magic
tech sky130A
timestamp 1616160187
<< nwell >>
rect 278 7469 1089 7619
rect 4103 7493 4914 7643
rect 1290 7288 2101 7438
rect 3090 7259 3901 7409
rect 277 7054 1088 7204
rect 4102 7078 4913 7228
rect 1345 6727 2156 6877
rect 3040 6839 3851 6989
rect 283 6488 1094 6638
rect 4108 6512 4919 6662
rect 1295 6307 2106 6457
rect 3095 6278 3906 6428
rect 282 6073 1093 6223
rect 4107 6097 4918 6247
rect 1510 5795 2321 5945
rect 2887 5811 3698 5961
rect 290 5509 1101 5659
rect 4115 5533 4926 5683
rect 1302 5328 2113 5478
rect 3102 5299 3913 5449
rect 289 5094 1100 5244
rect 4114 5118 4925 5268
rect 1357 4767 2168 4917
rect 3052 4879 3863 5029
rect 295 4528 1106 4678
rect 4120 4552 4931 4702
rect 1307 4347 2118 4497
rect 3107 4318 3918 4468
rect 294 4113 1105 4263
rect 4119 4137 4930 4287
rect 1605 3803 2416 3953
rect 2812 3886 3623 4036
rect 298 3552 1109 3702
rect 4123 3576 4934 3726
rect 1310 3371 2121 3521
rect 3110 3342 3921 3492
rect 297 3137 1108 3287
rect 4122 3161 4933 3311
rect 1365 2810 2176 2960
rect 3060 2922 3871 3072
rect 303 2571 1114 2721
rect 4128 2595 4939 2745
rect 1315 2390 2126 2540
rect 3115 2361 3926 2511
rect 302 2156 1113 2306
rect 4127 2180 4938 2330
rect 1530 1878 2341 2028
rect 2907 1894 3718 2044
rect 310 1592 1121 1742
rect 4135 1616 4946 1766
rect 1322 1411 2133 1561
rect 3122 1382 3933 1532
rect 309 1177 1120 1327
rect 4134 1201 4945 1351
rect 1377 850 2188 1000
rect 3072 962 3883 1112
rect 315 611 1126 761
rect 4140 635 4951 785
rect 1327 430 2138 580
rect 3127 401 3938 551
rect 314 196 1125 346
rect 4139 220 4950 370
rect 1717 -285 2528 -135
<< nmos >>
rect 4171 7702 4221 7744
rect 4379 7702 4429 7744
rect 4587 7702 4637 7744
rect 4800 7702 4850 7744
rect 3158 7468 3208 7510
rect 3366 7468 3416 7510
rect 3574 7468 3624 7510
rect 3787 7468 3837 7510
rect 342 7368 392 7410
rect 555 7368 605 7410
rect 763 7368 813 7410
rect 971 7368 1021 7410
rect 4170 7287 4220 7329
rect 4378 7287 4428 7329
rect 4586 7287 4636 7329
rect 4799 7287 4849 7329
rect 1354 7187 1404 7229
rect 1567 7187 1617 7229
rect 1775 7187 1825 7229
rect 1983 7187 2033 7229
rect 3108 7048 3158 7090
rect 3316 7048 3366 7090
rect 3524 7048 3574 7090
rect 3737 7048 3787 7090
rect 341 6953 391 6995
rect 554 6953 604 6995
rect 762 6953 812 6995
rect 970 6953 1020 6995
rect 4176 6721 4226 6763
rect 4384 6721 4434 6763
rect 4592 6721 4642 6763
rect 4805 6721 4855 6763
rect 1409 6626 1459 6668
rect 1622 6626 1672 6668
rect 1830 6626 1880 6668
rect 2038 6626 2088 6668
rect 3163 6487 3213 6529
rect 3371 6487 3421 6529
rect 3579 6487 3629 6529
rect 3792 6487 3842 6529
rect 347 6387 397 6429
rect 560 6387 610 6429
rect 768 6387 818 6429
rect 976 6387 1026 6429
rect 4175 6306 4225 6348
rect 4383 6306 4433 6348
rect 4591 6306 4641 6348
rect 4804 6306 4854 6348
rect 1359 6206 1409 6248
rect 1572 6206 1622 6248
rect 1780 6206 1830 6248
rect 1988 6206 2038 6248
rect 2955 6020 3005 6062
rect 3163 6020 3213 6062
rect 3371 6020 3421 6062
rect 3584 6020 3634 6062
rect 346 5972 396 6014
rect 559 5972 609 6014
rect 767 5972 817 6014
rect 975 5972 1025 6014
rect 4183 5742 4233 5784
rect 4391 5742 4441 5784
rect 4599 5742 4649 5784
rect 4812 5742 4862 5784
rect 1574 5694 1624 5736
rect 1787 5694 1837 5736
rect 1995 5694 2045 5736
rect 2203 5694 2253 5736
rect 3170 5508 3220 5550
rect 3378 5508 3428 5550
rect 3586 5508 3636 5550
rect 3799 5508 3849 5550
rect 354 5408 404 5450
rect 567 5408 617 5450
rect 775 5408 825 5450
rect 983 5408 1033 5450
rect 4182 5327 4232 5369
rect 4390 5327 4440 5369
rect 4598 5327 4648 5369
rect 4811 5327 4861 5369
rect 1366 5227 1416 5269
rect 1579 5227 1629 5269
rect 1787 5227 1837 5269
rect 1995 5227 2045 5269
rect 3120 5088 3170 5130
rect 3328 5088 3378 5130
rect 3536 5088 3586 5130
rect 3749 5088 3799 5130
rect 353 4993 403 5035
rect 566 4993 616 5035
rect 774 4993 824 5035
rect 982 4993 1032 5035
rect 4188 4761 4238 4803
rect 4396 4761 4446 4803
rect 4604 4761 4654 4803
rect 4817 4761 4867 4803
rect 1421 4666 1471 4708
rect 1634 4666 1684 4708
rect 1842 4666 1892 4708
rect 2050 4666 2100 4708
rect 3175 4527 3225 4569
rect 3383 4527 3433 4569
rect 3591 4527 3641 4569
rect 3804 4527 3854 4569
rect 359 4427 409 4469
rect 572 4427 622 4469
rect 780 4427 830 4469
rect 988 4427 1038 4469
rect 4187 4346 4237 4388
rect 4395 4346 4445 4388
rect 4603 4346 4653 4388
rect 4816 4346 4866 4388
rect 1371 4246 1421 4288
rect 1584 4246 1634 4288
rect 1792 4246 1842 4288
rect 2000 4246 2050 4288
rect 2880 4095 2930 4137
rect 3088 4095 3138 4137
rect 3296 4095 3346 4137
rect 3509 4095 3559 4137
rect 358 4012 408 4054
rect 571 4012 621 4054
rect 779 4012 829 4054
rect 987 4012 1037 4054
rect 4191 3785 4241 3827
rect 4399 3785 4449 3827
rect 4607 3785 4657 3827
rect 4820 3785 4870 3827
rect 1669 3702 1719 3744
rect 1882 3702 1932 3744
rect 2090 3702 2140 3744
rect 2298 3702 2348 3744
rect 3178 3551 3228 3593
rect 3386 3551 3436 3593
rect 3594 3551 3644 3593
rect 3807 3551 3857 3593
rect 362 3451 412 3493
rect 575 3451 625 3493
rect 783 3451 833 3493
rect 991 3451 1041 3493
rect 4190 3370 4240 3412
rect 4398 3370 4448 3412
rect 4606 3370 4656 3412
rect 4819 3370 4869 3412
rect 1374 3270 1424 3312
rect 1587 3270 1637 3312
rect 1795 3270 1845 3312
rect 2003 3270 2053 3312
rect 3128 3131 3178 3173
rect 3336 3131 3386 3173
rect 3544 3131 3594 3173
rect 3757 3131 3807 3173
rect 361 3036 411 3078
rect 574 3036 624 3078
rect 782 3036 832 3078
rect 990 3036 1040 3078
rect 4196 2804 4246 2846
rect 4404 2804 4454 2846
rect 4612 2804 4662 2846
rect 4825 2804 4875 2846
rect 1429 2709 1479 2751
rect 1642 2709 1692 2751
rect 1850 2709 1900 2751
rect 2058 2709 2108 2751
rect 3183 2570 3233 2612
rect 3391 2570 3441 2612
rect 3599 2570 3649 2612
rect 3812 2570 3862 2612
rect 367 2470 417 2512
rect 580 2470 630 2512
rect 788 2470 838 2512
rect 996 2470 1046 2512
rect 4195 2389 4245 2431
rect 4403 2389 4453 2431
rect 4611 2389 4661 2431
rect 4824 2389 4874 2431
rect 1379 2289 1429 2331
rect 1592 2289 1642 2331
rect 1800 2289 1850 2331
rect 2008 2289 2058 2331
rect 2975 2103 3025 2145
rect 3183 2103 3233 2145
rect 3391 2103 3441 2145
rect 3604 2103 3654 2145
rect 366 2055 416 2097
rect 579 2055 629 2097
rect 787 2055 837 2097
rect 995 2055 1045 2097
rect 4203 1825 4253 1867
rect 4411 1825 4461 1867
rect 4619 1825 4669 1867
rect 4832 1825 4882 1867
rect 1594 1777 1644 1819
rect 1807 1777 1857 1819
rect 2015 1777 2065 1819
rect 2223 1777 2273 1819
rect 3190 1591 3240 1633
rect 3398 1591 3448 1633
rect 3606 1591 3656 1633
rect 3819 1591 3869 1633
rect 374 1491 424 1533
rect 587 1491 637 1533
rect 795 1491 845 1533
rect 1003 1491 1053 1533
rect 4202 1410 4252 1452
rect 4410 1410 4460 1452
rect 4618 1410 4668 1452
rect 4831 1410 4881 1452
rect 1386 1310 1436 1352
rect 1599 1310 1649 1352
rect 1807 1310 1857 1352
rect 2015 1310 2065 1352
rect 3140 1171 3190 1213
rect 3348 1171 3398 1213
rect 3556 1171 3606 1213
rect 3769 1171 3819 1213
rect 373 1076 423 1118
rect 586 1076 636 1118
rect 794 1076 844 1118
rect 1002 1076 1052 1118
rect 4208 844 4258 886
rect 4416 844 4466 886
rect 4624 844 4674 886
rect 4837 844 4887 886
rect 1441 749 1491 791
rect 1654 749 1704 791
rect 1862 749 1912 791
rect 2070 749 2120 791
rect 3195 610 3245 652
rect 3403 610 3453 652
rect 3611 610 3661 652
rect 3824 610 3874 652
rect 379 510 429 552
rect 592 510 642 552
rect 800 510 850 552
rect 1008 510 1058 552
rect 4207 429 4257 471
rect 4415 429 4465 471
rect 4623 429 4673 471
rect 4836 429 4886 471
rect 1391 329 1441 371
rect 1604 329 1654 371
rect 1812 329 1862 371
rect 2020 329 2070 371
rect 378 95 428 137
rect 591 95 641 137
rect 799 95 849 137
rect 1007 95 1057 137
rect 1781 -386 1831 -344
rect 1994 -386 2044 -344
rect 2202 -386 2252 -344
rect 2410 -386 2460 -344
<< pmos >>
rect 342 7487 392 7587
rect 555 7487 605 7587
rect 763 7487 813 7587
rect 971 7487 1021 7587
rect 4171 7525 4221 7625
rect 4379 7525 4429 7625
rect 4587 7525 4637 7625
rect 4800 7525 4850 7625
rect 1354 7306 1404 7406
rect 1567 7306 1617 7406
rect 1775 7306 1825 7406
rect 1983 7306 2033 7406
rect 3158 7291 3208 7391
rect 3366 7291 3416 7391
rect 3574 7291 3624 7391
rect 3787 7291 3837 7391
rect 341 7072 391 7172
rect 554 7072 604 7172
rect 762 7072 812 7172
rect 970 7072 1020 7172
rect 4170 7110 4220 7210
rect 4378 7110 4428 7210
rect 4586 7110 4636 7210
rect 4799 7110 4849 7210
rect 3108 6871 3158 6971
rect 3316 6871 3366 6971
rect 3524 6871 3574 6971
rect 3737 6871 3787 6971
rect 1409 6745 1459 6845
rect 1622 6745 1672 6845
rect 1830 6745 1880 6845
rect 2038 6745 2088 6845
rect 347 6506 397 6606
rect 560 6506 610 6606
rect 768 6506 818 6606
rect 976 6506 1026 6606
rect 4176 6544 4226 6644
rect 4384 6544 4434 6644
rect 4592 6544 4642 6644
rect 4805 6544 4855 6644
rect 1359 6325 1409 6425
rect 1572 6325 1622 6425
rect 1780 6325 1830 6425
rect 1988 6325 2038 6425
rect 3163 6310 3213 6410
rect 3371 6310 3421 6410
rect 3579 6310 3629 6410
rect 3792 6310 3842 6410
rect 346 6091 396 6191
rect 559 6091 609 6191
rect 767 6091 817 6191
rect 975 6091 1025 6191
rect 4175 6129 4225 6229
rect 4383 6129 4433 6229
rect 4591 6129 4641 6229
rect 4804 6129 4854 6229
rect 1574 5813 1624 5913
rect 1787 5813 1837 5913
rect 1995 5813 2045 5913
rect 2203 5813 2253 5913
rect 2955 5843 3005 5943
rect 3163 5843 3213 5943
rect 3371 5843 3421 5943
rect 3584 5843 3634 5943
rect 354 5527 404 5627
rect 567 5527 617 5627
rect 775 5527 825 5627
rect 983 5527 1033 5627
rect 4183 5565 4233 5665
rect 4391 5565 4441 5665
rect 4599 5565 4649 5665
rect 4812 5565 4862 5665
rect 1366 5346 1416 5446
rect 1579 5346 1629 5446
rect 1787 5346 1837 5446
rect 1995 5346 2045 5446
rect 3170 5331 3220 5431
rect 3378 5331 3428 5431
rect 3586 5331 3636 5431
rect 3799 5331 3849 5431
rect 353 5112 403 5212
rect 566 5112 616 5212
rect 774 5112 824 5212
rect 982 5112 1032 5212
rect 4182 5150 4232 5250
rect 4390 5150 4440 5250
rect 4598 5150 4648 5250
rect 4811 5150 4861 5250
rect 3120 4911 3170 5011
rect 3328 4911 3378 5011
rect 3536 4911 3586 5011
rect 3749 4911 3799 5011
rect 1421 4785 1471 4885
rect 1634 4785 1684 4885
rect 1842 4785 1892 4885
rect 2050 4785 2100 4885
rect 359 4546 409 4646
rect 572 4546 622 4646
rect 780 4546 830 4646
rect 988 4546 1038 4646
rect 4188 4584 4238 4684
rect 4396 4584 4446 4684
rect 4604 4584 4654 4684
rect 4817 4584 4867 4684
rect 1371 4365 1421 4465
rect 1584 4365 1634 4465
rect 1792 4365 1842 4465
rect 2000 4365 2050 4465
rect 3175 4350 3225 4450
rect 3383 4350 3433 4450
rect 3591 4350 3641 4450
rect 3804 4350 3854 4450
rect 358 4131 408 4231
rect 571 4131 621 4231
rect 779 4131 829 4231
rect 987 4131 1037 4231
rect 4187 4169 4237 4269
rect 4395 4169 4445 4269
rect 4603 4169 4653 4269
rect 4816 4169 4866 4269
rect 1669 3821 1719 3921
rect 1882 3821 1932 3921
rect 2090 3821 2140 3921
rect 2298 3821 2348 3921
rect 2880 3918 2930 4018
rect 3088 3918 3138 4018
rect 3296 3918 3346 4018
rect 3509 3918 3559 4018
rect 362 3570 412 3670
rect 575 3570 625 3670
rect 783 3570 833 3670
rect 991 3570 1041 3670
rect 4191 3608 4241 3708
rect 4399 3608 4449 3708
rect 4607 3608 4657 3708
rect 4820 3608 4870 3708
rect 1374 3389 1424 3489
rect 1587 3389 1637 3489
rect 1795 3389 1845 3489
rect 2003 3389 2053 3489
rect 3178 3374 3228 3474
rect 3386 3374 3436 3474
rect 3594 3374 3644 3474
rect 3807 3374 3857 3474
rect 361 3155 411 3255
rect 574 3155 624 3255
rect 782 3155 832 3255
rect 990 3155 1040 3255
rect 4190 3193 4240 3293
rect 4398 3193 4448 3293
rect 4606 3193 4656 3293
rect 4819 3193 4869 3293
rect 3128 2954 3178 3054
rect 3336 2954 3386 3054
rect 3544 2954 3594 3054
rect 3757 2954 3807 3054
rect 1429 2828 1479 2928
rect 1642 2828 1692 2928
rect 1850 2828 1900 2928
rect 2058 2828 2108 2928
rect 367 2589 417 2689
rect 580 2589 630 2689
rect 788 2589 838 2689
rect 996 2589 1046 2689
rect 4196 2627 4246 2727
rect 4404 2627 4454 2727
rect 4612 2627 4662 2727
rect 4825 2627 4875 2727
rect 1379 2408 1429 2508
rect 1592 2408 1642 2508
rect 1800 2408 1850 2508
rect 2008 2408 2058 2508
rect 3183 2393 3233 2493
rect 3391 2393 3441 2493
rect 3599 2393 3649 2493
rect 3812 2393 3862 2493
rect 366 2174 416 2274
rect 579 2174 629 2274
rect 787 2174 837 2274
rect 995 2174 1045 2274
rect 4195 2212 4245 2312
rect 4403 2212 4453 2312
rect 4611 2212 4661 2312
rect 4824 2212 4874 2312
rect 1594 1896 1644 1996
rect 1807 1896 1857 1996
rect 2015 1896 2065 1996
rect 2223 1896 2273 1996
rect 2975 1926 3025 2026
rect 3183 1926 3233 2026
rect 3391 1926 3441 2026
rect 3604 1926 3654 2026
rect 374 1610 424 1710
rect 587 1610 637 1710
rect 795 1610 845 1710
rect 1003 1610 1053 1710
rect 4203 1648 4253 1748
rect 4411 1648 4461 1748
rect 4619 1648 4669 1748
rect 4832 1648 4882 1748
rect 1386 1429 1436 1529
rect 1599 1429 1649 1529
rect 1807 1429 1857 1529
rect 2015 1429 2065 1529
rect 3190 1414 3240 1514
rect 3398 1414 3448 1514
rect 3606 1414 3656 1514
rect 3819 1414 3869 1514
rect 373 1195 423 1295
rect 586 1195 636 1295
rect 794 1195 844 1295
rect 1002 1195 1052 1295
rect 4202 1233 4252 1333
rect 4410 1233 4460 1333
rect 4618 1233 4668 1333
rect 4831 1233 4881 1333
rect 3140 994 3190 1094
rect 3348 994 3398 1094
rect 3556 994 3606 1094
rect 3769 994 3819 1094
rect 1441 868 1491 968
rect 1654 868 1704 968
rect 1862 868 1912 968
rect 2070 868 2120 968
rect 379 629 429 729
rect 592 629 642 729
rect 800 629 850 729
rect 1008 629 1058 729
rect 4208 667 4258 767
rect 4416 667 4466 767
rect 4624 667 4674 767
rect 4837 667 4887 767
rect 1391 448 1441 548
rect 1604 448 1654 548
rect 1812 448 1862 548
rect 2020 448 2070 548
rect 3195 433 3245 533
rect 3403 433 3453 533
rect 3611 433 3661 533
rect 3824 433 3874 533
rect 378 214 428 314
rect 591 214 641 314
rect 799 214 849 314
rect 1007 214 1057 314
rect 4207 252 4257 352
rect 4415 252 4465 352
rect 4623 252 4673 352
rect 4836 252 4886 352
rect 1781 -267 1831 -167
rect 1994 -267 2044 -167
rect 2202 -267 2252 -167
rect 2410 -267 2460 -167
<< ndiff >>
rect 4122 7732 4171 7744
rect 4122 7712 4133 7732
rect 4153 7712 4171 7732
rect 4122 7702 4171 7712
rect 4221 7728 4265 7744
rect 4221 7708 4236 7728
rect 4256 7708 4265 7728
rect 4221 7702 4265 7708
rect 4335 7728 4379 7744
rect 4335 7708 4344 7728
rect 4364 7708 4379 7728
rect 4335 7702 4379 7708
rect 4429 7732 4478 7744
rect 4429 7712 4447 7732
rect 4467 7712 4478 7732
rect 4429 7702 4478 7712
rect 4543 7728 4587 7744
rect 4543 7708 4552 7728
rect 4572 7708 4587 7728
rect 4543 7702 4587 7708
rect 4637 7732 4686 7744
rect 4637 7712 4655 7732
rect 4675 7712 4686 7732
rect 4637 7702 4686 7712
rect 4756 7728 4800 7744
rect 4756 7708 4765 7728
rect 4785 7708 4800 7728
rect 4756 7702 4800 7708
rect 4850 7732 4899 7744
rect 4850 7712 4868 7732
rect 4888 7712 4899 7732
rect 4850 7702 4899 7712
rect 3109 7498 3158 7510
rect 3109 7478 3120 7498
rect 3140 7478 3158 7498
rect 3109 7468 3158 7478
rect 3208 7494 3252 7510
rect 3208 7474 3223 7494
rect 3243 7474 3252 7494
rect 3208 7468 3252 7474
rect 3322 7494 3366 7510
rect 3322 7474 3331 7494
rect 3351 7474 3366 7494
rect 3322 7468 3366 7474
rect 3416 7498 3465 7510
rect 3416 7478 3434 7498
rect 3454 7478 3465 7498
rect 3416 7468 3465 7478
rect 3530 7494 3574 7510
rect 3530 7474 3539 7494
rect 3559 7474 3574 7494
rect 3530 7468 3574 7474
rect 3624 7498 3673 7510
rect 3624 7478 3642 7498
rect 3662 7478 3673 7498
rect 3624 7468 3673 7478
rect 3743 7494 3787 7510
rect 3743 7474 3752 7494
rect 3772 7474 3787 7494
rect 3743 7468 3787 7474
rect 3837 7498 3886 7510
rect 3837 7478 3855 7498
rect 3875 7478 3886 7498
rect 3837 7468 3886 7478
rect 293 7400 342 7410
rect 293 7380 304 7400
rect 324 7380 342 7400
rect 293 7368 342 7380
rect 392 7404 436 7410
rect 392 7384 407 7404
rect 427 7384 436 7404
rect 392 7368 436 7384
rect 506 7400 555 7410
rect 506 7380 517 7400
rect 537 7380 555 7400
rect 506 7368 555 7380
rect 605 7404 649 7410
rect 605 7384 620 7404
rect 640 7384 649 7404
rect 605 7368 649 7384
rect 714 7400 763 7410
rect 714 7380 725 7400
rect 745 7380 763 7400
rect 714 7368 763 7380
rect 813 7404 857 7410
rect 813 7384 828 7404
rect 848 7384 857 7404
rect 813 7368 857 7384
rect 927 7404 971 7410
rect 927 7384 936 7404
rect 956 7384 971 7404
rect 927 7368 971 7384
rect 1021 7400 1070 7410
rect 1021 7380 1039 7400
rect 1059 7380 1070 7400
rect 1021 7368 1070 7380
rect 4121 7317 4170 7329
rect 4121 7297 4132 7317
rect 4152 7297 4170 7317
rect 4121 7287 4170 7297
rect 4220 7313 4264 7329
rect 4220 7293 4235 7313
rect 4255 7293 4264 7313
rect 4220 7287 4264 7293
rect 4334 7313 4378 7329
rect 4334 7293 4343 7313
rect 4363 7293 4378 7313
rect 4334 7287 4378 7293
rect 4428 7317 4477 7329
rect 4428 7297 4446 7317
rect 4466 7297 4477 7317
rect 4428 7287 4477 7297
rect 4542 7313 4586 7329
rect 4542 7293 4551 7313
rect 4571 7293 4586 7313
rect 4542 7287 4586 7293
rect 4636 7317 4685 7329
rect 4636 7297 4654 7317
rect 4674 7297 4685 7317
rect 4636 7287 4685 7297
rect 4755 7313 4799 7329
rect 4755 7293 4764 7313
rect 4784 7293 4799 7313
rect 4755 7287 4799 7293
rect 4849 7317 4898 7329
rect 4849 7297 4867 7317
rect 4887 7297 4898 7317
rect 4849 7287 4898 7297
rect 1305 7219 1354 7229
rect 1305 7199 1316 7219
rect 1336 7199 1354 7219
rect 1305 7187 1354 7199
rect 1404 7223 1448 7229
rect 1404 7203 1419 7223
rect 1439 7203 1448 7223
rect 1404 7187 1448 7203
rect 1518 7219 1567 7229
rect 1518 7199 1529 7219
rect 1549 7199 1567 7219
rect 1518 7187 1567 7199
rect 1617 7223 1661 7229
rect 1617 7203 1632 7223
rect 1652 7203 1661 7223
rect 1617 7187 1661 7203
rect 1726 7219 1775 7229
rect 1726 7199 1737 7219
rect 1757 7199 1775 7219
rect 1726 7187 1775 7199
rect 1825 7223 1869 7229
rect 1825 7203 1840 7223
rect 1860 7203 1869 7223
rect 1825 7187 1869 7203
rect 1939 7223 1983 7229
rect 1939 7203 1948 7223
rect 1968 7203 1983 7223
rect 1939 7187 1983 7203
rect 2033 7219 2082 7229
rect 2033 7199 2051 7219
rect 2071 7199 2082 7219
rect 2033 7187 2082 7199
rect 3059 7078 3108 7090
rect 3059 7058 3070 7078
rect 3090 7058 3108 7078
rect 3059 7048 3108 7058
rect 3158 7074 3202 7090
rect 3158 7054 3173 7074
rect 3193 7054 3202 7074
rect 3158 7048 3202 7054
rect 3272 7074 3316 7090
rect 3272 7054 3281 7074
rect 3301 7054 3316 7074
rect 3272 7048 3316 7054
rect 3366 7078 3415 7090
rect 3366 7058 3384 7078
rect 3404 7058 3415 7078
rect 3366 7048 3415 7058
rect 3480 7074 3524 7090
rect 3480 7054 3489 7074
rect 3509 7054 3524 7074
rect 3480 7048 3524 7054
rect 3574 7078 3623 7090
rect 3574 7058 3592 7078
rect 3612 7058 3623 7078
rect 3574 7048 3623 7058
rect 3693 7074 3737 7090
rect 3693 7054 3702 7074
rect 3722 7054 3737 7074
rect 3693 7048 3737 7054
rect 3787 7078 3836 7090
rect 3787 7058 3805 7078
rect 3825 7058 3836 7078
rect 3787 7048 3836 7058
rect 292 6985 341 6995
rect 292 6965 303 6985
rect 323 6965 341 6985
rect 292 6953 341 6965
rect 391 6989 435 6995
rect 391 6969 406 6989
rect 426 6969 435 6989
rect 391 6953 435 6969
rect 505 6985 554 6995
rect 505 6965 516 6985
rect 536 6965 554 6985
rect 505 6953 554 6965
rect 604 6989 648 6995
rect 604 6969 619 6989
rect 639 6969 648 6989
rect 604 6953 648 6969
rect 713 6985 762 6995
rect 713 6965 724 6985
rect 744 6965 762 6985
rect 713 6953 762 6965
rect 812 6989 856 6995
rect 812 6969 827 6989
rect 847 6969 856 6989
rect 812 6953 856 6969
rect 926 6989 970 6995
rect 926 6969 935 6989
rect 955 6969 970 6989
rect 926 6953 970 6969
rect 1020 6985 1069 6995
rect 1020 6965 1038 6985
rect 1058 6965 1069 6985
rect 1020 6953 1069 6965
rect 4127 6751 4176 6763
rect 4127 6731 4138 6751
rect 4158 6731 4176 6751
rect 4127 6721 4176 6731
rect 4226 6747 4270 6763
rect 4226 6727 4241 6747
rect 4261 6727 4270 6747
rect 4226 6721 4270 6727
rect 4340 6747 4384 6763
rect 4340 6727 4349 6747
rect 4369 6727 4384 6747
rect 4340 6721 4384 6727
rect 4434 6751 4483 6763
rect 4434 6731 4452 6751
rect 4472 6731 4483 6751
rect 4434 6721 4483 6731
rect 4548 6747 4592 6763
rect 4548 6727 4557 6747
rect 4577 6727 4592 6747
rect 4548 6721 4592 6727
rect 4642 6751 4691 6763
rect 4642 6731 4660 6751
rect 4680 6731 4691 6751
rect 4642 6721 4691 6731
rect 4761 6747 4805 6763
rect 4761 6727 4770 6747
rect 4790 6727 4805 6747
rect 4761 6721 4805 6727
rect 4855 6751 4904 6763
rect 4855 6731 4873 6751
rect 4893 6731 4904 6751
rect 4855 6721 4904 6731
rect 1360 6658 1409 6668
rect 1360 6638 1371 6658
rect 1391 6638 1409 6658
rect 1360 6626 1409 6638
rect 1459 6662 1503 6668
rect 1459 6642 1474 6662
rect 1494 6642 1503 6662
rect 1459 6626 1503 6642
rect 1573 6658 1622 6668
rect 1573 6638 1584 6658
rect 1604 6638 1622 6658
rect 1573 6626 1622 6638
rect 1672 6662 1716 6668
rect 1672 6642 1687 6662
rect 1707 6642 1716 6662
rect 1672 6626 1716 6642
rect 1781 6658 1830 6668
rect 1781 6638 1792 6658
rect 1812 6638 1830 6658
rect 1781 6626 1830 6638
rect 1880 6662 1924 6668
rect 1880 6642 1895 6662
rect 1915 6642 1924 6662
rect 1880 6626 1924 6642
rect 1994 6662 2038 6668
rect 1994 6642 2003 6662
rect 2023 6642 2038 6662
rect 1994 6626 2038 6642
rect 2088 6658 2137 6668
rect 2088 6638 2106 6658
rect 2126 6638 2137 6658
rect 2088 6626 2137 6638
rect 3114 6517 3163 6529
rect 3114 6497 3125 6517
rect 3145 6497 3163 6517
rect 3114 6487 3163 6497
rect 3213 6513 3257 6529
rect 3213 6493 3228 6513
rect 3248 6493 3257 6513
rect 3213 6487 3257 6493
rect 3327 6513 3371 6529
rect 3327 6493 3336 6513
rect 3356 6493 3371 6513
rect 3327 6487 3371 6493
rect 3421 6517 3470 6529
rect 3421 6497 3439 6517
rect 3459 6497 3470 6517
rect 3421 6487 3470 6497
rect 3535 6513 3579 6529
rect 3535 6493 3544 6513
rect 3564 6493 3579 6513
rect 3535 6487 3579 6493
rect 3629 6517 3678 6529
rect 3629 6497 3647 6517
rect 3667 6497 3678 6517
rect 3629 6487 3678 6497
rect 3748 6513 3792 6529
rect 3748 6493 3757 6513
rect 3777 6493 3792 6513
rect 3748 6487 3792 6493
rect 3842 6517 3891 6529
rect 3842 6497 3860 6517
rect 3880 6497 3891 6517
rect 3842 6487 3891 6497
rect 298 6419 347 6429
rect 298 6399 309 6419
rect 329 6399 347 6419
rect 298 6387 347 6399
rect 397 6423 441 6429
rect 397 6403 412 6423
rect 432 6403 441 6423
rect 397 6387 441 6403
rect 511 6419 560 6429
rect 511 6399 522 6419
rect 542 6399 560 6419
rect 511 6387 560 6399
rect 610 6423 654 6429
rect 610 6403 625 6423
rect 645 6403 654 6423
rect 610 6387 654 6403
rect 719 6419 768 6429
rect 719 6399 730 6419
rect 750 6399 768 6419
rect 719 6387 768 6399
rect 818 6423 862 6429
rect 818 6403 833 6423
rect 853 6403 862 6423
rect 818 6387 862 6403
rect 932 6423 976 6429
rect 932 6403 941 6423
rect 961 6403 976 6423
rect 932 6387 976 6403
rect 1026 6419 1075 6429
rect 1026 6399 1044 6419
rect 1064 6399 1075 6419
rect 1026 6387 1075 6399
rect 4126 6336 4175 6348
rect 4126 6316 4137 6336
rect 4157 6316 4175 6336
rect 4126 6306 4175 6316
rect 4225 6332 4269 6348
rect 4225 6312 4240 6332
rect 4260 6312 4269 6332
rect 4225 6306 4269 6312
rect 4339 6332 4383 6348
rect 4339 6312 4348 6332
rect 4368 6312 4383 6332
rect 4339 6306 4383 6312
rect 4433 6336 4482 6348
rect 4433 6316 4451 6336
rect 4471 6316 4482 6336
rect 4433 6306 4482 6316
rect 4547 6332 4591 6348
rect 4547 6312 4556 6332
rect 4576 6312 4591 6332
rect 4547 6306 4591 6312
rect 4641 6336 4690 6348
rect 4641 6316 4659 6336
rect 4679 6316 4690 6336
rect 4641 6306 4690 6316
rect 4760 6332 4804 6348
rect 4760 6312 4769 6332
rect 4789 6312 4804 6332
rect 4760 6306 4804 6312
rect 4854 6336 4903 6348
rect 4854 6316 4872 6336
rect 4892 6316 4903 6336
rect 4854 6306 4903 6316
rect 1310 6238 1359 6248
rect 1310 6218 1321 6238
rect 1341 6218 1359 6238
rect 1310 6206 1359 6218
rect 1409 6242 1453 6248
rect 1409 6222 1424 6242
rect 1444 6222 1453 6242
rect 1409 6206 1453 6222
rect 1523 6238 1572 6248
rect 1523 6218 1534 6238
rect 1554 6218 1572 6238
rect 1523 6206 1572 6218
rect 1622 6242 1666 6248
rect 1622 6222 1637 6242
rect 1657 6222 1666 6242
rect 1622 6206 1666 6222
rect 1731 6238 1780 6248
rect 1731 6218 1742 6238
rect 1762 6218 1780 6238
rect 1731 6206 1780 6218
rect 1830 6242 1874 6248
rect 1830 6222 1845 6242
rect 1865 6222 1874 6242
rect 1830 6206 1874 6222
rect 1944 6242 1988 6248
rect 1944 6222 1953 6242
rect 1973 6222 1988 6242
rect 1944 6206 1988 6222
rect 2038 6238 2087 6248
rect 2038 6218 2056 6238
rect 2076 6218 2087 6238
rect 2038 6206 2087 6218
rect 2906 6050 2955 6062
rect 2906 6030 2917 6050
rect 2937 6030 2955 6050
rect 2906 6020 2955 6030
rect 3005 6046 3049 6062
rect 3005 6026 3020 6046
rect 3040 6026 3049 6046
rect 3005 6020 3049 6026
rect 3119 6046 3163 6062
rect 3119 6026 3128 6046
rect 3148 6026 3163 6046
rect 3119 6020 3163 6026
rect 3213 6050 3262 6062
rect 3213 6030 3231 6050
rect 3251 6030 3262 6050
rect 3213 6020 3262 6030
rect 3327 6046 3371 6062
rect 3327 6026 3336 6046
rect 3356 6026 3371 6046
rect 3327 6020 3371 6026
rect 3421 6050 3470 6062
rect 3421 6030 3439 6050
rect 3459 6030 3470 6050
rect 3421 6020 3470 6030
rect 3540 6046 3584 6062
rect 3540 6026 3549 6046
rect 3569 6026 3584 6046
rect 3540 6020 3584 6026
rect 3634 6050 3683 6062
rect 3634 6030 3652 6050
rect 3672 6030 3683 6050
rect 3634 6020 3683 6030
rect 297 6004 346 6014
rect 297 5984 308 6004
rect 328 5984 346 6004
rect 297 5972 346 5984
rect 396 6008 440 6014
rect 396 5988 411 6008
rect 431 5988 440 6008
rect 396 5972 440 5988
rect 510 6004 559 6014
rect 510 5984 521 6004
rect 541 5984 559 6004
rect 510 5972 559 5984
rect 609 6008 653 6014
rect 609 5988 624 6008
rect 644 5988 653 6008
rect 609 5972 653 5988
rect 718 6004 767 6014
rect 718 5984 729 6004
rect 749 5984 767 6004
rect 718 5972 767 5984
rect 817 6008 861 6014
rect 817 5988 832 6008
rect 852 5988 861 6008
rect 817 5972 861 5988
rect 931 6008 975 6014
rect 931 5988 940 6008
rect 960 5988 975 6008
rect 931 5972 975 5988
rect 1025 6004 1074 6014
rect 1025 5984 1043 6004
rect 1063 5984 1074 6004
rect 1025 5972 1074 5984
rect 4134 5772 4183 5784
rect 4134 5752 4145 5772
rect 4165 5752 4183 5772
rect 4134 5742 4183 5752
rect 4233 5768 4277 5784
rect 4233 5748 4248 5768
rect 4268 5748 4277 5768
rect 4233 5742 4277 5748
rect 4347 5768 4391 5784
rect 4347 5748 4356 5768
rect 4376 5748 4391 5768
rect 4347 5742 4391 5748
rect 4441 5772 4490 5784
rect 4441 5752 4459 5772
rect 4479 5752 4490 5772
rect 4441 5742 4490 5752
rect 4555 5768 4599 5784
rect 4555 5748 4564 5768
rect 4584 5748 4599 5768
rect 4555 5742 4599 5748
rect 4649 5772 4698 5784
rect 4649 5752 4667 5772
rect 4687 5752 4698 5772
rect 4649 5742 4698 5752
rect 4768 5768 4812 5784
rect 4768 5748 4777 5768
rect 4797 5748 4812 5768
rect 4768 5742 4812 5748
rect 4862 5772 4911 5784
rect 4862 5752 4880 5772
rect 4900 5752 4911 5772
rect 4862 5742 4911 5752
rect 1525 5726 1574 5736
rect 1525 5706 1536 5726
rect 1556 5706 1574 5726
rect 1525 5694 1574 5706
rect 1624 5730 1668 5736
rect 1624 5710 1639 5730
rect 1659 5710 1668 5730
rect 1624 5694 1668 5710
rect 1738 5726 1787 5736
rect 1738 5706 1749 5726
rect 1769 5706 1787 5726
rect 1738 5694 1787 5706
rect 1837 5730 1881 5736
rect 1837 5710 1852 5730
rect 1872 5710 1881 5730
rect 1837 5694 1881 5710
rect 1946 5726 1995 5736
rect 1946 5706 1957 5726
rect 1977 5706 1995 5726
rect 1946 5694 1995 5706
rect 2045 5730 2089 5736
rect 2045 5710 2060 5730
rect 2080 5710 2089 5730
rect 2045 5694 2089 5710
rect 2159 5730 2203 5736
rect 2159 5710 2168 5730
rect 2188 5710 2203 5730
rect 2159 5694 2203 5710
rect 2253 5726 2302 5736
rect 2253 5706 2271 5726
rect 2291 5706 2302 5726
rect 2253 5694 2302 5706
rect 3121 5538 3170 5550
rect 3121 5518 3132 5538
rect 3152 5518 3170 5538
rect 3121 5508 3170 5518
rect 3220 5534 3264 5550
rect 3220 5514 3235 5534
rect 3255 5514 3264 5534
rect 3220 5508 3264 5514
rect 3334 5534 3378 5550
rect 3334 5514 3343 5534
rect 3363 5514 3378 5534
rect 3334 5508 3378 5514
rect 3428 5538 3477 5550
rect 3428 5518 3446 5538
rect 3466 5518 3477 5538
rect 3428 5508 3477 5518
rect 3542 5534 3586 5550
rect 3542 5514 3551 5534
rect 3571 5514 3586 5534
rect 3542 5508 3586 5514
rect 3636 5538 3685 5550
rect 3636 5518 3654 5538
rect 3674 5518 3685 5538
rect 3636 5508 3685 5518
rect 3755 5534 3799 5550
rect 3755 5514 3764 5534
rect 3784 5514 3799 5534
rect 3755 5508 3799 5514
rect 3849 5538 3898 5550
rect 3849 5518 3867 5538
rect 3887 5518 3898 5538
rect 3849 5508 3898 5518
rect 305 5440 354 5450
rect 305 5420 316 5440
rect 336 5420 354 5440
rect 305 5408 354 5420
rect 404 5444 448 5450
rect 404 5424 419 5444
rect 439 5424 448 5444
rect 404 5408 448 5424
rect 518 5440 567 5450
rect 518 5420 529 5440
rect 549 5420 567 5440
rect 518 5408 567 5420
rect 617 5444 661 5450
rect 617 5424 632 5444
rect 652 5424 661 5444
rect 617 5408 661 5424
rect 726 5440 775 5450
rect 726 5420 737 5440
rect 757 5420 775 5440
rect 726 5408 775 5420
rect 825 5444 869 5450
rect 825 5424 840 5444
rect 860 5424 869 5444
rect 825 5408 869 5424
rect 939 5444 983 5450
rect 939 5424 948 5444
rect 968 5424 983 5444
rect 939 5408 983 5424
rect 1033 5440 1082 5450
rect 1033 5420 1051 5440
rect 1071 5420 1082 5440
rect 1033 5408 1082 5420
rect 4133 5357 4182 5369
rect 4133 5337 4144 5357
rect 4164 5337 4182 5357
rect 4133 5327 4182 5337
rect 4232 5353 4276 5369
rect 4232 5333 4247 5353
rect 4267 5333 4276 5353
rect 4232 5327 4276 5333
rect 4346 5353 4390 5369
rect 4346 5333 4355 5353
rect 4375 5333 4390 5353
rect 4346 5327 4390 5333
rect 4440 5357 4489 5369
rect 4440 5337 4458 5357
rect 4478 5337 4489 5357
rect 4440 5327 4489 5337
rect 4554 5353 4598 5369
rect 4554 5333 4563 5353
rect 4583 5333 4598 5353
rect 4554 5327 4598 5333
rect 4648 5357 4697 5369
rect 4648 5337 4666 5357
rect 4686 5337 4697 5357
rect 4648 5327 4697 5337
rect 4767 5353 4811 5369
rect 4767 5333 4776 5353
rect 4796 5333 4811 5353
rect 4767 5327 4811 5333
rect 4861 5357 4910 5369
rect 4861 5337 4879 5357
rect 4899 5337 4910 5357
rect 4861 5327 4910 5337
rect 1317 5259 1366 5269
rect 1317 5239 1328 5259
rect 1348 5239 1366 5259
rect 1317 5227 1366 5239
rect 1416 5263 1460 5269
rect 1416 5243 1431 5263
rect 1451 5243 1460 5263
rect 1416 5227 1460 5243
rect 1530 5259 1579 5269
rect 1530 5239 1541 5259
rect 1561 5239 1579 5259
rect 1530 5227 1579 5239
rect 1629 5263 1673 5269
rect 1629 5243 1644 5263
rect 1664 5243 1673 5263
rect 1629 5227 1673 5243
rect 1738 5259 1787 5269
rect 1738 5239 1749 5259
rect 1769 5239 1787 5259
rect 1738 5227 1787 5239
rect 1837 5263 1881 5269
rect 1837 5243 1852 5263
rect 1872 5243 1881 5263
rect 1837 5227 1881 5243
rect 1951 5263 1995 5269
rect 1951 5243 1960 5263
rect 1980 5243 1995 5263
rect 1951 5227 1995 5243
rect 2045 5259 2094 5269
rect 2045 5239 2063 5259
rect 2083 5239 2094 5259
rect 2045 5227 2094 5239
rect 3071 5118 3120 5130
rect 3071 5098 3082 5118
rect 3102 5098 3120 5118
rect 3071 5088 3120 5098
rect 3170 5114 3214 5130
rect 3170 5094 3185 5114
rect 3205 5094 3214 5114
rect 3170 5088 3214 5094
rect 3284 5114 3328 5130
rect 3284 5094 3293 5114
rect 3313 5094 3328 5114
rect 3284 5088 3328 5094
rect 3378 5118 3427 5130
rect 3378 5098 3396 5118
rect 3416 5098 3427 5118
rect 3378 5088 3427 5098
rect 3492 5114 3536 5130
rect 3492 5094 3501 5114
rect 3521 5094 3536 5114
rect 3492 5088 3536 5094
rect 3586 5118 3635 5130
rect 3586 5098 3604 5118
rect 3624 5098 3635 5118
rect 3586 5088 3635 5098
rect 3705 5114 3749 5130
rect 3705 5094 3714 5114
rect 3734 5094 3749 5114
rect 3705 5088 3749 5094
rect 3799 5118 3848 5130
rect 3799 5098 3817 5118
rect 3837 5098 3848 5118
rect 3799 5088 3848 5098
rect 304 5025 353 5035
rect 304 5005 315 5025
rect 335 5005 353 5025
rect 304 4993 353 5005
rect 403 5029 447 5035
rect 403 5009 418 5029
rect 438 5009 447 5029
rect 403 4993 447 5009
rect 517 5025 566 5035
rect 517 5005 528 5025
rect 548 5005 566 5025
rect 517 4993 566 5005
rect 616 5029 660 5035
rect 616 5009 631 5029
rect 651 5009 660 5029
rect 616 4993 660 5009
rect 725 5025 774 5035
rect 725 5005 736 5025
rect 756 5005 774 5025
rect 725 4993 774 5005
rect 824 5029 868 5035
rect 824 5009 839 5029
rect 859 5009 868 5029
rect 824 4993 868 5009
rect 938 5029 982 5035
rect 938 5009 947 5029
rect 967 5009 982 5029
rect 938 4993 982 5009
rect 1032 5025 1081 5035
rect 1032 5005 1050 5025
rect 1070 5005 1081 5025
rect 1032 4993 1081 5005
rect 4139 4791 4188 4803
rect 4139 4771 4150 4791
rect 4170 4771 4188 4791
rect 4139 4761 4188 4771
rect 4238 4787 4282 4803
rect 4238 4767 4253 4787
rect 4273 4767 4282 4787
rect 4238 4761 4282 4767
rect 4352 4787 4396 4803
rect 4352 4767 4361 4787
rect 4381 4767 4396 4787
rect 4352 4761 4396 4767
rect 4446 4791 4495 4803
rect 4446 4771 4464 4791
rect 4484 4771 4495 4791
rect 4446 4761 4495 4771
rect 4560 4787 4604 4803
rect 4560 4767 4569 4787
rect 4589 4767 4604 4787
rect 4560 4761 4604 4767
rect 4654 4791 4703 4803
rect 4654 4771 4672 4791
rect 4692 4771 4703 4791
rect 4654 4761 4703 4771
rect 4773 4787 4817 4803
rect 4773 4767 4782 4787
rect 4802 4767 4817 4787
rect 4773 4761 4817 4767
rect 4867 4791 4916 4803
rect 4867 4771 4885 4791
rect 4905 4771 4916 4791
rect 4867 4761 4916 4771
rect 1372 4698 1421 4708
rect 1372 4678 1383 4698
rect 1403 4678 1421 4698
rect 1372 4666 1421 4678
rect 1471 4702 1515 4708
rect 1471 4682 1486 4702
rect 1506 4682 1515 4702
rect 1471 4666 1515 4682
rect 1585 4698 1634 4708
rect 1585 4678 1596 4698
rect 1616 4678 1634 4698
rect 1585 4666 1634 4678
rect 1684 4702 1728 4708
rect 1684 4682 1699 4702
rect 1719 4682 1728 4702
rect 1684 4666 1728 4682
rect 1793 4698 1842 4708
rect 1793 4678 1804 4698
rect 1824 4678 1842 4698
rect 1793 4666 1842 4678
rect 1892 4702 1936 4708
rect 1892 4682 1907 4702
rect 1927 4682 1936 4702
rect 1892 4666 1936 4682
rect 2006 4702 2050 4708
rect 2006 4682 2015 4702
rect 2035 4682 2050 4702
rect 2006 4666 2050 4682
rect 2100 4698 2149 4708
rect 2100 4678 2118 4698
rect 2138 4678 2149 4698
rect 2100 4666 2149 4678
rect 3126 4557 3175 4569
rect 3126 4537 3137 4557
rect 3157 4537 3175 4557
rect 3126 4527 3175 4537
rect 3225 4553 3269 4569
rect 3225 4533 3240 4553
rect 3260 4533 3269 4553
rect 3225 4527 3269 4533
rect 3339 4553 3383 4569
rect 3339 4533 3348 4553
rect 3368 4533 3383 4553
rect 3339 4527 3383 4533
rect 3433 4557 3482 4569
rect 3433 4537 3451 4557
rect 3471 4537 3482 4557
rect 3433 4527 3482 4537
rect 3547 4553 3591 4569
rect 3547 4533 3556 4553
rect 3576 4533 3591 4553
rect 3547 4527 3591 4533
rect 3641 4557 3690 4569
rect 3641 4537 3659 4557
rect 3679 4537 3690 4557
rect 3641 4527 3690 4537
rect 3760 4553 3804 4569
rect 3760 4533 3769 4553
rect 3789 4533 3804 4553
rect 3760 4527 3804 4533
rect 3854 4557 3903 4569
rect 3854 4537 3872 4557
rect 3892 4537 3903 4557
rect 3854 4527 3903 4537
rect 310 4459 359 4469
rect 310 4439 321 4459
rect 341 4439 359 4459
rect 310 4427 359 4439
rect 409 4463 453 4469
rect 409 4443 424 4463
rect 444 4443 453 4463
rect 409 4427 453 4443
rect 523 4459 572 4469
rect 523 4439 534 4459
rect 554 4439 572 4459
rect 523 4427 572 4439
rect 622 4463 666 4469
rect 622 4443 637 4463
rect 657 4443 666 4463
rect 622 4427 666 4443
rect 731 4459 780 4469
rect 731 4439 742 4459
rect 762 4439 780 4459
rect 731 4427 780 4439
rect 830 4463 874 4469
rect 830 4443 845 4463
rect 865 4443 874 4463
rect 830 4427 874 4443
rect 944 4463 988 4469
rect 944 4443 953 4463
rect 973 4443 988 4463
rect 944 4427 988 4443
rect 1038 4459 1087 4469
rect 1038 4439 1056 4459
rect 1076 4439 1087 4459
rect 1038 4427 1087 4439
rect 4138 4376 4187 4388
rect 4138 4356 4149 4376
rect 4169 4356 4187 4376
rect 4138 4346 4187 4356
rect 4237 4372 4281 4388
rect 4237 4352 4252 4372
rect 4272 4352 4281 4372
rect 4237 4346 4281 4352
rect 4351 4372 4395 4388
rect 4351 4352 4360 4372
rect 4380 4352 4395 4372
rect 4351 4346 4395 4352
rect 4445 4376 4494 4388
rect 4445 4356 4463 4376
rect 4483 4356 4494 4376
rect 4445 4346 4494 4356
rect 4559 4372 4603 4388
rect 4559 4352 4568 4372
rect 4588 4352 4603 4372
rect 4559 4346 4603 4352
rect 4653 4376 4702 4388
rect 4653 4356 4671 4376
rect 4691 4356 4702 4376
rect 4653 4346 4702 4356
rect 4772 4372 4816 4388
rect 4772 4352 4781 4372
rect 4801 4352 4816 4372
rect 4772 4346 4816 4352
rect 4866 4376 4915 4388
rect 4866 4356 4884 4376
rect 4904 4356 4915 4376
rect 4866 4346 4915 4356
rect 1322 4278 1371 4288
rect 1322 4258 1333 4278
rect 1353 4258 1371 4278
rect 1322 4246 1371 4258
rect 1421 4282 1465 4288
rect 1421 4262 1436 4282
rect 1456 4262 1465 4282
rect 1421 4246 1465 4262
rect 1535 4278 1584 4288
rect 1535 4258 1546 4278
rect 1566 4258 1584 4278
rect 1535 4246 1584 4258
rect 1634 4282 1678 4288
rect 1634 4262 1649 4282
rect 1669 4262 1678 4282
rect 1634 4246 1678 4262
rect 1743 4278 1792 4288
rect 1743 4258 1754 4278
rect 1774 4258 1792 4278
rect 1743 4246 1792 4258
rect 1842 4282 1886 4288
rect 1842 4262 1857 4282
rect 1877 4262 1886 4282
rect 1842 4246 1886 4262
rect 1956 4282 2000 4288
rect 1956 4262 1965 4282
rect 1985 4262 2000 4282
rect 1956 4246 2000 4262
rect 2050 4278 2099 4288
rect 2050 4258 2068 4278
rect 2088 4258 2099 4278
rect 2050 4246 2099 4258
rect 2831 4125 2880 4137
rect 2831 4105 2842 4125
rect 2862 4105 2880 4125
rect 2831 4095 2880 4105
rect 2930 4121 2974 4137
rect 2930 4101 2945 4121
rect 2965 4101 2974 4121
rect 2930 4095 2974 4101
rect 3044 4121 3088 4137
rect 3044 4101 3053 4121
rect 3073 4101 3088 4121
rect 3044 4095 3088 4101
rect 3138 4125 3187 4137
rect 3138 4105 3156 4125
rect 3176 4105 3187 4125
rect 3138 4095 3187 4105
rect 3252 4121 3296 4137
rect 3252 4101 3261 4121
rect 3281 4101 3296 4121
rect 3252 4095 3296 4101
rect 3346 4125 3395 4137
rect 3346 4105 3364 4125
rect 3384 4105 3395 4125
rect 3346 4095 3395 4105
rect 3465 4121 3509 4137
rect 3465 4101 3474 4121
rect 3494 4101 3509 4121
rect 3465 4095 3509 4101
rect 3559 4125 3608 4137
rect 3559 4105 3577 4125
rect 3597 4105 3608 4125
rect 3559 4095 3608 4105
rect 309 4044 358 4054
rect 309 4024 320 4044
rect 340 4024 358 4044
rect 309 4012 358 4024
rect 408 4048 452 4054
rect 408 4028 423 4048
rect 443 4028 452 4048
rect 408 4012 452 4028
rect 522 4044 571 4054
rect 522 4024 533 4044
rect 553 4024 571 4044
rect 522 4012 571 4024
rect 621 4048 665 4054
rect 621 4028 636 4048
rect 656 4028 665 4048
rect 621 4012 665 4028
rect 730 4044 779 4054
rect 730 4024 741 4044
rect 761 4024 779 4044
rect 730 4012 779 4024
rect 829 4048 873 4054
rect 829 4028 844 4048
rect 864 4028 873 4048
rect 829 4012 873 4028
rect 943 4048 987 4054
rect 943 4028 952 4048
rect 972 4028 987 4048
rect 943 4012 987 4028
rect 1037 4044 1086 4054
rect 1037 4024 1055 4044
rect 1075 4024 1086 4044
rect 1037 4012 1086 4024
rect 4142 3815 4191 3827
rect 4142 3795 4153 3815
rect 4173 3795 4191 3815
rect 4142 3785 4191 3795
rect 4241 3811 4285 3827
rect 4241 3791 4256 3811
rect 4276 3791 4285 3811
rect 4241 3785 4285 3791
rect 4355 3811 4399 3827
rect 4355 3791 4364 3811
rect 4384 3791 4399 3811
rect 4355 3785 4399 3791
rect 4449 3815 4498 3827
rect 4449 3795 4467 3815
rect 4487 3795 4498 3815
rect 4449 3785 4498 3795
rect 4563 3811 4607 3827
rect 4563 3791 4572 3811
rect 4592 3791 4607 3811
rect 4563 3785 4607 3791
rect 4657 3815 4706 3827
rect 4657 3795 4675 3815
rect 4695 3795 4706 3815
rect 4657 3785 4706 3795
rect 4776 3811 4820 3827
rect 4776 3791 4785 3811
rect 4805 3791 4820 3811
rect 4776 3785 4820 3791
rect 4870 3815 4919 3827
rect 4870 3795 4888 3815
rect 4908 3795 4919 3815
rect 4870 3785 4919 3795
rect 1620 3734 1669 3744
rect 1620 3714 1631 3734
rect 1651 3714 1669 3734
rect 1620 3702 1669 3714
rect 1719 3738 1763 3744
rect 1719 3718 1734 3738
rect 1754 3718 1763 3738
rect 1719 3702 1763 3718
rect 1833 3734 1882 3744
rect 1833 3714 1844 3734
rect 1864 3714 1882 3734
rect 1833 3702 1882 3714
rect 1932 3738 1976 3744
rect 1932 3718 1947 3738
rect 1967 3718 1976 3738
rect 1932 3702 1976 3718
rect 2041 3734 2090 3744
rect 2041 3714 2052 3734
rect 2072 3714 2090 3734
rect 2041 3702 2090 3714
rect 2140 3738 2184 3744
rect 2140 3718 2155 3738
rect 2175 3718 2184 3738
rect 2140 3702 2184 3718
rect 2254 3738 2298 3744
rect 2254 3718 2263 3738
rect 2283 3718 2298 3738
rect 2254 3702 2298 3718
rect 2348 3734 2397 3744
rect 2348 3714 2366 3734
rect 2386 3714 2397 3734
rect 2348 3702 2397 3714
rect 3129 3581 3178 3593
rect 3129 3561 3140 3581
rect 3160 3561 3178 3581
rect 3129 3551 3178 3561
rect 3228 3577 3272 3593
rect 3228 3557 3243 3577
rect 3263 3557 3272 3577
rect 3228 3551 3272 3557
rect 3342 3577 3386 3593
rect 3342 3557 3351 3577
rect 3371 3557 3386 3577
rect 3342 3551 3386 3557
rect 3436 3581 3485 3593
rect 3436 3561 3454 3581
rect 3474 3561 3485 3581
rect 3436 3551 3485 3561
rect 3550 3577 3594 3593
rect 3550 3557 3559 3577
rect 3579 3557 3594 3577
rect 3550 3551 3594 3557
rect 3644 3581 3693 3593
rect 3644 3561 3662 3581
rect 3682 3561 3693 3581
rect 3644 3551 3693 3561
rect 3763 3577 3807 3593
rect 3763 3557 3772 3577
rect 3792 3557 3807 3577
rect 3763 3551 3807 3557
rect 3857 3581 3906 3593
rect 3857 3561 3875 3581
rect 3895 3561 3906 3581
rect 3857 3551 3906 3561
rect 313 3483 362 3493
rect 313 3463 324 3483
rect 344 3463 362 3483
rect 313 3451 362 3463
rect 412 3487 456 3493
rect 412 3467 427 3487
rect 447 3467 456 3487
rect 412 3451 456 3467
rect 526 3483 575 3493
rect 526 3463 537 3483
rect 557 3463 575 3483
rect 526 3451 575 3463
rect 625 3487 669 3493
rect 625 3467 640 3487
rect 660 3467 669 3487
rect 625 3451 669 3467
rect 734 3483 783 3493
rect 734 3463 745 3483
rect 765 3463 783 3483
rect 734 3451 783 3463
rect 833 3487 877 3493
rect 833 3467 848 3487
rect 868 3467 877 3487
rect 833 3451 877 3467
rect 947 3487 991 3493
rect 947 3467 956 3487
rect 976 3467 991 3487
rect 947 3451 991 3467
rect 1041 3483 1090 3493
rect 1041 3463 1059 3483
rect 1079 3463 1090 3483
rect 1041 3451 1090 3463
rect 4141 3400 4190 3412
rect 4141 3380 4152 3400
rect 4172 3380 4190 3400
rect 4141 3370 4190 3380
rect 4240 3396 4284 3412
rect 4240 3376 4255 3396
rect 4275 3376 4284 3396
rect 4240 3370 4284 3376
rect 4354 3396 4398 3412
rect 4354 3376 4363 3396
rect 4383 3376 4398 3396
rect 4354 3370 4398 3376
rect 4448 3400 4497 3412
rect 4448 3380 4466 3400
rect 4486 3380 4497 3400
rect 4448 3370 4497 3380
rect 4562 3396 4606 3412
rect 4562 3376 4571 3396
rect 4591 3376 4606 3396
rect 4562 3370 4606 3376
rect 4656 3400 4705 3412
rect 4656 3380 4674 3400
rect 4694 3380 4705 3400
rect 4656 3370 4705 3380
rect 4775 3396 4819 3412
rect 4775 3376 4784 3396
rect 4804 3376 4819 3396
rect 4775 3370 4819 3376
rect 4869 3400 4918 3412
rect 4869 3380 4887 3400
rect 4907 3380 4918 3400
rect 4869 3370 4918 3380
rect 1325 3302 1374 3312
rect 1325 3282 1336 3302
rect 1356 3282 1374 3302
rect 1325 3270 1374 3282
rect 1424 3306 1468 3312
rect 1424 3286 1439 3306
rect 1459 3286 1468 3306
rect 1424 3270 1468 3286
rect 1538 3302 1587 3312
rect 1538 3282 1549 3302
rect 1569 3282 1587 3302
rect 1538 3270 1587 3282
rect 1637 3306 1681 3312
rect 1637 3286 1652 3306
rect 1672 3286 1681 3306
rect 1637 3270 1681 3286
rect 1746 3302 1795 3312
rect 1746 3282 1757 3302
rect 1777 3282 1795 3302
rect 1746 3270 1795 3282
rect 1845 3306 1889 3312
rect 1845 3286 1860 3306
rect 1880 3286 1889 3306
rect 1845 3270 1889 3286
rect 1959 3306 2003 3312
rect 1959 3286 1968 3306
rect 1988 3286 2003 3306
rect 1959 3270 2003 3286
rect 2053 3302 2102 3312
rect 2053 3282 2071 3302
rect 2091 3282 2102 3302
rect 2053 3270 2102 3282
rect 3079 3161 3128 3173
rect 3079 3141 3090 3161
rect 3110 3141 3128 3161
rect 3079 3131 3128 3141
rect 3178 3157 3222 3173
rect 3178 3137 3193 3157
rect 3213 3137 3222 3157
rect 3178 3131 3222 3137
rect 3292 3157 3336 3173
rect 3292 3137 3301 3157
rect 3321 3137 3336 3157
rect 3292 3131 3336 3137
rect 3386 3161 3435 3173
rect 3386 3141 3404 3161
rect 3424 3141 3435 3161
rect 3386 3131 3435 3141
rect 3500 3157 3544 3173
rect 3500 3137 3509 3157
rect 3529 3137 3544 3157
rect 3500 3131 3544 3137
rect 3594 3161 3643 3173
rect 3594 3141 3612 3161
rect 3632 3141 3643 3161
rect 3594 3131 3643 3141
rect 3713 3157 3757 3173
rect 3713 3137 3722 3157
rect 3742 3137 3757 3157
rect 3713 3131 3757 3137
rect 3807 3161 3856 3173
rect 3807 3141 3825 3161
rect 3845 3141 3856 3161
rect 3807 3131 3856 3141
rect 312 3068 361 3078
rect 312 3048 323 3068
rect 343 3048 361 3068
rect 312 3036 361 3048
rect 411 3072 455 3078
rect 411 3052 426 3072
rect 446 3052 455 3072
rect 411 3036 455 3052
rect 525 3068 574 3078
rect 525 3048 536 3068
rect 556 3048 574 3068
rect 525 3036 574 3048
rect 624 3072 668 3078
rect 624 3052 639 3072
rect 659 3052 668 3072
rect 624 3036 668 3052
rect 733 3068 782 3078
rect 733 3048 744 3068
rect 764 3048 782 3068
rect 733 3036 782 3048
rect 832 3072 876 3078
rect 832 3052 847 3072
rect 867 3052 876 3072
rect 832 3036 876 3052
rect 946 3072 990 3078
rect 946 3052 955 3072
rect 975 3052 990 3072
rect 946 3036 990 3052
rect 1040 3068 1089 3078
rect 1040 3048 1058 3068
rect 1078 3048 1089 3068
rect 1040 3036 1089 3048
rect 4147 2834 4196 2846
rect 4147 2814 4158 2834
rect 4178 2814 4196 2834
rect 4147 2804 4196 2814
rect 4246 2830 4290 2846
rect 4246 2810 4261 2830
rect 4281 2810 4290 2830
rect 4246 2804 4290 2810
rect 4360 2830 4404 2846
rect 4360 2810 4369 2830
rect 4389 2810 4404 2830
rect 4360 2804 4404 2810
rect 4454 2834 4503 2846
rect 4454 2814 4472 2834
rect 4492 2814 4503 2834
rect 4454 2804 4503 2814
rect 4568 2830 4612 2846
rect 4568 2810 4577 2830
rect 4597 2810 4612 2830
rect 4568 2804 4612 2810
rect 4662 2834 4711 2846
rect 4662 2814 4680 2834
rect 4700 2814 4711 2834
rect 4662 2804 4711 2814
rect 4781 2830 4825 2846
rect 4781 2810 4790 2830
rect 4810 2810 4825 2830
rect 4781 2804 4825 2810
rect 4875 2834 4924 2846
rect 4875 2814 4893 2834
rect 4913 2814 4924 2834
rect 4875 2804 4924 2814
rect 1380 2741 1429 2751
rect 1380 2721 1391 2741
rect 1411 2721 1429 2741
rect 1380 2709 1429 2721
rect 1479 2745 1523 2751
rect 1479 2725 1494 2745
rect 1514 2725 1523 2745
rect 1479 2709 1523 2725
rect 1593 2741 1642 2751
rect 1593 2721 1604 2741
rect 1624 2721 1642 2741
rect 1593 2709 1642 2721
rect 1692 2745 1736 2751
rect 1692 2725 1707 2745
rect 1727 2725 1736 2745
rect 1692 2709 1736 2725
rect 1801 2741 1850 2751
rect 1801 2721 1812 2741
rect 1832 2721 1850 2741
rect 1801 2709 1850 2721
rect 1900 2745 1944 2751
rect 1900 2725 1915 2745
rect 1935 2725 1944 2745
rect 1900 2709 1944 2725
rect 2014 2745 2058 2751
rect 2014 2725 2023 2745
rect 2043 2725 2058 2745
rect 2014 2709 2058 2725
rect 2108 2741 2157 2751
rect 2108 2721 2126 2741
rect 2146 2721 2157 2741
rect 2108 2709 2157 2721
rect 3134 2600 3183 2612
rect 3134 2580 3145 2600
rect 3165 2580 3183 2600
rect 3134 2570 3183 2580
rect 3233 2596 3277 2612
rect 3233 2576 3248 2596
rect 3268 2576 3277 2596
rect 3233 2570 3277 2576
rect 3347 2596 3391 2612
rect 3347 2576 3356 2596
rect 3376 2576 3391 2596
rect 3347 2570 3391 2576
rect 3441 2600 3490 2612
rect 3441 2580 3459 2600
rect 3479 2580 3490 2600
rect 3441 2570 3490 2580
rect 3555 2596 3599 2612
rect 3555 2576 3564 2596
rect 3584 2576 3599 2596
rect 3555 2570 3599 2576
rect 3649 2600 3698 2612
rect 3649 2580 3667 2600
rect 3687 2580 3698 2600
rect 3649 2570 3698 2580
rect 3768 2596 3812 2612
rect 3768 2576 3777 2596
rect 3797 2576 3812 2596
rect 3768 2570 3812 2576
rect 3862 2600 3911 2612
rect 3862 2580 3880 2600
rect 3900 2580 3911 2600
rect 3862 2570 3911 2580
rect 318 2502 367 2512
rect 318 2482 329 2502
rect 349 2482 367 2502
rect 318 2470 367 2482
rect 417 2506 461 2512
rect 417 2486 432 2506
rect 452 2486 461 2506
rect 417 2470 461 2486
rect 531 2502 580 2512
rect 531 2482 542 2502
rect 562 2482 580 2502
rect 531 2470 580 2482
rect 630 2506 674 2512
rect 630 2486 645 2506
rect 665 2486 674 2506
rect 630 2470 674 2486
rect 739 2502 788 2512
rect 739 2482 750 2502
rect 770 2482 788 2502
rect 739 2470 788 2482
rect 838 2506 882 2512
rect 838 2486 853 2506
rect 873 2486 882 2506
rect 838 2470 882 2486
rect 952 2506 996 2512
rect 952 2486 961 2506
rect 981 2486 996 2506
rect 952 2470 996 2486
rect 1046 2502 1095 2512
rect 1046 2482 1064 2502
rect 1084 2482 1095 2502
rect 1046 2470 1095 2482
rect 4146 2419 4195 2431
rect 4146 2399 4157 2419
rect 4177 2399 4195 2419
rect 4146 2389 4195 2399
rect 4245 2415 4289 2431
rect 4245 2395 4260 2415
rect 4280 2395 4289 2415
rect 4245 2389 4289 2395
rect 4359 2415 4403 2431
rect 4359 2395 4368 2415
rect 4388 2395 4403 2415
rect 4359 2389 4403 2395
rect 4453 2419 4502 2431
rect 4453 2399 4471 2419
rect 4491 2399 4502 2419
rect 4453 2389 4502 2399
rect 4567 2415 4611 2431
rect 4567 2395 4576 2415
rect 4596 2395 4611 2415
rect 4567 2389 4611 2395
rect 4661 2419 4710 2431
rect 4661 2399 4679 2419
rect 4699 2399 4710 2419
rect 4661 2389 4710 2399
rect 4780 2415 4824 2431
rect 4780 2395 4789 2415
rect 4809 2395 4824 2415
rect 4780 2389 4824 2395
rect 4874 2419 4923 2431
rect 4874 2399 4892 2419
rect 4912 2399 4923 2419
rect 4874 2389 4923 2399
rect 1330 2321 1379 2331
rect 1330 2301 1341 2321
rect 1361 2301 1379 2321
rect 1330 2289 1379 2301
rect 1429 2325 1473 2331
rect 1429 2305 1444 2325
rect 1464 2305 1473 2325
rect 1429 2289 1473 2305
rect 1543 2321 1592 2331
rect 1543 2301 1554 2321
rect 1574 2301 1592 2321
rect 1543 2289 1592 2301
rect 1642 2325 1686 2331
rect 1642 2305 1657 2325
rect 1677 2305 1686 2325
rect 1642 2289 1686 2305
rect 1751 2321 1800 2331
rect 1751 2301 1762 2321
rect 1782 2301 1800 2321
rect 1751 2289 1800 2301
rect 1850 2325 1894 2331
rect 1850 2305 1865 2325
rect 1885 2305 1894 2325
rect 1850 2289 1894 2305
rect 1964 2325 2008 2331
rect 1964 2305 1973 2325
rect 1993 2305 2008 2325
rect 1964 2289 2008 2305
rect 2058 2321 2107 2331
rect 2058 2301 2076 2321
rect 2096 2301 2107 2321
rect 2058 2289 2107 2301
rect 2926 2133 2975 2145
rect 2926 2113 2937 2133
rect 2957 2113 2975 2133
rect 2926 2103 2975 2113
rect 3025 2129 3069 2145
rect 3025 2109 3040 2129
rect 3060 2109 3069 2129
rect 3025 2103 3069 2109
rect 3139 2129 3183 2145
rect 3139 2109 3148 2129
rect 3168 2109 3183 2129
rect 3139 2103 3183 2109
rect 3233 2133 3282 2145
rect 3233 2113 3251 2133
rect 3271 2113 3282 2133
rect 3233 2103 3282 2113
rect 3347 2129 3391 2145
rect 3347 2109 3356 2129
rect 3376 2109 3391 2129
rect 3347 2103 3391 2109
rect 3441 2133 3490 2145
rect 3441 2113 3459 2133
rect 3479 2113 3490 2133
rect 3441 2103 3490 2113
rect 3560 2129 3604 2145
rect 3560 2109 3569 2129
rect 3589 2109 3604 2129
rect 3560 2103 3604 2109
rect 3654 2133 3703 2145
rect 3654 2113 3672 2133
rect 3692 2113 3703 2133
rect 3654 2103 3703 2113
rect 317 2087 366 2097
rect 317 2067 328 2087
rect 348 2067 366 2087
rect 317 2055 366 2067
rect 416 2091 460 2097
rect 416 2071 431 2091
rect 451 2071 460 2091
rect 416 2055 460 2071
rect 530 2087 579 2097
rect 530 2067 541 2087
rect 561 2067 579 2087
rect 530 2055 579 2067
rect 629 2091 673 2097
rect 629 2071 644 2091
rect 664 2071 673 2091
rect 629 2055 673 2071
rect 738 2087 787 2097
rect 738 2067 749 2087
rect 769 2067 787 2087
rect 738 2055 787 2067
rect 837 2091 881 2097
rect 837 2071 852 2091
rect 872 2071 881 2091
rect 837 2055 881 2071
rect 951 2091 995 2097
rect 951 2071 960 2091
rect 980 2071 995 2091
rect 951 2055 995 2071
rect 1045 2087 1094 2097
rect 1045 2067 1063 2087
rect 1083 2067 1094 2087
rect 1045 2055 1094 2067
rect 4154 1855 4203 1867
rect 4154 1835 4165 1855
rect 4185 1835 4203 1855
rect 4154 1825 4203 1835
rect 4253 1851 4297 1867
rect 4253 1831 4268 1851
rect 4288 1831 4297 1851
rect 4253 1825 4297 1831
rect 4367 1851 4411 1867
rect 4367 1831 4376 1851
rect 4396 1831 4411 1851
rect 4367 1825 4411 1831
rect 4461 1855 4510 1867
rect 4461 1835 4479 1855
rect 4499 1835 4510 1855
rect 4461 1825 4510 1835
rect 4575 1851 4619 1867
rect 4575 1831 4584 1851
rect 4604 1831 4619 1851
rect 4575 1825 4619 1831
rect 4669 1855 4718 1867
rect 4669 1835 4687 1855
rect 4707 1835 4718 1855
rect 4669 1825 4718 1835
rect 4788 1851 4832 1867
rect 4788 1831 4797 1851
rect 4817 1831 4832 1851
rect 4788 1825 4832 1831
rect 4882 1855 4931 1867
rect 4882 1835 4900 1855
rect 4920 1835 4931 1855
rect 4882 1825 4931 1835
rect 1545 1809 1594 1819
rect 1545 1789 1556 1809
rect 1576 1789 1594 1809
rect 1545 1777 1594 1789
rect 1644 1813 1688 1819
rect 1644 1793 1659 1813
rect 1679 1793 1688 1813
rect 1644 1777 1688 1793
rect 1758 1809 1807 1819
rect 1758 1789 1769 1809
rect 1789 1789 1807 1809
rect 1758 1777 1807 1789
rect 1857 1813 1901 1819
rect 1857 1793 1872 1813
rect 1892 1793 1901 1813
rect 1857 1777 1901 1793
rect 1966 1809 2015 1819
rect 1966 1789 1977 1809
rect 1997 1789 2015 1809
rect 1966 1777 2015 1789
rect 2065 1813 2109 1819
rect 2065 1793 2080 1813
rect 2100 1793 2109 1813
rect 2065 1777 2109 1793
rect 2179 1813 2223 1819
rect 2179 1793 2188 1813
rect 2208 1793 2223 1813
rect 2179 1777 2223 1793
rect 2273 1809 2322 1819
rect 2273 1789 2291 1809
rect 2311 1789 2322 1809
rect 2273 1777 2322 1789
rect 3141 1621 3190 1633
rect 3141 1601 3152 1621
rect 3172 1601 3190 1621
rect 3141 1591 3190 1601
rect 3240 1617 3284 1633
rect 3240 1597 3255 1617
rect 3275 1597 3284 1617
rect 3240 1591 3284 1597
rect 3354 1617 3398 1633
rect 3354 1597 3363 1617
rect 3383 1597 3398 1617
rect 3354 1591 3398 1597
rect 3448 1621 3497 1633
rect 3448 1601 3466 1621
rect 3486 1601 3497 1621
rect 3448 1591 3497 1601
rect 3562 1617 3606 1633
rect 3562 1597 3571 1617
rect 3591 1597 3606 1617
rect 3562 1591 3606 1597
rect 3656 1621 3705 1633
rect 3656 1601 3674 1621
rect 3694 1601 3705 1621
rect 3656 1591 3705 1601
rect 3775 1617 3819 1633
rect 3775 1597 3784 1617
rect 3804 1597 3819 1617
rect 3775 1591 3819 1597
rect 3869 1621 3918 1633
rect 3869 1601 3887 1621
rect 3907 1601 3918 1621
rect 3869 1591 3918 1601
rect 325 1523 374 1533
rect 325 1503 336 1523
rect 356 1503 374 1523
rect 325 1491 374 1503
rect 424 1527 468 1533
rect 424 1507 439 1527
rect 459 1507 468 1527
rect 424 1491 468 1507
rect 538 1523 587 1533
rect 538 1503 549 1523
rect 569 1503 587 1523
rect 538 1491 587 1503
rect 637 1527 681 1533
rect 637 1507 652 1527
rect 672 1507 681 1527
rect 637 1491 681 1507
rect 746 1523 795 1533
rect 746 1503 757 1523
rect 777 1503 795 1523
rect 746 1491 795 1503
rect 845 1527 889 1533
rect 845 1507 860 1527
rect 880 1507 889 1527
rect 845 1491 889 1507
rect 959 1527 1003 1533
rect 959 1507 968 1527
rect 988 1507 1003 1527
rect 959 1491 1003 1507
rect 1053 1523 1102 1533
rect 1053 1503 1071 1523
rect 1091 1503 1102 1523
rect 1053 1491 1102 1503
rect 4153 1440 4202 1452
rect 4153 1420 4164 1440
rect 4184 1420 4202 1440
rect 4153 1410 4202 1420
rect 4252 1436 4296 1452
rect 4252 1416 4267 1436
rect 4287 1416 4296 1436
rect 4252 1410 4296 1416
rect 4366 1436 4410 1452
rect 4366 1416 4375 1436
rect 4395 1416 4410 1436
rect 4366 1410 4410 1416
rect 4460 1440 4509 1452
rect 4460 1420 4478 1440
rect 4498 1420 4509 1440
rect 4460 1410 4509 1420
rect 4574 1436 4618 1452
rect 4574 1416 4583 1436
rect 4603 1416 4618 1436
rect 4574 1410 4618 1416
rect 4668 1440 4717 1452
rect 4668 1420 4686 1440
rect 4706 1420 4717 1440
rect 4668 1410 4717 1420
rect 4787 1436 4831 1452
rect 4787 1416 4796 1436
rect 4816 1416 4831 1436
rect 4787 1410 4831 1416
rect 4881 1440 4930 1452
rect 4881 1420 4899 1440
rect 4919 1420 4930 1440
rect 4881 1410 4930 1420
rect 1337 1342 1386 1352
rect 1337 1322 1348 1342
rect 1368 1322 1386 1342
rect 1337 1310 1386 1322
rect 1436 1346 1480 1352
rect 1436 1326 1451 1346
rect 1471 1326 1480 1346
rect 1436 1310 1480 1326
rect 1550 1342 1599 1352
rect 1550 1322 1561 1342
rect 1581 1322 1599 1342
rect 1550 1310 1599 1322
rect 1649 1346 1693 1352
rect 1649 1326 1664 1346
rect 1684 1326 1693 1346
rect 1649 1310 1693 1326
rect 1758 1342 1807 1352
rect 1758 1322 1769 1342
rect 1789 1322 1807 1342
rect 1758 1310 1807 1322
rect 1857 1346 1901 1352
rect 1857 1326 1872 1346
rect 1892 1326 1901 1346
rect 1857 1310 1901 1326
rect 1971 1346 2015 1352
rect 1971 1326 1980 1346
rect 2000 1326 2015 1346
rect 1971 1310 2015 1326
rect 2065 1342 2114 1352
rect 2065 1322 2083 1342
rect 2103 1322 2114 1342
rect 2065 1310 2114 1322
rect 3091 1201 3140 1213
rect 3091 1181 3102 1201
rect 3122 1181 3140 1201
rect 3091 1171 3140 1181
rect 3190 1197 3234 1213
rect 3190 1177 3205 1197
rect 3225 1177 3234 1197
rect 3190 1171 3234 1177
rect 3304 1197 3348 1213
rect 3304 1177 3313 1197
rect 3333 1177 3348 1197
rect 3304 1171 3348 1177
rect 3398 1201 3447 1213
rect 3398 1181 3416 1201
rect 3436 1181 3447 1201
rect 3398 1171 3447 1181
rect 3512 1197 3556 1213
rect 3512 1177 3521 1197
rect 3541 1177 3556 1197
rect 3512 1171 3556 1177
rect 3606 1201 3655 1213
rect 3606 1181 3624 1201
rect 3644 1181 3655 1201
rect 3606 1171 3655 1181
rect 3725 1197 3769 1213
rect 3725 1177 3734 1197
rect 3754 1177 3769 1197
rect 3725 1171 3769 1177
rect 3819 1201 3868 1213
rect 3819 1181 3837 1201
rect 3857 1181 3868 1201
rect 3819 1171 3868 1181
rect 324 1108 373 1118
rect 324 1088 335 1108
rect 355 1088 373 1108
rect 324 1076 373 1088
rect 423 1112 467 1118
rect 423 1092 438 1112
rect 458 1092 467 1112
rect 423 1076 467 1092
rect 537 1108 586 1118
rect 537 1088 548 1108
rect 568 1088 586 1108
rect 537 1076 586 1088
rect 636 1112 680 1118
rect 636 1092 651 1112
rect 671 1092 680 1112
rect 636 1076 680 1092
rect 745 1108 794 1118
rect 745 1088 756 1108
rect 776 1088 794 1108
rect 745 1076 794 1088
rect 844 1112 888 1118
rect 844 1092 859 1112
rect 879 1092 888 1112
rect 844 1076 888 1092
rect 958 1112 1002 1118
rect 958 1092 967 1112
rect 987 1092 1002 1112
rect 958 1076 1002 1092
rect 1052 1108 1101 1118
rect 1052 1088 1070 1108
rect 1090 1088 1101 1108
rect 1052 1076 1101 1088
rect 4159 874 4208 886
rect 4159 854 4170 874
rect 4190 854 4208 874
rect 4159 844 4208 854
rect 4258 870 4302 886
rect 4258 850 4273 870
rect 4293 850 4302 870
rect 4258 844 4302 850
rect 4372 870 4416 886
rect 4372 850 4381 870
rect 4401 850 4416 870
rect 4372 844 4416 850
rect 4466 874 4515 886
rect 4466 854 4484 874
rect 4504 854 4515 874
rect 4466 844 4515 854
rect 4580 870 4624 886
rect 4580 850 4589 870
rect 4609 850 4624 870
rect 4580 844 4624 850
rect 4674 874 4723 886
rect 4674 854 4692 874
rect 4712 854 4723 874
rect 4674 844 4723 854
rect 4793 870 4837 886
rect 4793 850 4802 870
rect 4822 850 4837 870
rect 4793 844 4837 850
rect 4887 874 4936 886
rect 4887 854 4905 874
rect 4925 854 4936 874
rect 4887 844 4936 854
rect 1392 781 1441 791
rect 1392 761 1403 781
rect 1423 761 1441 781
rect 1392 749 1441 761
rect 1491 785 1535 791
rect 1491 765 1506 785
rect 1526 765 1535 785
rect 1491 749 1535 765
rect 1605 781 1654 791
rect 1605 761 1616 781
rect 1636 761 1654 781
rect 1605 749 1654 761
rect 1704 785 1748 791
rect 1704 765 1719 785
rect 1739 765 1748 785
rect 1704 749 1748 765
rect 1813 781 1862 791
rect 1813 761 1824 781
rect 1844 761 1862 781
rect 1813 749 1862 761
rect 1912 785 1956 791
rect 1912 765 1927 785
rect 1947 765 1956 785
rect 1912 749 1956 765
rect 2026 785 2070 791
rect 2026 765 2035 785
rect 2055 765 2070 785
rect 2026 749 2070 765
rect 2120 781 2169 791
rect 2120 761 2138 781
rect 2158 761 2169 781
rect 2120 749 2169 761
rect 3146 640 3195 652
rect 3146 620 3157 640
rect 3177 620 3195 640
rect 3146 610 3195 620
rect 3245 636 3289 652
rect 3245 616 3260 636
rect 3280 616 3289 636
rect 3245 610 3289 616
rect 3359 636 3403 652
rect 3359 616 3368 636
rect 3388 616 3403 636
rect 3359 610 3403 616
rect 3453 640 3502 652
rect 3453 620 3471 640
rect 3491 620 3502 640
rect 3453 610 3502 620
rect 3567 636 3611 652
rect 3567 616 3576 636
rect 3596 616 3611 636
rect 3567 610 3611 616
rect 3661 640 3710 652
rect 3661 620 3679 640
rect 3699 620 3710 640
rect 3661 610 3710 620
rect 3780 636 3824 652
rect 3780 616 3789 636
rect 3809 616 3824 636
rect 3780 610 3824 616
rect 3874 640 3923 652
rect 3874 620 3892 640
rect 3912 620 3923 640
rect 3874 610 3923 620
rect 330 542 379 552
rect 330 522 341 542
rect 361 522 379 542
rect 330 510 379 522
rect 429 546 473 552
rect 429 526 444 546
rect 464 526 473 546
rect 429 510 473 526
rect 543 542 592 552
rect 543 522 554 542
rect 574 522 592 542
rect 543 510 592 522
rect 642 546 686 552
rect 642 526 657 546
rect 677 526 686 546
rect 642 510 686 526
rect 751 542 800 552
rect 751 522 762 542
rect 782 522 800 542
rect 751 510 800 522
rect 850 546 894 552
rect 850 526 865 546
rect 885 526 894 546
rect 850 510 894 526
rect 964 546 1008 552
rect 964 526 973 546
rect 993 526 1008 546
rect 964 510 1008 526
rect 1058 542 1107 552
rect 1058 522 1076 542
rect 1096 522 1107 542
rect 1058 510 1107 522
rect 4158 459 4207 471
rect 4158 439 4169 459
rect 4189 439 4207 459
rect 4158 429 4207 439
rect 4257 455 4301 471
rect 4257 435 4272 455
rect 4292 435 4301 455
rect 4257 429 4301 435
rect 4371 455 4415 471
rect 4371 435 4380 455
rect 4400 435 4415 455
rect 4371 429 4415 435
rect 4465 459 4514 471
rect 4465 439 4483 459
rect 4503 439 4514 459
rect 4465 429 4514 439
rect 4579 455 4623 471
rect 4579 435 4588 455
rect 4608 435 4623 455
rect 4579 429 4623 435
rect 4673 459 4722 471
rect 4673 439 4691 459
rect 4711 439 4722 459
rect 4673 429 4722 439
rect 4792 455 4836 471
rect 4792 435 4801 455
rect 4821 435 4836 455
rect 4792 429 4836 435
rect 4886 459 4935 471
rect 4886 439 4904 459
rect 4924 439 4935 459
rect 4886 429 4935 439
rect 1342 361 1391 371
rect 1342 341 1353 361
rect 1373 341 1391 361
rect 1342 329 1391 341
rect 1441 365 1485 371
rect 1441 345 1456 365
rect 1476 345 1485 365
rect 1441 329 1485 345
rect 1555 361 1604 371
rect 1555 341 1566 361
rect 1586 341 1604 361
rect 1555 329 1604 341
rect 1654 365 1698 371
rect 1654 345 1669 365
rect 1689 345 1698 365
rect 1654 329 1698 345
rect 1763 361 1812 371
rect 1763 341 1774 361
rect 1794 341 1812 361
rect 1763 329 1812 341
rect 1862 365 1906 371
rect 1862 345 1877 365
rect 1897 345 1906 365
rect 1862 329 1906 345
rect 1976 365 2020 371
rect 1976 345 1985 365
rect 2005 345 2020 365
rect 1976 329 2020 345
rect 2070 361 2119 371
rect 2070 341 2088 361
rect 2108 341 2119 361
rect 2070 329 2119 341
rect 329 127 378 137
rect 329 107 340 127
rect 360 107 378 127
rect 329 95 378 107
rect 428 131 472 137
rect 428 111 443 131
rect 463 111 472 131
rect 428 95 472 111
rect 542 127 591 137
rect 542 107 553 127
rect 573 107 591 127
rect 542 95 591 107
rect 641 131 685 137
rect 641 111 656 131
rect 676 111 685 131
rect 641 95 685 111
rect 750 127 799 137
rect 750 107 761 127
rect 781 107 799 127
rect 750 95 799 107
rect 849 131 893 137
rect 849 111 864 131
rect 884 111 893 131
rect 849 95 893 111
rect 963 131 1007 137
rect 963 111 972 131
rect 992 111 1007 131
rect 963 95 1007 111
rect 1057 127 1106 137
rect 1057 107 1075 127
rect 1095 107 1106 127
rect 1057 95 1106 107
rect 1732 -354 1781 -344
rect 1732 -374 1743 -354
rect 1763 -374 1781 -354
rect 1732 -386 1781 -374
rect 1831 -350 1875 -344
rect 1831 -370 1846 -350
rect 1866 -370 1875 -350
rect 1831 -386 1875 -370
rect 1945 -354 1994 -344
rect 1945 -374 1956 -354
rect 1976 -374 1994 -354
rect 1945 -386 1994 -374
rect 2044 -350 2088 -344
rect 2044 -370 2059 -350
rect 2079 -370 2088 -350
rect 2044 -386 2088 -370
rect 2153 -354 2202 -344
rect 2153 -374 2164 -354
rect 2184 -374 2202 -354
rect 2153 -386 2202 -374
rect 2252 -350 2296 -344
rect 2252 -370 2267 -350
rect 2287 -370 2296 -350
rect 2252 -386 2296 -370
rect 2366 -350 2410 -344
rect 2366 -370 2375 -350
rect 2395 -370 2410 -350
rect 2366 -386 2410 -370
rect 2460 -354 2509 -344
rect 2460 -374 2478 -354
rect 2498 -374 2509 -354
rect 2460 -386 2509 -374
<< pdiff >>
rect 298 7549 342 7587
rect 298 7529 310 7549
rect 330 7529 342 7549
rect 298 7487 342 7529
rect 392 7549 434 7587
rect 392 7529 406 7549
rect 426 7529 434 7549
rect 392 7487 434 7529
rect 511 7549 555 7587
rect 511 7529 523 7549
rect 543 7529 555 7549
rect 511 7487 555 7529
rect 605 7549 647 7587
rect 605 7529 619 7549
rect 639 7529 647 7549
rect 605 7487 647 7529
rect 719 7549 763 7587
rect 719 7529 731 7549
rect 751 7529 763 7549
rect 719 7487 763 7529
rect 813 7549 855 7587
rect 813 7529 827 7549
rect 847 7529 855 7549
rect 813 7487 855 7529
rect 929 7549 971 7587
rect 929 7529 937 7549
rect 957 7529 971 7549
rect 929 7487 971 7529
rect 1021 7556 1066 7587
rect 4127 7583 4171 7625
rect 4127 7563 4139 7583
rect 4159 7563 4171 7583
rect 4127 7556 4171 7563
rect 1021 7549 1065 7556
rect 1021 7529 1033 7549
rect 1053 7529 1065 7549
rect 1021 7487 1065 7529
rect 4126 7525 4171 7556
rect 4221 7583 4263 7625
rect 4221 7563 4235 7583
rect 4255 7563 4263 7583
rect 4221 7525 4263 7563
rect 4337 7583 4379 7625
rect 4337 7563 4345 7583
rect 4365 7563 4379 7583
rect 4337 7525 4379 7563
rect 4429 7583 4473 7625
rect 4429 7563 4441 7583
rect 4461 7563 4473 7583
rect 4429 7525 4473 7563
rect 4545 7583 4587 7625
rect 4545 7563 4553 7583
rect 4573 7563 4587 7583
rect 4545 7525 4587 7563
rect 4637 7583 4681 7625
rect 4637 7563 4649 7583
rect 4669 7563 4681 7583
rect 4637 7525 4681 7563
rect 4758 7583 4800 7625
rect 4758 7563 4766 7583
rect 4786 7563 4800 7583
rect 4758 7525 4800 7563
rect 4850 7583 4894 7625
rect 4850 7563 4862 7583
rect 4882 7563 4894 7583
rect 4850 7525 4894 7563
rect 1310 7368 1354 7406
rect 1310 7348 1322 7368
rect 1342 7348 1354 7368
rect 1310 7306 1354 7348
rect 1404 7368 1446 7406
rect 1404 7348 1418 7368
rect 1438 7348 1446 7368
rect 1404 7306 1446 7348
rect 1523 7368 1567 7406
rect 1523 7348 1535 7368
rect 1555 7348 1567 7368
rect 1523 7306 1567 7348
rect 1617 7368 1659 7406
rect 1617 7348 1631 7368
rect 1651 7348 1659 7368
rect 1617 7306 1659 7348
rect 1731 7368 1775 7406
rect 1731 7348 1743 7368
rect 1763 7348 1775 7368
rect 1731 7306 1775 7348
rect 1825 7368 1867 7406
rect 1825 7348 1839 7368
rect 1859 7348 1867 7368
rect 1825 7306 1867 7348
rect 1941 7368 1983 7406
rect 1941 7348 1949 7368
rect 1969 7348 1983 7368
rect 1941 7306 1983 7348
rect 2033 7375 2078 7406
rect 2033 7368 2077 7375
rect 2033 7348 2045 7368
rect 2065 7348 2077 7368
rect 2033 7306 2077 7348
rect 3114 7349 3158 7391
rect 3114 7329 3126 7349
rect 3146 7329 3158 7349
rect 3114 7322 3158 7329
rect 3113 7291 3158 7322
rect 3208 7349 3250 7391
rect 3208 7329 3222 7349
rect 3242 7329 3250 7349
rect 3208 7291 3250 7329
rect 3324 7349 3366 7391
rect 3324 7329 3332 7349
rect 3352 7329 3366 7349
rect 3324 7291 3366 7329
rect 3416 7349 3460 7391
rect 3416 7329 3428 7349
rect 3448 7329 3460 7349
rect 3416 7291 3460 7329
rect 3532 7349 3574 7391
rect 3532 7329 3540 7349
rect 3560 7329 3574 7349
rect 3532 7291 3574 7329
rect 3624 7349 3668 7391
rect 3624 7329 3636 7349
rect 3656 7329 3668 7349
rect 3624 7291 3668 7329
rect 3745 7349 3787 7391
rect 3745 7329 3753 7349
rect 3773 7329 3787 7349
rect 3745 7291 3787 7329
rect 3837 7349 3881 7391
rect 3837 7329 3849 7349
rect 3869 7329 3881 7349
rect 3837 7291 3881 7329
rect 297 7134 341 7172
rect 297 7114 309 7134
rect 329 7114 341 7134
rect 297 7072 341 7114
rect 391 7134 433 7172
rect 391 7114 405 7134
rect 425 7114 433 7134
rect 391 7072 433 7114
rect 510 7134 554 7172
rect 510 7114 522 7134
rect 542 7114 554 7134
rect 510 7072 554 7114
rect 604 7134 646 7172
rect 604 7114 618 7134
rect 638 7114 646 7134
rect 604 7072 646 7114
rect 718 7134 762 7172
rect 718 7114 730 7134
rect 750 7114 762 7134
rect 718 7072 762 7114
rect 812 7134 854 7172
rect 812 7114 826 7134
rect 846 7114 854 7134
rect 812 7072 854 7114
rect 928 7134 970 7172
rect 928 7114 936 7134
rect 956 7114 970 7134
rect 928 7072 970 7114
rect 1020 7141 1065 7172
rect 4126 7168 4170 7210
rect 4126 7148 4138 7168
rect 4158 7148 4170 7168
rect 4126 7141 4170 7148
rect 1020 7134 1064 7141
rect 1020 7114 1032 7134
rect 1052 7114 1064 7134
rect 1020 7072 1064 7114
rect 4125 7110 4170 7141
rect 4220 7168 4262 7210
rect 4220 7148 4234 7168
rect 4254 7148 4262 7168
rect 4220 7110 4262 7148
rect 4336 7168 4378 7210
rect 4336 7148 4344 7168
rect 4364 7148 4378 7168
rect 4336 7110 4378 7148
rect 4428 7168 4472 7210
rect 4428 7148 4440 7168
rect 4460 7148 4472 7168
rect 4428 7110 4472 7148
rect 4544 7168 4586 7210
rect 4544 7148 4552 7168
rect 4572 7148 4586 7168
rect 4544 7110 4586 7148
rect 4636 7168 4680 7210
rect 4636 7148 4648 7168
rect 4668 7148 4680 7168
rect 4636 7110 4680 7148
rect 4757 7168 4799 7210
rect 4757 7148 4765 7168
rect 4785 7148 4799 7168
rect 4757 7110 4799 7148
rect 4849 7168 4893 7210
rect 4849 7148 4861 7168
rect 4881 7148 4893 7168
rect 4849 7110 4893 7148
rect 3064 6929 3108 6971
rect 3064 6909 3076 6929
rect 3096 6909 3108 6929
rect 3064 6902 3108 6909
rect 3063 6871 3108 6902
rect 3158 6929 3200 6971
rect 3158 6909 3172 6929
rect 3192 6909 3200 6929
rect 3158 6871 3200 6909
rect 3274 6929 3316 6971
rect 3274 6909 3282 6929
rect 3302 6909 3316 6929
rect 3274 6871 3316 6909
rect 3366 6929 3410 6971
rect 3366 6909 3378 6929
rect 3398 6909 3410 6929
rect 3366 6871 3410 6909
rect 3482 6929 3524 6971
rect 3482 6909 3490 6929
rect 3510 6909 3524 6929
rect 3482 6871 3524 6909
rect 3574 6929 3618 6971
rect 3574 6909 3586 6929
rect 3606 6909 3618 6929
rect 3574 6871 3618 6909
rect 3695 6929 3737 6971
rect 3695 6909 3703 6929
rect 3723 6909 3737 6929
rect 3695 6871 3737 6909
rect 3787 6929 3831 6971
rect 3787 6909 3799 6929
rect 3819 6909 3831 6929
rect 3787 6871 3831 6909
rect 1365 6807 1409 6845
rect 1365 6787 1377 6807
rect 1397 6787 1409 6807
rect 1365 6745 1409 6787
rect 1459 6807 1501 6845
rect 1459 6787 1473 6807
rect 1493 6787 1501 6807
rect 1459 6745 1501 6787
rect 1578 6807 1622 6845
rect 1578 6787 1590 6807
rect 1610 6787 1622 6807
rect 1578 6745 1622 6787
rect 1672 6807 1714 6845
rect 1672 6787 1686 6807
rect 1706 6787 1714 6807
rect 1672 6745 1714 6787
rect 1786 6807 1830 6845
rect 1786 6787 1798 6807
rect 1818 6787 1830 6807
rect 1786 6745 1830 6787
rect 1880 6807 1922 6845
rect 1880 6787 1894 6807
rect 1914 6787 1922 6807
rect 1880 6745 1922 6787
rect 1996 6807 2038 6845
rect 1996 6787 2004 6807
rect 2024 6787 2038 6807
rect 1996 6745 2038 6787
rect 2088 6814 2133 6845
rect 2088 6807 2132 6814
rect 2088 6787 2100 6807
rect 2120 6787 2132 6807
rect 2088 6745 2132 6787
rect 303 6568 347 6606
rect 303 6548 315 6568
rect 335 6548 347 6568
rect 303 6506 347 6548
rect 397 6568 439 6606
rect 397 6548 411 6568
rect 431 6548 439 6568
rect 397 6506 439 6548
rect 516 6568 560 6606
rect 516 6548 528 6568
rect 548 6548 560 6568
rect 516 6506 560 6548
rect 610 6568 652 6606
rect 610 6548 624 6568
rect 644 6548 652 6568
rect 610 6506 652 6548
rect 724 6568 768 6606
rect 724 6548 736 6568
rect 756 6548 768 6568
rect 724 6506 768 6548
rect 818 6568 860 6606
rect 818 6548 832 6568
rect 852 6548 860 6568
rect 818 6506 860 6548
rect 934 6568 976 6606
rect 934 6548 942 6568
rect 962 6548 976 6568
rect 934 6506 976 6548
rect 1026 6575 1071 6606
rect 4132 6602 4176 6644
rect 4132 6582 4144 6602
rect 4164 6582 4176 6602
rect 4132 6575 4176 6582
rect 1026 6568 1070 6575
rect 1026 6548 1038 6568
rect 1058 6548 1070 6568
rect 1026 6506 1070 6548
rect 4131 6544 4176 6575
rect 4226 6602 4268 6644
rect 4226 6582 4240 6602
rect 4260 6582 4268 6602
rect 4226 6544 4268 6582
rect 4342 6602 4384 6644
rect 4342 6582 4350 6602
rect 4370 6582 4384 6602
rect 4342 6544 4384 6582
rect 4434 6602 4478 6644
rect 4434 6582 4446 6602
rect 4466 6582 4478 6602
rect 4434 6544 4478 6582
rect 4550 6602 4592 6644
rect 4550 6582 4558 6602
rect 4578 6582 4592 6602
rect 4550 6544 4592 6582
rect 4642 6602 4686 6644
rect 4642 6582 4654 6602
rect 4674 6582 4686 6602
rect 4642 6544 4686 6582
rect 4763 6602 4805 6644
rect 4763 6582 4771 6602
rect 4791 6582 4805 6602
rect 4763 6544 4805 6582
rect 4855 6602 4899 6644
rect 4855 6582 4867 6602
rect 4887 6582 4899 6602
rect 4855 6544 4899 6582
rect 1315 6387 1359 6425
rect 1315 6367 1327 6387
rect 1347 6367 1359 6387
rect 1315 6325 1359 6367
rect 1409 6387 1451 6425
rect 1409 6367 1423 6387
rect 1443 6367 1451 6387
rect 1409 6325 1451 6367
rect 1528 6387 1572 6425
rect 1528 6367 1540 6387
rect 1560 6367 1572 6387
rect 1528 6325 1572 6367
rect 1622 6387 1664 6425
rect 1622 6367 1636 6387
rect 1656 6367 1664 6387
rect 1622 6325 1664 6367
rect 1736 6387 1780 6425
rect 1736 6367 1748 6387
rect 1768 6367 1780 6387
rect 1736 6325 1780 6367
rect 1830 6387 1872 6425
rect 1830 6367 1844 6387
rect 1864 6367 1872 6387
rect 1830 6325 1872 6367
rect 1946 6387 1988 6425
rect 1946 6367 1954 6387
rect 1974 6367 1988 6387
rect 1946 6325 1988 6367
rect 2038 6394 2083 6425
rect 2038 6387 2082 6394
rect 2038 6367 2050 6387
rect 2070 6367 2082 6387
rect 2038 6325 2082 6367
rect 3119 6368 3163 6410
rect 3119 6348 3131 6368
rect 3151 6348 3163 6368
rect 3119 6341 3163 6348
rect 3118 6310 3163 6341
rect 3213 6368 3255 6410
rect 3213 6348 3227 6368
rect 3247 6348 3255 6368
rect 3213 6310 3255 6348
rect 3329 6368 3371 6410
rect 3329 6348 3337 6368
rect 3357 6348 3371 6368
rect 3329 6310 3371 6348
rect 3421 6368 3465 6410
rect 3421 6348 3433 6368
rect 3453 6348 3465 6368
rect 3421 6310 3465 6348
rect 3537 6368 3579 6410
rect 3537 6348 3545 6368
rect 3565 6348 3579 6368
rect 3537 6310 3579 6348
rect 3629 6368 3673 6410
rect 3629 6348 3641 6368
rect 3661 6348 3673 6368
rect 3629 6310 3673 6348
rect 3750 6368 3792 6410
rect 3750 6348 3758 6368
rect 3778 6348 3792 6368
rect 3750 6310 3792 6348
rect 3842 6368 3886 6410
rect 3842 6348 3854 6368
rect 3874 6348 3886 6368
rect 3842 6310 3886 6348
rect 302 6153 346 6191
rect 302 6133 314 6153
rect 334 6133 346 6153
rect 302 6091 346 6133
rect 396 6153 438 6191
rect 396 6133 410 6153
rect 430 6133 438 6153
rect 396 6091 438 6133
rect 515 6153 559 6191
rect 515 6133 527 6153
rect 547 6133 559 6153
rect 515 6091 559 6133
rect 609 6153 651 6191
rect 609 6133 623 6153
rect 643 6133 651 6153
rect 609 6091 651 6133
rect 723 6153 767 6191
rect 723 6133 735 6153
rect 755 6133 767 6153
rect 723 6091 767 6133
rect 817 6153 859 6191
rect 817 6133 831 6153
rect 851 6133 859 6153
rect 817 6091 859 6133
rect 933 6153 975 6191
rect 933 6133 941 6153
rect 961 6133 975 6153
rect 933 6091 975 6133
rect 1025 6160 1070 6191
rect 4131 6187 4175 6229
rect 4131 6167 4143 6187
rect 4163 6167 4175 6187
rect 4131 6160 4175 6167
rect 1025 6153 1069 6160
rect 1025 6133 1037 6153
rect 1057 6133 1069 6153
rect 1025 6091 1069 6133
rect 4130 6129 4175 6160
rect 4225 6187 4267 6229
rect 4225 6167 4239 6187
rect 4259 6167 4267 6187
rect 4225 6129 4267 6167
rect 4341 6187 4383 6229
rect 4341 6167 4349 6187
rect 4369 6167 4383 6187
rect 4341 6129 4383 6167
rect 4433 6187 4477 6229
rect 4433 6167 4445 6187
rect 4465 6167 4477 6187
rect 4433 6129 4477 6167
rect 4549 6187 4591 6229
rect 4549 6167 4557 6187
rect 4577 6167 4591 6187
rect 4549 6129 4591 6167
rect 4641 6187 4685 6229
rect 4641 6167 4653 6187
rect 4673 6167 4685 6187
rect 4641 6129 4685 6167
rect 4762 6187 4804 6229
rect 4762 6167 4770 6187
rect 4790 6167 4804 6187
rect 4762 6129 4804 6167
rect 4854 6187 4898 6229
rect 4854 6167 4866 6187
rect 4886 6167 4898 6187
rect 4854 6129 4898 6167
rect 1530 5875 1574 5913
rect 1530 5855 1542 5875
rect 1562 5855 1574 5875
rect 1530 5813 1574 5855
rect 1624 5875 1666 5913
rect 1624 5855 1638 5875
rect 1658 5855 1666 5875
rect 1624 5813 1666 5855
rect 1743 5875 1787 5913
rect 1743 5855 1755 5875
rect 1775 5855 1787 5875
rect 1743 5813 1787 5855
rect 1837 5875 1879 5913
rect 1837 5855 1851 5875
rect 1871 5855 1879 5875
rect 1837 5813 1879 5855
rect 1951 5875 1995 5913
rect 1951 5855 1963 5875
rect 1983 5855 1995 5875
rect 1951 5813 1995 5855
rect 2045 5875 2087 5913
rect 2045 5855 2059 5875
rect 2079 5855 2087 5875
rect 2045 5813 2087 5855
rect 2161 5875 2203 5913
rect 2161 5855 2169 5875
rect 2189 5855 2203 5875
rect 2161 5813 2203 5855
rect 2253 5882 2298 5913
rect 2911 5901 2955 5943
rect 2253 5875 2297 5882
rect 2253 5855 2265 5875
rect 2285 5855 2297 5875
rect 2911 5881 2923 5901
rect 2943 5881 2955 5901
rect 2911 5874 2955 5881
rect 2253 5813 2297 5855
rect 2910 5843 2955 5874
rect 3005 5901 3047 5943
rect 3005 5881 3019 5901
rect 3039 5881 3047 5901
rect 3005 5843 3047 5881
rect 3121 5901 3163 5943
rect 3121 5881 3129 5901
rect 3149 5881 3163 5901
rect 3121 5843 3163 5881
rect 3213 5901 3257 5943
rect 3213 5881 3225 5901
rect 3245 5881 3257 5901
rect 3213 5843 3257 5881
rect 3329 5901 3371 5943
rect 3329 5881 3337 5901
rect 3357 5881 3371 5901
rect 3329 5843 3371 5881
rect 3421 5901 3465 5943
rect 3421 5881 3433 5901
rect 3453 5881 3465 5901
rect 3421 5843 3465 5881
rect 3542 5901 3584 5943
rect 3542 5881 3550 5901
rect 3570 5881 3584 5901
rect 3542 5843 3584 5881
rect 3634 5901 3678 5943
rect 3634 5881 3646 5901
rect 3666 5881 3678 5901
rect 3634 5843 3678 5881
rect 310 5589 354 5627
rect 310 5569 322 5589
rect 342 5569 354 5589
rect 310 5527 354 5569
rect 404 5589 446 5627
rect 404 5569 418 5589
rect 438 5569 446 5589
rect 404 5527 446 5569
rect 523 5589 567 5627
rect 523 5569 535 5589
rect 555 5569 567 5589
rect 523 5527 567 5569
rect 617 5589 659 5627
rect 617 5569 631 5589
rect 651 5569 659 5589
rect 617 5527 659 5569
rect 731 5589 775 5627
rect 731 5569 743 5589
rect 763 5569 775 5589
rect 731 5527 775 5569
rect 825 5589 867 5627
rect 825 5569 839 5589
rect 859 5569 867 5589
rect 825 5527 867 5569
rect 941 5589 983 5627
rect 941 5569 949 5589
rect 969 5569 983 5589
rect 941 5527 983 5569
rect 1033 5596 1078 5627
rect 4139 5623 4183 5665
rect 4139 5603 4151 5623
rect 4171 5603 4183 5623
rect 4139 5596 4183 5603
rect 1033 5589 1077 5596
rect 1033 5569 1045 5589
rect 1065 5569 1077 5589
rect 1033 5527 1077 5569
rect 4138 5565 4183 5596
rect 4233 5623 4275 5665
rect 4233 5603 4247 5623
rect 4267 5603 4275 5623
rect 4233 5565 4275 5603
rect 4349 5623 4391 5665
rect 4349 5603 4357 5623
rect 4377 5603 4391 5623
rect 4349 5565 4391 5603
rect 4441 5623 4485 5665
rect 4441 5603 4453 5623
rect 4473 5603 4485 5623
rect 4441 5565 4485 5603
rect 4557 5623 4599 5665
rect 4557 5603 4565 5623
rect 4585 5603 4599 5623
rect 4557 5565 4599 5603
rect 4649 5623 4693 5665
rect 4649 5603 4661 5623
rect 4681 5603 4693 5623
rect 4649 5565 4693 5603
rect 4770 5623 4812 5665
rect 4770 5603 4778 5623
rect 4798 5603 4812 5623
rect 4770 5565 4812 5603
rect 4862 5623 4906 5665
rect 4862 5603 4874 5623
rect 4894 5603 4906 5623
rect 4862 5565 4906 5603
rect 1322 5408 1366 5446
rect 1322 5388 1334 5408
rect 1354 5388 1366 5408
rect 1322 5346 1366 5388
rect 1416 5408 1458 5446
rect 1416 5388 1430 5408
rect 1450 5388 1458 5408
rect 1416 5346 1458 5388
rect 1535 5408 1579 5446
rect 1535 5388 1547 5408
rect 1567 5388 1579 5408
rect 1535 5346 1579 5388
rect 1629 5408 1671 5446
rect 1629 5388 1643 5408
rect 1663 5388 1671 5408
rect 1629 5346 1671 5388
rect 1743 5408 1787 5446
rect 1743 5388 1755 5408
rect 1775 5388 1787 5408
rect 1743 5346 1787 5388
rect 1837 5408 1879 5446
rect 1837 5388 1851 5408
rect 1871 5388 1879 5408
rect 1837 5346 1879 5388
rect 1953 5408 1995 5446
rect 1953 5388 1961 5408
rect 1981 5388 1995 5408
rect 1953 5346 1995 5388
rect 2045 5415 2090 5446
rect 2045 5408 2089 5415
rect 2045 5388 2057 5408
rect 2077 5388 2089 5408
rect 2045 5346 2089 5388
rect 3126 5389 3170 5431
rect 3126 5369 3138 5389
rect 3158 5369 3170 5389
rect 3126 5362 3170 5369
rect 3125 5331 3170 5362
rect 3220 5389 3262 5431
rect 3220 5369 3234 5389
rect 3254 5369 3262 5389
rect 3220 5331 3262 5369
rect 3336 5389 3378 5431
rect 3336 5369 3344 5389
rect 3364 5369 3378 5389
rect 3336 5331 3378 5369
rect 3428 5389 3472 5431
rect 3428 5369 3440 5389
rect 3460 5369 3472 5389
rect 3428 5331 3472 5369
rect 3544 5389 3586 5431
rect 3544 5369 3552 5389
rect 3572 5369 3586 5389
rect 3544 5331 3586 5369
rect 3636 5389 3680 5431
rect 3636 5369 3648 5389
rect 3668 5369 3680 5389
rect 3636 5331 3680 5369
rect 3757 5389 3799 5431
rect 3757 5369 3765 5389
rect 3785 5369 3799 5389
rect 3757 5331 3799 5369
rect 3849 5389 3893 5431
rect 3849 5369 3861 5389
rect 3881 5369 3893 5389
rect 3849 5331 3893 5369
rect 309 5174 353 5212
rect 309 5154 321 5174
rect 341 5154 353 5174
rect 309 5112 353 5154
rect 403 5174 445 5212
rect 403 5154 417 5174
rect 437 5154 445 5174
rect 403 5112 445 5154
rect 522 5174 566 5212
rect 522 5154 534 5174
rect 554 5154 566 5174
rect 522 5112 566 5154
rect 616 5174 658 5212
rect 616 5154 630 5174
rect 650 5154 658 5174
rect 616 5112 658 5154
rect 730 5174 774 5212
rect 730 5154 742 5174
rect 762 5154 774 5174
rect 730 5112 774 5154
rect 824 5174 866 5212
rect 824 5154 838 5174
rect 858 5154 866 5174
rect 824 5112 866 5154
rect 940 5174 982 5212
rect 940 5154 948 5174
rect 968 5154 982 5174
rect 940 5112 982 5154
rect 1032 5181 1077 5212
rect 4138 5208 4182 5250
rect 4138 5188 4150 5208
rect 4170 5188 4182 5208
rect 4138 5181 4182 5188
rect 1032 5174 1076 5181
rect 1032 5154 1044 5174
rect 1064 5154 1076 5174
rect 1032 5112 1076 5154
rect 4137 5150 4182 5181
rect 4232 5208 4274 5250
rect 4232 5188 4246 5208
rect 4266 5188 4274 5208
rect 4232 5150 4274 5188
rect 4348 5208 4390 5250
rect 4348 5188 4356 5208
rect 4376 5188 4390 5208
rect 4348 5150 4390 5188
rect 4440 5208 4484 5250
rect 4440 5188 4452 5208
rect 4472 5188 4484 5208
rect 4440 5150 4484 5188
rect 4556 5208 4598 5250
rect 4556 5188 4564 5208
rect 4584 5188 4598 5208
rect 4556 5150 4598 5188
rect 4648 5208 4692 5250
rect 4648 5188 4660 5208
rect 4680 5188 4692 5208
rect 4648 5150 4692 5188
rect 4769 5208 4811 5250
rect 4769 5188 4777 5208
rect 4797 5188 4811 5208
rect 4769 5150 4811 5188
rect 4861 5208 4905 5250
rect 4861 5188 4873 5208
rect 4893 5188 4905 5208
rect 4861 5150 4905 5188
rect 3076 4969 3120 5011
rect 3076 4949 3088 4969
rect 3108 4949 3120 4969
rect 3076 4942 3120 4949
rect 3075 4911 3120 4942
rect 3170 4969 3212 5011
rect 3170 4949 3184 4969
rect 3204 4949 3212 4969
rect 3170 4911 3212 4949
rect 3286 4969 3328 5011
rect 3286 4949 3294 4969
rect 3314 4949 3328 4969
rect 3286 4911 3328 4949
rect 3378 4969 3422 5011
rect 3378 4949 3390 4969
rect 3410 4949 3422 4969
rect 3378 4911 3422 4949
rect 3494 4969 3536 5011
rect 3494 4949 3502 4969
rect 3522 4949 3536 4969
rect 3494 4911 3536 4949
rect 3586 4969 3630 5011
rect 3586 4949 3598 4969
rect 3618 4949 3630 4969
rect 3586 4911 3630 4949
rect 3707 4969 3749 5011
rect 3707 4949 3715 4969
rect 3735 4949 3749 4969
rect 3707 4911 3749 4949
rect 3799 4969 3843 5011
rect 3799 4949 3811 4969
rect 3831 4949 3843 4969
rect 3799 4911 3843 4949
rect 1377 4847 1421 4885
rect 1377 4827 1389 4847
rect 1409 4827 1421 4847
rect 1377 4785 1421 4827
rect 1471 4847 1513 4885
rect 1471 4827 1485 4847
rect 1505 4827 1513 4847
rect 1471 4785 1513 4827
rect 1590 4847 1634 4885
rect 1590 4827 1602 4847
rect 1622 4827 1634 4847
rect 1590 4785 1634 4827
rect 1684 4847 1726 4885
rect 1684 4827 1698 4847
rect 1718 4827 1726 4847
rect 1684 4785 1726 4827
rect 1798 4847 1842 4885
rect 1798 4827 1810 4847
rect 1830 4827 1842 4847
rect 1798 4785 1842 4827
rect 1892 4847 1934 4885
rect 1892 4827 1906 4847
rect 1926 4827 1934 4847
rect 1892 4785 1934 4827
rect 2008 4847 2050 4885
rect 2008 4827 2016 4847
rect 2036 4827 2050 4847
rect 2008 4785 2050 4827
rect 2100 4854 2145 4885
rect 2100 4847 2144 4854
rect 2100 4827 2112 4847
rect 2132 4827 2144 4847
rect 2100 4785 2144 4827
rect 315 4608 359 4646
rect 315 4588 327 4608
rect 347 4588 359 4608
rect 315 4546 359 4588
rect 409 4608 451 4646
rect 409 4588 423 4608
rect 443 4588 451 4608
rect 409 4546 451 4588
rect 528 4608 572 4646
rect 528 4588 540 4608
rect 560 4588 572 4608
rect 528 4546 572 4588
rect 622 4608 664 4646
rect 622 4588 636 4608
rect 656 4588 664 4608
rect 622 4546 664 4588
rect 736 4608 780 4646
rect 736 4588 748 4608
rect 768 4588 780 4608
rect 736 4546 780 4588
rect 830 4608 872 4646
rect 830 4588 844 4608
rect 864 4588 872 4608
rect 830 4546 872 4588
rect 946 4608 988 4646
rect 946 4588 954 4608
rect 974 4588 988 4608
rect 946 4546 988 4588
rect 1038 4615 1083 4646
rect 4144 4642 4188 4684
rect 4144 4622 4156 4642
rect 4176 4622 4188 4642
rect 4144 4615 4188 4622
rect 1038 4608 1082 4615
rect 1038 4588 1050 4608
rect 1070 4588 1082 4608
rect 1038 4546 1082 4588
rect 4143 4584 4188 4615
rect 4238 4642 4280 4684
rect 4238 4622 4252 4642
rect 4272 4622 4280 4642
rect 4238 4584 4280 4622
rect 4354 4642 4396 4684
rect 4354 4622 4362 4642
rect 4382 4622 4396 4642
rect 4354 4584 4396 4622
rect 4446 4642 4490 4684
rect 4446 4622 4458 4642
rect 4478 4622 4490 4642
rect 4446 4584 4490 4622
rect 4562 4642 4604 4684
rect 4562 4622 4570 4642
rect 4590 4622 4604 4642
rect 4562 4584 4604 4622
rect 4654 4642 4698 4684
rect 4654 4622 4666 4642
rect 4686 4622 4698 4642
rect 4654 4584 4698 4622
rect 4775 4642 4817 4684
rect 4775 4622 4783 4642
rect 4803 4622 4817 4642
rect 4775 4584 4817 4622
rect 4867 4642 4911 4684
rect 4867 4622 4879 4642
rect 4899 4622 4911 4642
rect 4867 4584 4911 4622
rect 1327 4427 1371 4465
rect 1327 4407 1339 4427
rect 1359 4407 1371 4427
rect 1327 4365 1371 4407
rect 1421 4427 1463 4465
rect 1421 4407 1435 4427
rect 1455 4407 1463 4427
rect 1421 4365 1463 4407
rect 1540 4427 1584 4465
rect 1540 4407 1552 4427
rect 1572 4407 1584 4427
rect 1540 4365 1584 4407
rect 1634 4427 1676 4465
rect 1634 4407 1648 4427
rect 1668 4407 1676 4427
rect 1634 4365 1676 4407
rect 1748 4427 1792 4465
rect 1748 4407 1760 4427
rect 1780 4407 1792 4427
rect 1748 4365 1792 4407
rect 1842 4427 1884 4465
rect 1842 4407 1856 4427
rect 1876 4407 1884 4427
rect 1842 4365 1884 4407
rect 1958 4427 2000 4465
rect 1958 4407 1966 4427
rect 1986 4407 2000 4427
rect 1958 4365 2000 4407
rect 2050 4434 2095 4465
rect 2050 4427 2094 4434
rect 2050 4407 2062 4427
rect 2082 4407 2094 4427
rect 2050 4365 2094 4407
rect 3131 4408 3175 4450
rect 3131 4388 3143 4408
rect 3163 4388 3175 4408
rect 3131 4381 3175 4388
rect 3130 4350 3175 4381
rect 3225 4408 3267 4450
rect 3225 4388 3239 4408
rect 3259 4388 3267 4408
rect 3225 4350 3267 4388
rect 3341 4408 3383 4450
rect 3341 4388 3349 4408
rect 3369 4388 3383 4408
rect 3341 4350 3383 4388
rect 3433 4408 3477 4450
rect 3433 4388 3445 4408
rect 3465 4388 3477 4408
rect 3433 4350 3477 4388
rect 3549 4408 3591 4450
rect 3549 4388 3557 4408
rect 3577 4388 3591 4408
rect 3549 4350 3591 4388
rect 3641 4408 3685 4450
rect 3641 4388 3653 4408
rect 3673 4388 3685 4408
rect 3641 4350 3685 4388
rect 3762 4408 3804 4450
rect 3762 4388 3770 4408
rect 3790 4388 3804 4408
rect 3762 4350 3804 4388
rect 3854 4408 3898 4450
rect 3854 4388 3866 4408
rect 3886 4388 3898 4408
rect 3854 4350 3898 4388
rect 314 4193 358 4231
rect 314 4173 326 4193
rect 346 4173 358 4193
rect 314 4131 358 4173
rect 408 4193 450 4231
rect 408 4173 422 4193
rect 442 4173 450 4193
rect 408 4131 450 4173
rect 527 4193 571 4231
rect 527 4173 539 4193
rect 559 4173 571 4193
rect 527 4131 571 4173
rect 621 4193 663 4231
rect 621 4173 635 4193
rect 655 4173 663 4193
rect 621 4131 663 4173
rect 735 4193 779 4231
rect 735 4173 747 4193
rect 767 4173 779 4193
rect 735 4131 779 4173
rect 829 4193 871 4231
rect 829 4173 843 4193
rect 863 4173 871 4193
rect 829 4131 871 4173
rect 945 4193 987 4231
rect 945 4173 953 4193
rect 973 4173 987 4193
rect 945 4131 987 4173
rect 1037 4200 1082 4231
rect 4143 4227 4187 4269
rect 4143 4207 4155 4227
rect 4175 4207 4187 4227
rect 4143 4200 4187 4207
rect 1037 4193 1081 4200
rect 1037 4173 1049 4193
rect 1069 4173 1081 4193
rect 1037 4131 1081 4173
rect 4142 4169 4187 4200
rect 4237 4227 4279 4269
rect 4237 4207 4251 4227
rect 4271 4207 4279 4227
rect 4237 4169 4279 4207
rect 4353 4227 4395 4269
rect 4353 4207 4361 4227
rect 4381 4207 4395 4227
rect 4353 4169 4395 4207
rect 4445 4227 4489 4269
rect 4445 4207 4457 4227
rect 4477 4207 4489 4227
rect 4445 4169 4489 4207
rect 4561 4227 4603 4269
rect 4561 4207 4569 4227
rect 4589 4207 4603 4227
rect 4561 4169 4603 4207
rect 4653 4227 4697 4269
rect 4653 4207 4665 4227
rect 4685 4207 4697 4227
rect 4653 4169 4697 4207
rect 4774 4227 4816 4269
rect 4774 4207 4782 4227
rect 4802 4207 4816 4227
rect 4774 4169 4816 4207
rect 4866 4227 4910 4269
rect 4866 4207 4878 4227
rect 4898 4207 4910 4227
rect 4866 4169 4910 4207
rect 2836 3976 2880 4018
rect 2836 3956 2848 3976
rect 2868 3956 2880 3976
rect 2836 3949 2880 3956
rect 1625 3883 1669 3921
rect 1625 3863 1637 3883
rect 1657 3863 1669 3883
rect 1625 3821 1669 3863
rect 1719 3883 1761 3921
rect 1719 3863 1733 3883
rect 1753 3863 1761 3883
rect 1719 3821 1761 3863
rect 1838 3883 1882 3921
rect 1838 3863 1850 3883
rect 1870 3863 1882 3883
rect 1838 3821 1882 3863
rect 1932 3883 1974 3921
rect 1932 3863 1946 3883
rect 1966 3863 1974 3883
rect 1932 3821 1974 3863
rect 2046 3883 2090 3921
rect 2046 3863 2058 3883
rect 2078 3863 2090 3883
rect 2046 3821 2090 3863
rect 2140 3883 2182 3921
rect 2140 3863 2154 3883
rect 2174 3863 2182 3883
rect 2140 3821 2182 3863
rect 2256 3883 2298 3921
rect 2256 3863 2264 3883
rect 2284 3863 2298 3883
rect 2256 3821 2298 3863
rect 2348 3890 2393 3921
rect 2835 3918 2880 3949
rect 2930 3976 2972 4018
rect 2930 3956 2944 3976
rect 2964 3956 2972 3976
rect 2930 3918 2972 3956
rect 3046 3976 3088 4018
rect 3046 3956 3054 3976
rect 3074 3956 3088 3976
rect 3046 3918 3088 3956
rect 3138 3976 3182 4018
rect 3138 3956 3150 3976
rect 3170 3956 3182 3976
rect 3138 3918 3182 3956
rect 3254 3976 3296 4018
rect 3254 3956 3262 3976
rect 3282 3956 3296 3976
rect 3254 3918 3296 3956
rect 3346 3976 3390 4018
rect 3346 3956 3358 3976
rect 3378 3956 3390 3976
rect 3346 3918 3390 3956
rect 3467 3976 3509 4018
rect 3467 3956 3475 3976
rect 3495 3956 3509 3976
rect 3467 3918 3509 3956
rect 3559 3976 3603 4018
rect 3559 3956 3571 3976
rect 3591 3956 3603 3976
rect 3559 3918 3603 3956
rect 2348 3883 2392 3890
rect 2348 3863 2360 3883
rect 2380 3863 2392 3883
rect 2348 3821 2392 3863
rect 318 3632 362 3670
rect 318 3612 330 3632
rect 350 3612 362 3632
rect 318 3570 362 3612
rect 412 3632 454 3670
rect 412 3612 426 3632
rect 446 3612 454 3632
rect 412 3570 454 3612
rect 531 3632 575 3670
rect 531 3612 543 3632
rect 563 3612 575 3632
rect 531 3570 575 3612
rect 625 3632 667 3670
rect 625 3612 639 3632
rect 659 3612 667 3632
rect 625 3570 667 3612
rect 739 3632 783 3670
rect 739 3612 751 3632
rect 771 3612 783 3632
rect 739 3570 783 3612
rect 833 3632 875 3670
rect 833 3612 847 3632
rect 867 3612 875 3632
rect 833 3570 875 3612
rect 949 3632 991 3670
rect 949 3612 957 3632
rect 977 3612 991 3632
rect 949 3570 991 3612
rect 1041 3639 1086 3670
rect 4147 3666 4191 3708
rect 4147 3646 4159 3666
rect 4179 3646 4191 3666
rect 4147 3639 4191 3646
rect 1041 3632 1085 3639
rect 1041 3612 1053 3632
rect 1073 3612 1085 3632
rect 1041 3570 1085 3612
rect 4146 3608 4191 3639
rect 4241 3666 4283 3708
rect 4241 3646 4255 3666
rect 4275 3646 4283 3666
rect 4241 3608 4283 3646
rect 4357 3666 4399 3708
rect 4357 3646 4365 3666
rect 4385 3646 4399 3666
rect 4357 3608 4399 3646
rect 4449 3666 4493 3708
rect 4449 3646 4461 3666
rect 4481 3646 4493 3666
rect 4449 3608 4493 3646
rect 4565 3666 4607 3708
rect 4565 3646 4573 3666
rect 4593 3646 4607 3666
rect 4565 3608 4607 3646
rect 4657 3666 4701 3708
rect 4657 3646 4669 3666
rect 4689 3646 4701 3666
rect 4657 3608 4701 3646
rect 4778 3666 4820 3708
rect 4778 3646 4786 3666
rect 4806 3646 4820 3666
rect 4778 3608 4820 3646
rect 4870 3666 4914 3708
rect 4870 3646 4882 3666
rect 4902 3646 4914 3666
rect 4870 3608 4914 3646
rect 1330 3451 1374 3489
rect 1330 3431 1342 3451
rect 1362 3431 1374 3451
rect 1330 3389 1374 3431
rect 1424 3451 1466 3489
rect 1424 3431 1438 3451
rect 1458 3431 1466 3451
rect 1424 3389 1466 3431
rect 1543 3451 1587 3489
rect 1543 3431 1555 3451
rect 1575 3431 1587 3451
rect 1543 3389 1587 3431
rect 1637 3451 1679 3489
rect 1637 3431 1651 3451
rect 1671 3431 1679 3451
rect 1637 3389 1679 3431
rect 1751 3451 1795 3489
rect 1751 3431 1763 3451
rect 1783 3431 1795 3451
rect 1751 3389 1795 3431
rect 1845 3451 1887 3489
rect 1845 3431 1859 3451
rect 1879 3431 1887 3451
rect 1845 3389 1887 3431
rect 1961 3451 2003 3489
rect 1961 3431 1969 3451
rect 1989 3431 2003 3451
rect 1961 3389 2003 3431
rect 2053 3458 2098 3489
rect 2053 3451 2097 3458
rect 2053 3431 2065 3451
rect 2085 3431 2097 3451
rect 2053 3389 2097 3431
rect 3134 3432 3178 3474
rect 3134 3412 3146 3432
rect 3166 3412 3178 3432
rect 3134 3405 3178 3412
rect 3133 3374 3178 3405
rect 3228 3432 3270 3474
rect 3228 3412 3242 3432
rect 3262 3412 3270 3432
rect 3228 3374 3270 3412
rect 3344 3432 3386 3474
rect 3344 3412 3352 3432
rect 3372 3412 3386 3432
rect 3344 3374 3386 3412
rect 3436 3432 3480 3474
rect 3436 3412 3448 3432
rect 3468 3412 3480 3432
rect 3436 3374 3480 3412
rect 3552 3432 3594 3474
rect 3552 3412 3560 3432
rect 3580 3412 3594 3432
rect 3552 3374 3594 3412
rect 3644 3432 3688 3474
rect 3644 3412 3656 3432
rect 3676 3412 3688 3432
rect 3644 3374 3688 3412
rect 3765 3432 3807 3474
rect 3765 3412 3773 3432
rect 3793 3412 3807 3432
rect 3765 3374 3807 3412
rect 3857 3432 3901 3474
rect 3857 3412 3869 3432
rect 3889 3412 3901 3432
rect 3857 3374 3901 3412
rect 317 3217 361 3255
rect 317 3197 329 3217
rect 349 3197 361 3217
rect 317 3155 361 3197
rect 411 3217 453 3255
rect 411 3197 425 3217
rect 445 3197 453 3217
rect 411 3155 453 3197
rect 530 3217 574 3255
rect 530 3197 542 3217
rect 562 3197 574 3217
rect 530 3155 574 3197
rect 624 3217 666 3255
rect 624 3197 638 3217
rect 658 3197 666 3217
rect 624 3155 666 3197
rect 738 3217 782 3255
rect 738 3197 750 3217
rect 770 3197 782 3217
rect 738 3155 782 3197
rect 832 3217 874 3255
rect 832 3197 846 3217
rect 866 3197 874 3217
rect 832 3155 874 3197
rect 948 3217 990 3255
rect 948 3197 956 3217
rect 976 3197 990 3217
rect 948 3155 990 3197
rect 1040 3224 1085 3255
rect 4146 3251 4190 3293
rect 4146 3231 4158 3251
rect 4178 3231 4190 3251
rect 4146 3224 4190 3231
rect 1040 3217 1084 3224
rect 1040 3197 1052 3217
rect 1072 3197 1084 3217
rect 1040 3155 1084 3197
rect 4145 3193 4190 3224
rect 4240 3251 4282 3293
rect 4240 3231 4254 3251
rect 4274 3231 4282 3251
rect 4240 3193 4282 3231
rect 4356 3251 4398 3293
rect 4356 3231 4364 3251
rect 4384 3231 4398 3251
rect 4356 3193 4398 3231
rect 4448 3251 4492 3293
rect 4448 3231 4460 3251
rect 4480 3231 4492 3251
rect 4448 3193 4492 3231
rect 4564 3251 4606 3293
rect 4564 3231 4572 3251
rect 4592 3231 4606 3251
rect 4564 3193 4606 3231
rect 4656 3251 4700 3293
rect 4656 3231 4668 3251
rect 4688 3231 4700 3251
rect 4656 3193 4700 3231
rect 4777 3251 4819 3293
rect 4777 3231 4785 3251
rect 4805 3231 4819 3251
rect 4777 3193 4819 3231
rect 4869 3251 4913 3293
rect 4869 3231 4881 3251
rect 4901 3231 4913 3251
rect 4869 3193 4913 3231
rect 3084 3012 3128 3054
rect 3084 2992 3096 3012
rect 3116 2992 3128 3012
rect 3084 2985 3128 2992
rect 3083 2954 3128 2985
rect 3178 3012 3220 3054
rect 3178 2992 3192 3012
rect 3212 2992 3220 3012
rect 3178 2954 3220 2992
rect 3294 3012 3336 3054
rect 3294 2992 3302 3012
rect 3322 2992 3336 3012
rect 3294 2954 3336 2992
rect 3386 3012 3430 3054
rect 3386 2992 3398 3012
rect 3418 2992 3430 3012
rect 3386 2954 3430 2992
rect 3502 3012 3544 3054
rect 3502 2992 3510 3012
rect 3530 2992 3544 3012
rect 3502 2954 3544 2992
rect 3594 3012 3638 3054
rect 3594 2992 3606 3012
rect 3626 2992 3638 3012
rect 3594 2954 3638 2992
rect 3715 3012 3757 3054
rect 3715 2992 3723 3012
rect 3743 2992 3757 3012
rect 3715 2954 3757 2992
rect 3807 3012 3851 3054
rect 3807 2992 3819 3012
rect 3839 2992 3851 3012
rect 3807 2954 3851 2992
rect 1385 2890 1429 2928
rect 1385 2870 1397 2890
rect 1417 2870 1429 2890
rect 1385 2828 1429 2870
rect 1479 2890 1521 2928
rect 1479 2870 1493 2890
rect 1513 2870 1521 2890
rect 1479 2828 1521 2870
rect 1598 2890 1642 2928
rect 1598 2870 1610 2890
rect 1630 2870 1642 2890
rect 1598 2828 1642 2870
rect 1692 2890 1734 2928
rect 1692 2870 1706 2890
rect 1726 2870 1734 2890
rect 1692 2828 1734 2870
rect 1806 2890 1850 2928
rect 1806 2870 1818 2890
rect 1838 2870 1850 2890
rect 1806 2828 1850 2870
rect 1900 2890 1942 2928
rect 1900 2870 1914 2890
rect 1934 2870 1942 2890
rect 1900 2828 1942 2870
rect 2016 2890 2058 2928
rect 2016 2870 2024 2890
rect 2044 2870 2058 2890
rect 2016 2828 2058 2870
rect 2108 2897 2153 2928
rect 2108 2890 2152 2897
rect 2108 2870 2120 2890
rect 2140 2870 2152 2890
rect 2108 2828 2152 2870
rect 323 2651 367 2689
rect 323 2631 335 2651
rect 355 2631 367 2651
rect 323 2589 367 2631
rect 417 2651 459 2689
rect 417 2631 431 2651
rect 451 2631 459 2651
rect 417 2589 459 2631
rect 536 2651 580 2689
rect 536 2631 548 2651
rect 568 2631 580 2651
rect 536 2589 580 2631
rect 630 2651 672 2689
rect 630 2631 644 2651
rect 664 2631 672 2651
rect 630 2589 672 2631
rect 744 2651 788 2689
rect 744 2631 756 2651
rect 776 2631 788 2651
rect 744 2589 788 2631
rect 838 2651 880 2689
rect 838 2631 852 2651
rect 872 2631 880 2651
rect 838 2589 880 2631
rect 954 2651 996 2689
rect 954 2631 962 2651
rect 982 2631 996 2651
rect 954 2589 996 2631
rect 1046 2658 1091 2689
rect 4152 2685 4196 2727
rect 4152 2665 4164 2685
rect 4184 2665 4196 2685
rect 4152 2658 4196 2665
rect 1046 2651 1090 2658
rect 1046 2631 1058 2651
rect 1078 2631 1090 2651
rect 1046 2589 1090 2631
rect 4151 2627 4196 2658
rect 4246 2685 4288 2727
rect 4246 2665 4260 2685
rect 4280 2665 4288 2685
rect 4246 2627 4288 2665
rect 4362 2685 4404 2727
rect 4362 2665 4370 2685
rect 4390 2665 4404 2685
rect 4362 2627 4404 2665
rect 4454 2685 4498 2727
rect 4454 2665 4466 2685
rect 4486 2665 4498 2685
rect 4454 2627 4498 2665
rect 4570 2685 4612 2727
rect 4570 2665 4578 2685
rect 4598 2665 4612 2685
rect 4570 2627 4612 2665
rect 4662 2685 4706 2727
rect 4662 2665 4674 2685
rect 4694 2665 4706 2685
rect 4662 2627 4706 2665
rect 4783 2685 4825 2727
rect 4783 2665 4791 2685
rect 4811 2665 4825 2685
rect 4783 2627 4825 2665
rect 4875 2685 4919 2727
rect 4875 2665 4887 2685
rect 4907 2665 4919 2685
rect 4875 2627 4919 2665
rect 1335 2470 1379 2508
rect 1335 2450 1347 2470
rect 1367 2450 1379 2470
rect 1335 2408 1379 2450
rect 1429 2470 1471 2508
rect 1429 2450 1443 2470
rect 1463 2450 1471 2470
rect 1429 2408 1471 2450
rect 1548 2470 1592 2508
rect 1548 2450 1560 2470
rect 1580 2450 1592 2470
rect 1548 2408 1592 2450
rect 1642 2470 1684 2508
rect 1642 2450 1656 2470
rect 1676 2450 1684 2470
rect 1642 2408 1684 2450
rect 1756 2470 1800 2508
rect 1756 2450 1768 2470
rect 1788 2450 1800 2470
rect 1756 2408 1800 2450
rect 1850 2470 1892 2508
rect 1850 2450 1864 2470
rect 1884 2450 1892 2470
rect 1850 2408 1892 2450
rect 1966 2470 2008 2508
rect 1966 2450 1974 2470
rect 1994 2450 2008 2470
rect 1966 2408 2008 2450
rect 2058 2477 2103 2508
rect 2058 2470 2102 2477
rect 2058 2450 2070 2470
rect 2090 2450 2102 2470
rect 2058 2408 2102 2450
rect 3139 2451 3183 2493
rect 3139 2431 3151 2451
rect 3171 2431 3183 2451
rect 3139 2424 3183 2431
rect 3138 2393 3183 2424
rect 3233 2451 3275 2493
rect 3233 2431 3247 2451
rect 3267 2431 3275 2451
rect 3233 2393 3275 2431
rect 3349 2451 3391 2493
rect 3349 2431 3357 2451
rect 3377 2431 3391 2451
rect 3349 2393 3391 2431
rect 3441 2451 3485 2493
rect 3441 2431 3453 2451
rect 3473 2431 3485 2451
rect 3441 2393 3485 2431
rect 3557 2451 3599 2493
rect 3557 2431 3565 2451
rect 3585 2431 3599 2451
rect 3557 2393 3599 2431
rect 3649 2451 3693 2493
rect 3649 2431 3661 2451
rect 3681 2431 3693 2451
rect 3649 2393 3693 2431
rect 3770 2451 3812 2493
rect 3770 2431 3778 2451
rect 3798 2431 3812 2451
rect 3770 2393 3812 2431
rect 3862 2451 3906 2493
rect 3862 2431 3874 2451
rect 3894 2431 3906 2451
rect 3862 2393 3906 2431
rect 322 2236 366 2274
rect 322 2216 334 2236
rect 354 2216 366 2236
rect 322 2174 366 2216
rect 416 2236 458 2274
rect 416 2216 430 2236
rect 450 2216 458 2236
rect 416 2174 458 2216
rect 535 2236 579 2274
rect 535 2216 547 2236
rect 567 2216 579 2236
rect 535 2174 579 2216
rect 629 2236 671 2274
rect 629 2216 643 2236
rect 663 2216 671 2236
rect 629 2174 671 2216
rect 743 2236 787 2274
rect 743 2216 755 2236
rect 775 2216 787 2236
rect 743 2174 787 2216
rect 837 2236 879 2274
rect 837 2216 851 2236
rect 871 2216 879 2236
rect 837 2174 879 2216
rect 953 2236 995 2274
rect 953 2216 961 2236
rect 981 2216 995 2236
rect 953 2174 995 2216
rect 1045 2243 1090 2274
rect 4151 2270 4195 2312
rect 4151 2250 4163 2270
rect 4183 2250 4195 2270
rect 4151 2243 4195 2250
rect 1045 2236 1089 2243
rect 1045 2216 1057 2236
rect 1077 2216 1089 2236
rect 1045 2174 1089 2216
rect 4150 2212 4195 2243
rect 4245 2270 4287 2312
rect 4245 2250 4259 2270
rect 4279 2250 4287 2270
rect 4245 2212 4287 2250
rect 4361 2270 4403 2312
rect 4361 2250 4369 2270
rect 4389 2250 4403 2270
rect 4361 2212 4403 2250
rect 4453 2270 4497 2312
rect 4453 2250 4465 2270
rect 4485 2250 4497 2270
rect 4453 2212 4497 2250
rect 4569 2270 4611 2312
rect 4569 2250 4577 2270
rect 4597 2250 4611 2270
rect 4569 2212 4611 2250
rect 4661 2270 4705 2312
rect 4661 2250 4673 2270
rect 4693 2250 4705 2270
rect 4661 2212 4705 2250
rect 4782 2270 4824 2312
rect 4782 2250 4790 2270
rect 4810 2250 4824 2270
rect 4782 2212 4824 2250
rect 4874 2270 4918 2312
rect 4874 2250 4886 2270
rect 4906 2250 4918 2270
rect 4874 2212 4918 2250
rect 1550 1958 1594 1996
rect 1550 1938 1562 1958
rect 1582 1938 1594 1958
rect 1550 1896 1594 1938
rect 1644 1958 1686 1996
rect 1644 1938 1658 1958
rect 1678 1938 1686 1958
rect 1644 1896 1686 1938
rect 1763 1958 1807 1996
rect 1763 1938 1775 1958
rect 1795 1938 1807 1958
rect 1763 1896 1807 1938
rect 1857 1958 1899 1996
rect 1857 1938 1871 1958
rect 1891 1938 1899 1958
rect 1857 1896 1899 1938
rect 1971 1958 2015 1996
rect 1971 1938 1983 1958
rect 2003 1938 2015 1958
rect 1971 1896 2015 1938
rect 2065 1958 2107 1996
rect 2065 1938 2079 1958
rect 2099 1938 2107 1958
rect 2065 1896 2107 1938
rect 2181 1958 2223 1996
rect 2181 1938 2189 1958
rect 2209 1938 2223 1958
rect 2181 1896 2223 1938
rect 2273 1965 2318 1996
rect 2931 1984 2975 2026
rect 2273 1958 2317 1965
rect 2273 1938 2285 1958
rect 2305 1938 2317 1958
rect 2931 1964 2943 1984
rect 2963 1964 2975 1984
rect 2931 1957 2975 1964
rect 2273 1896 2317 1938
rect 2930 1926 2975 1957
rect 3025 1984 3067 2026
rect 3025 1964 3039 1984
rect 3059 1964 3067 1984
rect 3025 1926 3067 1964
rect 3141 1984 3183 2026
rect 3141 1964 3149 1984
rect 3169 1964 3183 1984
rect 3141 1926 3183 1964
rect 3233 1984 3277 2026
rect 3233 1964 3245 1984
rect 3265 1964 3277 1984
rect 3233 1926 3277 1964
rect 3349 1984 3391 2026
rect 3349 1964 3357 1984
rect 3377 1964 3391 1984
rect 3349 1926 3391 1964
rect 3441 1984 3485 2026
rect 3441 1964 3453 1984
rect 3473 1964 3485 1984
rect 3441 1926 3485 1964
rect 3562 1984 3604 2026
rect 3562 1964 3570 1984
rect 3590 1964 3604 1984
rect 3562 1926 3604 1964
rect 3654 1984 3698 2026
rect 3654 1964 3666 1984
rect 3686 1964 3698 1984
rect 3654 1926 3698 1964
rect 330 1672 374 1710
rect 330 1652 342 1672
rect 362 1652 374 1672
rect 330 1610 374 1652
rect 424 1672 466 1710
rect 424 1652 438 1672
rect 458 1652 466 1672
rect 424 1610 466 1652
rect 543 1672 587 1710
rect 543 1652 555 1672
rect 575 1652 587 1672
rect 543 1610 587 1652
rect 637 1672 679 1710
rect 637 1652 651 1672
rect 671 1652 679 1672
rect 637 1610 679 1652
rect 751 1672 795 1710
rect 751 1652 763 1672
rect 783 1652 795 1672
rect 751 1610 795 1652
rect 845 1672 887 1710
rect 845 1652 859 1672
rect 879 1652 887 1672
rect 845 1610 887 1652
rect 961 1672 1003 1710
rect 961 1652 969 1672
rect 989 1652 1003 1672
rect 961 1610 1003 1652
rect 1053 1679 1098 1710
rect 4159 1706 4203 1748
rect 4159 1686 4171 1706
rect 4191 1686 4203 1706
rect 4159 1679 4203 1686
rect 1053 1672 1097 1679
rect 1053 1652 1065 1672
rect 1085 1652 1097 1672
rect 1053 1610 1097 1652
rect 4158 1648 4203 1679
rect 4253 1706 4295 1748
rect 4253 1686 4267 1706
rect 4287 1686 4295 1706
rect 4253 1648 4295 1686
rect 4369 1706 4411 1748
rect 4369 1686 4377 1706
rect 4397 1686 4411 1706
rect 4369 1648 4411 1686
rect 4461 1706 4505 1748
rect 4461 1686 4473 1706
rect 4493 1686 4505 1706
rect 4461 1648 4505 1686
rect 4577 1706 4619 1748
rect 4577 1686 4585 1706
rect 4605 1686 4619 1706
rect 4577 1648 4619 1686
rect 4669 1706 4713 1748
rect 4669 1686 4681 1706
rect 4701 1686 4713 1706
rect 4669 1648 4713 1686
rect 4790 1706 4832 1748
rect 4790 1686 4798 1706
rect 4818 1686 4832 1706
rect 4790 1648 4832 1686
rect 4882 1706 4926 1748
rect 4882 1686 4894 1706
rect 4914 1686 4926 1706
rect 4882 1648 4926 1686
rect 1342 1491 1386 1529
rect 1342 1471 1354 1491
rect 1374 1471 1386 1491
rect 1342 1429 1386 1471
rect 1436 1491 1478 1529
rect 1436 1471 1450 1491
rect 1470 1471 1478 1491
rect 1436 1429 1478 1471
rect 1555 1491 1599 1529
rect 1555 1471 1567 1491
rect 1587 1471 1599 1491
rect 1555 1429 1599 1471
rect 1649 1491 1691 1529
rect 1649 1471 1663 1491
rect 1683 1471 1691 1491
rect 1649 1429 1691 1471
rect 1763 1491 1807 1529
rect 1763 1471 1775 1491
rect 1795 1471 1807 1491
rect 1763 1429 1807 1471
rect 1857 1491 1899 1529
rect 1857 1471 1871 1491
rect 1891 1471 1899 1491
rect 1857 1429 1899 1471
rect 1973 1491 2015 1529
rect 1973 1471 1981 1491
rect 2001 1471 2015 1491
rect 1973 1429 2015 1471
rect 2065 1498 2110 1529
rect 2065 1491 2109 1498
rect 2065 1471 2077 1491
rect 2097 1471 2109 1491
rect 2065 1429 2109 1471
rect 3146 1472 3190 1514
rect 3146 1452 3158 1472
rect 3178 1452 3190 1472
rect 3146 1445 3190 1452
rect 3145 1414 3190 1445
rect 3240 1472 3282 1514
rect 3240 1452 3254 1472
rect 3274 1452 3282 1472
rect 3240 1414 3282 1452
rect 3356 1472 3398 1514
rect 3356 1452 3364 1472
rect 3384 1452 3398 1472
rect 3356 1414 3398 1452
rect 3448 1472 3492 1514
rect 3448 1452 3460 1472
rect 3480 1452 3492 1472
rect 3448 1414 3492 1452
rect 3564 1472 3606 1514
rect 3564 1452 3572 1472
rect 3592 1452 3606 1472
rect 3564 1414 3606 1452
rect 3656 1472 3700 1514
rect 3656 1452 3668 1472
rect 3688 1452 3700 1472
rect 3656 1414 3700 1452
rect 3777 1472 3819 1514
rect 3777 1452 3785 1472
rect 3805 1452 3819 1472
rect 3777 1414 3819 1452
rect 3869 1472 3913 1514
rect 3869 1452 3881 1472
rect 3901 1452 3913 1472
rect 3869 1414 3913 1452
rect 329 1257 373 1295
rect 329 1237 341 1257
rect 361 1237 373 1257
rect 329 1195 373 1237
rect 423 1257 465 1295
rect 423 1237 437 1257
rect 457 1237 465 1257
rect 423 1195 465 1237
rect 542 1257 586 1295
rect 542 1237 554 1257
rect 574 1237 586 1257
rect 542 1195 586 1237
rect 636 1257 678 1295
rect 636 1237 650 1257
rect 670 1237 678 1257
rect 636 1195 678 1237
rect 750 1257 794 1295
rect 750 1237 762 1257
rect 782 1237 794 1257
rect 750 1195 794 1237
rect 844 1257 886 1295
rect 844 1237 858 1257
rect 878 1237 886 1257
rect 844 1195 886 1237
rect 960 1257 1002 1295
rect 960 1237 968 1257
rect 988 1237 1002 1257
rect 960 1195 1002 1237
rect 1052 1264 1097 1295
rect 4158 1291 4202 1333
rect 4158 1271 4170 1291
rect 4190 1271 4202 1291
rect 4158 1264 4202 1271
rect 1052 1257 1096 1264
rect 1052 1237 1064 1257
rect 1084 1237 1096 1257
rect 1052 1195 1096 1237
rect 4157 1233 4202 1264
rect 4252 1291 4294 1333
rect 4252 1271 4266 1291
rect 4286 1271 4294 1291
rect 4252 1233 4294 1271
rect 4368 1291 4410 1333
rect 4368 1271 4376 1291
rect 4396 1271 4410 1291
rect 4368 1233 4410 1271
rect 4460 1291 4504 1333
rect 4460 1271 4472 1291
rect 4492 1271 4504 1291
rect 4460 1233 4504 1271
rect 4576 1291 4618 1333
rect 4576 1271 4584 1291
rect 4604 1271 4618 1291
rect 4576 1233 4618 1271
rect 4668 1291 4712 1333
rect 4668 1271 4680 1291
rect 4700 1271 4712 1291
rect 4668 1233 4712 1271
rect 4789 1291 4831 1333
rect 4789 1271 4797 1291
rect 4817 1271 4831 1291
rect 4789 1233 4831 1271
rect 4881 1291 4925 1333
rect 4881 1271 4893 1291
rect 4913 1271 4925 1291
rect 4881 1233 4925 1271
rect 3096 1052 3140 1094
rect 3096 1032 3108 1052
rect 3128 1032 3140 1052
rect 3096 1025 3140 1032
rect 3095 994 3140 1025
rect 3190 1052 3232 1094
rect 3190 1032 3204 1052
rect 3224 1032 3232 1052
rect 3190 994 3232 1032
rect 3306 1052 3348 1094
rect 3306 1032 3314 1052
rect 3334 1032 3348 1052
rect 3306 994 3348 1032
rect 3398 1052 3442 1094
rect 3398 1032 3410 1052
rect 3430 1032 3442 1052
rect 3398 994 3442 1032
rect 3514 1052 3556 1094
rect 3514 1032 3522 1052
rect 3542 1032 3556 1052
rect 3514 994 3556 1032
rect 3606 1052 3650 1094
rect 3606 1032 3618 1052
rect 3638 1032 3650 1052
rect 3606 994 3650 1032
rect 3727 1052 3769 1094
rect 3727 1032 3735 1052
rect 3755 1032 3769 1052
rect 3727 994 3769 1032
rect 3819 1052 3863 1094
rect 3819 1032 3831 1052
rect 3851 1032 3863 1052
rect 3819 994 3863 1032
rect 1397 930 1441 968
rect 1397 910 1409 930
rect 1429 910 1441 930
rect 1397 868 1441 910
rect 1491 930 1533 968
rect 1491 910 1505 930
rect 1525 910 1533 930
rect 1491 868 1533 910
rect 1610 930 1654 968
rect 1610 910 1622 930
rect 1642 910 1654 930
rect 1610 868 1654 910
rect 1704 930 1746 968
rect 1704 910 1718 930
rect 1738 910 1746 930
rect 1704 868 1746 910
rect 1818 930 1862 968
rect 1818 910 1830 930
rect 1850 910 1862 930
rect 1818 868 1862 910
rect 1912 930 1954 968
rect 1912 910 1926 930
rect 1946 910 1954 930
rect 1912 868 1954 910
rect 2028 930 2070 968
rect 2028 910 2036 930
rect 2056 910 2070 930
rect 2028 868 2070 910
rect 2120 937 2165 968
rect 2120 930 2164 937
rect 2120 910 2132 930
rect 2152 910 2164 930
rect 2120 868 2164 910
rect 335 691 379 729
rect 335 671 347 691
rect 367 671 379 691
rect 335 629 379 671
rect 429 691 471 729
rect 429 671 443 691
rect 463 671 471 691
rect 429 629 471 671
rect 548 691 592 729
rect 548 671 560 691
rect 580 671 592 691
rect 548 629 592 671
rect 642 691 684 729
rect 642 671 656 691
rect 676 671 684 691
rect 642 629 684 671
rect 756 691 800 729
rect 756 671 768 691
rect 788 671 800 691
rect 756 629 800 671
rect 850 691 892 729
rect 850 671 864 691
rect 884 671 892 691
rect 850 629 892 671
rect 966 691 1008 729
rect 966 671 974 691
rect 994 671 1008 691
rect 966 629 1008 671
rect 1058 698 1103 729
rect 4164 725 4208 767
rect 4164 705 4176 725
rect 4196 705 4208 725
rect 4164 698 4208 705
rect 1058 691 1102 698
rect 1058 671 1070 691
rect 1090 671 1102 691
rect 1058 629 1102 671
rect 4163 667 4208 698
rect 4258 725 4300 767
rect 4258 705 4272 725
rect 4292 705 4300 725
rect 4258 667 4300 705
rect 4374 725 4416 767
rect 4374 705 4382 725
rect 4402 705 4416 725
rect 4374 667 4416 705
rect 4466 725 4510 767
rect 4466 705 4478 725
rect 4498 705 4510 725
rect 4466 667 4510 705
rect 4582 725 4624 767
rect 4582 705 4590 725
rect 4610 705 4624 725
rect 4582 667 4624 705
rect 4674 725 4718 767
rect 4674 705 4686 725
rect 4706 705 4718 725
rect 4674 667 4718 705
rect 4795 725 4837 767
rect 4795 705 4803 725
rect 4823 705 4837 725
rect 4795 667 4837 705
rect 4887 725 4931 767
rect 4887 705 4899 725
rect 4919 705 4931 725
rect 4887 667 4931 705
rect 1347 510 1391 548
rect 1347 490 1359 510
rect 1379 490 1391 510
rect 1347 448 1391 490
rect 1441 510 1483 548
rect 1441 490 1455 510
rect 1475 490 1483 510
rect 1441 448 1483 490
rect 1560 510 1604 548
rect 1560 490 1572 510
rect 1592 490 1604 510
rect 1560 448 1604 490
rect 1654 510 1696 548
rect 1654 490 1668 510
rect 1688 490 1696 510
rect 1654 448 1696 490
rect 1768 510 1812 548
rect 1768 490 1780 510
rect 1800 490 1812 510
rect 1768 448 1812 490
rect 1862 510 1904 548
rect 1862 490 1876 510
rect 1896 490 1904 510
rect 1862 448 1904 490
rect 1978 510 2020 548
rect 1978 490 1986 510
rect 2006 490 2020 510
rect 1978 448 2020 490
rect 2070 517 2115 548
rect 2070 510 2114 517
rect 2070 490 2082 510
rect 2102 490 2114 510
rect 2070 448 2114 490
rect 3151 491 3195 533
rect 3151 471 3163 491
rect 3183 471 3195 491
rect 3151 464 3195 471
rect 3150 433 3195 464
rect 3245 491 3287 533
rect 3245 471 3259 491
rect 3279 471 3287 491
rect 3245 433 3287 471
rect 3361 491 3403 533
rect 3361 471 3369 491
rect 3389 471 3403 491
rect 3361 433 3403 471
rect 3453 491 3497 533
rect 3453 471 3465 491
rect 3485 471 3497 491
rect 3453 433 3497 471
rect 3569 491 3611 533
rect 3569 471 3577 491
rect 3597 471 3611 491
rect 3569 433 3611 471
rect 3661 491 3705 533
rect 3661 471 3673 491
rect 3693 471 3705 491
rect 3661 433 3705 471
rect 3782 491 3824 533
rect 3782 471 3790 491
rect 3810 471 3824 491
rect 3782 433 3824 471
rect 3874 491 3918 533
rect 3874 471 3886 491
rect 3906 471 3918 491
rect 3874 433 3918 471
rect 334 276 378 314
rect 334 256 346 276
rect 366 256 378 276
rect 334 214 378 256
rect 428 276 470 314
rect 428 256 442 276
rect 462 256 470 276
rect 428 214 470 256
rect 547 276 591 314
rect 547 256 559 276
rect 579 256 591 276
rect 547 214 591 256
rect 641 276 683 314
rect 641 256 655 276
rect 675 256 683 276
rect 641 214 683 256
rect 755 276 799 314
rect 755 256 767 276
rect 787 256 799 276
rect 755 214 799 256
rect 849 276 891 314
rect 849 256 863 276
rect 883 256 891 276
rect 849 214 891 256
rect 965 276 1007 314
rect 965 256 973 276
rect 993 256 1007 276
rect 965 214 1007 256
rect 1057 283 1102 314
rect 4163 310 4207 352
rect 4163 290 4175 310
rect 4195 290 4207 310
rect 4163 283 4207 290
rect 1057 276 1101 283
rect 1057 256 1069 276
rect 1089 256 1101 276
rect 1057 214 1101 256
rect 4162 252 4207 283
rect 4257 310 4299 352
rect 4257 290 4271 310
rect 4291 290 4299 310
rect 4257 252 4299 290
rect 4373 310 4415 352
rect 4373 290 4381 310
rect 4401 290 4415 310
rect 4373 252 4415 290
rect 4465 310 4509 352
rect 4465 290 4477 310
rect 4497 290 4509 310
rect 4465 252 4509 290
rect 4581 310 4623 352
rect 4581 290 4589 310
rect 4609 290 4623 310
rect 4581 252 4623 290
rect 4673 310 4717 352
rect 4673 290 4685 310
rect 4705 290 4717 310
rect 4673 252 4717 290
rect 4794 310 4836 352
rect 4794 290 4802 310
rect 4822 290 4836 310
rect 4794 252 4836 290
rect 4886 310 4930 352
rect 4886 290 4898 310
rect 4918 290 4930 310
rect 4886 252 4930 290
rect 1737 -205 1781 -167
rect 1737 -225 1749 -205
rect 1769 -225 1781 -205
rect 1737 -267 1781 -225
rect 1831 -205 1873 -167
rect 1831 -225 1845 -205
rect 1865 -225 1873 -205
rect 1831 -267 1873 -225
rect 1950 -205 1994 -167
rect 1950 -225 1962 -205
rect 1982 -225 1994 -205
rect 1950 -267 1994 -225
rect 2044 -205 2086 -167
rect 2044 -225 2058 -205
rect 2078 -225 2086 -205
rect 2044 -267 2086 -225
rect 2158 -205 2202 -167
rect 2158 -225 2170 -205
rect 2190 -225 2202 -205
rect 2158 -267 2202 -225
rect 2252 -205 2294 -167
rect 2252 -225 2266 -205
rect 2286 -225 2294 -205
rect 2252 -267 2294 -225
rect 2368 -205 2410 -167
rect 2368 -225 2376 -205
rect 2396 -225 2410 -205
rect 2368 -267 2410 -225
rect 2460 -198 2505 -167
rect 2460 -205 2504 -198
rect 2460 -225 2472 -205
rect 2492 -225 2504 -205
rect 2460 -267 2504 -225
<< ndiffc >>
rect 118 7764 136 7782
rect 4133 7712 4153 7732
rect 4236 7708 4256 7728
rect 4344 7708 4364 7728
rect 4447 7712 4467 7732
rect 4552 7708 4572 7728
rect 4655 7712 4675 7732
rect 4765 7708 4785 7728
rect 4868 7712 4888 7732
rect 5048 7711 5066 7729
rect 120 7665 138 7683
rect 116 7550 134 7568
rect 5050 7612 5068 7630
rect 5055 7510 5073 7528
rect 118 7451 136 7469
rect 3120 7478 3140 7498
rect 3223 7474 3243 7494
rect 3331 7474 3351 7494
rect 3434 7478 3454 7498
rect 3539 7474 3559 7494
rect 3642 7478 3662 7498
rect 3752 7474 3772 7494
rect 3855 7478 3875 7498
rect 304 7380 324 7400
rect 407 7384 427 7404
rect 517 7380 537 7400
rect 620 7384 640 7404
rect 725 7380 745 7400
rect 828 7384 848 7404
rect 936 7384 956 7404
rect 1039 7380 1059 7400
rect 5057 7411 5075 7429
rect 116 7268 134 7286
rect 4132 7297 4152 7317
rect 4235 7293 4255 7313
rect 4343 7293 4363 7313
rect 4446 7297 4466 7317
rect 4551 7293 4571 7313
rect 4654 7297 4674 7317
rect 4764 7293 4784 7313
rect 4867 7297 4887 7317
rect 1316 7199 1336 7219
rect 1419 7203 1439 7223
rect 1529 7199 1549 7219
rect 1632 7203 1652 7223
rect 1737 7199 1757 7219
rect 1840 7203 1860 7223
rect 1948 7203 1968 7223
rect 2051 7199 2071 7219
rect 5055 7228 5073 7246
rect 118 7169 136 7187
rect 123 7067 141 7085
rect 5057 7129 5075 7147
rect 3070 7058 3090 7078
rect 3173 7054 3193 7074
rect 3281 7054 3301 7074
rect 3384 7058 3404 7078
rect 3489 7054 3509 7074
rect 3592 7058 3612 7078
rect 3702 7054 3722 7074
rect 3805 7058 3825 7078
rect 125 6968 143 6986
rect 303 6965 323 6985
rect 406 6969 426 6989
rect 516 6965 536 6985
rect 619 6969 639 6989
rect 724 6965 744 6985
rect 827 6969 847 6989
rect 935 6969 955 6989
rect 1038 6965 1058 6985
rect 5053 7014 5071 7032
rect 5055 6915 5073 6933
rect 123 6783 141 6801
rect 125 6684 143 6702
rect 4138 6731 4158 6751
rect 4241 6727 4261 6747
rect 4349 6727 4369 6747
rect 4452 6731 4472 6751
rect 4557 6727 4577 6747
rect 4660 6731 4680 6751
rect 4770 6727 4790 6747
rect 4873 6731 4893 6751
rect 5053 6730 5071 6748
rect 1371 6638 1391 6658
rect 1474 6642 1494 6662
rect 1584 6638 1604 6658
rect 1687 6642 1707 6662
rect 1792 6638 1812 6658
rect 1895 6642 1915 6662
rect 2003 6642 2023 6662
rect 2106 6638 2126 6658
rect 121 6569 139 6587
rect 5055 6631 5073 6649
rect 5060 6529 5078 6547
rect 123 6470 141 6488
rect 3125 6497 3145 6517
rect 3228 6493 3248 6513
rect 3336 6493 3356 6513
rect 3439 6497 3459 6517
rect 3544 6493 3564 6513
rect 3647 6497 3667 6517
rect 3757 6493 3777 6513
rect 3860 6497 3880 6517
rect 309 6399 329 6419
rect 412 6403 432 6423
rect 522 6399 542 6419
rect 625 6403 645 6423
rect 730 6399 750 6419
rect 833 6403 853 6423
rect 941 6403 961 6423
rect 1044 6399 1064 6419
rect 5062 6430 5080 6448
rect 121 6287 139 6305
rect 4137 6316 4157 6336
rect 4240 6312 4260 6332
rect 4348 6312 4368 6332
rect 4451 6316 4471 6336
rect 4556 6312 4576 6332
rect 4659 6316 4679 6336
rect 4769 6312 4789 6332
rect 4872 6316 4892 6336
rect 1321 6218 1341 6238
rect 1424 6222 1444 6242
rect 1534 6218 1554 6238
rect 1637 6222 1657 6242
rect 1742 6218 1762 6238
rect 1845 6222 1865 6242
rect 1953 6222 1973 6242
rect 2056 6218 2076 6238
rect 5060 6247 5078 6265
rect 123 6188 141 6206
rect 128 6086 146 6104
rect 5062 6148 5080 6166
rect 2917 6030 2937 6050
rect 3020 6026 3040 6046
rect 3128 6026 3148 6046
rect 3231 6030 3251 6050
rect 3336 6026 3356 6046
rect 3439 6030 3459 6050
rect 3549 6026 3569 6046
rect 3652 6030 3672 6050
rect 5058 6033 5076 6051
rect 130 5987 148 6005
rect 308 5984 328 6004
rect 411 5988 431 6008
rect 521 5984 541 6004
rect 624 5988 644 6008
rect 729 5984 749 6004
rect 832 5988 852 6008
rect 940 5988 960 6008
rect 1043 5984 1063 6004
rect 130 5804 148 5822
rect 5060 5934 5078 5952
rect 4145 5752 4165 5772
rect 4248 5748 4268 5768
rect 4356 5748 4376 5768
rect 4459 5752 4479 5772
rect 4564 5748 4584 5768
rect 4667 5752 4687 5772
rect 4777 5748 4797 5768
rect 4880 5752 4900 5772
rect 5060 5751 5078 5769
rect 132 5705 150 5723
rect 1536 5706 1556 5726
rect 1639 5710 1659 5730
rect 1749 5706 1769 5726
rect 1852 5710 1872 5730
rect 1957 5706 1977 5726
rect 2060 5710 2080 5730
rect 2168 5710 2188 5730
rect 2271 5706 2291 5726
rect 128 5590 146 5608
rect 5062 5652 5080 5670
rect 5067 5550 5085 5568
rect 130 5491 148 5509
rect 3132 5518 3152 5538
rect 3235 5514 3255 5534
rect 3343 5514 3363 5534
rect 3446 5518 3466 5538
rect 3551 5514 3571 5534
rect 3654 5518 3674 5538
rect 3764 5514 3784 5534
rect 3867 5518 3887 5538
rect 316 5420 336 5440
rect 419 5424 439 5444
rect 529 5420 549 5440
rect 632 5424 652 5444
rect 737 5420 757 5440
rect 840 5424 860 5444
rect 948 5424 968 5444
rect 1051 5420 1071 5440
rect 5069 5451 5087 5469
rect 128 5308 146 5326
rect 4144 5337 4164 5357
rect 4247 5333 4267 5353
rect 4355 5333 4375 5353
rect 4458 5337 4478 5357
rect 4563 5333 4583 5353
rect 4666 5337 4686 5357
rect 4776 5333 4796 5353
rect 4879 5337 4899 5357
rect 1328 5239 1348 5259
rect 1431 5243 1451 5263
rect 1541 5239 1561 5259
rect 1644 5243 1664 5263
rect 1749 5239 1769 5259
rect 1852 5243 1872 5263
rect 1960 5243 1980 5263
rect 2063 5239 2083 5259
rect 5067 5268 5085 5286
rect 130 5209 148 5227
rect 135 5107 153 5125
rect 5069 5169 5087 5187
rect 3082 5098 3102 5118
rect 3185 5094 3205 5114
rect 3293 5094 3313 5114
rect 3396 5098 3416 5118
rect 3501 5094 3521 5114
rect 3604 5098 3624 5118
rect 3714 5094 3734 5114
rect 3817 5098 3837 5118
rect 137 5008 155 5026
rect 315 5005 335 5025
rect 418 5009 438 5029
rect 528 5005 548 5025
rect 631 5009 651 5029
rect 736 5005 756 5025
rect 839 5009 859 5029
rect 947 5009 967 5029
rect 1050 5005 1070 5025
rect 5065 5054 5083 5072
rect 5067 4955 5085 4973
rect 135 4823 153 4841
rect 137 4724 155 4742
rect 4150 4771 4170 4791
rect 4253 4767 4273 4787
rect 4361 4767 4381 4787
rect 4464 4771 4484 4791
rect 4569 4767 4589 4787
rect 4672 4771 4692 4791
rect 4782 4767 4802 4787
rect 4885 4771 4905 4791
rect 5065 4770 5083 4788
rect 1383 4678 1403 4698
rect 1486 4682 1506 4702
rect 1596 4678 1616 4698
rect 1699 4682 1719 4702
rect 1804 4678 1824 4698
rect 1907 4682 1927 4702
rect 2015 4682 2035 4702
rect 2118 4678 2138 4698
rect 133 4609 151 4627
rect 5067 4671 5085 4689
rect 5072 4569 5090 4587
rect 135 4510 153 4528
rect 3137 4537 3157 4557
rect 3240 4533 3260 4553
rect 3348 4533 3368 4553
rect 3451 4537 3471 4557
rect 3556 4533 3576 4553
rect 3659 4537 3679 4557
rect 3769 4533 3789 4553
rect 3872 4537 3892 4557
rect 321 4439 341 4459
rect 424 4443 444 4463
rect 534 4439 554 4459
rect 637 4443 657 4463
rect 742 4439 762 4459
rect 845 4443 865 4463
rect 953 4443 973 4463
rect 1056 4439 1076 4459
rect 5074 4470 5092 4488
rect 133 4327 151 4345
rect 4149 4356 4169 4376
rect 4252 4352 4272 4372
rect 4360 4352 4380 4372
rect 4463 4356 4483 4376
rect 4568 4352 4588 4372
rect 4671 4356 4691 4376
rect 4781 4352 4801 4372
rect 4884 4356 4904 4376
rect 1333 4258 1353 4278
rect 1436 4262 1456 4282
rect 1546 4258 1566 4278
rect 1649 4262 1669 4282
rect 1754 4258 1774 4278
rect 1857 4262 1877 4282
rect 1965 4262 1985 4282
rect 2068 4258 2088 4278
rect 5072 4287 5090 4305
rect 135 4228 153 4246
rect 140 4126 158 4144
rect 5074 4188 5092 4206
rect 2842 4105 2862 4125
rect 2945 4101 2965 4121
rect 3053 4101 3073 4121
rect 3156 4105 3176 4125
rect 3261 4101 3281 4121
rect 3364 4105 3384 4125
rect 3474 4101 3494 4121
rect 3577 4105 3597 4125
rect 142 4027 160 4045
rect 320 4024 340 4044
rect 423 4028 443 4048
rect 533 4024 553 4044
rect 636 4028 656 4048
rect 741 4024 761 4044
rect 844 4028 864 4048
rect 952 4028 972 4048
rect 1055 4024 1075 4044
rect 5070 4073 5088 4091
rect 138 3847 156 3865
rect 5072 3974 5090 3992
rect 140 3748 158 3766
rect 4153 3795 4173 3815
rect 4256 3791 4276 3811
rect 4364 3791 4384 3811
rect 4467 3795 4487 3815
rect 4572 3791 4592 3811
rect 4675 3795 4695 3815
rect 4785 3791 4805 3811
rect 4888 3795 4908 3815
rect 5068 3794 5086 3812
rect 1631 3714 1651 3734
rect 1734 3718 1754 3738
rect 1844 3714 1864 3734
rect 1947 3718 1967 3738
rect 2052 3714 2072 3734
rect 2155 3718 2175 3738
rect 2263 3718 2283 3738
rect 2366 3714 2386 3734
rect 136 3633 154 3651
rect 5070 3695 5088 3713
rect 5075 3593 5093 3611
rect 138 3534 156 3552
rect 3140 3561 3160 3581
rect 3243 3557 3263 3577
rect 3351 3557 3371 3577
rect 3454 3561 3474 3581
rect 3559 3557 3579 3577
rect 3662 3561 3682 3581
rect 3772 3557 3792 3577
rect 3875 3561 3895 3581
rect 324 3463 344 3483
rect 427 3467 447 3487
rect 537 3463 557 3483
rect 640 3467 660 3487
rect 745 3463 765 3483
rect 848 3467 868 3487
rect 956 3467 976 3487
rect 1059 3463 1079 3483
rect 5077 3494 5095 3512
rect 136 3351 154 3369
rect 4152 3380 4172 3400
rect 4255 3376 4275 3396
rect 4363 3376 4383 3396
rect 4466 3380 4486 3400
rect 4571 3376 4591 3396
rect 4674 3380 4694 3400
rect 4784 3376 4804 3396
rect 4887 3380 4907 3400
rect 1336 3282 1356 3302
rect 1439 3286 1459 3306
rect 1549 3282 1569 3302
rect 1652 3286 1672 3306
rect 1757 3282 1777 3302
rect 1860 3286 1880 3306
rect 1968 3286 1988 3306
rect 2071 3282 2091 3302
rect 5075 3311 5093 3329
rect 138 3252 156 3270
rect 143 3150 161 3168
rect 5077 3212 5095 3230
rect 3090 3141 3110 3161
rect 3193 3137 3213 3157
rect 3301 3137 3321 3157
rect 3404 3141 3424 3161
rect 3509 3137 3529 3157
rect 3612 3141 3632 3161
rect 3722 3137 3742 3157
rect 3825 3141 3845 3161
rect 145 3051 163 3069
rect 323 3048 343 3068
rect 426 3052 446 3072
rect 536 3048 556 3068
rect 639 3052 659 3072
rect 744 3048 764 3068
rect 847 3052 867 3072
rect 955 3052 975 3072
rect 1058 3048 1078 3068
rect 5073 3097 5091 3115
rect 5075 2998 5093 3016
rect 143 2866 161 2884
rect 145 2767 163 2785
rect 4158 2814 4178 2834
rect 4261 2810 4281 2830
rect 4369 2810 4389 2830
rect 4472 2814 4492 2834
rect 4577 2810 4597 2830
rect 4680 2814 4700 2834
rect 4790 2810 4810 2830
rect 4893 2814 4913 2834
rect 5073 2813 5091 2831
rect 1391 2721 1411 2741
rect 1494 2725 1514 2745
rect 1604 2721 1624 2741
rect 1707 2725 1727 2745
rect 1812 2721 1832 2741
rect 1915 2725 1935 2745
rect 2023 2725 2043 2745
rect 2126 2721 2146 2741
rect 141 2652 159 2670
rect 5075 2714 5093 2732
rect 5080 2612 5098 2630
rect 143 2553 161 2571
rect 3145 2580 3165 2600
rect 3248 2576 3268 2596
rect 3356 2576 3376 2596
rect 3459 2580 3479 2600
rect 3564 2576 3584 2596
rect 3667 2580 3687 2600
rect 3777 2576 3797 2596
rect 3880 2580 3900 2600
rect 329 2482 349 2502
rect 432 2486 452 2506
rect 542 2482 562 2502
rect 645 2486 665 2506
rect 750 2482 770 2502
rect 853 2486 873 2506
rect 961 2486 981 2506
rect 1064 2482 1084 2502
rect 5082 2513 5100 2531
rect 141 2370 159 2388
rect 4157 2399 4177 2419
rect 4260 2395 4280 2415
rect 4368 2395 4388 2415
rect 4471 2399 4491 2419
rect 4576 2395 4596 2415
rect 4679 2399 4699 2419
rect 4789 2395 4809 2415
rect 4892 2399 4912 2419
rect 1341 2301 1361 2321
rect 1444 2305 1464 2325
rect 1554 2301 1574 2321
rect 1657 2305 1677 2325
rect 1762 2301 1782 2321
rect 1865 2305 1885 2325
rect 1973 2305 1993 2325
rect 2076 2301 2096 2321
rect 5080 2330 5098 2348
rect 143 2271 161 2289
rect 148 2169 166 2187
rect 5082 2231 5100 2249
rect 2937 2113 2957 2133
rect 3040 2109 3060 2129
rect 3148 2109 3168 2129
rect 3251 2113 3271 2133
rect 3356 2109 3376 2129
rect 3459 2113 3479 2133
rect 3569 2109 3589 2129
rect 3672 2113 3692 2133
rect 5078 2116 5096 2134
rect 150 2070 168 2088
rect 328 2067 348 2087
rect 431 2071 451 2091
rect 541 2067 561 2087
rect 644 2071 664 2091
rect 749 2067 769 2087
rect 852 2071 872 2091
rect 960 2071 980 2091
rect 1063 2067 1083 2087
rect 150 1887 168 1905
rect 5080 2017 5098 2035
rect 4165 1835 4185 1855
rect 4268 1831 4288 1851
rect 4376 1831 4396 1851
rect 4479 1835 4499 1855
rect 4584 1831 4604 1851
rect 4687 1835 4707 1855
rect 4797 1831 4817 1851
rect 4900 1835 4920 1855
rect 5080 1834 5098 1852
rect 152 1788 170 1806
rect 1556 1789 1576 1809
rect 1659 1793 1679 1813
rect 1769 1789 1789 1809
rect 1872 1793 1892 1813
rect 1977 1789 1997 1809
rect 2080 1793 2100 1813
rect 2188 1793 2208 1813
rect 2291 1789 2311 1809
rect 148 1673 166 1691
rect 5082 1735 5100 1753
rect 5087 1633 5105 1651
rect 150 1574 168 1592
rect 3152 1601 3172 1621
rect 3255 1597 3275 1617
rect 3363 1597 3383 1617
rect 3466 1601 3486 1621
rect 3571 1597 3591 1617
rect 3674 1601 3694 1621
rect 3784 1597 3804 1617
rect 3887 1601 3907 1621
rect 336 1503 356 1523
rect 439 1507 459 1527
rect 549 1503 569 1523
rect 652 1507 672 1527
rect 757 1503 777 1523
rect 860 1507 880 1527
rect 968 1507 988 1527
rect 1071 1503 1091 1523
rect 5089 1534 5107 1552
rect 148 1391 166 1409
rect 4164 1420 4184 1440
rect 4267 1416 4287 1436
rect 4375 1416 4395 1436
rect 4478 1420 4498 1440
rect 4583 1416 4603 1436
rect 4686 1420 4706 1440
rect 4796 1416 4816 1436
rect 4899 1420 4919 1440
rect 1348 1322 1368 1342
rect 1451 1326 1471 1346
rect 1561 1322 1581 1342
rect 1664 1326 1684 1346
rect 1769 1322 1789 1342
rect 1872 1326 1892 1346
rect 1980 1326 2000 1346
rect 2083 1322 2103 1342
rect 5087 1351 5105 1369
rect 150 1292 168 1310
rect 155 1190 173 1208
rect 5089 1252 5107 1270
rect 3102 1181 3122 1201
rect 3205 1177 3225 1197
rect 3313 1177 3333 1197
rect 3416 1181 3436 1201
rect 3521 1177 3541 1197
rect 3624 1181 3644 1201
rect 3734 1177 3754 1197
rect 3837 1181 3857 1201
rect 157 1091 175 1109
rect 335 1088 355 1108
rect 438 1092 458 1112
rect 548 1088 568 1108
rect 651 1092 671 1112
rect 756 1088 776 1108
rect 859 1092 879 1112
rect 967 1092 987 1112
rect 1070 1088 1090 1108
rect 5085 1137 5103 1155
rect 5087 1038 5105 1056
rect 155 906 173 924
rect 157 807 175 825
rect 4170 854 4190 874
rect 4273 850 4293 870
rect 4381 850 4401 870
rect 4484 854 4504 874
rect 4589 850 4609 870
rect 4692 854 4712 874
rect 4802 850 4822 870
rect 4905 854 4925 874
rect 5085 853 5103 871
rect 1403 761 1423 781
rect 1506 765 1526 785
rect 1616 761 1636 781
rect 1719 765 1739 785
rect 1824 761 1844 781
rect 1927 765 1947 785
rect 2035 765 2055 785
rect 2138 761 2158 781
rect 153 692 171 710
rect 5087 754 5105 772
rect 5092 652 5110 670
rect 155 593 173 611
rect 3157 620 3177 640
rect 3260 616 3280 636
rect 3368 616 3388 636
rect 3471 620 3491 640
rect 3576 616 3596 636
rect 3679 620 3699 640
rect 3789 616 3809 636
rect 3892 620 3912 640
rect 341 522 361 542
rect 444 526 464 546
rect 554 522 574 542
rect 657 526 677 546
rect 762 522 782 542
rect 865 526 885 546
rect 973 526 993 546
rect 1076 522 1096 542
rect 5094 553 5112 571
rect 153 410 171 428
rect 4169 439 4189 459
rect 4272 435 4292 455
rect 4380 435 4400 455
rect 4483 439 4503 459
rect 4588 435 4608 455
rect 4691 439 4711 459
rect 4801 435 4821 455
rect 4904 439 4924 459
rect 1353 341 1373 361
rect 1456 345 1476 365
rect 1566 341 1586 361
rect 1669 345 1689 365
rect 1774 341 1794 361
rect 1877 345 1897 365
rect 1985 345 2005 365
rect 2088 341 2108 361
rect 5092 370 5110 388
rect 155 311 173 329
rect 160 209 178 227
rect 5094 271 5112 289
rect 5090 156 5108 174
rect 162 110 180 128
rect 340 107 360 127
rect 443 111 463 131
rect 553 107 573 127
rect 656 111 676 131
rect 761 107 781 127
rect 864 111 884 131
rect 972 111 992 131
rect 1075 107 1095 127
rect 5092 57 5110 75
rect 1743 -374 1763 -354
rect 1846 -370 1866 -350
rect 1956 -374 1976 -354
rect 2059 -370 2079 -350
rect 2164 -374 2184 -354
rect 2267 -370 2287 -350
rect 2375 -370 2395 -350
rect 2478 -374 2498 -354
<< pdiffc >>
rect 310 7529 330 7549
rect 406 7529 426 7549
rect 523 7529 543 7549
rect 619 7529 639 7549
rect 731 7529 751 7549
rect 827 7529 847 7549
rect 937 7529 957 7549
rect 4139 7563 4159 7583
rect 1033 7529 1053 7549
rect 4235 7563 4255 7583
rect 4345 7563 4365 7583
rect 4441 7563 4461 7583
rect 4553 7563 4573 7583
rect 4649 7563 4669 7583
rect 4766 7563 4786 7583
rect 4862 7563 4882 7583
rect 1322 7348 1342 7368
rect 1418 7348 1438 7368
rect 1535 7348 1555 7368
rect 1631 7348 1651 7368
rect 1743 7348 1763 7368
rect 1839 7348 1859 7368
rect 1949 7348 1969 7368
rect 2045 7348 2065 7368
rect 3126 7329 3146 7349
rect 3222 7329 3242 7349
rect 3332 7329 3352 7349
rect 3428 7329 3448 7349
rect 3540 7329 3560 7349
rect 3636 7329 3656 7349
rect 3753 7329 3773 7349
rect 3849 7329 3869 7349
rect 309 7114 329 7134
rect 405 7114 425 7134
rect 522 7114 542 7134
rect 618 7114 638 7134
rect 730 7114 750 7134
rect 826 7114 846 7134
rect 936 7114 956 7134
rect 4138 7148 4158 7168
rect 1032 7114 1052 7134
rect 4234 7148 4254 7168
rect 4344 7148 4364 7168
rect 4440 7148 4460 7168
rect 4552 7148 4572 7168
rect 4648 7148 4668 7168
rect 4765 7148 4785 7168
rect 4861 7148 4881 7168
rect 3076 6909 3096 6929
rect 3172 6909 3192 6929
rect 3282 6909 3302 6929
rect 3378 6909 3398 6929
rect 3490 6909 3510 6929
rect 3586 6909 3606 6929
rect 3703 6909 3723 6929
rect 3799 6909 3819 6929
rect 1377 6787 1397 6807
rect 1473 6787 1493 6807
rect 1590 6787 1610 6807
rect 1686 6787 1706 6807
rect 1798 6787 1818 6807
rect 1894 6787 1914 6807
rect 2004 6787 2024 6807
rect 2100 6787 2120 6807
rect 315 6548 335 6568
rect 411 6548 431 6568
rect 528 6548 548 6568
rect 624 6548 644 6568
rect 736 6548 756 6568
rect 832 6548 852 6568
rect 942 6548 962 6568
rect 4144 6582 4164 6602
rect 1038 6548 1058 6568
rect 4240 6582 4260 6602
rect 4350 6582 4370 6602
rect 4446 6582 4466 6602
rect 4558 6582 4578 6602
rect 4654 6582 4674 6602
rect 4771 6582 4791 6602
rect 4867 6582 4887 6602
rect 1327 6367 1347 6387
rect 1423 6367 1443 6387
rect 1540 6367 1560 6387
rect 1636 6367 1656 6387
rect 1748 6367 1768 6387
rect 1844 6367 1864 6387
rect 1954 6367 1974 6387
rect 2050 6367 2070 6387
rect 3131 6348 3151 6368
rect 3227 6348 3247 6368
rect 3337 6348 3357 6368
rect 3433 6348 3453 6368
rect 3545 6348 3565 6368
rect 3641 6348 3661 6368
rect 3758 6348 3778 6368
rect 3854 6348 3874 6368
rect 314 6133 334 6153
rect 410 6133 430 6153
rect 527 6133 547 6153
rect 623 6133 643 6153
rect 735 6133 755 6153
rect 831 6133 851 6153
rect 941 6133 961 6153
rect 4143 6167 4163 6187
rect 1037 6133 1057 6153
rect 4239 6167 4259 6187
rect 4349 6167 4369 6187
rect 4445 6167 4465 6187
rect 4557 6167 4577 6187
rect 4653 6167 4673 6187
rect 4770 6167 4790 6187
rect 4866 6167 4886 6187
rect 1542 5855 1562 5875
rect 1638 5855 1658 5875
rect 1755 5855 1775 5875
rect 1851 5855 1871 5875
rect 1963 5855 1983 5875
rect 2059 5855 2079 5875
rect 2169 5855 2189 5875
rect 2265 5855 2285 5875
rect 2923 5881 2943 5901
rect 3019 5881 3039 5901
rect 3129 5881 3149 5901
rect 3225 5881 3245 5901
rect 3337 5881 3357 5901
rect 3433 5881 3453 5901
rect 3550 5881 3570 5901
rect 3646 5881 3666 5901
rect 322 5569 342 5589
rect 418 5569 438 5589
rect 535 5569 555 5589
rect 631 5569 651 5589
rect 743 5569 763 5589
rect 839 5569 859 5589
rect 949 5569 969 5589
rect 4151 5603 4171 5623
rect 1045 5569 1065 5589
rect 4247 5603 4267 5623
rect 4357 5603 4377 5623
rect 4453 5603 4473 5623
rect 4565 5603 4585 5623
rect 4661 5603 4681 5623
rect 4778 5603 4798 5623
rect 4874 5603 4894 5623
rect 1334 5388 1354 5408
rect 1430 5388 1450 5408
rect 1547 5388 1567 5408
rect 1643 5388 1663 5408
rect 1755 5388 1775 5408
rect 1851 5388 1871 5408
rect 1961 5388 1981 5408
rect 2057 5388 2077 5408
rect 3138 5369 3158 5389
rect 3234 5369 3254 5389
rect 3344 5369 3364 5389
rect 3440 5369 3460 5389
rect 3552 5369 3572 5389
rect 3648 5369 3668 5389
rect 3765 5369 3785 5389
rect 3861 5369 3881 5389
rect 321 5154 341 5174
rect 417 5154 437 5174
rect 534 5154 554 5174
rect 630 5154 650 5174
rect 742 5154 762 5174
rect 838 5154 858 5174
rect 948 5154 968 5174
rect 4150 5188 4170 5208
rect 1044 5154 1064 5174
rect 4246 5188 4266 5208
rect 4356 5188 4376 5208
rect 4452 5188 4472 5208
rect 4564 5188 4584 5208
rect 4660 5188 4680 5208
rect 4777 5188 4797 5208
rect 4873 5188 4893 5208
rect 3088 4949 3108 4969
rect 3184 4949 3204 4969
rect 3294 4949 3314 4969
rect 3390 4949 3410 4969
rect 3502 4949 3522 4969
rect 3598 4949 3618 4969
rect 3715 4949 3735 4969
rect 3811 4949 3831 4969
rect 1389 4827 1409 4847
rect 1485 4827 1505 4847
rect 1602 4827 1622 4847
rect 1698 4827 1718 4847
rect 1810 4827 1830 4847
rect 1906 4827 1926 4847
rect 2016 4827 2036 4847
rect 2112 4827 2132 4847
rect 327 4588 347 4608
rect 423 4588 443 4608
rect 540 4588 560 4608
rect 636 4588 656 4608
rect 748 4588 768 4608
rect 844 4588 864 4608
rect 954 4588 974 4608
rect 4156 4622 4176 4642
rect 1050 4588 1070 4608
rect 4252 4622 4272 4642
rect 4362 4622 4382 4642
rect 4458 4622 4478 4642
rect 4570 4622 4590 4642
rect 4666 4622 4686 4642
rect 4783 4622 4803 4642
rect 4879 4622 4899 4642
rect 1339 4407 1359 4427
rect 1435 4407 1455 4427
rect 1552 4407 1572 4427
rect 1648 4407 1668 4427
rect 1760 4407 1780 4427
rect 1856 4407 1876 4427
rect 1966 4407 1986 4427
rect 2062 4407 2082 4427
rect 3143 4388 3163 4408
rect 3239 4388 3259 4408
rect 3349 4388 3369 4408
rect 3445 4388 3465 4408
rect 3557 4388 3577 4408
rect 3653 4388 3673 4408
rect 3770 4388 3790 4408
rect 3866 4388 3886 4408
rect 326 4173 346 4193
rect 422 4173 442 4193
rect 539 4173 559 4193
rect 635 4173 655 4193
rect 747 4173 767 4193
rect 843 4173 863 4193
rect 953 4173 973 4193
rect 4155 4207 4175 4227
rect 1049 4173 1069 4193
rect 4251 4207 4271 4227
rect 4361 4207 4381 4227
rect 4457 4207 4477 4227
rect 4569 4207 4589 4227
rect 4665 4207 4685 4227
rect 4782 4207 4802 4227
rect 4878 4207 4898 4227
rect 2848 3956 2868 3976
rect 1637 3863 1657 3883
rect 1733 3863 1753 3883
rect 1850 3863 1870 3883
rect 1946 3863 1966 3883
rect 2058 3863 2078 3883
rect 2154 3863 2174 3883
rect 2264 3863 2284 3883
rect 2944 3956 2964 3976
rect 3054 3956 3074 3976
rect 3150 3956 3170 3976
rect 3262 3956 3282 3976
rect 3358 3956 3378 3976
rect 3475 3956 3495 3976
rect 3571 3956 3591 3976
rect 2360 3863 2380 3883
rect 330 3612 350 3632
rect 426 3612 446 3632
rect 543 3612 563 3632
rect 639 3612 659 3632
rect 751 3612 771 3632
rect 847 3612 867 3632
rect 957 3612 977 3632
rect 4159 3646 4179 3666
rect 1053 3612 1073 3632
rect 4255 3646 4275 3666
rect 4365 3646 4385 3666
rect 4461 3646 4481 3666
rect 4573 3646 4593 3666
rect 4669 3646 4689 3666
rect 4786 3646 4806 3666
rect 4882 3646 4902 3666
rect 1342 3431 1362 3451
rect 1438 3431 1458 3451
rect 1555 3431 1575 3451
rect 1651 3431 1671 3451
rect 1763 3431 1783 3451
rect 1859 3431 1879 3451
rect 1969 3431 1989 3451
rect 2065 3431 2085 3451
rect 3146 3412 3166 3432
rect 3242 3412 3262 3432
rect 3352 3412 3372 3432
rect 3448 3412 3468 3432
rect 3560 3412 3580 3432
rect 3656 3412 3676 3432
rect 3773 3412 3793 3432
rect 3869 3412 3889 3432
rect 329 3197 349 3217
rect 425 3197 445 3217
rect 542 3197 562 3217
rect 638 3197 658 3217
rect 750 3197 770 3217
rect 846 3197 866 3217
rect 956 3197 976 3217
rect 4158 3231 4178 3251
rect 1052 3197 1072 3217
rect 4254 3231 4274 3251
rect 4364 3231 4384 3251
rect 4460 3231 4480 3251
rect 4572 3231 4592 3251
rect 4668 3231 4688 3251
rect 4785 3231 4805 3251
rect 4881 3231 4901 3251
rect 3096 2992 3116 3012
rect 3192 2992 3212 3012
rect 3302 2992 3322 3012
rect 3398 2992 3418 3012
rect 3510 2992 3530 3012
rect 3606 2992 3626 3012
rect 3723 2992 3743 3012
rect 3819 2992 3839 3012
rect 1397 2870 1417 2890
rect 1493 2870 1513 2890
rect 1610 2870 1630 2890
rect 1706 2870 1726 2890
rect 1818 2870 1838 2890
rect 1914 2870 1934 2890
rect 2024 2870 2044 2890
rect 2120 2870 2140 2890
rect 335 2631 355 2651
rect 431 2631 451 2651
rect 548 2631 568 2651
rect 644 2631 664 2651
rect 756 2631 776 2651
rect 852 2631 872 2651
rect 962 2631 982 2651
rect 4164 2665 4184 2685
rect 1058 2631 1078 2651
rect 4260 2665 4280 2685
rect 4370 2665 4390 2685
rect 4466 2665 4486 2685
rect 4578 2665 4598 2685
rect 4674 2665 4694 2685
rect 4791 2665 4811 2685
rect 4887 2665 4907 2685
rect 1347 2450 1367 2470
rect 1443 2450 1463 2470
rect 1560 2450 1580 2470
rect 1656 2450 1676 2470
rect 1768 2450 1788 2470
rect 1864 2450 1884 2470
rect 1974 2450 1994 2470
rect 2070 2450 2090 2470
rect 3151 2431 3171 2451
rect 3247 2431 3267 2451
rect 3357 2431 3377 2451
rect 3453 2431 3473 2451
rect 3565 2431 3585 2451
rect 3661 2431 3681 2451
rect 3778 2431 3798 2451
rect 3874 2431 3894 2451
rect 334 2216 354 2236
rect 430 2216 450 2236
rect 547 2216 567 2236
rect 643 2216 663 2236
rect 755 2216 775 2236
rect 851 2216 871 2236
rect 961 2216 981 2236
rect 4163 2250 4183 2270
rect 1057 2216 1077 2236
rect 4259 2250 4279 2270
rect 4369 2250 4389 2270
rect 4465 2250 4485 2270
rect 4577 2250 4597 2270
rect 4673 2250 4693 2270
rect 4790 2250 4810 2270
rect 4886 2250 4906 2270
rect 1562 1938 1582 1958
rect 1658 1938 1678 1958
rect 1775 1938 1795 1958
rect 1871 1938 1891 1958
rect 1983 1938 2003 1958
rect 2079 1938 2099 1958
rect 2189 1938 2209 1958
rect 2285 1938 2305 1958
rect 2943 1964 2963 1984
rect 3039 1964 3059 1984
rect 3149 1964 3169 1984
rect 3245 1964 3265 1984
rect 3357 1964 3377 1984
rect 3453 1964 3473 1984
rect 3570 1964 3590 1984
rect 3666 1964 3686 1984
rect 342 1652 362 1672
rect 438 1652 458 1672
rect 555 1652 575 1672
rect 651 1652 671 1672
rect 763 1652 783 1672
rect 859 1652 879 1672
rect 969 1652 989 1672
rect 4171 1686 4191 1706
rect 1065 1652 1085 1672
rect 4267 1686 4287 1706
rect 4377 1686 4397 1706
rect 4473 1686 4493 1706
rect 4585 1686 4605 1706
rect 4681 1686 4701 1706
rect 4798 1686 4818 1706
rect 4894 1686 4914 1706
rect 1354 1471 1374 1491
rect 1450 1471 1470 1491
rect 1567 1471 1587 1491
rect 1663 1471 1683 1491
rect 1775 1471 1795 1491
rect 1871 1471 1891 1491
rect 1981 1471 2001 1491
rect 2077 1471 2097 1491
rect 3158 1452 3178 1472
rect 3254 1452 3274 1472
rect 3364 1452 3384 1472
rect 3460 1452 3480 1472
rect 3572 1452 3592 1472
rect 3668 1452 3688 1472
rect 3785 1452 3805 1472
rect 3881 1452 3901 1472
rect 341 1237 361 1257
rect 437 1237 457 1257
rect 554 1237 574 1257
rect 650 1237 670 1257
rect 762 1237 782 1257
rect 858 1237 878 1257
rect 968 1237 988 1257
rect 4170 1271 4190 1291
rect 1064 1237 1084 1257
rect 4266 1271 4286 1291
rect 4376 1271 4396 1291
rect 4472 1271 4492 1291
rect 4584 1271 4604 1291
rect 4680 1271 4700 1291
rect 4797 1271 4817 1291
rect 4893 1271 4913 1291
rect 3108 1032 3128 1052
rect 3204 1032 3224 1052
rect 3314 1032 3334 1052
rect 3410 1032 3430 1052
rect 3522 1032 3542 1052
rect 3618 1032 3638 1052
rect 3735 1032 3755 1052
rect 3831 1032 3851 1052
rect 1409 910 1429 930
rect 1505 910 1525 930
rect 1622 910 1642 930
rect 1718 910 1738 930
rect 1830 910 1850 930
rect 1926 910 1946 930
rect 2036 910 2056 930
rect 2132 910 2152 930
rect 347 671 367 691
rect 443 671 463 691
rect 560 671 580 691
rect 656 671 676 691
rect 768 671 788 691
rect 864 671 884 691
rect 974 671 994 691
rect 4176 705 4196 725
rect 1070 671 1090 691
rect 4272 705 4292 725
rect 4382 705 4402 725
rect 4478 705 4498 725
rect 4590 705 4610 725
rect 4686 705 4706 725
rect 4803 705 4823 725
rect 4899 705 4919 725
rect 1359 490 1379 510
rect 1455 490 1475 510
rect 1572 490 1592 510
rect 1668 490 1688 510
rect 1780 490 1800 510
rect 1876 490 1896 510
rect 1986 490 2006 510
rect 2082 490 2102 510
rect 3163 471 3183 491
rect 3259 471 3279 491
rect 3369 471 3389 491
rect 3465 471 3485 491
rect 3577 471 3597 491
rect 3673 471 3693 491
rect 3790 471 3810 491
rect 3886 471 3906 491
rect 346 256 366 276
rect 442 256 462 276
rect 559 256 579 276
rect 655 256 675 276
rect 767 256 787 276
rect 863 256 883 276
rect 973 256 993 276
rect 4175 290 4195 310
rect 1069 256 1089 276
rect 4271 290 4291 310
rect 4381 290 4401 310
rect 4477 290 4497 310
rect 4589 290 4609 310
rect 4685 290 4705 310
rect 4802 290 4822 310
rect 4898 290 4918 310
rect 1749 -225 1769 -205
rect 1845 -225 1865 -205
rect 1962 -225 1982 -205
rect 2058 -225 2078 -205
rect 2170 -225 2190 -205
rect 2266 -225 2286 -205
rect 2376 -225 2396 -205
rect 2472 -225 2492 -205
<< poly >>
rect 4171 7744 4221 7760
rect 4379 7744 4429 7760
rect 4587 7744 4637 7760
rect 4800 7744 4850 7760
rect 4171 7677 4221 7702
rect 4171 7651 4177 7677
rect 4203 7651 4221 7677
rect 4171 7625 4221 7651
rect 4379 7673 4429 7702
rect 4379 7649 4393 7673
rect 4417 7649 4429 7673
rect 4379 7625 4429 7649
rect 4587 7678 4637 7702
rect 4587 7654 4602 7678
rect 4626 7654 4637 7678
rect 4587 7625 4637 7654
rect 4800 7673 4850 7702
rect 4800 7653 4817 7673
rect 4837 7653 4850 7673
rect 4800 7625 4850 7653
rect 342 7587 392 7600
rect 555 7587 605 7600
rect 763 7587 813 7600
rect 971 7587 1021 7600
rect 3158 7510 3208 7526
rect 3366 7510 3416 7526
rect 3574 7510 3624 7526
rect 3787 7510 3837 7526
rect 4171 7512 4221 7525
rect 4379 7512 4429 7525
rect 4587 7512 4637 7525
rect 4800 7512 4850 7525
rect 342 7459 392 7487
rect 342 7439 355 7459
rect 375 7439 392 7459
rect 342 7410 392 7439
rect 555 7458 605 7487
rect 555 7434 566 7458
rect 590 7434 605 7458
rect 555 7410 605 7434
rect 763 7463 813 7487
rect 763 7439 775 7463
rect 799 7439 813 7463
rect 763 7410 813 7439
rect 971 7461 1021 7487
rect 971 7435 989 7461
rect 1015 7435 1021 7461
rect 971 7410 1021 7435
rect 3158 7443 3208 7468
rect 1354 7406 1404 7419
rect 1567 7406 1617 7419
rect 1775 7406 1825 7419
rect 1983 7406 2033 7419
rect 3158 7417 3164 7443
rect 3190 7417 3208 7443
rect 342 7352 392 7368
rect 555 7352 605 7368
rect 763 7352 813 7368
rect 971 7352 1021 7368
rect 3158 7391 3208 7417
rect 3366 7439 3416 7468
rect 3366 7415 3380 7439
rect 3404 7415 3416 7439
rect 3366 7391 3416 7415
rect 3574 7444 3624 7468
rect 3574 7420 3589 7444
rect 3613 7420 3624 7444
rect 3574 7391 3624 7420
rect 3787 7439 3837 7468
rect 3787 7419 3804 7439
rect 3824 7419 3837 7439
rect 3787 7391 3837 7419
rect 1354 7278 1404 7306
rect 1354 7258 1367 7278
rect 1387 7258 1404 7278
rect 1354 7229 1404 7258
rect 1567 7277 1617 7306
rect 1567 7253 1578 7277
rect 1602 7253 1617 7277
rect 1567 7229 1617 7253
rect 1775 7282 1825 7306
rect 1775 7258 1787 7282
rect 1811 7258 1825 7282
rect 1775 7229 1825 7258
rect 1983 7280 2033 7306
rect 4170 7329 4220 7345
rect 4378 7329 4428 7345
rect 4586 7329 4636 7345
rect 4799 7329 4849 7345
rect 1983 7254 2001 7280
rect 2027 7254 2033 7280
rect 3158 7278 3208 7291
rect 3366 7278 3416 7291
rect 3574 7278 3624 7291
rect 3787 7278 3837 7291
rect 1983 7229 2033 7254
rect 4170 7262 4220 7287
rect 4170 7236 4176 7262
rect 4202 7236 4220 7262
rect 4170 7210 4220 7236
rect 4378 7258 4428 7287
rect 4378 7234 4392 7258
rect 4416 7234 4428 7258
rect 4378 7210 4428 7234
rect 4586 7263 4636 7287
rect 4586 7239 4601 7263
rect 4625 7239 4636 7263
rect 4586 7210 4636 7239
rect 4799 7258 4849 7287
rect 4799 7238 4816 7258
rect 4836 7238 4849 7258
rect 4799 7210 4849 7238
rect 341 7172 391 7185
rect 554 7172 604 7185
rect 762 7172 812 7185
rect 970 7172 1020 7185
rect 1354 7171 1404 7187
rect 1567 7171 1617 7187
rect 1775 7171 1825 7187
rect 1983 7171 2033 7187
rect 3108 7090 3158 7106
rect 3316 7090 3366 7106
rect 3524 7090 3574 7106
rect 3737 7090 3787 7106
rect 4170 7097 4220 7110
rect 4378 7097 4428 7110
rect 4586 7097 4636 7110
rect 4799 7097 4849 7110
rect 341 7044 391 7072
rect 341 7024 354 7044
rect 374 7024 391 7044
rect 341 6995 391 7024
rect 554 7043 604 7072
rect 554 7019 565 7043
rect 589 7019 604 7043
rect 554 6995 604 7019
rect 762 7048 812 7072
rect 762 7024 774 7048
rect 798 7024 812 7048
rect 762 6995 812 7024
rect 970 7046 1020 7072
rect 970 7020 988 7046
rect 1014 7020 1020 7046
rect 970 6995 1020 7020
rect 3108 7023 3158 7048
rect 3108 6997 3114 7023
rect 3140 6997 3158 7023
rect 3108 6971 3158 6997
rect 3316 7019 3366 7048
rect 3316 6995 3330 7019
rect 3354 6995 3366 7019
rect 3316 6971 3366 6995
rect 3524 7024 3574 7048
rect 3524 7000 3539 7024
rect 3563 7000 3574 7024
rect 3524 6971 3574 7000
rect 3737 7019 3787 7048
rect 3737 6999 3754 7019
rect 3774 6999 3787 7019
rect 3737 6971 3787 6999
rect 341 6937 391 6953
rect 554 6937 604 6953
rect 762 6937 812 6953
rect 970 6937 1020 6953
rect 3108 6858 3158 6871
rect 3316 6858 3366 6871
rect 3524 6858 3574 6871
rect 3737 6858 3787 6871
rect 1409 6845 1459 6858
rect 1622 6845 1672 6858
rect 1830 6845 1880 6858
rect 2038 6845 2088 6858
rect 4176 6763 4226 6779
rect 4384 6763 4434 6779
rect 4592 6763 4642 6779
rect 4805 6763 4855 6779
rect 1409 6717 1459 6745
rect 1409 6697 1422 6717
rect 1442 6697 1459 6717
rect 1409 6668 1459 6697
rect 1622 6716 1672 6745
rect 1622 6692 1633 6716
rect 1657 6692 1672 6716
rect 1622 6668 1672 6692
rect 1830 6721 1880 6745
rect 1830 6697 1842 6721
rect 1866 6697 1880 6721
rect 1830 6668 1880 6697
rect 2038 6719 2088 6745
rect 2038 6693 2056 6719
rect 2082 6693 2088 6719
rect 2038 6668 2088 6693
rect 4176 6696 4226 6721
rect 4176 6670 4182 6696
rect 4208 6670 4226 6696
rect 4176 6644 4226 6670
rect 4384 6692 4434 6721
rect 4384 6668 4398 6692
rect 4422 6668 4434 6692
rect 4384 6644 4434 6668
rect 4592 6697 4642 6721
rect 4592 6673 4607 6697
rect 4631 6673 4642 6697
rect 4592 6644 4642 6673
rect 4805 6692 4855 6721
rect 4805 6672 4822 6692
rect 4842 6672 4855 6692
rect 4805 6644 4855 6672
rect 347 6606 397 6619
rect 560 6606 610 6619
rect 768 6606 818 6619
rect 976 6606 1026 6619
rect 1409 6610 1459 6626
rect 1622 6610 1672 6626
rect 1830 6610 1880 6626
rect 2038 6610 2088 6626
rect 3163 6529 3213 6545
rect 3371 6529 3421 6545
rect 3579 6529 3629 6545
rect 3792 6529 3842 6545
rect 4176 6531 4226 6544
rect 4384 6531 4434 6544
rect 4592 6531 4642 6544
rect 4805 6531 4855 6544
rect 347 6478 397 6506
rect 347 6458 360 6478
rect 380 6458 397 6478
rect 347 6429 397 6458
rect 560 6477 610 6506
rect 560 6453 571 6477
rect 595 6453 610 6477
rect 560 6429 610 6453
rect 768 6482 818 6506
rect 768 6458 780 6482
rect 804 6458 818 6482
rect 768 6429 818 6458
rect 976 6480 1026 6506
rect 976 6454 994 6480
rect 1020 6454 1026 6480
rect 976 6429 1026 6454
rect 3163 6462 3213 6487
rect 1359 6425 1409 6438
rect 1572 6425 1622 6438
rect 1780 6425 1830 6438
rect 1988 6425 2038 6438
rect 3163 6436 3169 6462
rect 3195 6436 3213 6462
rect 347 6371 397 6387
rect 560 6371 610 6387
rect 768 6371 818 6387
rect 976 6371 1026 6387
rect 3163 6410 3213 6436
rect 3371 6458 3421 6487
rect 3371 6434 3385 6458
rect 3409 6434 3421 6458
rect 3371 6410 3421 6434
rect 3579 6463 3629 6487
rect 3579 6439 3594 6463
rect 3618 6439 3629 6463
rect 3579 6410 3629 6439
rect 3792 6458 3842 6487
rect 3792 6438 3809 6458
rect 3829 6438 3842 6458
rect 3792 6410 3842 6438
rect 1359 6297 1409 6325
rect 1359 6277 1372 6297
rect 1392 6277 1409 6297
rect 1359 6248 1409 6277
rect 1572 6296 1622 6325
rect 1572 6272 1583 6296
rect 1607 6272 1622 6296
rect 1572 6248 1622 6272
rect 1780 6301 1830 6325
rect 1780 6277 1792 6301
rect 1816 6277 1830 6301
rect 1780 6248 1830 6277
rect 1988 6299 2038 6325
rect 4175 6348 4225 6364
rect 4383 6348 4433 6364
rect 4591 6348 4641 6364
rect 4804 6348 4854 6364
rect 1988 6273 2006 6299
rect 2032 6273 2038 6299
rect 3163 6297 3213 6310
rect 3371 6297 3421 6310
rect 3579 6297 3629 6310
rect 3792 6297 3842 6310
rect 1988 6248 2038 6273
rect 4175 6281 4225 6306
rect 4175 6255 4181 6281
rect 4207 6255 4225 6281
rect 4175 6229 4225 6255
rect 4383 6277 4433 6306
rect 4383 6253 4397 6277
rect 4421 6253 4433 6277
rect 4383 6229 4433 6253
rect 4591 6282 4641 6306
rect 4591 6258 4606 6282
rect 4630 6258 4641 6282
rect 4591 6229 4641 6258
rect 4804 6277 4854 6306
rect 4804 6257 4821 6277
rect 4841 6257 4854 6277
rect 4804 6229 4854 6257
rect 346 6191 396 6204
rect 559 6191 609 6204
rect 767 6191 817 6204
rect 975 6191 1025 6204
rect 1359 6190 1409 6206
rect 1572 6190 1622 6206
rect 1780 6190 1830 6206
rect 1988 6190 2038 6206
rect 4175 6116 4225 6129
rect 4383 6116 4433 6129
rect 4591 6116 4641 6129
rect 4804 6116 4854 6129
rect 346 6063 396 6091
rect 346 6043 359 6063
rect 379 6043 396 6063
rect 346 6014 396 6043
rect 559 6062 609 6091
rect 559 6038 570 6062
rect 594 6038 609 6062
rect 559 6014 609 6038
rect 767 6067 817 6091
rect 767 6043 779 6067
rect 803 6043 817 6067
rect 767 6014 817 6043
rect 975 6065 1025 6091
rect 975 6039 993 6065
rect 1019 6039 1025 6065
rect 2955 6062 3005 6078
rect 3163 6062 3213 6078
rect 3371 6062 3421 6078
rect 3584 6062 3634 6078
rect 975 6014 1025 6039
rect 2955 5995 3005 6020
rect 346 5956 396 5972
rect 559 5956 609 5972
rect 767 5956 817 5972
rect 975 5956 1025 5972
rect 2955 5969 2961 5995
rect 2987 5969 3005 5995
rect 2955 5943 3005 5969
rect 3163 5991 3213 6020
rect 3163 5967 3177 5991
rect 3201 5967 3213 5991
rect 3163 5943 3213 5967
rect 3371 5996 3421 6020
rect 3371 5972 3386 5996
rect 3410 5972 3421 5996
rect 3371 5943 3421 5972
rect 3584 5991 3634 6020
rect 3584 5971 3601 5991
rect 3621 5971 3634 5991
rect 3584 5943 3634 5971
rect 1574 5913 1624 5926
rect 1787 5913 1837 5926
rect 1995 5913 2045 5926
rect 2203 5913 2253 5926
rect 2955 5830 3005 5843
rect 3163 5830 3213 5843
rect 3371 5830 3421 5843
rect 3584 5830 3634 5843
rect 1574 5785 1624 5813
rect 1574 5765 1587 5785
rect 1607 5765 1624 5785
rect 1574 5736 1624 5765
rect 1787 5784 1837 5813
rect 1787 5760 1798 5784
rect 1822 5760 1837 5784
rect 1787 5736 1837 5760
rect 1995 5789 2045 5813
rect 1995 5765 2007 5789
rect 2031 5765 2045 5789
rect 1995 5736 2045 5765
rect 2203 5787 2253 5813
rect 2203 5761 2221 5787
rect 2247 5761 2253 5787
rect 4183 5784 4233 5800
rect 4391 5784 4441 5800
rect 4599 5784 4649 5800
rect 4812 5784 4862 5800
rect 2203 5736 2253 5761
rect 4183 5717 4233 5742
rect 1574 5678 1624 5694
rect 1787 5678 1837 5694
rect 1995 5678 2045 5694
rect 2203 5678 2253 5694
rect 4183 5691 4189 5717
rect 4215 5691 4233 5717
rect 4183 5665 4233 5691
rect 4391 5713 4441 5742
rect 4391 5689 4405 5713
rect 4429 5689 4441 5713
rect 4391 5665 4441 5689
rect 4599 5718 4649 5742
rect 4599 5694 4614 5718
rect 4638 5694 4649 5718
rect 4599 5665 4649 5694
rect 4812 5713 4862 5742
rect 4812 5693 4829 5713
rect 4849 5693 4862 5713
rect 4812 5665 4862 5693
rect 354 5627 404 5640
rect 567 5627 617 5640
rect 775 5627 825 5640
rect 983 5627 1033 5640
rect 3170 5550 3220 5566
rect 3378 5550 3428 5566
rect 3586 5550 3636 5566
rect 3799 5550 3849 5566
rect 4183 5552 4233 5565
rect 4391 5552 4441 5565
rect 4599 5552 4649 5565
rect 4812 5552 4862 5565
rect 354 5499 404 5527
rect 354 5479 367 5499
rect 387 5479 404 5499
rect 354 5450 404 5479
rect 567 5498 617 5527
rect 567 5474 578 5498
rect 602 5474 617 5498
rect 567 5450 617 5474
rect 775 5503 825 5527
rect 775 5479 787 5503
rect 811 5479 825 5503
rect 775 5450 825 5479
rect 983 5501 1033 5527
rect 983 5475 1001 5501
rect 1027 5475 1033 5501
rect 983 5450 1033 5475
rect 3170 5483 3220 5508
rect 1366 5446 1416 5459
rect 1579 5446 1629 5459
rect 1787 5446 1837 5459
rect 1995 5446 2045 5459
rect 3170 5457 3176 5483
rect 3202 5457 3220 5483
rect 354 5392 404 5408
rect 567 5392 617 5408
rect 775 5392 825 5408
rect 983 5392 1033 5408
rect 3170 5431 3220 5457
rect 3378 5479 3428 5508
rect 3378 5455 3392 5479
rect 3416 5455 3428 5479
rect 3378 5431 3428 5455
rect 3586 5484 3636 5508
rect 3586 5460 3601 5484
rect 3625 5460 3636 5484
rect 3586 5431 3636 5460
rect 3799 5479 3849 5508
rect 3799 5459 3816 5479
rect 3836 5459 3849 5479
rect 3799 5431 3849 5459
rect 1366 5318 1416 5346
rect 1366 5298 1379 5318
rect 1399 5298 1416 5318
rect 1366 5269 1416 5298
rect 1579 5317 1629 5346
rect 1579 5293 1590 5317
rect 1614 5293 1629 5317
rect 1579 5269 1629 5293
rect 1787 5322 1837 5346
rect 1787 5298 1799 5322
rect 1823 5298 1837 5322
rect 1787 5269 1837 5298
rect 1995 5320 2045 5346
rect 4182 5369 4232 5385
rect 4390 5369 4440 5385
rect 4598 5369 4648 5385
rect 4811 5369 4861 5385
rect 1995 5294 2013 5320
rect 2039 5294 2045 5320
rect 3170 5318 3220 5331
rect 3378 5318 3428 5331
rect 3586 5318 3636 5331
rect 3799 5318 3849 5331
rect 1995 5269 2045 5294
rect 4182 5302 4232 5327
rect 4182 5276 4188 5302
rect 4214 5276 4232 5302
rect 4182 5250 4232 5276
rect 4390 5298 4440 5327
rect 4390 5274 4404 5298
rect 4428 5274 4440 5298
rect 4390 5250 4440 5274
rect 4598 5303 4648 5327
rect 4598 5279 4613 5303
rect 4637 5279 4648 5303
rect 4598 5250 4648 5279
rect 4811 5298 4861 5327
rect 4811 5278 4828 5298
rect 4848 5278 4861 5298
rect 4811 5250 4861 5278
rect 353 5212 403 5225
rect 566 5212 616 5225
rect 774 5212 824 5225
rect 982 5212 1032 5225
rect 1366 5211 1416 5227
rect 1579 5211 1629 5227
rect 1787 5211 1837 5227
rect 1995 5211 2045 5227
rect 3120 5130 3170 5146
rect 3328 5130 3378 5146
rect 3536 5130 3586 5146
rect 3749 5130 3799 5146
rect 4182 5137 4232 5150
rect 4390 5137 4440 5150
rect 4598 5137 4648 5150
rect 4811 5137 4861 5150
rect 353 5084 403 5112
rect 353 5064 366 5084
rect 386 5064 403 5084
rect 353 5035 403 5064
rect 566 5083 616 5112
rect 566 5059 577 5083
rect 601 5059 616 5083
rect 566 5035 616 5059
rect 774 5088 824 5112
rect 774 5064 786 5088
rect 810 5064 824 5088
rect 774 5035 824 5064
rect 982 5086 1032 5112
rect 982 5060 1000 5086
rect 1026 5060 1032 5086
rect 982 5035 1032 5060
rect 3120 5063 3170 5088
rect 3120 5037 3126 5063
rect 3152 5037 3170 5063
rect 3120 5011 3170 5037
rect 3328 5059 3378 5088
rect 3328 5035 3342 5059
rect 3366 5035 3378 5059
rect 3328 5011 3378 5035
rect 3536 5064 3586 5088
rect 3536 5040 3551 5064
rect 3575 5040 3586 5064
rect 3536 5011 3586 5040
rect 3749 5059 3799 5088
rect 3749 5039 3766 5059
rect 3786 5039 3799 5059
rect 3749 5011 3799 5039
rect 353 4977 403 4993
rect 566 4977 616 4993
rect 774 4977 824 4993
rect 982 4977 1032 4993
rect 3120 4898 3170 4911
rect 3328 4898 3378 4911
rect 3536 4898 3586 4911
rect 3749 4898 3799 4911
rect 1421 4885 1471 4898
rect 1634 4885 1684 4898
rect 1842 4885 1892 4898
rect 2050 4885 2100 4898
rect 4188 4803 4238 4819
rect 4396 4803 4446 4819
rect 4604 4803 4654 4819
rect 4817 4803 4867 4819
rect 1421 4757 1471 4785
rect 1421 4737 1434 4757
rect 1454 4737 1471 4757
rect 1421 4708 1471 4737
rect 1634 4756 1684 4785
rect 1634 4732 1645 4756
rect 1669 4732 1684 4756
rect 1634 4708 1684 4732
rect 1842 4761 1892 4785
rect 1842 4737 1854 4761
rect 1878 4737 1892 4761
rect 1842 4708 1892 4737
rect 2050 4759 2100 4785
rect 2050 4733 2068 4759
rect 2094 4733 2100 4759
rect 2050 4708 2100 4733
rect 4188 4736 4238 4761
rect 4188 4710 4194 4736
rect 4220 4710 4238 4736
rect 4188 4684 4238 4710
rect 4396 4732 4446 4761
rect 4396 4708 4410 4732
rect 4434 4708 4446 4732
rect 4396 4684 4446 4708
rect 4604 4737 4654 4761
rect 4604 4713 4619 4737
rect 4643 4713 4654 4737
rect 4604 4684 4654 4713
rect 4817 4732 4867 4761
rect 4817 4712 4834 4732
rect 4854 4712 4867 4732
rect 4817 4684 4867 4712
rect 359 4646 409 4659
rect 572 4646 622 4659
rect 780 4646 830 4659
rect 988 4646 1038 4659
rect 1421 4650 1471 4666
rect 1634 4650 1684 4666
rect 1842 4650 1892 4666
rect 2050 4650 2100 4666
rect 3175 4569 3225 4585
rect 3383 4569 3433 4585
rect 3591 4569 3641 4585
rect 3804 4569 3854 4585
rect 4188 4571 4238 4584
rect 4396 4571 4446 4584
rect 4604 4571 4654 4584
rect 4817 4571 4867 4584
rect 359 4518 409 4546
rect 359 4498 372 4518
rect 392 4498 409 4518
rect 359 4469 409 4498
rect 572 4517 622 4546
rect 572 4493 583 4517
rect 607 4493 622 4517
rect 572 4469 622 4493
rect 780 4522 830 4546
rect 780 4498 792 4522
rect 816 4498 830 4522
rect 780 4469 830 4498
rect 988 4520 1038 4546
rect 988 4494 1006 4520
rect 1032 4494 1038 4520
rect 988 4469 1038 4494
rect 3175 4502 3225 4527
rect 1371 4465 1421 4478
rect 1584 4465 1634 4478
rect 1792 4465 1842 4478
rect 2000 4465 2050 4478
rect 3175 4476 3181 4502
rect 3207 4476 3225 4502
rect 359 4411 409 4427
rect 572 4411 622 4427
rect 780 4411 830 4427
rect 988 4411 1038 4427
rect 3175 4450 3225 4476
rect 3383 4498 3433 4527
rect 3383 4474 3397 4498
rect 3421 4474 3433 4498
rect 3383 4450 3433 4474
rect 3591 4503 3641 4527
rect 3591 4479 3606 4503
rect 3630 4479 3641 4503
rect 3591 4450 3641 4479
rect 3804 4498 3854 4527
rect 3804 4478 3821 4498
rect 3841 4478 3854 4498
rect 3804 4450 3854 4478
rect 1371 4337 1421 4365
rect 1371 4317 1384 4337
rect 1404 4317 1421 4337
rect 1371 4288 1421 4317
rect 1584 4336 1634 4365
rect 1584 4312 1595 4336
rect 1619 4312 1634 4336
rect 1584 4288 1634 4312
rect 1792 4341 1842 4365
rect 1792 4317 1804 4341
rect 1828 4317 1842 4341
rect 1792 4288 1842 4317
rect 2000 4339 2050 4365
rect 4187 4388 4237 4404
rect 4395 4388 4445 4404
rect 4603 4388 4653 4404
rect 4816 4388 4866 4404
rect 2000 4313 2018 4339
rect 2044 4313 2050 4339
rect 3175 4337 3225 4350
rect 3383 4337 3433 4350
rect 3591 4337 3641 4350
rect 3804 4337 3854 4350
rect 2000 4288 2050 4313
rect 4187 4321 4237 4346
rect 4187 4295 4193 4321
rect 4219 4295 4237 4321
rect 4187 4269 4237 4295
rect 4395 4317 4445 4346
rect 4395 4293 4409 4317
rect 4433 4293 4445 4317
rect 4395 4269 4445 4293
rect 4603 4322 4653 4346
rect 4603 4298 4618 4322
rect 4642 4298 4653 4322
rect 4603 4269 4653 4298
rect 4816 4317 4866 4346
rect 4816 4297 4833 4317
rect 4853 4297 4866 4317
rect 4816 4269 4866 4297
rect 358 4231 408 4244
rect 571 4231 621 4244
rect 779 4231 829 4244
rect 987 4231 1037 4244
rect 1371 4230 1421 4246
rect 1584 4230 1634 4246
rect 1792 4230 1842 4246
rect 2000 4230 2050 4246
rect 4187 4156 4237 4169
rect 4395 4156 4445 4169
rect 4603 4156 4653 4169
rect 4816 4156 4866 4169
rect 2880 4137 2930 4153
rect 3088 4137 3138 4153
rect 3296 4137 3346 4153
rect 3509 4137 3559 4153
rect 358 4103 408 4131
rect 358 4083 371 4103
rect 391 4083 408 4103
rect 358 4054 408 4083
rect 571 4102 621 4131
rect 571 4078 582 4102
rect 606 4078 621 4102
rect 571 4054 621 4078
rect 779 4107 829 4131
rect 779 4083 791 4107
rect 815 4083 829 4107
rect 779 4054 829 4083
rect 987 4105 1037 4131
rect 987 4079 1005 4105
rect 1031 4079 1037 4105
rect 987 4054 1037 4079
rect 2880 4070 2930 4095
rect 2880 4044 2886 4070
rect 2912 4044 2930 4070
rect 2880 4018 2930 4044
rect 3088 4066 3138 4095
rect 3088 4042 3102 4066
rect 3126 4042 3138 4066
rect 3088 4018 3138 4042
rect 3296 4071 3346 4095
rect 3296 4047 3311 4071
rect 3335 4047 3346 4071
rect 3296 4018 3346 4047
rect 3509 4066 3559 4095
rect 3509 4046 3526 4066
rect 3546 4046 3559 4066
rect 3509 4018 3559 4046
rect 358 3996 408 4012
rect 571 3996 621 4012
rect 779 3996 829 4012
rect 987 3996 1037 4012
rect 1669 3921 1719 3934
rect 1882 3921 1932 3934
rect 2090 3921 2140 3934
rect 2298 3921 2348 3934
rect 2880 3905 2930 3918
rect 3088 3905 3138 3918
rect 3296 3905 3346 3918
rect 3509 3905 3559 3918
rect 4191 3827 4241 3843
rect 4399 3827 4449 3843
rect 4607 3827 4657 3843
rect 4820 3827 4870 3843
rect 1669 3793 1719 3821
rect 1669 3773 1682 3793
rect 1702 3773 1719 3793
rect 1669 3744 1719 3773
rect 1882 3792 1932 3821
rect 1882 3768 1893 3792
rect 1917 3768 1932 3792
rect 1882 3744 1932 3768
rect 2090 3797 2140 3821
rect 2090 3773 2102 3797
rect 2126 3773 2140 3797
rect 2090 3744 2140 3773
rect 2298 3795 2348 3821
rect 2298 3769 2316 3795
rect 2342 3769 2348 3795
rect 2298 3744 2348 3769
rect 4191 3760 4241 3785
rect 4191 3734 4197 3760
rect 4223 3734 4241 3760
rect 4191 3708 4241 3734
rect 4399 3756 4449 3785
rect 4399 3732 4413 3756
rect 4437 3732 4449 3756
rect 4399 3708 4449 3732
rect 4607 3761 4657 3785
rect 4607 3737 4622 3761
rect 4646 3737 4657 3761
rect 4607 3708 4657 3737
rect 4820 3756 4870 3785
rect 4820 3736 4837 3756
rect 4857 3736 4870 3756
rect 4820 3708 4870 3736
rect 1669 3686 1719 3702
rect 1882 3686 1932 3702
rect 2090 3686 2140 3702
rect 2298 3686 2348 3702
rect 362 3670 412 3683
rect 575 3670 625 3683
rect 783 3670 833 3683
rect 991 3670 1041 3683
rect 3178 3593 3228 3609
rect 3386 3593 3436 3609
rect 3594 3593 3644 3609
rect 3807 3593 3857 3609
rect 4191 3595 4241 3608
rect 4399 3595 4449 3608
rect 4607 3595 4657 3608
rect 4820 3595 4870 3608
rect 362 3542 412 3570
rect 362 3522 375 3542
rect 395 3522 412 3542
rect 362 3493 412 3522
rect 575 3541 625 3570
rect 575 3517 586 3541
rect 610 3517 625 3541
rect 575 3493 625 3517
rect 783 3546 833 3570
rect 783 3522 795 3546
rect 819 3522 833 3546
rect 783 3493 833 3522
rect 991 3544 1041 3570
rect 991 3518 1009 3544
rect 1035 3518 1041 3544
rect 991 3493 1041 3518
rect 3178 3526 3228 3551
rect 1374 3489 1424 3502
rect 1587 3489 1637 3502
rect 1795 3489 1845 3502
rect 2003 3489 2053 3502
rect 3178 3500 3184 3526
rect 3210 3500 3228 3526
rect 362 3435 412 3451
rect 575 3435 625 3451
rect 783 3435 833 3451
rect 991 3435 1041 3451
rect 3178 3474 3228 3500
rect 3386 3522 3436 3551
rect 3386 3498 3400 3522
rect 3424 3498 3436 3522
rect 3386 3474 3436 3498
rect 3594 3527 3644 3551
rect 3594 3503 3609 3527
rect 3633 3503 3644 3527
rect 3594 3474 3644 3503
rect 3807 3522 3857 3551
rect 3807 3502 3824 3522
rect 3844 3502 3857 3522
rect 3807 3474 3857 3502
rect 1374 3361 1424 3389
rect 1374 3341 1387 3361
rect 1407 3341 1424 3361
rect 1374 3312 1424 3341
rect 1587 3360 1637 3389
rect 1587 3336 1598 3360
rect 1622 3336 1637 3360
rect 1587 3312 1637 3336
rect 1795 3365 1845 3389
rect 1795 3341 1807 3365
rect 1831 3341 1845 3365
rect 1795 3312 1845 3341
rect 2003 3363 2053 3389
rect 4190 3412 4240 3428
rect 4398 3412 4448 3428
rect 4606 3412 4656 3428
rect 4819 3412 4869 3428
rect 2003 3337 2021 3363
rect 2047 3337 2053 3363
rect 3178 3361 3228 3374
rect 3386 3361 3436 3374
rect 3594 3361 3644 3374
rect 3807 3361 3857 3374
rect 2003 3312 2053 3337
rect 4190 3345 4240 3370
rect 4190 3319 4196 3345
rect 4222 3319 4240 3345
rect 4190 3293 4240 3319
rect 4398 3341 4448 3370
rect 4398 3317 4412 3341
rect 4436 3317 4448 3341
rect 4398 3293 4448 3317
rect 4606 3346 4656 3370
rect 4606 3322 4621 3346
rect 4645 3322 4656 3346
rect 4606 3293 4656 3322
rect 4819 3341 4869 3370
rect 4819 3321 4836 3341
rect 4856 3321 4869 3341
rect 4819 3293 4869 3321
rect 361 3255 411 3268
rect 574 3255 624 3268
rect 782 3255 832 3268
rect 990 3255 1040 3268
rect 1374 3254 1424 3270
rect 1587 3254 1637 3270
rect 1795 3254 1845 3270
rect 2003 3254 2053 3270
rect 3128 3173 3178 3189
rect 3336 3173 3386 3189
rect 3544 3173 3594 3189
rect 3757 3173 3807 3189
rect 4190 3180 4240 3193
rect 4398 3180 4448 3193
rect 4606 3180 4656 3193
rect 4819 3180 4869 3193
rect 361 3127 411 3155
rect 361 3107 374 3127
rect 394 3107 411 3127
rect 361 3078 411 3107
rect 574 3126 624 3155
rect 574 3102 585 3126
rect 609 3102 624 3126
rect 574 3078 624 3102
rect 782 3131 832 3155
rect 782 3107 794 3131
rect 818 3107 832 3131
rect 782 3078 832 3107
rect 990 3129 1040 3155
rect 990 3103 1008 3129
rect 1034 3103 1040 3129
rect 990 3078 1040 3103
rect 3128 3106 3178 3131
rect 3128 3080 3134 3106
rect 3160 3080 3178 3106
rect 3128 3054 3178 3080
rect 3336 3102 3386 3131
rect 3336 3078 3350 3102
rect 3374 3078 3386 3102
rect 3336 3054 3386 3078
rect 3544 3107 3594 3131
rect 3544 3083 3559 3107
rect 3583 3083 3594 3107
rect 3544 3054 3594 3083
rect 3757 3102 3807 3131
rect 3757 3082 3774 3102
rect 3794 3082 3807 3102
rect 3757 3054 3807 3082
rect 361 3020 411 3036
rect 574 3020 624 3036
rect 782 3020 832 3036
rect 990 3020 1040 3036
rect 3128 2941 3178 2954
rect 3336 2941 3386 2954
rect 3544 2941 3594 2954
rect 3757 2941 3807 2954
rect 1429 2928 1479 2941
rect 1642 2928 1692 2941
rect 1850 2928 1900 2941
rect 2058 2928 2108 2941
rect 4196 2846 4246 2862
rect 4404 2846 4454 2862
rect 4612 2846 4662 2862
rect 4825 2846 4875 2862
rect 1429 2800 1479 2828
rect 1429 2780 1442 2800
rect 1462 2780 1479 2800
rect 1429 2751 1479 2780
rect 1642 2799 1692 2828
rect 1642 2775 1653 2799
rect 1677 2775 1692 2799
rect 1642 2751 1692 2775
rect 1850 2804 1900 2828
rect 1850 2780 1862 2804
rect 1886 2780 1900 2804
rect 1850 2751 1900 2780
rect 2058 2802 2108 2828
rect 2058 2776 2076 2802
rect 2102 2776 2108 2802
rect 2058 2751 2108 2776
rect 4196 2779 4246 2804
rect 4196 2753 4202 2779
rect 4228 2753 4246 2779
rect 4196 2727 4246 2753
rect 4404 2775 4454 2804
rect 4404 2751 4418 2775
rect 4442 2751 4454 2775
rect 4404 2727 4454 2751
rect 4612 2780 4662 2804
rect 4612 2756 4627 2780
rect 4651 2756 4662 2780
rect 4612 2727 4662 2756
rect 4825 2775 4875 2804
rect 4825 2755 4842 2775
rect 4862 2755 4875 2775
rect 4825 2727 4875 2755
rect 367 2689 417 2702
rect 580 2689 630 2702
rect 788 2689 838 2702
rect 996 2689 1046 2702
rect 1429 2693 1479 2709
rect 1642 2693 1692 2709
rect 1850 2693 1900 2709
rect 2058 2693 2108 2709
rect 3183 2612 3233 2628
rect 3391 2612 3441 2628
rect 3599 2612 3649 2628
rect 3812 2612 3862 2628
rect 4196 2614 4246 2627
rect 4404 2614 4454 2627
rect 4612 2614 4662 2627
rect 4825 2614 4875 2627
rect 367 2561 417 2589
rect 367 2541 380 2561
rect 400 2541 417 2561
rect 367 2512 417 2541
rect 580 2560 630 2589
rect 580 2536 591 2560
rect 615 2536 630 2560
rect 580 2512 630 2536
rect 788 2565 838 2589
rect 788 2541 800 2565
rect 824 2541 838 2565
rect 788 2512 838 2541
rect 996 2563 1046 2589
rect 996 2537 1014 2563
rect 1040 2537 1046 2563
rect 996 2512 1046 2537
rect 3183 2545 3233 2570
rect 1379 2508 1429 2521
rect 1592 2508 1642 2521
rect 1800 2508 1850 2521
rect 2008 2508 2058 2521
rect 3183 2519 3189 2545
rect 3215 2519 3233 2545
rect 367 2454 417 2470
rect 580 2454 630 2470
rect 788 2454 838 2470
rect 996 2454 1046 2470
rect 3183 2493 3233 2519
rect 3391 2541 3441 2570
rect 3391 2517 3405 2541
rect 3429 2517 3441 2541
rect 3391 2493 3441 2517
rect 3599 2546 3649 2570
rect 3599 2522 3614 2546
rect 3638 2522 3649 2546
rect 3599 2493 3649 2522
rect 3812 2541 3862 2570
rect 3812 2521 3829 2541
rect 3849 2521 3862 2541
rect 3812 2493 3862 2521
rect 1379 2380 1429 2408
rect 1379 2360 1392 2380
rect 1412 2360 1429 2380
rect 1379 2331 1429 2360
rect 1592 2379 1642 2408
rect 1592 2355 1603 2379
rect 1627 2355 1642 2379
rect 1592 2331 1642 2355
rect 1800 2384 1850 2408
rect 1800 2360 1812 2384
rect 1836 2360 1850 2384
rect 1800 2331 1850 2360
rect 2008 2382 2058 2408
rect 4195 2431 4245 2447
rect 4403 2431 4453 2447
rect 4611 2431 4661 2447
rect 4824 2431 4874 2447
rect 2008 2356 2026 2382
rect 2052 2356 2058 2382
rect 3183 2380 3233 2393
rect 3391 2380 3441 2393
rect 3599 2380 3649 2393
rect 3812 2380 3862 2393
rect 2008 2331 2058 2356
rect 4195 2364 4245 2389
rect 4195 2338 4201 2364
rect 4227 2338 4245 2364
rect 4195 2312 4245 2338
rect 4403 2360 4453 2389
rect 4403 2336 4417 2360
rect 4441 2336 4453 2360
rect 4403 2312 4453 2336
rect 4611 2365 4661 2389
rect 4611 2341 4626 2365
rect 4650 2341 4661 2365
rect 4611 2312 4661 2341
rect 4824 2360 4874 2389
rect 4824 2340 4841 2360
rect 4861 2340 4874 2360
rect 4824 2312 4874 2340
rect 366 2274 416 2287
rect 579 2274 629 2287
rect 787 2274 837 2287
rect 995 2274 1045 2287
rect 1379 2273 1429 2289
rect 1592 2273 1642 2289
rect 1800 2273 1850 2289
rect 2008 2273 2058 2289
rect 4195 2199 4245 2212
rect 4403 2199 4453 2212
rect 4611 2199 4661 2212
rect 4824 2199 4874 2212
rect 366 2146 416 2174
rect 366 2126 379 2146
rect 399 2126 416 2146
rect 366 2097 416 2126
rect 579 2145 629 2174
rect 579 2121 590 2145
rect 614 2121 629 2145
rect 579 2097 629 2121
rect 787 2150 837 2174
rect 787 2126 799 2150
rect 823 2126 837 2150
rect 787 2097 837 2126
rect 995 2148 1045 2174
rect 995 2122 1013 2148
rect 1039 2122 1045 2148
rect 2975 2145 3025 2161
rect 3183 2145 3233 2161
rect 3391 2145 3441 2161
rect 3604 2145 3654 2161
rect 995 2097 1045 2122
rect 2975 2078 3025 2103
rect 366 2039 416 2055
rect 579 2039 629 2055
rect 787 2039 837 2055
rect 995 2039 1045 2055
rect 2975 2052 2981 2078
rect 3007 2052 3025 2078
rect 2975 2026 3025 2052
rect 3183 2074 3233 2103
rect 3183 2050 3197 2074
rect 3221 2050 3233 2074
rect 3183 2026 3233 2050
rect 3391 2079 3441 2103
rect 3391 2055 3406 2079
rect 3430 2055 3441 2079
rect 3391 2026 3441 2055
rect 3604 2074 3654 2103
rect 3604 2054 3621 2074
rect 3641 2054 3654 2074
rect 3604 2026 3654 2054
rect 1594 1996 1644 2009
rect 1807 1996 1857 2009
rect 2015 1996 2065 2009
rect 2223 1996 2273 2009
rect 2975 1913 3025 1926
rect 3183 1913 3233 1926
rect 3391 1913 3441 1926
rect 3604 1913 3654 1926
rect 1594 1868 1644 1896
rect 1594 1848 1607 1868
rect 1627 1848 1644 1868
rect 1594 1819 1644 1848
rect 1807 1867 1857 1896
rect 1807 1843 1818 1867
rect 1842 1843 1857 1867
rect 1807 1819 1857 1843
rect 2015 1872 2065 1896
rect 2015 1848 2027 1872
rect 2051 1848 2065 1872
rect 2015 1819 2065 1848
rect 2223 1870 2273 1896
rect 2223 1844 2241 1870
rect 2267 1844 2273 1870
rect 4203 1867 4253 1883
rect 4411 1867 4461 1883
rect 4619 1867 4669 1883
rect 4832 1867 4882 1883
rect 2223 1819 2273 1844
rect 4203 1800 4253 1825
rect 1594 1761 1644 1777
rect 1807 1761 1857 1777
rect 2015 1761 2065 1777
rect 2223 1761 2273 1777
rect 4203 1774 4209 1800
rect 4235 1774 4253 1800
rect 4203 1748 4253 1774
rect 4411 1796 4461 1825
rect 4411 1772 4425 1796
rect 4449 1772 4461 1796
rect 4411 1748 4461 1772
rect 4619 1801 4669 1825
rect 4619 1777 4634 1801
rect 4658 1777 4669 1801
rect 4619 1748 4669 1777
rect 4832 1796 4882 1825
rect 4832 1776 4849 1796
rect 4869 1776 4882 1796
rect 4832 1748 4882 1776
rect 374 1710 424 1723
rect 587 1710 637 1723
rect 795 1710 845 1723
rect 1003 1710 1053 1723
rect 3190 1633 3240 1649
rect 3398 1633 3448 1649
rect 3606 1633 3656 1649
rect 3819 1633 3869 1649
rect 4203 1635 4253 1648
rect 4411 1635 4461 1648
rect 4619 1635 4669 1648
rect 4832 1635 4882 1648
rect 374 1582 424 1610
rect 374 1562 387 1582
rect 407 1562 424 1582
rect 374 1533 424 1562
rect 587 1581 637 1610
rect 587 1557 598 1581
rect 622 1557 637 1581
rect 587 1533 637 1557
rect 795 1586 845 1610
rect 795 1562 807 1586
rect 831 1562 845 1586
rect 795 1533 845 1562
rect 1003 1584 1053 1610
rect 1003 1558 1021 1584
rect 1047 1558 1053 1584
rect 1003 1533 1053 1558
rect 3190 1566 3240 1591
rect 1386 1529 1436 1542
rect 1599 1529 1649 1542
rect 1807 1529 1857 1542
rect 2015 1529 2065 1542
rect 3190 1540 3196 1566
rect 3222 1540 3240 1566
rect 374 1475 424 1491
rect 587 1475 637 1491
rect 795 1475 845 1491
rect 1003 1475 1053 1491
rect 3190 1514 3240 1540
rect 3398 1562 3448 1591
rect 3398 1538 3412 1562
rect 3436 1538 3448 1562
rect 3398 1514 3448 1538
rect 3606 1567 3656 1591
rect 3606 1543 3621 1567
rect 3645 1543 3656 1567
rect 3606 1514 3656 1543
rect 3819 1562 3869 1591
rect 3819 1542 3836 1562
rect 3856 1542 3869 1562
rect 3819 1514 3869 1542
rect 1386 1401 1436 1429
rect 1386 1381 1399 1401
rect 1419 1381 1436 1401
rect 1386 1352 1436 1381
rect 1599 1400 1649 1429
rect 1599 1376 1610 1400
rect 1634 1376 1649 1400
rect 1599 1352 1649 1376
rect 1807 1405 1857 1429
rect 1807 1381 1819 1405
rect 1843 1381 1857 1405
rect 1807 1352 1857 1381
rect 2015 1403 2065 1429
rect 4202 1452 4252 1468
rect 4410 1452 4460 1468
rect 4618 1452 4668 1468
rect 4831 1452 4881 1468
rect 2015 1377 2033 1403
rect 2059 1377 2065 1403
rect 3190 1401 3240 1414
rect 3398 1401 3448 1414
rect 3606 1401 3656 1414
rect 3819 1401 3869 1414
rect 2015 1352 2065 1377
rect 4202 1385 4252 1410
rect 4202 1359 4208 1385
rect 4234 1359 4252 1385
rect 4202 1333 4252 1359
rect 4410 1381 4460 1410
rect 4410 1357 4424 1381
rect 4448 1357 4460 1381
rect 4410 1333 4460 1357
rect 4618 1386 4668 1410
rect 4618 1362 4633 1386
rect 4657 1362 4668 1386
rect 4618 1333 4668 1362
rect 4831 1381 4881 1410
rect 4831 1361 4848 1381
rect 4868 1361 4881 1381
rect 4831 1333 4881 1361
rect 373 1295 423 1308
rect 586 1295 636 1308
rect 794 1295 844 1308
rect 1002 1295 1052 1308
rect 1386 1294 1436 1310
rect 1599 1294 1649 1310
rect 1807 1294 1857 1310
rect 2015 1294 2065 1310
rect 3140 1213 3190 1229
rect 3348 1213 3398 1229
rect 3556 1213 3606 1229
rect 3769 1213 3819 1229
rect 4202 1220 4252 1233
rect 4410 1220 4460 1233
rect 4618 1220 4668 1233
rect 4831 1220 4881 1233
rect 373 1167 423 1195
rect 373 1147 386 1167
rect 406 1147 423 1167
rect 373 1118 423 1147
rect 586 1166 636 1195
rect 586 1142 597 1166
rect 621 1142 636 1166
rect 586 1118 636 1142
rect 794 1171 844 1195
rect 794 1147 806 1171
rect 830 1147 844 1171
rect 794 1118 844 1147
rect 1002 1169 1052 1195
rect 1002 1143 1020 1169
rect 1046 1143 1052 1169
rect 1002 1118 1052 1143
rect 3140 1146 3190 1171
rect 3140 1120 3146 1146
rect 3172 1120 3190 1146
rect 3140 1094 3190 1120
rect 3348 1142 3398 1171
rect 3348 1118 3362 1142
rect 3386 1118 3398 1142
rect 3348 1094 3398 1118
rect 3556 1147 3606 1171
rect 3556 1123 3571 1147
rect 3595 1123 3606 1147
rect 3556 1094 3606 1123
rect 3769 1142 3819 1171
rect 3769 1122 3786 1142
rect 3806 1122 3819 1142
rect 3769 1094 3819 1122
rect 373 1060 423 1076
rect 586 1060 636 1076
rect 794 1060 844 1076
rect 1002 1060 1052 1076
rect 3140 981 3190 994
rect 3348 981 3398 994
rect 3556 981 3606 994
rect 3769 981 3819 994
rect 1441 968 1491 981
rect 1654 968 1704 981
rect 1862 968 1912 981
rect 2070 968 2120 981
rect 4208 886 4258 902
rect 4416 886 4466 902
rect 4624 886 4674 902
rect 4837 886 4887 902
rect 1441 840 1491 868
rect 1441 820 1454 840
rect 1474 820 1491 840
rect 1441 791 1491 820
rect 1654 839 1704 868
rect 1654 815 1665 839
rect 1689 815 1704 839
rect 1654 791 1704 815
rect 1862 844 1912 868
rect 1862 820 1874 844
rect 1898 820 1912 844
rect 1862 791 1912 820
rect 2070 842 2120 868
rect 2070 816 2088 842
rect 2114 816 2120 842
rect 2070 791 2120 816
rect 4208 819 4258 844
rect 4208 793 4214 819
rect 4240 793 4258 819
rect 4208 767 4258 793
rect 4416 815 4466 844
rect 4416 791 4430 815
rect 4454 791 4466 815
rect 4416 767 4466 791
rect 4624 820 4674 844
rect 4624 796 4639 820
rect 4663 796 4674 820
rect 4624 767 4674 796
rect 4837 815 4887 844
rect 4837 795 4854 815
rect 4874 795 4887 815
rect 4837 767 4887 795
rect 379 729 429 742
rect 592 729 642 742
rect 800 729 850 742
rect 1008 729 1058 742
rect 1441 733 1491 749
rect 1654 733 1704 749
rect 1862 733 1912 749
rect 2070 733 2120 749
rect 3195 652 3245 668
rect 3403 652 3453 668
rect 3611 652 3661 668
rect 3824 652 3874 668
rect 4208 654 4258 667
rect 4416 654 4466 667
rect 4624 654 4674 667
rect 4837 654 4887 667
rect 379 601 429 629
rect 379 581 392 601
rect 412 581 429 601
rect 379 552 429 581
rect 592 600 642 629
rect 592 576 603 600
rect 627 576 642 600
rect 592 552 642 576
rect 800 605 850 629
rect 800 581 812 605
rect 836 581 850 605
rect 800 552 850 581
rect 1008 603 1058 629
rect 1008 577 1026 603
rect 1052 577 1058 603
rect 1008 552 1058 577
rect 3195 585 3245 610
rect 1391 548 1441 561
rect 1604 548 1654 561
rect 1812 548 1862 561
rect 2020 548 2070 561
rect 3195 559 3201 585
rect 3227 559 3245 585
rect 379 494 429 510
rect 592 494 642 510
rect 800 494 850 510
rect 1008 494 1058 510
rect 3195 533 3245 559
rect 3403 581 3453 610
rect 3403 557 3417 581
rect 3441 557 3453 581
rect 3403 533 3453 557
rect 3611 586 3661 610
rect 3611 562 3626 586
rect 3650 562 3661 586
rect 3611 533 3661 562
rect 3824 581 3874 610
rect 3824 561 3841 581
rect 3861 561 3874 581
rect 3824 533 3874 561
rect 1391 420 1441 448
rect 1391 400 1404 420
rect 1424 400 1441 420
rect 1391 371 1441 400
rect 1604 419 1654 448
rect 1604 395 1615 419
rect 1639 395 1654 419
rect 1604 371 1654 395
rect 1812 424 1862 448
rect 1812 400 1824 424
rect 1848 400 1862 424
rect 1812 371 1862 400
rect 2020 422 2070 448
rect 4207 471 4257 487
rect 4415 471 4465 487
rect 4623 471 4673 487
rect 4836 471 4886 487
rect 2020 396 2038 422
rect 2064 396 2070 422
rect 3195 420 3245 433
rect 3403 420 3453 433
rect 3611 420 3661 433
rect 3824 420 3874 433
rect 2020 371 2070 396
rect 4207 404 4257 429
rect 4207 378 4213 404
rect 4239 378 4257 404
rect 4207 352 4257 378
rect 4415 400 4465 429
rect 4415 376 4429 400
rect 4453 376 4465 400
rect 4415 352 4465 376
rect 4623 405 4673 429
rect 4623 381 4638 405
rect 4662 381 4673 405
rect 4623 352 4673 381
rect 4836 400 4886 429
rect 4836 380 4853 400
rect 4873 380 4886 400
rect 4836 352 4886 380
rect 378 314 428 327
rect 591 314 641 327
rect 799 314 849 327
rect 1007 314 1057 327
rect 1391 313 1441 329
rect 1604 313 1654 329
rect 1812 313 1862 329
rect 2020 313 2070 329
rect 4207 239 4257 252
rect 4415 239 4465 252
rect 4623 239 4673 252
rect 4836 239 4886 252
rect 378 186 428 214
rect 378 166 391 186
rect 411 166 428 186
rect 378 137 428 166
rect 591 185 641 214
rect 591 161 602 185
rect 626 161 641 185
rect 591 137 641 161
rect 799 190 849 214
rect 799 166 811 190
rect 835 166 849 190
rect 799 137 849 166
rect 1007 188 1057 214
rect 1007 162 1025 188
rect 1051 162 1057 188
rect 1007 137 1057 162
rect 378 79 428 95
rect 591 79 641 95
rect 799 79 849 95
rect 1007 79 1057 95
rect 1781 -167 1831 -154
rect 1994 -167 2044 -154
rect 2202 -167 2252 -154
rect 2410 -167 2460 -154
rect 1781 -295 1831 -267
rect 1781 -315 1794 -295
rect 1814 -315 1831 -295
rect 1781 -344 1831 -315
rect 1994 -296 2044 -267
rect 1994 -320 2005 -296
rect 2029 -320 2044 -296
rect 1994 -344 2044 -320
rect 2202 -291 2252 -267
rect 2202 -315 2214 -291
rect 2238 -315 2252 -291
rect 2202 -344 2252 -315
rect 2410 -293 2460 -267
rect 2410 -319 2428 -293
rect 2454 -319 2460 -293
rect 2410 -344 2460 -319
rect 1781 -402 1831 -386
rect 1994 -402 2044 -386
rect 2202 -402 2252 -386
rect 2410 -402 2460 -386
<< polycont >>
rect 4177 7651 4203 7677
rect 4393 7649 4417 7673
rect 4602 7654 4626 7678
rect 4817 7653 4837 7673
rect 355 7439 375 7459
rect 566 7434 590 7458
rect 775 7439 799 7463
rect 989 7435 1015 7461
rect 3164 7417 3190 7443
rect 3380 7415 3404 7439
rect 3589 7420 3613 7444
rect 3804 7419 3824 7439
rect 1367 7258 1387 7278
rect 1578 7253 1602 7277
rect 1787 7258 1811 7282
rect 2001 7254 2027 7280
rect 4176 7236 4202 7262
rect 4392 7234 4416 7258
rect 4601 7239 4625 7263
rect 4816 7238 4836 7258
rect 354 7024 374 7044
rect 565 7019 589 7043
rect 774 7024 798 7048
rect 988 7020 1014 7046
rect 3114 6997 3140 7023
rect 3330 6995 3354 7019
rect 3539 7000 3563 7024
rect 3754 6999 3774 7019
rect 1422 6697 1442 6717
rect 1633 6692 1657 6716
rect 1842 6697 1866 6721
rect 2056 6693 2082 6719
rect 4182 6670 4208 6696
rect 4398 6668 4422 6692
rect 4607 6673 4631 6697
rect 4822 6672 4842 6692
rect 360 6458 380 6478
rect 571 6453 595 6477
rect 780 6458 804 6482
rect 994 6454 1020 6480
rect 3169 6436 3195 6462
rect 3385 6434 3409 6458
rect 3594 6439 3618 6463
rect 3809 6438 3829 6458
rect 1372 6277 1392 6297
rect 1583 6272 1607 6296
rect 1792 6277 1816 6301
rect 2006 6273 2032 6299
rect 4181 6255 4207 6281
rect 4397 6253 4421 6277
rect 4606 6258 4630 6282
rect 4821 6257 4841 6277
rect 359 6043 379 6063
rect 570 6038 594 6062
rect 779 6043 803 6067
rect 993 6039 1019 6065
rect 2961 5969 2987 5995
rect 3177 5967 3201 5991
rect 3386 5972 3410 5996
rect 3601 5971 3621 5991
rect 1587 5765 1607 5785
rect 1798 5760 1822 5784
rect 2007 5765 2031 5789
rect 2221 5761 2247 5787
rect 4189 5691 4215 5717
rect 4405 5689 4429 5713
rect 4614 5694 4638 5718
rect 4829 5693 4849 5713
rect 367 5479 387 5499
rect 578 5474 602 5498
rect 787 5479 811 5503
rect 1001 5475 1027 5501
rect 3176 5457 3202 5483
rect 3392 5455 3416 5479
rect 3601 5460 3625 5484
rect 3816 5459 3836 5479
rect 1379 5298 1399 5318
rect 1590 5293 1614 5317
rect 1799 5298 1823 5322
rect 2013 5294 2039 5320
rect 4188 5276 4214 5302
rect 4404 5274 4428 5298
rect 4613 5279 4637 5303
rect 4828 5278 4848 5298
rect 366 5064 386 5084
rect 577 5059 601 5083
rect 786 5064 810 5088
rect 1000 5060 1026 5086
rect 3126 5037 3152 5063
rect 3342 5035 3366 5059
rect 3551 5040 3575 5064
rect 3766 5039 3786 5059
rect 1434 4737 1454 4757
rect 1645 4732 1669 4756
rect 1854 4737 1878 4761
rect 2068 4733 2094 4759
rect 4194 4710 4220 4736
rect 4410 4708 4434 4732
rect 4619 4713 4643 4737
rect 4834 4712 4854 4732
rect 372 4498 392 4518
rect 583 4493 607 4517
rect 792 4498 816 4522
rect 1006 4494 1032 4520
rect 3181 4476 3207 4502
rect 3397 4474 3421 4498
rect 3606 4479 3630 4503
rect 3821 4478 3841 4498
rect 1384 4317 1404 4337
rect 1595 4312 1619 4336
rect 1804 4317 1828 4341
rect 2018 4313 2044 4339
rect 4193 4295 4219 4321
rect 4409 4293 4433 4317
rect 4618 4298 4642 4322
rect 4833 4297 4853 4317
rect 371 4083 391 4103
rect 582 4078 606 4102
rect 791 4083 815 4107
rect 1005 4079 1031 4105
rect 2886 4044 2912 4070
rect 3102 4042 3126 4066
rect 3311 4047 3335 4071
rect 3526 4046 3546 4066
rect 1682 3773 1702 3793
rect 1893 3768 1917 3792
rect 2102 3773 2126 3797
rect 2316 3769 2342 3795
rect 4197 3734 4223 3760
rect 4413 3732 4437 3756
rect 4622 3737 4646 3761
rect 4837 3736 4857 3756
rect 375 3522 395 3542
rect 586 3517 610 3541
rect 795 3522 819 3546
rect 1009 3518 1035 3544
rect 3184 3500 3210 3526
rect 3400 3498 3424 3522
rect 3609 3503 3633 3527
rect 3824 3502 3844 3522
rect 1387 3341 1407 3361
rect 1598 3336 1622 3360
rect 1807 3341 1831 3365
rect 2021 3337 2047 3363
rect 4196 3319 4222 3345
rect 4412 3317 4436 3341
rect 4621 3322 4645 3346
rect 4836 3321 4856 3341
rect 374 3107 394 3127
rect 585 3102 609 3126
rect 794 3107 818 3131
rect 1008 3103 1034 3129
rect 3134 3080 3160 3106
rect 3350 3078 3374 3102
rect 3559 3083 3583 3107
rect 3774 3082 3794 3102
rect 1442 2780 1462 2800
rect 1653 2775 1677 2799
rect 1862 2780 1886 2804
rect 2076 2776 2102 2802
rect 4202 2753 4228 2779
rect 4418 2751 4442 2775
rect 4627 2756 4651 2780
rect 4842 2755 4862 2775
rect 380 2541 400 2561
rect 591 2536 615 2560
rect 800 2541 824 2565
rect 1014 2537 1040 2563
rect 3189 2519 3215 2545
rect 3405 2517 3429 2541
rect 3614 2522 3638 2546
rect 3829 2521 3849 2541
rect 1392 2360 1412 2380
rect 1603 2355 1627 2379
rect 1812 2360 1836 2384
rect 2026 2356 2052 2382
rect 4201 2338 4227 2364
rect 4417 2336 4441 2360
rect 4626 2341 4650 2365
rect 4841 2340 4861 2360
rect 379 2126 399 2146
rect 590 2121 614 2145
rect 799 2126 823 2150
rect 1013 2122 1039 2148
rect 2981 2052 3007 2078
rect 3197 2050 3221 2074
rect 3406 2055 3430 2079
rect 3621 2054 3641 2074
rect 1607 1848 1627 1868
rect 1818 1843 1842 1867
rect 2027 1848 2051 1872
rect 2241 1844 2267 1870
rect 4209 1774 4235 1800
rect 4425 1772 4449 1796
rect 4634 1777 4658 1801
rect 4849 1776 4869 1796
rect 387 1562 407 1582
rect 598 1557 622 1581
rect 807 1562 831 1586
rect 1021 1558 1047 1584
rect 3196 1540 3222 1566
rect 3412 1538 3436 1562
rect 3621 1543 3645 1567
rect 3836 1542 3856 1562
rect 1399 1381 1419 1401
rect 1610 1376 1634 1400
rect 1819 1381 1843 1405
rect 2033 1377 2059 1403
rect 4208 1359 4234 1385
rect 4424 1357 4448 1381
rect 4633 1362 4657 1386
rect 4848 1361 4868 1381
rect 386 1147 406 1167
rect 597 1142 621 1166
rect 806 1147 830 1171
rect 1020 1143 1046 1169
rect 3146 1120 3172 1146
rect 3362 1118 3386 1142
rect 3571 1123 3595 1147
rect 3786 1122 3806 1142
rect 1454 820 1474 840
rect 1665 815 1689 839
rect 1874 820 1898 844
rect 2088 816 2114 842
rect 4214 793 4240 819
rect 4430 791 4454 815
rect 4639 796 4663 820
rect 4854 795 4874 815
rect 392 581 412 601
rect 603 576 627 600
rect 812 581 836 605
rect 1026 577 1052 603
rect 3201 559 3227 585
rect 3417 557 3441 581
rect 3626 562 3650 586
rect 3841 561 3861 581
rect 1404 400 1424 420
rect 1615 395 1639 419
rect 1824 400 1848 424
rect 2038 396 2064 422
rect 4213 378 4239 404
rect 4429 376 4453 400
rect 4638 381 4662 405
rect 4853 380 4873 400
rect 391 166 411 186
rect 602 161 626 185
rect 811 166 835 190
rect 1025 162 1051 188
rect 1794 -315 1814 -295
rect 2005 -320 2029 -296
rect 2214 -315 2238 -291
rect 2428 -319 2454 -293
<< ndiffres >>
rect 97 7782 154 7801
rect 97 7779 118 7782
rect 3 7764 118 7779
rect 136 7764 154 7782
rect 3 7741 154 7764
rect 3 7705 45 7741
rect 2 7704 102 7705
rect 2 7683 158 7704
rect 5028 7733 5089 7749
rect 5028 7729 5184 7733
rect 5028 7711 5048 7729
rect 5066 7711 5184 7729
rect 2 7665 120 7683
rect 138 7665 158 7683
rect 2 7661 158 7665
rect 97 7645 158 7661
rect 5028 7690 5184 7711
rect 5084 7689 5184 7690
rect 5141 7653 5183 7689
rect 5032 7630 5183 7653
rect 95 7568 152 7587
rect 95 7565 116 7568
rect 1 7550 116 7565
rect 134 7550 152 7568
rect 1 7527 152 7550
rect 1 7491 43 7527
rect 0 7490 100 7491
rect 0 7469 156 7490
rect 5032 7612 5050 7630
rect 5068 7615 5183 7630
rect 5068 7612 5089 7615
rect 5032 7593 5089 7612
rect 5035 7532 5096 7548
rect 5035 7528 5191 7532
rect 5035 7510 5055 7528
rect 5073 7510 5191 7528
rect 0 7451 118 7469
rect 136 7451 156 7469
rect 0 7447 156 7451
rect 95 7431 156 7447
rect 5035 7489 5191 7510
rect 5091 7488 5191 7489
rect 5148 7452 5190 7488
rect 5039 7429 5190 7452
rect 5039 7411 5057 7429
rect 5075 7414 5190 7429
rect 5075 7411 5096 7414
rect 5039 7392 5096 7411
rect 95 7286 152 7305
rect 95 7283 116 7286
rect 1 7268 116 7283
rect 134 7268 152 7286
rect 1 7245 152 7268
rect 1 7209 43 7245
rect 0 7208 100 7209
rect 0 7187 156 7208
rect 5035 7250 5096 7266
rect 5035 7246 5191 7250
rect 5035 7228 5055 7246
rect 5073 7228 5191 7246
rect 0 7169 118 7187
rect 136 7169 156 7187
rect 0 7165 156 7169
rect 95 7149 156 7165
rect 102 7085 159 7104
rect 102 7082 123 7085
rect 8 7067 123 7082
rect 141 7067 159 7085
rect 5035 7207 5191 7228
rect 5091 7206 5191 7207
rect 5148 7170 5190 7206
rect 5039 7147 5190 7170
rect 5039 7129 5057 7147
rect 5075 7132 5190 7147
rect 5075 7129 5096 7132
rect 5039 7110 5096 7129
rect 8 7044 159 7067
rect 8 7008 50 7044
rect 7 7007 107 7008
rect 7 6986 163 7007
rect 7 6968 125 6986
rect 143 6968 163 6986
rect 7 6964 163 6968
rect 102 6948 163 6964
rect 5033 7036 5094 7052
rect 5033 7032 5189 7036
rect 5033 7014 5053 7032
rect 5071 7014 5189 7032
rect 5033 6993 5189 7014
rect 5089 6992 5189 6993
rect 5146 6956 5188 6992
rect 5037 6933 5188 6956
rect 5037 6915 5055 6933
rect 5073 6918 5188 6933
rect 5073 6915 5094 6918
rect 5037 6896 5094 6915
rect 102 6801 159 6820
rect 102 6798 123 6801
rect 8 6783 123 6798
rect 141 6783 159 6801
rect 8 6760 159 6783
rect 8 6724 50 6760
rect 7 6723 107 6724
rect 7 6702 163 6723
rect 7 6684 125 6702
rect 143 6684 163 6702
rect 7 6680 163 6684
rect 102 6664 163 6680
rect 5033 6752 5094 6768
rect 5033 6748 5189 6752
rect 5033 6730 5053 6748
rect 5071 6730 5189 6748
rect 5033 6709 5189 6730
rect 5089 6708 5189 6709
rect 5146 6672 5188 6708
rect 5037 6649 5188 6672
rect 100 6587 157 6606
rect 100 6584 121 6587
rect 6 6569 121 6584
rect 139 6569 157 6587
rect 6 6546 157 6569
rect 6 6510 48 6546
rect 5 6509 105 6510
rect 5 6488 161 6509
rect 5037 6631 5055 6649
rect 5073 6634 5188 6649
rect 5073 6631 5094 6634
rect 5037 6612 5094 6631
rect 5040 6551 5101 6567
rect 5040 6547 5196 6551
rect 5040 6529 5060 6547
rect 5078 6529 5196 6547
rect 5 6470 123 6488
rect 141 6470 161 6488
rect 5 6466 161 6470
rect 100 6450 161 6466
rect 5040 6508 5196 6529
rect 5096 6507 5196 6508
rect 5153 6471 5195 6507
rect 5044 6448 5195 6471
rect 5044 6430 5062 6448
rect 5080 6433 5195 6448
rect 5080 6430 5101 6433
rect 5044 6411 5101 6430
rect 100 6305 157 6324
rect 100 6302 121 6305
rect 6 6287 121 6302
rect 139 6287 157 6305
rect 6 6264 157 6287
rect 6 6228 48 6264
rect 5 6227 105 6228
rect 5 6206 161 6227
rect 5040 6269 5101 6285
rect 5040 6265 5196 6269
rect 5040 6247 5060 6265
rect 5078 6247 5196 6265
rect 5 6188 123 6206
rect 141 6188 161 6206
rect 5 6184 161 6188
rect 100 6168 161 6184
rect 107 6104 164 6123
rect 107 6101 128 6104
rect 13 6086 128 6101
rect 146 6086 164 6104
rect 5040 6226 5196 6247
rect 5096 6225 5196 6226
rect 5153 6189 5195 6225
rect 5044 6166 5195 6189
rect 5044 6148 5062 6166
rect 5080 6151 5195 6166
rect 5080 6148 5101 6151
rect 5044 6129 5101 6148
rect 13 6063 164 6086
rect 13 6027 55 6063
rect 12 6026 112 6027
rect 12 6005 168 6026
rect 5038 6055 5099 6071
rect 5038 6051 5194 6055
rect 5038 6033 5058 6051
rect 5076 6033 5194 6051
rect 12 5987 130 6005
rect 148 5987 168 6005
rect 12 5983 168 5987
rect 107 5967 168 5983
rect 5038 6012 5194 6033
rect 5094 6011 5194 6012
rect 5151 5975 5193 6011
rect 5042 5952 5193 5975
rect 109 5822 166 5841
rect 109 5819 130 5822
rect 15 5804 130 5819
rect 148 5804 166 5822
rect 5042 5934 5060 5952
rect 5078 5937 5193 5952
rect 5078 5934 5099 5937
rect 5042 5915 5099 5934
rect 15 5781 166 5804
rect 15 5745 57 5781
rect 14 5744 114 5745
rect 14 5723 170 5744
rect 5040 5773 5101 5789
rect 5040 5769 5196 5773
rect 5040 5751 5060 5769
rect 5078 5751 5196 5769
rect 14 5705 132 5723
rect 150 5705 170 5723
rect 14 5701 170 5705
rect 109 5685 170 5701
rect 5040 5730 5196 5751
rect 5096 5729 5196 5730
rect 5153 5693 5195 5729
rect 5044 5670 5195 5693
rect 107 5608 164 5627
rect 107 5605 128 5608
rect 13 5590 128 5605
rect 146 5590 164 5608
rect 13 5567 164 5590
rect 13 5531 55 5567
rect 12 5530 112 5531
rect 12 5509 168 5530
rect 5044 5652 5062 5670
rect 5080 5655 5195 5670
rect 5080 5652 5101 5655
rect 5044 5633 5101 5652
rect 5047 5572 5108 5588
rect 5047 5568 5203 5572
rect 5047 5550 5067 5568
rect 5085 5550 5203 5568
rect 12 5491 130 5509
rect 148 5491 168 5509
rect 12 5487 168 5491
rect 107 5471 168 5487
rect 5047 5529 5203 5550
rect 5103 5528 5203 5529
rect 5160 5492 5202 5528
rect 5051 5469 5202 5492
rect 5051 5451 5069 5469
rect 5087 5454 5202 5469
rect 5087 5451 5108 5454
rect 5051 5432 5108 5451
rect 107 5326 164 5345
rect 107 5323 128 5326
rect 13 5308 128 5323
rect 146 5308 164 5326
rect 13 5285 164 5308
rect 13 5249 55 5285
rect 12 5248 112 5249
rect 12 5227 168 5248
rect 5047 5290 5108 5306
rect 5047 5286 5203 5290
rect 5047 5268 5067 5286
rect 5085 5268 5203 5286
rect 12 5209 130 5227
rect 148 5209 168 5227
rect 12 5205 168 5209
rect 107 5189 168 5205
rect 114 5125 171 5144
rect 114 5122 135 5125
rect 20 5107 135 5122
rect 153 5107 171 5125
rect 5047 5247 5203 5268
rect 5103 5246 5203 5247
rect 5160 5210 5202 5246
rect 5051 5187 5202 5210
rect 5051 5169 5069 5187
rect 5087 5172 5202 5187
rect 5087 5169 5108 5172
rect 5051 5150 5108 5169
rect 20 5084 171 5107
rect 20 5048 62 5084
rect 19 5047 119 5048
rect 19 5026 175 5047
rect 19 5008 137 5026
rect 155 5008 175 5026
rect 19 5004 175 5008
rect 114 4988 175 5004
rect 5045 5076 5106 5092
rect 5045 5072 5201 5076
rect 5045 5054 5065 5072
rect 5083 5054 5201 5072
rect 5045 5033 5201 5054
rect 5101 5032 5201 5033
rect 5158 4996 5200 5032
rect 5049 4973 5200 4996
rect 5049 4955 5067 4973
rect 5085 4958 5200 4973
rect 5085 4955 5106 4958
rect 5049 4936 5106 4955
rect 114 4841 171 4860
rect 114 4838 135 4841
rect 20 4823 135 4838
rect 153 4823 171 4841
rect 20 4800 171 4823
rect 20 4764 62 4800
rect 19 4763 119 4764
rect 19 4742 175 4763
rect 19 4724 137 4742
rect 155 4724 175 4742
rect 19 4720 175 4724
rect 114 4704 175 4720
rect 5045 4792 5106 4808
rect 5045 4788 5201 4792
rect 5045 4770 5065 4788
rect 5083 4770 5201 4788
rect 5045 4749 5201 4770
rect 5101 4748 5201 4749
rect 5158 4712 5200 4748
rect 5049 4689 5200 4712
rect 112 4627 169 4646
rect 112 4624 133 4627
rect 18 4609 133 4624
rect 151 4609 169 4627
rect 18 4586 169 4609
rect 18 4550 60 4586
rect 17 4549 117 4550
rect 17 4528 173 4549
rect 5049 4671 5067 4689
rect 5085 4674 5200 4689
rect 5085 4671 5106 4674
rect 5049 4652 5106 4671
rect 5052 4591 5113 4607
rect 5052 4587 5208 4591
rect 5052 4569 5072 4587
rect 5090 4569 5208 4587
rect 17 4510 135 4528
rect 153 4510 173 4528
rect 17 4506 173 4510
rect 112 4490 173 4506
rect 5052 4548 5208 4569
rect 5108 4547 5208 4548
rect 5165 4511 5207 4547
rect 5056 4488 5207 4511
rect 5056 4470 5074 4488
rect 5092 4473 5207 4488
rect 5092 4470 5113 4473
rect 5056 4451 5113 4470
rect 112 4345 169 4364
rect 112 4342 133 4345
rect 18 4327 133 4342
rect 151 4327 169 4345
rect 18 4304 169 4327
rect 18 4268 60 4304
rect 17 4267 117 4268
rect 17 4246 173 4267
rect 5052 4309 5113 4325
rect 5052 4305 5208 4309
rect 5052 4287 5072 4305
rect 5090 4287 5208 4305
rect 17 4228 135 4246
rect 153 4228 173 4246
rect 17 4224 173 4228
rect 112 4208 173 4224
rect 119 4144 176 4163
rect 119 4141 140 4144
rect 25 4126 140 4141
rect 158 4126 176 4144
rect 5052 4266 5208 4287
rect 5108 4265 5208 4266
rect 5165 4229 5207 4265
rect 5056 4206 5207 4229
rect 5056 4188 5074 4206
rect 5092 4191 5207 4206
rect 5092 4188 5113 4191
rect 5056 4169 5113 4188
rect 25 4103 176 4126
rect 25 4067 67 4103
rect 24 4066 124 4067
rect 24 4045 180 4066
rect 5050 4095 5111 4111
rect 24 4027 142 4045
rect 160 4027 180 4045
rect 24 4023 180 4027
rect 119 4007 180 4023
rect 5050 4091 5206 4095
rect 5050 4073 5070 4091
rect 5088 4073 5206 4091
rect 5050 4052 5206 4073
rect 5106 4051 5206 4052
rect 117 3865 174 3884
rect 117 3862 138 3865
rect 23 3847 138 3862
rect 156 3847 174 3865
rect 23 3824 174 3847
rect 23 3788 65 3824
rect 5163 4015 5205 4051
rect 5054 3992 5205 4015
rect 5054 3974 5072 3992
rect 5090 3977 5205 3992
rect 5090 3974 5111 3977
rect 5054 3955 5111 3974
rect 22 3787 122 3788
rect 22 3766 178 3787
rect 22 3748 140 3766
rect 158 3748 178 3766
rect 22 3744 178 3748
rect 5048 3816 5109 3832
rect 5048 3812 5204 3816
rect 5048 3794 5068 3812
rect 5086 3794 5204 3812
rect 117 3728 178 3744
rect 5048 3773 5204 3794
rect 5104 3772 5204 3773
rect 5161 3736 5203 3772
rect 5052 3713 5203 3736
rect 115 3651 172 3670
rect 115 3648 136 3651
rect 21 3633 136 3648
rect 154 3633 172 3651
rect 21 3610 172 3633
rect 21 3574 63 3610
rect 20 3573 120 3574
rect 20 3552 176 3573
rect 5052 3695 5070 3713
rect 5088 3698 5203 3713
rect 5088 3695 5109 3698
rect 5052 3676 5109 3695
rect 5055 3615 5116 3631
rect 5055 3611 5211 3615
rect 5055 3593 5075 3611
rect 5093 3593 5211 3611
rect 20 3534 138 3552
rect 156 3534 176 3552
rect 20 3530 176 3534
rect 115 3514 176 3530
rect 5055 3572 5211 3593
rect 5111 3571 5211 3572
rect 5168 3535 5210 3571
rect 5059 3512 5210 3535
rect 5059 3494 5077 3512
rect 5095 3497 5210 3512
rect 5095 3494 5116 3497
rect 5059 3475 5116 3494
rect 115 3369 172 3388
rect 115 3366 136 3369
rect 21 3351 136 3366
rect 154 3351 172 3369
rect 21 3328 172 3351
rect 21 3292 63 3328
rect 20 3291 120 3292
rect 20 3270 176 3291
rect 5055 3333 5116 3349
rect 5055 3329 5211 3333
rect 5055 3311 5075 3329
rect 5093 3311 5211 3329
rect 20 3252 138 3270
rect 156 3252 176 3270
rect 20 3248 176 3252
rect 115 3232 176 3248
rect 122 3168 179 3187
rect 122 3165 143 3168
rect 28 3150 143 3165
rect 161 3150 179 3168
rect 5055 3290 5211 3311
rect 5111 3289 5211 3290
rect 5168 3253 5210 3289
rect 5059 3230 5210 3253
rect 5059 3212 5077 3230
rect 5095 3215 5210 3230
rect 5095 3212 5116 3215
rect 5059 3193 5116 3212
rect 28 3127 179 3150
rect 28 3091 70 3127
rect 27 3090 127 3091
rect 27 3069 183 3090
rect 27 3051 145 3069
rect 163 3051 183 3069
rect 27 3047 183 3051
rect 122 3031 183 3047
rect 5053 3119 5114 3135
rect 5053 3115 5209 3119
rect 5053 3097 5073 3115
rect 5091 3097 5209 3115
rect 5053 3076 5209 3097
rect 5109 3075 5209 3076
rect 5166 3039 5208 3075
rect 5057 3016 5208 3039
rect 5057 2998 5075 3016
rect 5093 3001 5208 3016
rect 5093 2998 5114 3001
rect 5057 2979 5114 2998
rect 122 2884 179 2903
rect 122 2881 143 2884
rect 28 2866 143 2881
rect 161 2866 179 2884
rect 28 2843 179 2866
rect 28 2807 70 2843
rect 27 2806 127 2807
rect 27 2785 183 2806
rect 27 2767 145 2785
rect 163 2767 183 2785
rect 27 2763 183 2767
rect 122 2747 183 2763
rect 5053 2835 5114 2851
rect 5053 2831 5209 2835
rect 5053 2813 5073 2831
rect 5091 2813 5209 2831
rect 5053 2792 5209 2813
rect 5109 2791 5209 2792
rect 5166 2755 5208 2791
rect 5057 2732 5208 2755
rect 120 2670 177 2689
rect 120 2667 141 2670
rect 26 2652 141 2667
rect 159 2652 177 2670
rect 26 2629 177 2652
rect 26 2593 68 2629
rect 25 2592 125 2593
rect 25 2571 181 2592
rect 5057 2714 5075 2732
rect 5093 2717 5208 2732
rect 5093 2714 5114 2717
rect 5057 2695 5114 2714
rect 5060 2634 5121 2650
rect 5060 2630 5216 2634
rect 5060 2612 5080 2630
rect 5098 2612 5216 2630
rect 25 2553 143 2571
rect 161 2553 181 2571
rect 25 2549 181 2553
rect 120 2533 181 2549
rect 5060 2591 5216 2612
rect 5116 2590 5216 2591
rect 5173 2554 5215 2590
rect 5064 2531 5215 2554
rect 5064 2513 5082 2531
rect 5100 2516 5215 2531
rect 5100 2513 5121 2516
rect 5064 2494 5121 2513
rect 120 2388 177 2407
rect 120 2385 141 2388
rect 26 2370 141 2385
rect 159 2370 177 2388
rect 26 2347 177 2370
rect 26 2311 68 2347
rect 25 2310 125 2311
rect 25 2289 181 2310
rect 5060 2352 5121 2368
rect 5060 2348 5216 2352
rect 5060 2330 5080 2348
rect 5098 2330 5216 2348
rect 25 2271 143 2289
rect 161 2271 181 2289
rect 25 2267 181 2271
rect 120 2251 181 2267
rect 127 2187 184 2206
rect 127 2184 148 2187
rect 33 2169 148 2184
rect 166 2169 184 2187
rect 5060 2309 5216 2330
rect 5116 2308 5216 2309
rect 5173 2272 5215 2308
rect 5064 2249 5215 2272
rect 5064 2231 5082 2249
rect 5100 2234 5215 2249
rect 5100 2231 5121 2234
rect 5064 2212 5121 2231
rect 33 2146 184 2169
rect 33 2110 75 2146
rect 32 2109 132 2110
rect 32 2088 188 2109
rect 5058 2138 5119 2154
rect 5058 2134 5214 2138
rect 5058 2116 5078 2134
rect 5096 2116 5214 2134
rect 32 2070 150 2088
rect 168 2070 188 2088
rect 32 2066 188 2070
rect 127 2050 188 2066
rect 5058 2095 5214 2116
rect 5114 2094 5214 2095
rect 5171 2058 5213 2094
rect 5062 2035 5213 2058
rect 129 1905 186 1924
rect 129 1902 150 1905
rect 35 1887 150 1902
rect 168 1887 186 1905
rect 5062 2017 5080 2035
rect 5098 2020 5213 2035
rect 5098 2017 5119 2020
rect 5062 1998 5119 2017
rect 35 1864 186 1887
rect 35 1828 77 1864
rect 34 1827 134 1828
rect 34 1806 190 1827
rect 5060 1856 5121 1872
rect 5060 1852 5216 1856
rect 5060 1834 5080 1852
rect 5098 1834 5216 1852
rect 34 1788 152 1806
rect 170 1788 190 1806
rect 34 1784 190 1788
rect 129 1768 190 1784
rect 5060 1813 5216 1834
rect 5116 1812 5216 1813
rect 5173 1776 5215 1812
rect 5064 1753 5215 1776
rect 127 1691 184 1710
rect 127 1688 148 1691
rect 33 1673 148 1688
rect 166 1673 184 1691
rect 33 1650 184 1673
rect 33 1614 75 1650
rect 32 1613 132 1614
rect 32 1592 188 1613
rect 5064 1735 5082 1753
rect 5100 1738 5215 1753
rect 5100 1735 5121 1738
rect 5064 1716 5121 1735
rect 5067 1655 5128 1671
rect 5067 1651 5223 1655
rect 5067 1633 5087 1651
rect 5105 1633 5223 1651
rect 32 1574 150 1592
rect 168 1574 188 1592
rect 32 1570 188 1574
rect 127 1554 188 1570
rect 5067 1612 5223 1633
rect 5123 1611 5223 1612
rect 5180 1575 5222 1611
rect 5071 1552 5222 1575
rect 5071 1534 5089 1552
rect 5107 1537 5222 1552
rect 5107 1534 5128 1537
rect 5071 1515 5128 1534
rect 127 1409 184 1428
rect 127 1406 148 1409
rect 33 1391 148 1406
rect 166 1391 184 1409
rect 33 1368 184 1391
rect 33 1332 75 1368
rect 32 1331 132 1332
rect 32 1310 188 1331
rect 5067 1373 5128 1389
rect 5067 1369 5223 1373
rect 5067 1351 5087 1369
rect 5105 1351 5223 1369
rect 32 1292 150 1310
rect 168 1292 188 1310
rect 32 1288 188 1292
rect 127 1272 188 1288
rect 134 1208 191 1227
rect 134 1205 155 1208
rect 40 1190 155 1205
rect 173 1190 191 1208
rect 5067 1330 5223 1351
rect 5123 1329 5223 1330
rect 5180 1293 5222 1329
rect 5071 1270 5222 1293
rect 5071 1252 5089 1270
rect 5107 1255 5222 1270
rect 5107 1252 5128 1255
rect 5071 1233 5128 1252
rect 40 1167 191 1190
rect 40 1131 82 1167
rect 39 1130 139 1131
rect 39 1109 195 1130
rect 39 1091 157 1109
rect 175 1091 195 1109
rect 39 1087 195 1091
rect 134 1071 195 1087
rect 5065 1159 5126 1175
rect 5065 1155 5221 1159
rect 5065 1137 5085 1155
rect 5103 1137 5221 1155
rect 5065 1116 5221 1137
rect 5121 1115 5221 1116
rect 5178 1079 5220 1115
rect 5069 1056 5220 1079
rect 5069 1038 5087 1056
rect 5105 1041 5220 1056
rect 5105 1038 5126 1041
rect 5069 1019 5126 1038
rect 134 924 191 943
rect 134 921 155 924
rect 40 906 155 921
rect 173 906 191 924
rect 40 883 191 906
rect 40 847 82 883
rect 39 846 139 847
rect 39 825 195 846
rect 39 807 157 825
rect 175 807 195 825
rect 39 803 195 807
rect 134 787 195 803
rect 5065 875 5126 891
rect 5065 871 5221 875
rect 5065 853 5085 871
rect 5103 853 5221 871
rect 5065 832 5221 853
rect 5121 831 5221 832
rect 5178 795 5220 831
rect 5069 772 5220 795
rect 132 710 189 729
rect 132 707 153 710
rect 38 692 153 707
rect 171 692 189 710
rect 38 669 189 692
rect 38 633 80 669
rect 37 632 137 633
rect 37 611 193 632
rect 5069 754 5087 772
rect 5105 757 5220 772
rect 5105 754 5126 757
rect 5069 735 5126 754
rect 5072 674 5133 690
rect 5072 670 5228 674
rect 5072 652 5092 670
rect 5110 652 5228 670
rect 37 593 155 611
rect 173 593 193 611
rect 37 589 193 593
rect 132 573 193 589
rect 5072 631 5228 652
rect 5128 630 5228 631
rect 5185 594 5227 630
rect 5076 571 5227 594
rect 5076 553 5094 571
rect 5112 556 5227 571
rect 5112 553 5133 556
rect 5076 534 5133 553
rect 132 428 189 447
rect 132 425 153 428
rect 38 410 153 425
rect 171 410 189 428
rect 38 387 189 410
rect 38 351 80 387
rect 37 350 137 351
rect 37 329 193 350
rect 5072 392 5133 408
rect 5072 388 5228 392
rect 5072 370 5092 388
rect 5110 370 5228 388
rect 37 311 155 329
rect 173 311 193 329
rect 37 307 193 311
rect 132 291 193 307
rect 139 227 196 246
rect 139 224 160 227
rect 45 209 160 224
rect 178 209 196 227
rect 5072 349 5228 370
rect 5128 348 5228 349
rect 5185 312 5227 348
rect 5076 289 5227 312
rect 5076 271 5094 289
rect 5112 274 5227 289
rect 5112 271 5133 274
rect 5076 252 5133 271
rect 45 186 196 209
rect 45 150 87 186
rect 44 149 144 150
rect 44 128 200 149
rect 5070 178 5131 194
rect 5070 174 5226 178
rect 5070 156 5090 174
rect 5108 156 5226 174
rect 44 110 162 128
rect 180 110 200 128
rect 44 106 200 110
rect 139 90 200 106
rect 5070 135 5226 156
rect 5126 134 5226 135
rect 5183 98 5225 134
rect 5074 75 5225 98
rect 5074 57 5092 75
rect 5110 60 5225 75
rect 5110 57 5131 60
rect 5074 38 5131 57
<< locali >>
rect 110 7791 145 7839
rect 5038 7833 5076 7839
rect 4449 7815 5076 7833
rect 108 7782 145 7791
rect 108 7764 118 7782
rect 136 7764 145 7782
rect 108 7754 145 7764
rect 4031 7798 4199 7799
rect 4450 7798 4474 7815
rect 4031 7772 4475 7798
rect 4031 7770 4199 7772
rect 111 7690 148 7692
rect 111 7689 759 7690
rect 110 7683 759 7689
rect 110 7665 120 7683
rect 138 7669 759 7683
rect 138 7665 148 7669
rect 589 7668 759 7669
rect 110 7655 148 7665
rect 110 7577 145 7655
rect 722 7645 759 7668
rect 106 7568 145 7577
rect 106 7550 116 7568
rect 134 7550 145 7568
rect 106 7544 145 7550
rect 301 7620 551 7644
rect 301 7549 338 7620
rect 453 7559 484 7560
rect 106 7540 143 7544
rect 301 7529 310 7549
rect 330 7529 338 7549
rect 301 7519 338 7529
rect 397 7549 484 7559
rect 397 7529 406 7549
rect 426 7529 484 7549
rect 397 7520 484 7529
rect 397 7519 434 7520
rect 109 7469 146 7478
rect 107 7451 118 7469
rect 136 7451 146 7469
rect 453 7467 484 7520
rect 514 7549 551 7620
rect 722 7625 1115 7645
rect 1135 7625 1138 7645
rect 722 7620 1138 7625
rect 722 7619 1063 7620
rect 666 7559 697 7560
rect 514 7529 523 7549
rect 543 7529 551 7549
rect 514 7519 551 7529
rect 610 7552 697 7559
rect 610 7549 671 7552
rect 610 7529 619 7549
rect 639 7532 671 7549
rect 692 7532 697 7552
rect 639 7529 697 7532
rect 610 7522 697 7529
rect 722 7549 759 7619
rect 1025 7618 1062 7619
rect 4031 7592 4058 7770
rect 4098 7732 4162 7744
rect 4438 7740 4475 7772
rect 4646 7771 4895 7793
rect 4646 7740 4683 7771
rect 4859 7769 4895 7771
rect 5038 7774 5076 7815
rect 4859 7740 4896 7769
rect 4098 7731 4133 7732
rect 4075 7726 4133 7731
rect 4075 7706 4078 7726
rect 4098 7712 4133 7726
rect 4153 7712 4162 7732
rect 4098 7704 4162 7712
rect 4124 7703 4162 7704
rect 4125 7702 4162 7703
rect 4228 7736 4264 7737
rect 4336 7736 4372 7737
rect 4228 7730 4372 7736
rect 4228 7728 4294 7730
rect 4228 7708 4236 7728
rect 4256 7709 4294 7728
rect 4316 7728 4372 7730
rect 4316 7709 4344 7728
rect 4256 7708 4344 7709
rect 4364 7708 4372 7728
rect 4228 7702 4372 7708
rect 4438 7732 4476 7740
rect 4544 7736 4580 7737
rect 4438 7712 4447 7732
rect 4467 7712 4476 7732
rect 4438 7703 4476 7712
rect 4495 7729 4580 7736
rect 4495 7709 4502 7729
rect 4523 7728 4580 7729
rect 4523 7709 4552 7728
rect 4495 7708 4552 7709
rect 4572 7708 4580 7728
rect 4438 7702 4475 7703
rect 4495 7702 4580 7708
rect 4646 7732 4684 7740
rect 4757 7736 4793 7737
rect 4646 7712 4655 7732
rect 4675 7712 4684 7732
rect 4646 7703 4684 7712
rect 4708 7728 4793 7736
rect 4708 7708 4765 7728
rect 4785 7708 4793 7728
rect 4646 7702 4683 7703
rect 4708 7702 4793 7708
rect 4859 7732 4897 7740
rect 4859 7712 4868 7732
rect 4888 7712 4897 7732
rect 4859 7703 4897 7712
rect 5038 7739 5074 7774
rect 5038 7729 5075 7739
rect 5038 7711 5048 7729
rect 5066 7711 5075 7729
rect 4859 7702 4896 7703
rect 5038 7702 5075 7711
rect 4282 7681 4318 7702
rect 4708 7681 4739 7702
rect 4115 7677 4215 7681
rect 4115 7673 4177 7677
rect 4115 7647 4122 7673
rect 4148 7651 4177 7673
rect 4203 7651 4215 7677
rect 4148 7647 4215 7651
rect 4115 7644 4215 7647
rect 4283 7644 4318 7681
rect 4380 7678 4739 7681
rect 4380 7673 4602 7678
rect 4380 7649 4393 7673
rect 4417 7654 4602 7673
rect 4626 7654 4739 7678
rect 4417 7649 4739 7654
rect 4380 7645 4739 7649
rect 4806 7673 4955 7681
rect 4806 7653 4817 7673
rect 4837 7653 4955 7673
rect 4806 7646 4955 7653
rect 4806 7645 4847 7646
rect 4130 7592 4167 7593
rect 4226 7592 4263 7593
rect 4282 7592 4318 7644
rect 4337 7592 4374 7593
rect 4030 7583 4168 7592
rect 2966 7565 2997 7568
rect 874 7559 910 7560
rect 722 7529 731 7549
rect 751 7529 759 7549
rect 610 7520 666 7522
rect 610 7519 647 7520
rect 722 7519 759 7529
rect 818 7549 966 7559
rect 1066 7556 1162 7558
rect 818 7529 827 7549
rect 847 7529 937 7549
rect 957 7529 966 7549
rect 818 7520 966 7529
rect 1024 7549 1162 7556
rect 1024 7529 1033 7549
rect 1053 7529 1162 7549
rect 1024 7520 1162 7529
rect 2966 7539 2973 7565
rect 2992 7539 2997 7565
rect 818 7519 855 7520
rect 874 7468 910 7520
rect 929 7519 966 7520
rect 1025 7519 1062 7520
rect 345 7466 386 7467
rect 107 7302 146 7451
rect 237 7459 386 7466
rect 237 7439 355 7459
rect 375 7439 386 7459
rect 237 7431 386 7439
rect 453 7463 812 7467
rect 453 7458 775 7463
rect 453 7434 566 7458
rect 590 7439 775 7458
rect 799 7439 812 7463
rect 590 7434 812 7439
rect 453 7431 812 7434
rect 874 7431 909 7468
rect 977 7465 1077 7468
rect 977 7461 1044 7465
rect 977 7435 989 7461
rect 1015 7439 1044 7461
rect 1070 7439 1077 7465
rect 1015 7435 1077 7439
rect 977 7431 1077 7435
rect 453 7410 484 7431
rect 874 7410 910 7431
rect 296 7409 333 7410
rect 295 7400 333 7409
rect 295 7380 304 7400
rect 324 7380 333 7400
rect 295 7372 333 7380
rect 399 7404 484 7410
rect 509 7409 546 7410
rect 399 7384 407 7404
rect 427 7384 484 7404
rect 399 7376 484 7384
rect 508 7400 546 7409
rect 508 7380 517 7400
rect 537 7380 546 7400
rect 399 7375 435 7376
rect 508 7372 546 7380
rect 612 7404 697 7410
rect 717 7409 754 7410
rect 612 7384 620 7404
rect 640 7403 697 7404
rect 640 7384 669 7403
rect 612 7383 669 7384
rect 690 7383 697 7403
rect 612 7376 697 7383
rect 716 7400 754 7409
rect 716 7380 725 7400
rect 745 7380 754 7400
rect 612 7375 648 7376
rect 716 7372 754 7380
rect 820 7405 964 7410
rect 820 7404 885 7405
rect 820 7384 828 7404
rect 848 7384 885 7404
rect 907 7404 964 7405
rect 907 7384 936 7404
rect 956 7384 964 7404
rect 820 7376 964 7384
rect 820 7375 856 7376
rect 928 7375 964 7376
rect 1030 7409 1067 7410
rect 1030 7408 1068 7409
rect 1030 7400 1094 7408
rect 1030 7380 1039 7400
rect 1059 7386 1094 7400
rect 1114 7386 1117 7406
rect 1059 7381 1117 7386
rect 1059 7380 1094 7381
rect 296 7343 333 7372
rect 297 7341 333 7343
rect 509 7341 546 7372
rect 297 7319 546 7341
rect 717 7340 754 7372
rect 1030 7368 1094 7380
rect 1134 7342 1161 7520
rect 993 7340 1161 7342
rect 717 7314 1161 7340
rect 1313 7439 1563 7463
rect 1313 7368 1350 7439
rect 1465 7378 1496 7379
rect 1313 7348 1322 7368
rect 1342 7348 1350 7368
rect 1313 7338 1350 7348
rect 1409 7368 1496 7378
rect 1409 7348 1418 7368
rect 1438 7348 1496 7368
rect 1409 7339 1496 7348
rect 1409 7338 1446 7339
rect 717 7304 739 7314
rect 993 7313 1161 7314
rect 677 7302 739 7304
rect 107 7295 739 7302
rect 106 7286 739 7295
rect 1465 7286 1496 7339
rect 1526 7368 1563 7439
rect 1734 7444 2127 7464
rect 2147 7444 2150 7464
rect 1734 7439 2150 7444
rect 1734 7438 2075 7439
rect 1678 7378 1709 7379
rect 1526 7348 1535 7368
rect 1555 7348 1563 7368
rect 1526 7338 1563 7348
rect 1622 7371 1709 7378
rect 1622 7368 1683 7371
rect 1622 7348 1631 7368
rect 1651 7351 1683 7368
rect 1704 7351 1709 7371
rect 1651 7348 1709 7351
rect 1622 7341 1709 7348
rect 1734 7368 1771 7438
rect 2037 7437 2074 7438
rect 1886 7378 1922 7379
rect 1734 7348 1743 7368
rect 1763 7348 1771 7368
rect 1622 7339 1678 7341
rect 1622 7338 1659 7339
rect 1734 7338 1771 7348
rect 1830 7368 1978 7378
rect 2078 7375 2174 7377
rect 1830 7348 1839 7368
rect 1859 7348 1949 7368
rect 1969 7348 1978 7368
rect 1830 7339 1978 7348
rect 2036 7368 2174 7375
rect 2036 7348 2045 7368
rect 2065 7348 2174 7368
rect 2036 7339 2174 7348
rect 1830 7338 1867 7339
rect 1886 7287 1922 7339
rect 1941 7338 1978 7339
rect 2037 7338 2074 7339
rect 106 7268 116 7286
rect 134 7285 739 7286
rect 1357 7285 1398 7286
rect 134 7280 155 7285
rect 134 7268 146 7280
rect 1249 7278 1398 7285
rect 106 7260 146 7268
rect 189 7267 215 7268
rect 106 7258 143 7260
rect 189 7249 743 7267
rect 1249 7258 1367 7278
rect 1387 7258 1398 7278
rect 1249 7250 1398 7258
rect 1465 7282 1824 7286
rect 1465 7277 1787 7282
rect 1465 7253 1578 7277
rect 1602 7258 1787 7277
rect 1811 7258 1824 7282
rect 1602 7253 1824 7258
rect 1465 7250 1824 7253
rect 1886 7250 1921 7287
rect 1989 7284 2089 7287
rect 1989 7280 2056 7284
rect 1989 7254 2001 7280
rect 2027 7258 2056 7280
rect 2082 7258 2089 7284
rect 2027 7254 2089 7258
rect 1989 7250 2089 7254
rect 109 7190 146 7196
rect 189 7190 215 7249
rect 722 7230 743 7249
rect 109 7187 215 7190
rect 109 7169 118 7187
rect 136 7173 215 7187
rect 300 7205 550 7229
rect 136 7171 212 7173
rect 136 7169 146 7171
rect 109 7159 146 7169
rect 114 7094 145 7159
rect 300 7134 337 7205
rect 452 7144 483 7145
rect 300 7114 309 7134
rect 329 7114 337 7134
rect 300 7104 337 7114
rect 396 7134 483 7144
rect 396 7114 405 7134
rect 425 7114 483 7134
rect 396 7105 483 7114
rect 396 7104 433 7105
rect 113 7085 150 7094
rect 113 7067 123 7085
rect 141 7067 150 7085
rect 113 7057 150 7067
rect 452 7052 483 7105
rect 513 7134 550 7205
rect 721 7210 1114 7230
rect 1134 7210 1137 7230
rect 1465 7229 1496 7250
rect 1886 7229 1922 7250
rect 1308 7228 1345 7229
rect 721 7205 1137 7210
rect 1307 7219 1345 7228
rect 721 7204 1062 7205
rect 665 7144 696 7145
rect 513 7114 522 7134
rect 542 7114 550 7134
rect 513 7104 550 7114
rect 609 7137 696 7144
rect 609 7134 670 7137
rect 609 7114 618 7134
rect 638 7117 670 7134
rect 691 7117 696 7137
rect 638 7114 696 7117
rect 609 7107 696 7114
rect 721 7134 758 7204
rect 1024 7203 1061 7204
rect 1307 7199 1316 7219
rect 1336 7199 1345 7219
rect 1307 7191 1345 7199
rect 1411 7223 1496 7229
rect 1521 7228 1558 7229
rect 1411 7203 1419 7223
rect 1439 7203 1496 7223
rect 1411 7195 1496 7203
rect 1520 7219 1558 7228
rect 1520 7199 1529 7219
rect 1549 7199 1558 7219
rect 1411 7194 1447 7195
rect 1520 7191 1558 7199
rect 1624 7223 1709 7229
rect 1729 7228 1766 7229
rect 1624 7203 1632 7223
rect 1652 7222 1709 7223
rect 1652 7203 1681 7222
rect 1624 7202 1681 7203
rect 1702 7202 1709 7222
rect 1624 7195 1709 7202
rect 1728 7219 1766 7228
rect 1728 7199 1737 7219
rect 1757 7199 1766 7219
rect 1624 7194 1660 7195
rect 1728 7191 1766 7199
rect 1832 7223 1976 7229
rect 1832 7203 1840 7223
rect 1860 7203 1892 7223
rect 1916 7203 1948 7223
rect 1968 7203 1976 7223
rect 1832 7195 1976 7203
rect 1832 7194 1868 7195
rect 1940 7194 1976 7195
rect 2042 7228 2079 7229
rect 2042 7227 2080 7228
rect 2042 7219 2106 7227
rect 2042 7199 2051 7219
rect 2071 7205 2106 7219
rect 2126 7205 2129 7225
rect 2071 7200 2129 7205
rect 2071 7199 2106 7200
rect 1308 7162 1345 7191
rect 1309 7160 1345 7162
rect 1521 7160 1558 7191
rect 873 7144 909 7145
rect 721 7114 730 7134
rect 750 7114 758 7134
rect 609 7105 665 7107
rect 609 7104 646 7105
rect 721 7104 758 7114
rect 817 7134 965 7144
rect 1065 7141 1161 7143
rect 817 7114 826 7134
rect 846 7114 936 7134
rect 956 7114 965 7134
rect 817 7105 965 7114
rect 1023 7134 1161 7141
rect 1309 7138 1558 7160
rect 1729 7159 1766 7191
rect 2042 7187 2106 7199
rect 2146 7161 2173 7339
rect 2005 7159 2173 7161
rect 1729 7155 2173 7159
rect 1023 7114 1032 7134
rect 1052 7114 1161 7134
rect 1729 7136 1778 7155
rect 1798 7136 2173 7155
rect 1729 7133 2173 7136
rect 2005 7132 2173 7133
rect 2873 7146 2902 7148
rect 2873 7141 2905 7146
rect 2873 7123 2880 7141
rect 2900 7123 2905 7141
rect 2966 7145 2997 7539
rect 3018 7564 3186 7565
rect 3018 7561 3462 7564
rect 3018 7542 3393 7561
rect 3413 7542 3462 7561
rect 4030 7563 4139 7583
rect 4159 7563 4168 7583
rect 3018 7538 3462 7542
rect 3018 7536 3186 7538
rect 3018 7358 3045 7536
rect 3085 7498 3149 7510
rect 3425 7506 3462 7538
rect 3633 7537 3882 7559
rect 4030 7556 4168 7563
rect 4226 7583 4374 7592
rect 4226 7563 4235 7583
rect 4255 7563 4345 7583
rect 4365 7563 4374 7583
rect 4030 7554 4126 7556
rect 4226 7553 4374 7563
rect 4433 7583 4470 7593
rect 4545 7592 4582 7593
rect 4526 7590 4582 7592
rect 4433 7563 4441 7583
rect 4461 7563 4470 7583
rect 4282 7552 4318 7553
rect 3633 7506 3670 7537
rect 3846 7535 3882 7537
rect 3846 7506 3883 7535
rect 3085 7497 3120 7498
rect 3062 7492 3120 7497
rect 3062 7472 3065 7492
rect 3085 7478 3120 7492
rect 3140 7478 3149 7498
rect 3085 7470 3149 7478
rect 3111 7469 3149 7470
rect 3112 7468 3149 7469
rect 3215 7502 3251 7503
rect 3323 7502 3359 7503
rect 3215 7494 3359 7502
rect 3215 7474 3223 7494
rect 3243 7493 3331 7494
rect 3243 7474 3276 7493
rect 3215 7473 3276 7474
rect 3300 7474 3331 7493
rect 3351 7474 3359 7494
rect 3300 7473 3359 7474
rect 3215 7468 3359 7473
rect 3425 7498 3463 7506
rect 3531 7502 3567 7503
rect 3425 7478 3434 7498
rect 3454 7478 3463 7498
rect 3425 7469 3463 7478
rect 3482 7495 3567 7502
rect 3482 7475 3489 7495
rect 3510 7494 3567 7495
rect 3510 7475 3539 7494
rect 3482 7474 3539 7475
rect 3559 7474 3567 7494
rect 3425 7468 3462 7469
rect 3482 7468 3567 7474
rect 3633 7498 3671 7506
rect 3744 7502 3780 7503
rect 3633 7478 3642 7498
rect 3662 7478 3671 7498
rect 3633 7469 3671 7478
rect 3695 7494 3780 7502
rect 3695 7474 3752 7494
rect 3772 7474 3780 7494
rect 3633 7468 3670 7469
rect 3695 7468 3780 7474
rect 3846 7498 3884 7506
rect 3846 7478 3855 7498
rect 3875 7478 3884 7498
rect 4130 7493 4167 7494
rect 4433 7493 4470 7563
rect 4495 7583 4582 7590
rect 4495 7580 4553 7583
rect 4495 7560 4500 7580
rect 4521 7563 4553 7580
rect 4573 7563 4582 7583
rect 4521 7560 4582 7563
rect 4495 7553 4582 7560
rect 4641 7583 4678 7593
rect 4641 7563 4649 7583
rect 4669 7563 4678 7583
rect 4495 7552 4526 7553
rect 4129 7492 4470 7493
rect 3846 7469 3884 7478
rect 4054 7487 4470 7492
rect 3846 7468 3883 7469
rect 3269 7447 3305 7468
rect 3695 7447 3726 7468
rect 4054 7467 4057 7487
rect 4077 7467 4470 7487
rect 4641 7492 4678 7563
rect 4708 7592 4739 7645
rect 5041 7630 5078 7640
rect 5041 7612 5050 7630
rect 5068 7612 5078 7630
rect 5041 7603 5078 7612
rect 4758 7592 4795 7593
rect 4708 7583 4795 7592
rect 4708 7563 4766 7583
rect 4786 7563 4795 7583
rect 4708 7553 4795 7563
rect 4854 7583 4891 7593
rect 4854 7563 4862 7583
rect 4882 7563 4891 7583
rect 4708 7552 4739 7553
rect 4854 7492 4891 7563
rect 5046 7538 5077 7603
rect 5045 7528 5082 7538
rect 5045 7526 5055 7528
rect 4979 7524 5055 7526
rect 4641 7468 4891 7492
rect 4976 7510 5055 7524
rect 5073 7510 5082 7528
rect 4976 7507 5082 7510
rect 4448 7448 4469 7467
rect 4976 7448 5002 7507
rect 5045 7501 5082 7507
rect 3102 7443 3202 7447
rect 3102 7439 3164 7443
rect 3102 7413 3109 7439
rect 3135 7417 3164 7439
rect 3190 7417 3202 7443
rect 3135 7413 3202 7417
rect 3102 7410 3202 7413
rect 3270 7410 3305 7447
rect 3367 7444 3726 7447
rect 3367 7439 3589 7444
rect 3367 7415 3380 7439
rect 3404 7420 3589 7439
rect 3613 7420 3726 7444
rect 3404 7415 3726 7420
rect 3367 7411 3726 7415
rect 3793 7439 3942 7447
rect 3793 7419 3804 7439
rect 3824 7419 3942 7439
rect 4448 7430 5002 7448
rect 5048 7437 5085 7439
rect 4976 7429 5002 7430
rect 5045 7429 5085 7437
rect 3793 7412 3942 7419
rect 5045 7417 5057 7429
rect 5036 7412 5057 7417
rect 3793 7411 3834 7412
rect 4452 7411 5057 7412
rect 5075 7411 5085 7429
rect 3117 7358 3154 7359
rect 3213 7358 3250 7359
rect 3269 7358 3305 7410
rect 3324 7358 3361 7359
rect 3017 7349 3155 7358
rect 3017 7329 3126 7349
rect 3146 7329 3155 7349
rect 3017 7322 3155 7329
rect 3213 7349 3361 7358
rect 3213 7329 3222 7349
rect 3242 7329 3332 7349
rect 3352 7329 3361 7349
rect 3017 7320 3113 7322
rect 3213 7319 3361 7329
rect 3420 7349 3457 7359
rect 3532 7358 3569 7359
rect 3513 7356 3569 7358
rect 3420 7329 3428 7349
rect 3448 7329 3457 7349
rect 3269 7318 3305 7319
rect 3117 7259 3154 7260
rect 3420 7259 3457 7329
rect 3482 7349 3569 7356
rect 3482 7346 3540 7349
rect 3482 7326 3487 7346
rect 3508 7329 3540 7346
rect 3560 7329 3569 7349
rect 3508 7326 3569 7329
rect 3482 7319 3569 7326
rect 3628 7349 3665 7359
rect 3628 7329 3636 7349
rect 3656 7329 3665 7349
rect 3482 7318 3513 7319
rect 3116 7258 3457 7259
rect 3041 7253 3457 7258
rect 3041 7233 3044 7253
rect 3064 7233 3457 7253
rect 3628 7258 3665 7329
rect 3695 7358 3726 7411
rect 4452 7402 5085 7411
rect 4452 7395 5084 7402
rect 4452 7393 4514 7395
rect 4030 7383 4198 7384
rect 4452 7383 4474 7393
rect 3745 7358 3782 7359
rect 3695 7349 3782 7358
rect 3695 7329 3753 7349
rect 3773 7329 3782 7349
rect 3695 7319 3782 7329
rect 3841 7349 3878 7359
rect 3841 7329 3849 7349
rect 3869 7329 3878 7349
rect 3695 7318 3726 7319
rect 3841 7258 3878 7329
rect 3628 7234 3878 7258
rect 4030 7357 4474 7383
rect 4030 7355 4198 7357
rect 4030 7177 4057 7355
rect 4097 7317 4161 7329
rect 4437 7325 4474 7357
rect 4645 7356 4894 7378
rect 4645 7325 4682 7356
rect 4858 7354 4894 7356
rect 4858 7325 4895 7354
rect 4097 7316 4132 7317
rect 4074 7311 4132 7316
rect 4074 7291 4077 7311
rect 4097 7297 4132 7311
rect 4152 7297 4161 7317
rect 4097 7289 4161 7297
rect 4123 7288 4161 7289
rect 4124 7287 4161 7288
rect 4227 7321 4263 7322
rect 4335 7321 4371 7322
rect 4227 7313 4371 7321
rect 4227 7293 4235 7313
rect 4255 7293 4284 7313
rect 4227 7292 4284 7293
rect 4306 7293 4343 7313
rect 4363 7293 4371 7313
rect 4306 7292 4371 7293
rect 4227 7287 4371 7292
rect 4437 7317 4475 7325
rect 4543 7321 4579 7322
rect 4437 7297 4446 7317
rect 4466 7297 4475 7317
rect 4437 7288 4475 7297
rect 4494 7314 4579 7321
rect 4494 7294 4501 7314
rect 4522 7313 4579 7314
rect 4522 7294 4551 7313
rect 4494 7293 4551 7294
rect 4571 7293 4579 7313
rect 4437 7287 4474 7288
rect 4494 7287 4579 7293
rect 4645 7317 4683 7325
rect 4756 7321 4792 7322
rect 4645 7297 4654 7317
rect 4674 7297 4683 7317
rect 4645 7288 4683 7297
rect 4707 7313 4792 7321
rect 4707 7293 4764 7313
rect 4784 7293 4792 7313
rect 4645 7287 4682 7288
rect 4707 7287 4792 7293
rect 4858 7317 4896 7325
rect 4858 7297 4867 7317
rect 4887 7297 4896 7317
rect 4858 7288 4896 7297
rect 4858 7287 4895 7288
rect 4281 7266 4317 7287
rect 4707 7266 4738 7287
rect 4114 7262 4214 7266
rect 4114 7258 4176 7262
rect 4114 7232 4121 7258
rect 4147 7236 4176 7258
rect 4202 7236 4214 7262
rect 4147 7232 4214 7236
rect 4114 7229 4214 7232
rect 4282 7229 4317 7266
rect 4379 7263 4738 7266
rect 4379 7258 4601 7263
rect 4379 7234 4392 7258
rect 4416 7239 4601 7258
rect 4625 7239 4738 7263
rect 4416 7234 4738 7239
rect 4379 7230 4738 7234
rect 4805 7258 4954 7266
rect 4805 7238 4816 7258
rect 4836 7238 4954 7258
rect 4805 7231 4954 7238
rect 5045 7246 5084 7395
rect 4805 7230 4846 7231
rect 4129 7177 4166 7178
rect 4225 7177 4262 7178
rect 4281 7177 4317 7229
rect 4336 7177 4373 7178
rect 4029 7168 4167 7177
rect 4029 7148 4138 7168
rect 4158 7148 4167 7168
rect 2966 7144 3136 7145
rect 2966 7129 3412 7144
rect 4029 7141 4167 7148
rect 4225 7168 4373 7177
rect 4225 7148 4234 7168
rect 4254 7148 4344 7168
rect 4364 7148 4373 7168
rect 4029 7139 4125 7141
rect 2873 7118 2905 7123
rect 1023 7105 1161 7114
rect 817 7104 854 7105
rect 873 7053 909 7105
rect 928 7104 965 7105
rect 1024 7104 1061 7105
rect 344 7051 385 7052
rect 236 7044 385 7051
rect 236 7024 354 7044
rect 374 7024 385 7044
rect 236 7016 385 7024
rect 452 7048 811 7052
rect 452 7043 774 7048
rect 452 7019 565 7043
rect 589 7024 774 7043
rect 798 7024 811 7048
rect 589 7019 811 7024
rect 452 7016 811 7019
rect 873 7016 908 7053
rect 976 7050 1076 7053
rect 976 7046 1043 7050
rect 976 7020 988 7046
rect 1014 7024 1043 7046
rect 1069 7024 1076 7050
rect 1014 7020 1076 7024
rect 976 7016 1076 7020
rect 452 6995 483 7016
rect 873 6995 909 7016
rect 116 6986 153 6995
rect 295 6994 332 6995
rect 116 6968 125 6986
rect 143 6968 153 6986
rect 116 6958 153 6968
rect 117 6923 153 6958
rect 294 6985 332 6994
rect 294 6965 303 6985
rect 323 6965 332 6985
rect 294 6957 332 6965
rect 398 6989 483 6995
rect 508 6994 545 6995
rect 398 6969 406 6989
rect 426 6969 483 6989
rect 398 6961 483 6969
rect 507 6985 545 6994
rect 507 6965 516 6985
rect 536 6965 545 6985
rect 398 6960 434 6961
rect 507 6957 545 6965
rect 611 6989 696 6995
rect 716 6994 753 6995
rect 611 6969 619 6989
rect 639 6988 696 6989
rect 639 6969 668 6988
rect 611 6968 668 6969
rect 689 6968 696 6988
rect 611 6961 696 6968
rect 715 6985 753 6994
rect 715 6965 724 6985
rect 744 6965 753 6985
rect 611 6960 647 6961
rect 715 6957 753 6965
rect 819 6989 963 6995
rect 819 6969 827 6989
rect 847 6988 935 6989
rect 847 6969 875 6988
rect 819 6967 875 6969
rect 897 6969 935 6988
rect 955 6969 963 6989
rect 897 6967 963 6969
rect 819 6961 963 6967
rect 819 6960 855 6961
rect 927 6960 963 6961
rect 1029 6994 1066 6995
rect 1029 6993 1067 6994
rect 1029 6985 1093 6993
rect 1029 6965 1038 6985
rect 1058 6971 1093 6985
rect 1113 6971 1116 6991
rect 1058 6966 1116 6971
rect 1058 6965 1093 6966
rect 295 6928 332 6957
rect 115 6882 153 6923
rect 296 6926 332 6928
rect 508 6926 545 6957
rect 296 6904 545 6926
rect 716 6925 753 6957
rect 1029 6953 1093 6965
rect 1133 6927 1160 7105
rect 992 6925 1160 6927
rect 716 6899 1160 6925
rect 717 6882 741 6899
rect 992 6898 1160 6899
rect 115 6864 742 6882
rect 1368 6878 1618 6902
rect 115 6858 153 6864
rect 115 6834 152 6858
rect 115 6810 150 6834
rect 113 6801 150 6810
rect 113 6783 123 6801
rect 141 6783 150 6801
rect 113 6773 150 6783
rect 1368 6807 1405 6878
rect 1520 6817 1551 6818
rect 1368 6787 1377 6807
rect 1397 6787 1405 6807
rect 1368 6777 1405 6787
rect 1464 6807 1551 6817
rect 1464 6787 1473 6807
rect 1493 6787 1551 6807
rect 1464 6778 1551 6787
rect 1464 6777 1501 6778
rect 1520 6725 1551 6778
rect 1581 6807 1618 6878
rect 1789 6883 2182 6903
rect 2202 6883 2205 6903
rect 1789 6878 2205 6883
rect 1789 6877 2130 6878
rect 1733 6817 1764 6818
rect 1581 6787 1590 6807
rect 1610 6787 1618 6807
rect 1581 6777 1618 6787
rect 1677 6810 1764 6817
rect 1677 6807 1738 6810
rect 1677 6787 1686 6807
rect 1706 6790 1738 6807
rect 1759 6790 1764 6810
rect 1706 6787 1764 6790
rect 1677 6780 1764 6787
rect 1789 6807 1826 6877
rect 2092 6876 2129 6877
rect 1941 6817 1977 6818
rect 1789 6787 1798 6807
rect 1818 6787 1826 6807
rect 1677 6778 1733 6780
rect 1677 6777 1714 6778
rect 1789 6777 1826 6787
rect 1885 6807 2033 6817
rect 2133 6814 2229 6816
rect 1885 6787 1894 6807
rect 1914 6787 2004 6807
rect 2024 6787 2033 6807
rect 1885 6778 2033 6787
rect 2091 6807 2229 6814
rect 2091 6787 2100 6807
rect 2120 6787 2229 6807
rect 2091 6778 2229 6787
rect 1885 6777 1922 6778
rect 1941 6726 1977 6778
rect 1996 6777 2033 6778
rect 2092 6777 2129 6778
rect 1412 6724 1453 6725
rect 1304 6717 1453 6724
rect 116 6709 153 6711
rect 116 6708 764 6709
rect 115 6702 764 6708
rect 115 6684 125 6702
rect 143 6688 764 6702
rect 1304 6697 1422 6717
rect 1442 6697 1453 6717
rect 1304 6689 1453 6697
rect 1520 6721 1879 6725
rect 1520 6716 1842 6721
rect 1520 6692 1633 6716
rect 1657 6697 1842 6716
rect 1866 6697 1879 6721
rect 1657 6692 1879 6697
rect 1520 6689 1879 6692
rect 1941 6689 1976 6726
rect 2044 6723 2144 6726
rect 2044 6719 2111 6723
rect 2044 6693 2056 6719
rect 2082 6697 2111 6719
rect 2137 6697 2144 6723
rect 2082 6693 2144 6697
rect 2044 6689 2144 6693
rect 143 6684 153 6688
rect 594 6687 764 6688
rect 115 6674 153 6684
rect 115 6596 150 6674
rect 727 6664 764 6687
rect 1520 6668 1551 6689
rect 1941 6668 1977 6689
rect 1363 6667 1400 6668
rect 111 6587 150 6596
rect 111 6569 121 6587
rect 139 6569 150 6587
rect 111 6563 150 6569
rect 306 6639 556 6663
rect 306 6568 343 6639
rect 458 6578 489 6579
rect 111 6559 148 6563
rect 306 6548 315 6568
rect 335 6548 343 6568
rect 306 6538 343 6548
rect 402 6568 489 6578
rect 402 6548 411 6568
rect 431 6548 489 6568
rect 402 6539 489 6548
rect 402 6538 439 6539
rect 114 6488 151 6497
rect 112 6470 123 6488
rect 141 6470 151 6488
rect 458 6486 489 6539
rect 519 6568 556 6639
rect 727 6644 1120 6664
rect 1140 6644 1143 6664
rect 727 6639 1143 6644
rect 1362 6658 1400 6667
rect 727 6638 1068 6639
rect 1362 6638 1371 6658
rect 1391 6638 1400 6658
rect 671 6578 702 6579
rect 519 6548 528 6568
rect 548 6548 556 6568
rect 519 6538 556 6548
rect 615 6571 702 6578
rect 615 6568 676 6571
rect 615 6548 624 6568
rect 644 6551 676 6568
rect 697 6551 702 6571
rect 644 6548 702 6551
rect 615 6541 702 6548
rect 727 6568 764 6638
rect 1030 6637 1067 6638
rect 1362 6630 1400 6638
rect 1466 6662 1551 6668
rect 1576 6667 1613 6668
rect 1466 6642 1474 6662
rect 1494 6642 1551 6662
rect 1466 6634 1551 6642
rect 1575 6658 1613 6667
rect 1575 6638 1584 6658
rect 1604 6638 1613 6658
rect 1466 6633 1502 6634
rect 1575 6630 1613 6638
rect 1679 6662 1764 6668
rect 1784 6667 1821 6668
rect 1679 6642 1687 6662
rect 1707 6661 1764 6662
rect 1707 6642 1736 6661
rect 1679 6641 1736 6642
rect 1757 6641 1764 6661
rect 1679 6634 1764 6641
rect 1783 6658 1821 6667
rect 1783 6638 1792 6658
rect 1812 6638 1821 6658
rect 1679 6633 1715 6634
rect 1783 6630 1821 6638
rect 1887 6662 2031 6668
rect 1887 6642 1895 6662
rect 1915 6660 2003 6662
rect 1915 6643 1951 6660
rect 1975 6643 2003 6660
rect 1915 6642 2003 6643
rect 2023 6642 2031 6662
rect 1887 6634 2031 6642
rect 1887 6633 1923 6634
rect 1995 6633 2031 6634
rect 2097 6667 2134 6668
rect 2097 6666 2135 6667
rect 2097 6658 2161 6666
rect 2097 6638 2106 6658
rect 2126 6644 2161 6658
rect 2181 6644 2184 6664
rect 2126 6639 2184 6644
rect 2126 6638 2161 6639
rect 1363 6601 1400 6630
rect 1364 6599 1400 6601
rect 1576 6599 1613 6630
rect 879 6578 915 6579
rect 727 6548 736 6568
rect 756 6548 764 6568
rect 615 6539 671 6541
rect 615 6538 652 6539
rect 727 6538 764 6548
rect 823 6568 971 6578
rect 1364 6577 1613 6599
rect 1784 6598 1821 6630
rect 2097 6626 2161 6638
rect 2201 6600 2228 6778
rect 2060 6598 2228 6600
rect 1784 6587 2228 6598
rect 1071 6575 1167 6577
rect 823 6548 832 6568
rect 852 6548 942 6568
rect 962 6548 971 6568
rect 823 6539 971 6548
rect 1029 6568 1167 6575
rect 1784 6572 2230 6587
rect 2060 6571 2230 6572
rect 1029 6548 1038 6568
rect 1058 6548 1167 6568
rect 1029 6539 1167 6548
rect 823 6538 860 6539
rect 879 6487 915 6539
rect 934 6538 971 6539
rect 1030 6538 1067 6539
rect 350 6485 391 6486
rect 112 6321 151 6470
rect 242 6478 391 6485
rect 242 6458 360 6478
rect 380 6458 391 6478
rect 242 6450 391 6458
rect 458 6482 817 6486
rect 458 6477 780 6482
rect 458 6453 571 6477
rect 595 6458 780 6477
rect 804 6458 817 6482
rect 595 6453 817 6458
rect 458 6450 817 6453
rect 879 6450 914 6487
rect 982 6484 1082 6487
rect 982 6480 1049 6484
rect 982 6454 994 6480
rect 1020 6458 1049 6480
rect 1075 6458 1082 6484
rect 1020 6454 1082 6458
rect 982 6450 1082 6454
rect 458 6429 489 6450
rect 879 6429 915 6450
rect 301 6428 338 6429
rect 300 6419 338 6428
rect 300 6399 309 6419
rect 329 6399 338 6419
rect 300 6391 338 6399
rect 404 6423 489 6429
rect 514 6428 551 6429
rect 404 6403 412 6423
rect 432 6403 489 6423
rect 404 6395 489 6403
rect 513 6419 551 6428
rect 513 6399 522 6419
rect 542 6399 551 6419
rect 404 6394 440 6395
rect 513 6391 551 6399
rect 617 6423 702 6429
rect 722 6428 759 6429
rect 617 6403 625 6423
rect 645 6422 702 6423
rect 645 6403 674 6422
rect 617 6402 674 6403
rect 695 6402 702 6422
rect 617 6395 702 6402
rect 721 6419 759 6428
rect 721 6399 730 6419
rect 750 6399 759 6419
rect 617 6394 653 6395
rect 721 6391 759 6399
rect 825 6424 969 6429
rect 825 6423 890 6424
rect 825 6403 833 6423
rect 853 6403 890 6423
rect 912 6423 969 6424
rect 912 6403 941 6423
rect 961 6403 969 6423
rect 825 6395 969 6403
rect 825 6394 861 6395
rect 933 6394 969 6395
rect 1035 6428 1072 6429
rect 1035 6427 1073 6428
rect 1035 6419 1099 6427
rect 1035 6399 1044 6419
rect 1064 6405 1099 6419
rect 1119 6405 1122 6425
rect 1064 6400 1122 6405
rect 1064 6399 1099 6400
rect 301 6362 338 6391
rect 302 6360 338 6362
rect 514 6360 551 6391
rect 302 6338 551 6360
rect 722 6359 759 6391
rect 1035 6387 1099 6399
rect 1139 6361 1166 6539
rect 998 6359 1166 6361
rect 722 6333 1166 6359
rect 1318 6458 1568 6482
rect 1318 6387 1355 6458
rect 1470 6397 1501 6398
rect 1318 6367 1327 6387
rect 1347 6367 1355 6387
rect 1318 6357 1355 6367
rect 1414 6387 1501 6397
rect 1414 6367 1423 6387
rect 1443 6367 1501 6387
rect 1414 6358 1501 6367
rect 1414 6357 1451 6358
rect 722 6323 744 6333
rect 998 6332 1166 6333
rect 682 6321 744 6323
rect 112 6314 744 6321
rect 111 6305 744 6314
rect 1470 6305 1501 6358
rect 1531 6387 1568 6458
rect 1739 6463 2132 6483
rect 2152 6463 2155 6483
rect 1739 6458 2155 6463
rect 1739 6457 2080 6458
rect 1683 6397 1714 6398
rect 1531 6367 1540 6387
rect 1560 6367 1568 6387
rect 1531 6357 1568 6367
rect 1627 6390 1714 6397
rect 1627 6387 1688 6390
rect 1627 6367 1636 6387
rect 1656 6370 1688 6387
rect 1709 6370 1714 6390
rect 1656 6367 1714 6370
rect 1627 6360 1714 6367
rect 1739 6387 1776 6457
rect 2042 6456 2079 6457
rect 1891 6397 1927 6398
rect 1739 6367 1748 6387
rect 1768 6367 1776 6387
rect 1627 6358 1683 6360
rect 1627 6357 1664 6358
rect 1739 6357 1776 6367
rect 1835 6387 1983 6397
rect 2083 6394 2179 6396
rect 1835 6367 1844 6387
rect 1864 6367 1954 6387
rect 1974 6367 1983 6387
rect 1835 6358 1983 6367
rect 2041 6387 2179 6394
rect 2041 6367 2050 6387
rect 2070 6367 2179 6387
rect 2041 6358 2179 6367
rect 1835 6357 1872 6358
rect 1891 6306 1927 6358
rect 1946 6357 1983 6358
rect 2042 6357 2079 6358
rect 111 6287 121 6305
rect 139 6304 744 6305
rect 1362 6304 1403 6305
rect 139 6299 160 6304
rect 139 6287 151 6299
rect 1254 6297 1403 6304
rect 111 6279 151 6287
rect 194 6286 220 6287
rect 111 6277 148 6279
rect 194 6268 748 6286
rect 1254 6277 1372 6297
rect 1392 6277 1403 6297
rect 1254 6269 1403 6277
rect 1470 6301 1829 6305
rect 1470 6296 1792 6301
rect 1470 6272 1583 6296
rect 1607 6277 1792 6296
rect 1816 6277 1829 6301
rect 1607 6272 1829 6277
rect 1470 6269 1829 6272
rect 1891 6269 1926 6306
rect 1994 6303 2094 6306
rect 1994 6299 2061 6303
rect 1994 6273 2006 6299
rect 2032 6277 2061 6299
rect 2087 6277 2094 6303
rect 2032 6273 2094 6277
rect 1994 6269 2094 6273
rect 114 6209 151 6215
rect 194 6209 220 6268
rect 727 6249 748 6268
rect 114 6206 220 6209
rect 114 6188 123 6206
rect 141 6192 220 6206
rect 305 6224 555 6248
rect 141 6190 217 6192
rect 141 6188 151 6190
rect 114 6178 151 6188
rect 119 6113 150 6178
rect 305 6153 342 6224
rect 457 6163 488 6164
rect 305 6133 314 6153
rect 334 6133 342 6153
rect 305 6123 342 6133
rect 401 6153 488 6163
rect 401 6133 410 6153
rect 430 6133 488 6153
rect 401 6124 488 6133
rect 401 6123 438 6124
rect 118 6104 155 6113
rect 118 6086 128 6104
rect 146 6086 155 6104
rect 118 6076 155 6086
rect 457 6071 488 6124
rect 518 6153 555 6224
rect 726 6229 1119 6249
rect 1139 6229 1142 6249
rect 1470 6248 1501 6269
rect 1891 6248 1927 6269
rect 1313 6247 1350 6248
rect 726 6224 1142 6229
rect 1312 6238 1350 6247
rect 726 6223 1067 6224
rect 670 6163 701 6164
rect 518 6133 527 6153
rect 547 6133 555 6153
rect 518 6123 555 6133
rect 614 6156 701 6163
rect 614 6153 675 6156
rect 614 6133 623 6153
rect 643 6136 675 6153
rect 696 6136 701 6156
rect 643 6133 701 6136
rect 614 6126 701 6133
rect 726 6153 763 6223
rect 1029 6222 1066 6223
rect 1312 6218 1321 6238
rect 1341 6218 1350 6238
rect 1312 6210 1350 6218
rect 1416 6242 1501 6248
rect 1526 6247 1563 6248
rect 1416 6222 1424 6242
rect 1444 6222 1501 6242
rect 1416 6214 1501 6222
rect 1525 6238 1563 6247
rect 1525 6218 1534 6238
rect 1554 6218 1563 6238
rect 1416 6213 1452 6214
rect 1525 6210 1563 6218
rect 1629 6242 1714 6248
rect 1734 6247 1771 6248
rect 1629 6222 1637 6242
rect 1657 6241 1714 6242
rect 1657 6222 1686 6241
rect 1629 6221 1686 6222
rect 1707 6221 1714 6241
rect 1629 6214 1714 6221
rect 1733 6238 1771 6247
rect 1733 6218 1742 6238
rect 1762 6218 1771 6238
rect 1629 6213 1665 6214
rect 1733 6210 1771 6218
rect 1837 6243 1981 6248
rect 1837 6242 1896 6243
rect 1837 6222 1845 6242
rect 1865 6223 1896 6242
rect 1920 6242 1981 6243
rect 1920 6223 1953 6242
rect 1865 6222 1953 6223
rect 1973 6222 1981 6242
rect 1837 6214 1981 6222
rect 1837 6213 1873 6214
rect 1945 6213 1981 6214
rect 2047 6247 2084 6248
rect 2047 6246 2085 6247
rect 2047 6238 2111 6246
rect 2047 6218 2056 6238
rect 2076 6224 2111 6238
rect 2131 6224 2134 6244
rect 2076 6219 2134 6224
rect 2076 6218 2111 6219
rect 1313 6181 1350 6210
rect 1314 6179 1350 6181
rect 1526 6179 1563 6210
rect 878 6163 914 6164
rect 726 6133 735 6153
rect 755 6133 763 6153
rect 614 6124 670 6126
rect 614 6123 651 6124
rect 726 6123 763 6133
rect 822 6153 970 6163
rect 1070 6160 1166 6162
rect 822 6133 831 6153
rect 851 6133 941 6153
rect 961 6133 970 6153
rect 822 6124 970 6133
rect 1028 6153 1166 6160
rect 1314 6157 1563 6179
rect 1734 6178 1771 6210
rect 2047 6206 2111 6218
rect 2151 6180 2178 6358
rect 2010 6178 2178 6180
rect 1734 6174 2178 6178
rect 1028 6133 1037 6153
rect 1057 6133 1166 6153
rect 1734 6155 1783 6174
rect 1803 6155 2178 6174
rect 1734 6152 2178 6155
rect 2010 6151 2178 6152
rect 2199 6177 2230 6571
rect 2199 6151 2204 6177
rect 2223 6151 2230 6177
rect 2199 6148 2230 6151
rect 1028 6124 1166 6133
rect 822 6123 859 6124
rect 878 6072 914 6124
rect 933 6123 970 6124
rect 1029 6123 1066 6124
rect 349 6070 390 6071
rect 241 6063 390 6070
rect 241 6043 359 6063
rect 379 6043 390 6063
rect 241 6035 390 6043
rect 457 6067 816 6071
rect 457 6062 779 6067
rect 457 6038 570 6062
rect 594 6043 779 6062
rect 803 6043 816 6067
rect 594 6038 816 6043
rect 457 6035 816 6038
rect 878 6035 913 6072
rect 981 6069 1081 6072
rect 981 6065 1048 6069
rect 981 6039 993 6065
rect 1019 6043 1048 6065
rect 1074 6043 1081 6069
rect 1019 6039 1081 6043
rect 981 6035 1081 6039
rect 457 6014 488 6035
rect 878 6014 914 6035
rect 121 6005 158 6014
rect 300 6013 337 6014
rect 121 5987 130 6005
rect 148 5987 158 6005
rect 121 5977 158 5987
rect 122 5942 158 5977
rect 299 6004 337 6013
rect 299 5984 308 6004
rect 328 5984 337 6004
rect 299 5976 337 5984
rect 403 6008 488 6014
rect 513 6013 550 6014
rect 403 5988 411 6008
rect 431 5988 488 6008
rect 403 5980 488 5988
rect 512 6004 550 6013
rect 512 5984 521 6004
rect 541 5984 550 6004
rect 403 5979 439 5980
rect 512 5976 550 5984
rect 616 6008 701 6014
rect 721 6013 758 6014
rect 616 5988 624 6008
rect 644 6007 701 6008
rect 644 5988 673 6007
rect 616 5987 673 5988
rect 694 5987 701 6007
rect 616 5980 701 5987
rect 720 6004 758 6013
rect 720 5984 729 6004
rect 749 5984 758 6004
rect 616 5979 652 5980
rect 720 5976 758 5984
rect 824 6008 968 6014
rect 824 5988 832 6008
rect 852 6007 940 6008
rect 852 5988 880 6007
rect 824 5986 880 5988
rect 902 5988 940 6007
rect 960 5988 968 6008
rect 902 5986 968 5988
rect 824 5980 968 5986
rect 824 5979 860 5980
rect 932 5979 968 5980
rect 1034 6013 1071 6014
rect 1034 6012 1072 6013
rect 1034 6004 1098 6012
rect 1034 5984 1043 6004
rect 1063 5990 1098 6004
rect 1118 5990 1121 6010
rect 1063 5985 1121 5990
rect 1063 5984 1098 5985
rect 300 5947 337 5976
rect 120 5901 158 5942
rect 301 5945 337 5947
rect 513 5945 550 5976
rect 301 5923 550 5945
rect 721 5944 758 5976
rect 1034 5972 1098 5984
rect 1138 5946 1165 6124
rect 2749 6113 2786 6124
rect 2875 6117 2905 7118
rect 2968 7118 3412 7129
rect 2968 7116 3136 7118
rect 2968 6938 2995 7116
rect 3035 7078 3099 7090
rect 3375 7086 3412 7118
rect 3583 7117 3832 7139
rect 4225 7138 4373 7148
rect 4432 7168 4469 7178
rect 4544 7177 4581 7178
rect 4525 7175 4581 7177
rect 4432 7148 4440 7168
rect 4460 7148 4469 7168
rect 4281 7137 4317 7138
rect 3583 7086 3620 7117
rect 3796 7115 3832 7117
rect 3796 7086 3833 7115
rect 3035 7077 3070 7078
rect 3012 7072 3070 7077
rect 3012 7052 3015 7072
rect 3035 7058 3070 7072
rect 3090 7058 3099 7078
rect 3035 7050 3099 7058
rect 3061 7049 3099 7050
rect 3062 7048 3099 7049
rect 3165 7082 3201 7083
rect 3273 7082 3309 7083
rect 3165 7074 3309 7082
rect 3165 7054 3173 7074
rect 3193 7055 3225 7074
rect 3248 7055 3281 7074
rect 3193 7054 3281 7055
rect 3301 7054 3309 7074
rect 3165 7048 3309 7054
rect 3375 7078 3413 7086
rect 3481 7082 3517 7083
rect 3375 7058 3384 7078
rect 3404 7058 3413 7078
rect 3375 7049 3413 7058
rect 3432 7075 3517 7082
rect 3432 7055 3439 7075
rect 3460 7074 3517 7075
rect 3460 7055 3489 7074
rect 3432 7054 3489 7055
rect 3509 7054 3517 7074
rect 3375 7048 3412 7049
rect 3432 7048 3517 7054
rect 3583 7078 3621 7086
rect 3694 7082 3730 7083
rect 3583 7058 3592 7078
rect 3612 7058 3621 7078
rect 3583 7049 3621 7058
rect 3645 7074 3730 7082
rect 3645 7054 3702 7074
rect 3722 7054 3730 7074
rect 3583 7048 3620 7049
rect 3645 7048 3730 7054
rect 3796 7078 3834 7086
rect 4129 7078 4166 7079
rect 4432 7078 4469 7148
rect 4494 7168 4581 7175
rect 4494 7165 4552 7168
rect 4494 7145 4499 7165
rect 4520 7148 4552 7165
rect 4572 7148 4581 7168
rect 4520 7145 4581 7148
rect 4494 7138 4581 7145
rect 4640 7168 4677 7178
rect 4640 7148 4648 7168
rect 4668 7148 4677 7168
rect 4494 7137 4525 7138
rect 3796 7058 3805 7078
rect 3825 7058 3834 7078
rect 4128 7077 4469 7078
rect 3796 7049 3834 7058
rect 4053 7072 4469 7077
rect 4053 7052 4056 7072
rect 4076 7052 4469 7072
rect 4640 7077 4677 7148
rect 4707 7177 4738 7230
rect 5045 7228 5055 7246
rect 5073 7228 5084 7246
rect 5045 7219 5082 7228
rect 4757 7177 4794 7178
rect 4707 7168 4794 7177
rect 4707 7148 4765 7168
rect 4785 7148 4794 7168
rect 4707 7138 4794 7148
rect 4853 7168 4890 7178
rect 4853 7148 4861 7168
rect 4881 7148 4890 7168
rect 5048 7153 5085 7157
rect 4707 7137 4738 7138
rect 4853 7077 4890 7148
rect 4640 7053 4890 7077
rect 5046 7147 5085 7153
rect 5046 7129 5057 7147
rect 5075 7129 5085 7147
rect 5046 7120 5085 7129
rect 3796 7048 3833 7049
rect 3219 7027 3255 7048
rect 3645 7027 3676 7048
rect 4432 7029 4469 7052
rect 5046 7042 5081 7120
rect 5043 7032 5081 7042
rect 4432 7028 4602 7029
rect 5043 7028 5053 7032
rect 3052 7023 3152 7027
rect 3052 7019 3114 7023
rect 3052 6993 3059 7019
rect 3085 6997 3114 7019
rect 3140 6997 3152 7023
rect 3085 6993 3152 6997
rect 3052 6990 3152 6993
rect 3220 6990 3255 7027
rect 3317 7024 3676 7027
rect 3317 7019 3539 7024
rect 3317 6995 3330 7019
rect 3354 7000 3539 7019
rect 3563 7000 3676 7024
rect 3354 6995 3676 7000
rect 3317 6991 3676 6995
rect 3743 7019 3892 7027
rect 3743 6999 3754 7019
rect 3774 6999 3892 7019
rect 4432 7014 5053 7028
rect 5071 7014 5081 7032
rect 4432 7008 5081 7014
rect 4432 7007 5080 7008
rect 5043 7005 5080 7007
rect 3743 6992 3892 6999
rect 3743 6991 3784 6992
rect 3067 6938 3104 6939
rect 3163 6938 3200 6939
rect 3219 6938 3255 6990
rect 3274 6938 3311 6939
rect 2967 6929 3105 6938
rect 2967 6909 3076 6929
rect 3096 6909 3105 6929
rect 2967 6902 3105 6909
rect 3163 6929 3311 6938
rect 3163 6909 3172 6929
rect 3192 6909 3282 6929
rect 3302 6909 3311 6929
rect 2967 6900 3063 6902
rect 3163 6899 3311 6909
rect 3370 6929 3407 6939
rect 3482 6938 3519 6939
rect 3463 6936 3519 6938
rect 3370 6909 3378 6929
rect 3398 6909 3407 6929
rect 3219 6898 3255 6899
rect 3067 6839 3104 6840
rect 3370 6839 3407 6909
rect 3432 6929 3519 6936
rect 3432 6926 3490 6929
rect 3432 6906 3437 6926
rect 3458 6909 3490 6926
rect 3510 6909 3519 6929
rect 3458 6906 3519 6909
rect 3432 6899 3519 6906
rect 3578 6929 3615 6939
rect 3578 6909 3586 6929
rect 3606 6909 3615 6929
rect 3432 6898 3463 6899
rect 3066 6838 3407 6839
rect 2991 6833 3407 6838
rect 2991 6813 2994 6833
rect 3014 6813 3407 6833
rect 3578 6838 3615 6909
rect 3645 6938 3676 6991
rect 3695 6938 3732 6939
rect 3645 6929 3732 6938
rect 3645 6909 3703 6929
rect 3723 6909 3732 6929
rect 3645 6899 3732 6909
rect 3791 6929 3828 6939
rect 3791 6909 3799 6929
rect 3819 6909 3828 6929
rect 3645 6898 3676 6899
rect 3791 6838 3828 6909
rect 5046 6933 5083 6943
rect 5046 6915 5055 6933
rect 5073 6915 5083 6933
rect 5046 6906 5083 6915
rect 5046 6882 5081 6906
rect 5044 6858 5081 6882
rect 5043 6852 5081 6858
rect 3578 6814 3828 6838
rect 4454 6834 5081 6852
rect 4036 6817 4204 6818
rect 4455 6817 4479 6834
rect 4036 6791 4480 6817
rect 4036 6789 4204 6791
rect 4036 6611 4063 6789
rect 4103 6751 4167 6763
rect 4443 6759 4480 6791
rect 4651 6790 4900 6812
rect 4651 6759 4688 6790
rect 4864 6788 4900 6790
rect 5043 6793 5081 6834
rect 4864 6759 4901 6788
rect 4103 6750 4138 6751
rect 4080 6745 4138 6750
rect 4080 6725 4083 6745
rect 4103 6731 4138 6745
rect 4158 6731 4167 6751
rect 4103 6723 4167 6731
rect 4129 6722 4167 6723
rect 4130 6721 4167 6722
rect 4233 6755 4269 6756
rect 4341 6755 4377 6756
rect 4233 6749 4377 6755
rect 4233 6747 4299 6749
rect 4233 6727 4241 6747
rect 4261 6728 4299 6747
rect 4321 6747 4377 6749
rect 4321 6728 4349 6747
rect 4261 6727 4349 6728
rect 4369 6727 4377 6747
rect 4233 6721 4377 6727
rect 4443 6751 4481 6759
rect 4549 6755 4585 6756
rect 4443 6731 4452 6751
rect 4472 6731 4481 6751
rect 4443 6722 4481 6731
rect 4500 6748 4585 6755
rect 4500 6728 4507 6748
rect 4528 6747 4585 6748
rect 4528 6728 4557 6747
rect 4500 6727 4557 6728
rect 4577 6727 4585 6747
rect 4443 6721 4480 6722
rect 4500 6721 4585 6727
rect 4651 6751 4689 6759
rect 4762 6755 4798 6756
rect 4651 6731 4660 6751
rect 4680 6731 4689 6751
rect 4651 6722 4689 6731
rect 4713 6747 4798 6755
rect 4713 6727 4770 6747
rect 4790 6727 4798 6747
rect 4651 6721 4688 6722
rect 4713 6721 4798 6727
rect 4864 6751 4902 6759
rect 4864 6731 4873 6751
rect 4893 6731 4902 6751
rect 4864 6722 4902 6731
rect 5043 6758 5079 6793
rect 5043 6748 5080 6758
rect 5043 6730 5053 6748
rect 5071 6730 5080 6748
rect 4864 6721 4901 6722
rect 5043 6721 5080 6730
rect 4287 6700 4323 6721
rect 4713 6700 4744 6721
rect 4120 6696 4220 6700
rect 4120 6692 4182 6696
rect 4120 6666 4127 6692
rect 4153 6670 4182 6692
rect 4208 6670 4220 6696
rect 4153 6666 4220 6670
rect 4120 6663 4220 6666
rect 4288 6663 4323 6700
rect 4385 6697 4744 6700
rect 4385 6692 4607 6697
rect 4385 6668 4398 6692
rect 4422 6673 4607 6692
rect 4631 6673 4744 6697
rect 4422 6668 4744 6673
rect 4385 6664 4744 6668
rect 4811 6692 4960 6700
rect 4811 6672 4822 6692
rect 4842 6672 4960 6692
rect 4811 6665 4960 6672
rect 4811 6664 4852 6665
rect 4135 6611 4172 6612
rect 4231 6611 4268 6612
rect 4287 6611 4323 6663
rect 4342 6611 4379 6612
rect 4035 6602 4173 6611
rect 3023 6583 3191 6584
rect 3023 6580 3467 6583
rect 3023 6561 3398 6580
rect 3418 6561 3467 6580
rect 4035 6582 4144 6602
rect 4164 6582 4173 6602
rect 3023 6557 3467 6561
rect 3023 6555 3191 6557
rect 3023 6377 3050 6555
rect 3090 6517 3154 6529
rect 3430 6525 3467 6557
rect 3638 6556 3887 6578
rect 4035 6575 4173 6582
rect 4231 6602 4379 6611
rect 4231 6582 4240 6602
rect 4260 6582 4350 6602
rect 4370 6582 4379 6602
rect 4035 6573 4131 6575
rect 4231 6572 4379 6582
rect 4438 6602 4475 6612
rect 4550 6611 4587 6612
rect 4531 6609 4587 6611
rect 4438 6582 4446 6602
rect 4466 6582 4475 6602
rect 4287 6571 4323 6572
rect 3638 6525 3675 6556
rect 3851 6554 3887 6556
rect 3851 6525 3888 6554
rect 3090 6516 3125 6517
rect 3067 6511 3125 6516
rect 3067 6491 3070 6511
rect 3090 6497 3125 6511
rect 3145 6497 3154 6517
rect 3090 6489 3154 6497
rect 3116 6488 3154 6489
rect 3117 6487 3154 6488
rect 3220 6521 3256 6522
rect 3328 6521 3364 6522
rect 3220 6513 3364 6521
rect 3220 6493 3228 6513
rect 3248 6493 3280 6513
rect 3304 6493 3336 6513
rect 3356 6493 3364 6513
rect 3220 6487 3364 6493
rect 3430 6517 3468 6525
rect 3536 6521 3572 6522
rect 3430 6497 3439 6517
rect 3459 6497 3468 6517
rect 3430 6488 3468 6497
rect 3487 6514 3572 6521
rect 3487 6494 3494 6514
rect 3515 6513 3572 6514
rect 3515 6494 3544 6513
rect 3487 6493 3544 6494
rect 3564 6493 3572 6513
rect 3430 6487 3467 6488
rect 3487 6487 3572 6493
rect 3638 6517 3676 6525
rect 3749 6521 3785 6522
rect 3638 6497 3647 6517
rect 3667 6497 3676 6517
rect 3638 6488 3676 6497
rect 3700 6513 3785 6521
rect 3700 6493 3757 6513
rect 3777 6493 3785 6513
rect 3638 6487 3675 6488
rect 3700 6487 3785 6493
rect 3851 6517 3889 6525
rect 3851 6497 3860 6517
rect 3880 6497 3889 6517
rect 4135 6512 4172 6513
rect 4438 6512 4475 6582
rect 4500 6602 4587 6609
rect 4500 6599 4558 6602
rect 4500 6579 4505 6599
rect 4526 6582 4558 6599
rect 4578 6582 4587 6602
rect 4526 6579 4587 6582
rect 4500 6572 4587 6579
rect 4646 6602 4683 6612
rect 4646 6582 4654 6602
rect 4674 6582 4683 6602
rect 4500 6571 4531 6572
rect 4134 6511 4475 6512
rect 3851 6488 3889 6497
rect 4059 6506 4475 6511
rect 3851 6487 3888 6488
rect 3274 6466 3310 6487
rect 3700 6466 3731 6487
rect 4059 6486 4062 6506
rect 4082 6486 4475 6506
rect 4646 6511 4683 6582
rect 4713 6611 4744 6664
rect 5046 6649 5083 6659
rect 5046 6631 5055 6649
rect 5073 6631 5083 6649
rect 5046 6622 5083 6631
rect 4763 6611 4800 6612
rect 4713 6602 4800 6611
rect 4713 6582 4771 6602
rect 4791 6582 4800 6602
rect 4713 6572 4800 6582
rect 4859 6602 4896 6612
rect 4859 6582 4867 6602
rect 4887 6582 4896 6602
rect 4713 6571 4744 6572
rect 4859 6511 4896 6582
rect 5051 6557 5082 6622
rect 5050 6547 5087 6557
rect 5050 6545 5060 6547
rect 4984 6543 5060 6545
rect 4646 6487 4896 6511
rect 4981 6529 5060 6543
rect 5078 6529 5087 6547
rect 4981 6526 5087 6529
rect 4453 6467 4474 6486
rect 4981 6467 5007 6526
rect 5050 6520 5087 6526
rect 3107 6462 3207 6466
rect 3107 6458 3169 6462
rect 3107 6432 3114 6458
rect 3140 6436 3169 6458
rect 3195 6436 3207 6462
rect 3140 6432 3207 6436
rect 3107 6429 3207 6432
rect 3275 6429 3310 6466
rect 3372 6463 3731 6466
rect 3372 6458 3594 6463
rect 3372 6434 3385 6458
rect 3409 6439 3594 6458
rect 3618 6439 3731 6463
rect 3409 6434 3731 6439
rect 3372 6430 3731 6434
rect 3798 6458 3947 6466
rect 3798 6438 3809 6458
rect 3829 6438 3947 6458
rect 4453 6449 5007 6467
rect 5053 6456 5090 6458
rect 4981 6448 5007 6449
rect 5050 6448 5090 6456
rect 3798 6431 3947 6438
rect 5050 6436 5062 6448
rect 5041 6431 5062 6436
rect 3798 6430 3839 6431
rect 4457 6430 5062 6431
rect 5080 6430 5090 6448
rect 3122 6377 3159 6378
rect 3218 6377 3255 6378
rect 3274 6377 3310 6429
rect 3329 6377 3366 6378
rect 3022 6368 3160 6377
rect 3022 6348 3131 6368
rect 3151 6348 3160 6368
rect 3022 6341 3160 6348
rect 3218 6368 3366 6377
rect 3218 6348 3227 6368
rect 3247 6348 3337 6368
rect 3357 6348 3366 6368
rect 3022 6339 3118 6341
rect 3218 6338 3366 6348
rect 3425 6368 3462 6378
rect 3537 6377 3574 6378
rect 3518 6375 3574 6377
rect 3425 6348 3433 6368
rect 3453 6348 3462 6368
rect 3274 6337 3310 6338
rect 3122 6278 3159 6279
rect 3425 6278 3462 6348
rect 3487 6368 3574 6375
rect 3487 6365 3545 6368
rect 3487 6345 3492 6365
rect 3513 6348 3545 6365
rect 3565 6348 3574 6368
rect 3513 6345 3574 6348
rect 3487 6338 3574 6345
rect 3633 6368 3670 6378
rect 3633 6348 3641 6368
rect 3661 6348 3670 6368
rect 3487 6337 3518 6338
rect 3121 6277 3462 6278
rect 3046 6272 3462 6277
rect 3046 6252 3049 6272
rect 3069 6252 3462 6272
rect 3633 6277 3670 6348
rect 3700 6377 3731 6430
rect 4457 6421 5090 6430
rect 4457 6414 5089 6421
rect 4457 6412 4519 6414
rect 4035 6402 4203 6403
rect 4457 6402 4479 6412
rect 3750 6377 3787 6378
rect 3700 6368 3787 6377
rect 3700 6348 3758 6368
rect 3778 6348 3787 6368
rect 3700 6338 3787 6348
rect 3846 6368 3883 6378
rect 3846 6348 3854 6368
rect 3874 6348 3883 6368
rect 3700 6337 3731 6338
rect 3846 6277 3883 6348
rect 3633 6253 3883 6277
rect 4035 6376 4479 6402
rect 4035 6374 4203 6376
rect 4035 6196 4062 6374
rect 4102 6336 4166 6348
rect 4442 6344 4479 6376
rect 4650 6375 4899 6397
rect 4650 6344 4687 6375
rect 4863 6373 4899 6375
rect 4863 6344 4900 6373
rect 4102 6335 4137 6336
rect 4079 6330 4137 6335
rect 4079 6310 4082 6330
rect 4102 6316 4137 6330
rect 4157 6316 4166 6336
rect 4102 6308 4166 6316
rect 4128 6307 4166 6308
rect 4129 6306 4166 6307
rect 4232 6340 4268 6341
rect 4340 6340 4376 6341
rect 4232 6332 4376 6340
rect 4232 6312 4240 6332
rect 4260 6312 4289 6332
rect 4232 6311 4289 6312
rect 4311 6312 4348 6332
rect 4368 6312 4376 6332
rect 4311 6311 4376 6312
rect 4232 6306 4376 6311
rect 4442 6336 4480 6344
rect 4548 6340 4584 6341
rect 4442 6316 4451 6336
rect 4471 6316 4480 6336
rect 4442 6307 4480 6316
rect 4499 6333 4584 6340
rect 4499 6313 4506 6333
rect 4527 6332 4584 6333
rect 4527 6313 4556 6332
rect 4499 6312 4556 6313
rect 4576 6312 4584 6332
rect 4442 6306 4479 6307
rect 4499 6306 4584 6312
rect 4650 6336 4688 6344
rect 4761 6340 4797 6341
rect 4650 6316 4659 6336
rect 4679 6316 4688 6336
rect 4650 6307 4688 6316
rect 4712 6332 4797 6340
rect 4712 6312 4769 6332
rect 4789 6312 4797 6332
rect 4650 6306 4687 6307
rect 4712 6306 4797 6312
rect 4863 6336 4901 6344
rect 4863 6316 4872 6336
rect 4892 6316 4901 6336
rect 4863 6307 4901 6316
rect 4863 6306 4900 6307
rect 4286 6285 4322 6306
rect 4712 6285 4743 6306
rect 4119 6281 4219 6285
rect 4119 6277 4181 6281
rect 4119 6251 4126 6277
rect 4152 6255 4181 6277
rect 4207 6255 4219 6281
rect 4152 6251 4219 6255
rect 4119 6248 4219 6251
rect 4287 6248 4322 6285
rect 4384 6282 4743 6285
rect 4384 6277 4606 6282
rect 4384 6253 4397 6277
rect 4421 6258 4606 6277
rect 4630 6258 4743 6282
rect 4421 6253 4743 6258
rect 4384 6249 4743 6253
rect 4810 6277 4959 6285
rect 4810 6257 4821 6277
rect 4841 6257 4959 6277
rect 4810 6250 4959 6257
rect 5050 6265 5089 6414
rect 4810 6249 4851 6250
rect 4134 6196 4171 6197
rect 4230 6196 4267 6197
rect 4286 6196 4322 6248
rect 4341 6196 4378 6197
rect 4034 6187 4172 6196
rect 4034 6167 4143 6187
rect 4163 6167 4172 6187
rect 4034 6160 4172 6167
rect 4230 6187 4378 6196
rect 4230 6167 4239 6187
rect 4259 6167 4349 6187
rect 4369 6167 4378 6187
rect 4034 6158 4130 6160
rect 4230 6157 4378 6167
rect 4437 6187 4474 6197
rect 4549 6196 4586 6197
rect 4530 6194 4586 6196
rect 4437 6167 4445 6187
rect 4465 6167 4474 6187
rect 4286 6156 4322 6157
rect 2749 6094 2757 6113
rect 2780 6094 2786 6113
rect 2749 6083 2786 6094
rect 2815 6116 2983 6117
rect 2815 6090 3259 6116
rect 2815 6088 2983 6090
rect 2752 6023 2785 6083
rect 997 5944 1165 5946
rect 721 5918 1165 5944
rect 722 5901 746 5918
rect 997 5917 1165 5918
rect 1533 5946 1783 5970
rect 120 5883 747 5901
rect 120 5877 158 5883
rect 122 5831 157 5877
rect 1533 5875 1570 5946
rect 1685 5885 1716 5886
rect 1533 5855 1542 5875
rect 1562 5855 1570 5875
rect 1533 5845 1570 5855
rect 1629 5875 1716 5885
rect 1629 5855 1638 5875
rect 1658 5855 1716 5875
rect 1629 5846 1716 5855
rect 1629 5845 1666 5846
rect 120 5822 157 5831
rect 120 5804 130 5822
rect 148 5804 157 5822
rect 120 5794 157 5804
rect 1685 5793 1716 5846
rect 1746 5875 1783 5946
rect 1954 5951 2347 5971
rect 2367 5951 2370 5971
rect 1954 5946 2370 5951
rect 1954 5945 2295 5946
rect 1898 5885 1929 5886
rect 1746 5855 1755 5875
rect 1775 5855 1783 5875
rect 1746 5845 1783 5855
rect 1842 5878 1929 5885
rect 1842 5875 1903 5878
rect 1842 5855 1851 5875
rect 1871 5858 1903 5875
rect 1924 5858 1929 5878
rect 1871 5855 1929 5858
rect 1842 5848 1929 5855
rect 1954 5875 1991 5945
rect 2257 5944 2294 5945
rect 2106 5885 2142 5886
rect 1954 5855 1963 5875
rect 1983 5855 1991 5875
rect 1842 5846 1898 5848
rect 1842 5845 1879 5846
rect 1954 5845 1991 5855
rect 2050 5875 2198 5885
rect 2298 5882 2394 5884
rect 2050 5855 2059 5875
rect 2079 5855 2169 5875
rect 2189 5855 2198 5875
rect 2050 5846 2198 5855
rect 2256 5875 2394 5882
rect 2256 5855 2265 5875
rect 2285 5855 2394 5875
rect 2256 5846 2394 5855
rect 2050 5845 2087 5846
rect 2106 5794 2142 5846
rect 2161 5845 2198 5846
rect 2257 5845 2294 5846
rect 1577 5792 1618 5793
rect 1469 5785 1618 5792
rect 1469 5765 1587 5785
rect 1607 5765 1618 5785
rect 1469 5757 1618 5765
rect 1685 5789 2044 5793
rect 1685 5784 2007 5789
rect 1685 5760 1798 5784
rect 1822 5765 2007 5784
rect 2031 5765 2044 5789
rect 1822 5760 2044 5765
rect 1685 5757 2044 5760
rect 2106 5757 2141 5794
rect 2209 5791 2309 5794
rect 2209 5787 2276 5791
rect 2209 5761 2221 5787
rect 2247 5765 2276 5787
rect 2302 5765 2309 5791
rect 2247 5761 2309 5765
rect 2209 5757 2309 5761
rect 1685 5736 1716 5757
rect 2106 5736 2142 5757
rect 1528 5735 1565 5736
rect 123 5730 160 5732
rect 123 5729 771 5730
rect 122 5723 771 5729
rect 122 5705 132 5723
rect 150 5709 771 5723
rect 150 5705 160 5709
rect 601 5708 771 5709
rect 122 5695 160 5705
rect 122 5617 157 5695
rect 734 5685 771 5708
rect 1527 5726 1565 5735
rect 1527 5706 1536 5726
rect 1556 5706 1565 5726
rect 1527 5698 1565 5706
rect 1631 5730 1716 5736
rect 1741 5735 1778 5736
rect 1631 5710 1639 5730
rect 1659 5710 1716 5730
rect 1631 5702 1716 5710
rect 1740 5726 1778 5735
rect 1740 5706 1749 5726
rect 1769 5706 1778 5726
rect 1631 5701 1667 5702
rect 1740 5698 1778 5706
rect 1844 5730 1929 5736
rect 1949 5735 1986 5736
rect 1844 5710 1852 5730
rect 1872 5729 1929 5730
rect 1872 5710 1901 5729
rect 1844 5709 1901 5710
rect 1922 5709 1929 5729
rect 1844 5702 1929 5709
rect 1948 5726 1986 5735
rect 1948 5706 1957 5726
rect 1977 5706 1986 5726
rect 1844 5701 1880 5702
rect 1948 5698 1986 5706
rect 2052 5734 2196 5736
rect 2052 5730 2110 5734
rect 2052 5710 2060 5730
rect 2080 5710 2110 5730
rect 2052 5708 2110 5710
rect 2135 5730 2196 5734
rect 2135 5710 2168 5730
rect 2188 5710 2196 5730
rect 2135 5708 2196 5710
rect 2052 5702 2196 5708
rect 2052 5701 2088 5702
rect 2160 5701 2196 5702
rect 2262 5735 2299 5736
rect 2262 5734 2300 5735
rect 2262 5726 2326 5734
rect 2262 5706 2271 5726
rect 2291 5712 2326 5726
rect 2346 5712 2349 5732
rect 2291 5707 2349 5712
rect 2291 5706 2326 5707
rect 118 5608 157 5617
rect 118 5590 128 5608
rect 146 5590 157 5608
rect 118 5584 157 5590
rect 313 5660 563 5684
rect 313 5589 350 5660
rect 465 5599 496 5600
rect 118 5580 155 5584
rect 313 5569 322 5589
rect 342 5569 350 5589
rect 313 5559 350 5569
rect 409 5589 496 5599
rect 409 5569 418 5589
rect 438 5569 496 5589
rect 409 5560 496 5569
rect 409 5559 446 5560
rect 121 5509 158 5518
rect 119 5491 130 5509
rect 148 5491 158 5509
rect 465 5507 496 5560
rect 526 5589 563 5660
rect 734 5665 1127 5685
rect 1147 5665 1150 5685
rect 1528 5669 1565 5698
rect 734 5660 1150 5665
rect 1529 5667 1565 5669
rect 1741 5667 1778 5698
rect 734 5659 1075 5660
rect 678 5599 709 5600
rect 526 5569 535 5589
rect 555 5569 563 5589
rect 526 5559 563 5569
rect 622 5592 709 5599
rect 622 5589 683 5592
rect 622 5569 631 5589
rect 651 5572 683 5589
rect 704 5572 709 5592
rect 651 5569 709 5572
rect 622 5562 709 5569
rect 734 5589 771 5659
rect 1037 5658 1074 5659
rect 1529 5645 1778 5667
rect 1949 5666 1986 5698
rect 2262 5694 2326 5706
rect 2366 5668 2393 5846
rect 2225 5666 2393 5668
rect 1949 5640 2393 5666
rect 2225 5639 2393 5640
rect 886 5599 922 5600
rect 734 5569 743 5589
rect 763 5569 771 5589
rect 622 5560 678 5562
rect 622 5559 659 5560
rect 734 5559 771 5569
rect 830 5589 978 5599
rect 1078 5596 1174 5598
rect 830 5569 839 5589
rect 859 5569 949 5589
rect 969 5569 978 5589
rect 830 5560 978 5569
rect 1036 5589 1174 5596
rect 1036 5569 1045 5589
rect 1065 5569 1174 5589
rect 1036 5560 1174 5569
rect 830 5559 867 5560
rect 886 5508 922 5560
rect 941 5559 978 5560
rect 1037 5559 1074 5560
rect 357 5506 398 5507
rect 119 5342 158 5491
rect 249 5499 398 5506
rect 249 5479 367 5499
rect 387 5479 398 5499
rect 249 5471 398 5479
rect 465 5503 824 5507
rect 465 5498 787 5503
rect 465 5474 578 5498
rect 602 5479 787 5498
rect 811 5479 824 5503
rect 602 5474 824 5479
rect 465 5471 824 5474
rect 886 5471 921 5508
rect 989 5505 1089 5508
rect 989 5501 1056 5505
rect 989 5475 1001 5501
rect 1027 5479 1056 5501
rect 1082 5479 1089 5505
rect 1027 5475 1089 5479
rect 989 5471 1089 5475
rect 465 5450 496 5471
rect 886 5450 922 5471
rect 308 5449 345 5450
rect 307 5440 345 5449
rect 307 5420 316 5440
rect 336 5420 345 5440
rect 307 5412 345 5420
rect 411 5444 496 5450
rect 521 5449 558 5450
rect 411 5424 419 5444
rect 439 5424 496 5444
rect 411 5416 496 5424
rect 520 5440 558 5449
rect 520 5420 529 5440
rect 549 5420 558 5440
rect 411 5415 447 5416
rect 520 5412 558 5420
rect 624 5444 709 5450
rect 729 5449 766 5450
rect 624 5424 632 5444
rect 652 5443 709 5444
rect 652 5424 681 5443
rect 624 5423 681 5424
rect 702 5423 709 5443
rect 624 5416 709 5423
rect 728 5440 766 5449
rect 728 5420 737 5440
rect 757 5420 766 5440
rect 624 5415 660 5416
rect 728 5412 766 5420
rect 832 5445 976 5450
rect 832 5444 897 5445
rect 832 5424 840 5444
rect 860 5424 897 5444
rect 919 5444 976 5445
rect 919 5424 948 5444
rect 968 5424 976 5444
rect 832 5416 976 5424
rect 832 5415 868 5416
rect 940 5415 976 5416
rect 1042 5449 1079 5450
rect 1042 5448 1080 5449
rect 1042 5440 1106 5448
rect 1042 5420 1051 5440
rect 1071 5426 1106 5440
rect 1126 5426 1129 5446
rect 1071 5421 1129 5426
rect 1071 5420 1106 5421
rect 308 5383 345 5412
rect 309 5381 345 5383
rect 521 5381 558 5412
rect 309 5359 558 5381
rect 729 5380 766 5412
rect 1042 5408 1106 5420
rect 1146 5382 1173 5560
rect 1005 5380 1173 5382
rect 729 5354 1173 5380
rect 1325 5479 1575 5503
rect 1325 5408 1362 5479
rect 1477 5418 1508 5419
rect 1325 5388 1334 5408
rect 1354 5388 1362 5408
rect 1325 5378 1362 5388
rect 1421 5408 1508 5418
rect 1421 5388 1430 5408
rect 1450 5388 1508 5408
rect 1421 5379 1508 5388
rect 1421 5378 1458 5379
rect 729 5344 751 5354
rect 1005 5353 1173 5354
rect 689 5342 751 5344
rect 119 5335 751 5342
rect 118 5326 751 5335
rect 1477 5326 1508 5379
rect 1538 5408 1575 5479
rect 1746 5484 2139 5504
rect 2159 5484 2162 5504
rect 1746 5479 2162 5484
rect 1746 5478 2087 5479
rect 1690 5418 1721 5419
rect 1538 5388 1547 5408
rect 1567 5388 1575 5408
rect 1538 5378 1575 5388
rect 1634 5411 1721 5418
rect 1634 5408 1695 5411
rect 1634 5388 1643 5408
rect 1663 5391 1695 5408
rect 1716 5391 1721 5411
rect 1663 5388 1721 5391
rect 1634 5381 1721 5388
rect 1746 5408 1783 5478
rect 2049 5477 2086 5478
rect 1898 5418 1934 5419
rect 1746 5388 1755 5408
rect 1775 5388 1783 5408
rect 1634 5379 1690 5381
rect 1634 5378 1671 5379
rect 1746 5378 1783 5388
rect 1842 5408 1990 5418
rect 2090 5415 2186 5417
rect 1842 5388 1851 5408
rect 1871 5388 1961 5408
rect 1981 5388 1990 5408
rect 1842 5379 1990 5388
rect 2048 5408 2186 5415
rect 2048 5388 2057 5408
rect 2077 5388 2186 5408
rect 2048 5379 2186 5388
rect 1842 5378 1879 5379
rect 1898 5327 1934 5379
rect 1953 5378 1990 5379
rect 2049 5378 2086 5379
rect 118 5308 128 5326
rect 146 5325 751 5326
rect 1369 5325 1410 5326
rect 146 5320 167 5325
rect 146 5308 158 5320
rect 1261 5318 1410 5325
rect 118 5300 158 5308
rect 201 5307 227 5308
rect 118 5298 155 5300
rect 201 5289 755 5307
rect 1261 5298 1379 5318
rect 1399 5298 1410 5318
rect 1261 5290 1410 5298
rect 1477 5322 1836 5326
rect 1477 5317 1799 5322
rect 1477 5293 1590 5317
rect 1614 5298 1799 5317
rect 1823 5298 1836 5322
rect 1614 5293 1836 5298
rect 1477 5290 1836 5293
rect 1898 5290 1933 5327
rect 2001 5324 2101 5327
rect 2001 5320 2068 5324
rect 2001 5294 2013 5320
rect 2039 5298 2068 5320
rect 2094 5298 2101 5324
rect 2039 5294 2101 5298
rect 2001 5290 2101 5294
rect 121 5230 158 5236
rect 201 5230 227 5289
rect 734 5270 755 5289
rect 121 5227 227 5230
rect 121 5209 130 5227
rect 148 5213 227 5227
rect 312 5245 562 5269
rect 148 5211 224 5213
rect 148 5209 158 5211
rect 121 5199 158 5209
rect 126 5134 157 5199
rect 312 5174 349 5245
rect 464 5184 495 5185
rect 312 5154 321 5174
rect 341 5154 349 5174
rect 312 5144 349 5154
rect 408 5174 495 5184
rect 408 5154 417 5174
rect 437 5154 495 5174
rect 408 5145 495 5154
rect 408 5144 445 5145
rect 125 5125 162 5134
rect 125 5107 135 5125
rect 153 5107 162 5125
rect 125 5097 162 5107
rect 464 5092 495 5145
rect 525 5174 562 5245
rect 733 5250 1126 5270
rect 1146 5250 1149 5270
rect 1477 5269 1508 5290
rect 1898 5269 1934 5290
rect 1320 5268 1357 5269
rect 733 5245 1149 5250
rect 1319 5259 1357 5268
rect 733 5244 1074 5245
rect 677 5184 708 5185
rect 525 5154 534 5174
rect 554 5154 562 5174
rect 525 5144 562 5154
rect 621 5177 708 5184
rect 621 5174 682 5177
rect 621 5154 630 5174
rect 650 5157 682 5174
rect 703 5157 708 5177
rect 650 5154 708 5157
rect 621 5147 708 5154
rect 733 5174 770 5244
rect 1036 5243 1073 5244
rect 1319 5239 1328 5259
rect 1348 5239 1357 5259
rect 1319 5231 1357 5239
rect 1423 5263 1508 5269
rect 1533 5268 1570 5269
rect 1423 5243 1431 5263
rect 1451 5243 1508 5263
rect 1423 5235 1508 5243
rect 1532 5259 1570 5268
rect 1532 5239 1541 5259
rect 1561 5239 1570 5259
rect 1423 5234 1459 5235
rect 1532 5231 1570 5239
rect 1636 5263 1721 5269
rect 1741 5268 1778 5269
rect 1636 5243 1644 5263
rect 1664 5262 1721 5263
rect 1664 5243 1693 5262
rect 1636 5242 1693 5243
rect 1714 5242 1721 5262
rect 1636 5235 1721 5242
rect 1740 5259 1778 5268
rect 1740 5239 1749 5259
rect 1769 5239 1778 5259
rect 1636 5234 1672 5235
rect 1740 5231 1778 5239
rect 1844 5263 1988 5269
rect 1844 5243 1852 5263
rect 1872 5243 1904 5263
rect 1928 5243 1960 5263
rect 1980 5243 1988 5263
rect 1844 5235 1988 5243
rect 1844 5234 1880 5235
rect 1952 5234 1988 5235
rect 2054 5268 2091 5269
rect 2054 5267 2092 5268
rect 2054 5259 2118 5267
rect 2054 5239 2063 5259
rect 2083 5245 2118 5259
rect 2138 5245 2141 5265
rect 2083 5240 2141 5245
rect 2083 5239 2118 5240
rect 1320 5202 1357 5231
rect 1321 5200 1357 5202
rect 1533 5200 1570 5231
rect 885 5184 921 5185
rect 733 5154 742 5174
rect 762 5154 770 5174
rect 621 5145 677 5147
rect 621 5144 658 5145
rect 733 5144 770 5154
rect 829 5174 977 5184
rect 1077 5181 1173 5183
rect 829 5154 838 5174
rect 858 5154 948 5174
rect 968 5154 977 5174
rect 829 5145 977 5154
rect 1035 5174 1173 5181
rect 1321 5178 1570 5200
rect 1741 5199 1778 5231
rect 2054 5227 2118 5239
rect 2158 5201 2185 5379
rect 2017 5199 2185 5201
rect 1741 5195 2185 5199
rect 1035 5154 1044 5174
rect 1064 5154 1173 5174
rect 1741 5176 1790 5195
rect 1810 5176 2185 5195
rect 1741 5173 2185 5176
rect 2017 5172 2185 5173
rect 1035 5145 1173 5154
rect 829 5144 866 5145
rect 885 5093 921 5145
rect 940 5144 977 5145
rect 1036 5144 1073 5145
rect 356 5091 397 5092
rect 248 5084 397 5091
rect 248 5064 366 5084
rect 386 5064 397 5084
rect 248 5056 397 5064
rect 464 5088 823 5092
rect 464 5083 786 5088
rect 464 5059 577 5083
rect 601 5064 786 5083
rect 810 5064 823 5088
rect 601 5059 823 5064
rect 464 5056 823 5059
rect 885 5056 920 5093
rect 988 5090 1088 5093
rect 988 5086 1055 5090
rect 988 5060 1000 5086
rect 1026 5064 1055 5086
rect 1081 5064 1088 5090
rect 1026 5060 1088 5064
rect 988 5056 1088 5060
rect 464 5035 495 5056
rect 885 5035 921 5056
rect 128 5026 165 5035
rect 307 5034 344 5035
rect 128 5008 137 5026
rect 155 5008 165 5026
rect 128 4998 165 5008
rect 129 4963 165 4998
rect 306 5025 344 5034
rect 306 5005 315 5025
rect 335 5005 344 5025
rect 306 4997 344 5005
rect 410 5029 495 5035
rect 520 5034 557 5035
rect 410 5009 418 5029
rect 438 5009 495 5029
rect 410 5001 495 5009
rect 519 5025 557 5034
rect 519 5005 528 5025
rect 548 5005 557 5025
rect 410 5000 446 5001
rect 519 4997 557 5005
rect 623 5029 708 5035
rect 728 5034 765 5035
rect 623 5009 631 5029
rect 651 5028 708 5029
rect 651 5009 680 5028
rect 623 5008 680 5009
rect 701 5008 708 5028
rect 623 5001 708 5008
rect 727 5025 765 5034
rect 727 5005 736 5025
rect 756 5005 765 5025
rect 623 5000 659 5001
rect 727 4997 765 5005
rect 831 5029 975 5035
rect 831 5009 839 5029
rect 859 5028 947 5029
rect 859 5009 887 5028
rect 831 5007 887 5009
rect 909 5009 947 5028
rect 967 5009 975 5029
rect 909 5007 975 5009
rect 831 5001 975 5007
rect 831 5000 867 5001
rect 939 5000 975 5001
rect 1041 5034 1078 5035
rect 1041 5033 1079 5034
rect 1041 5025 1105 5033
rect 1041 5005 1050 5025
rect 1070 5011 1105 5025
rect 1125 5011 1128 5031
rect 1070 5006 1128 5011
rect 1070 5005 1105 5006
rect 307 4968 344 4997
rect 127 4922 165 4963
rect 308 4966 344 4968
rect 520 4966 557 4997
rect 308 4944 557 4966
rect 728 4965 765 4997
rect 1041 4993 1105 5005
rect 1145 4967 1172 5145
rect 1004 4965 1172 4967
rect 728 4939 1172 4965
rect 729 4922 753 4939
rect 1004 4938 1172 4939
rect 127 4904 754 4922
rect 1380 4918 1630 4942
rect 127 4898 165 4904
rect 127 4874 164 4898
rect 127 4850 162 4874
rect 125 4841 162 4850
rect 125 4823 135 4841
rect 153 4823 162 4841
rect 125 4813 162 4823
rect 1380 4847 1417 4918
rect 1532 4857 1563 4858
rect 1380 4827 1389 4847
rect 1409 4827 1417 4847
rect 1380 4817 1417 4827
rect 1476 4847 1563 4857
rect 1476 4827 1485 4847
rect 1505 4827 1563 4847
rect 1476 4818 1563 4827
rect 1476 4817 1513 4818
rect 1532 4765 1563 4818
rect 1593 4847 1630 4918
rect 1801 4923 2194 4943
rect 2214 4923 2217 4943
rect 1801 4918 2217 4923
rect 1801 4917 2142 4918
rect 1745 4857 1776 4858
rect 1593 4827 1602 4847
rect 1622 4827 1630 4847
rect 1593 4817 1630 4827
rect 1689 4850 1776 4857
rect 1689 4847 1750 4850
rect 1689 4827 1698 4847
rect 1718 4830 1750 4847
rect 1771 4830 1776 4850
rect 1718 4827 1776 4830
rect 1689 4820 1776 4827
rect 1801 4847 1838 4917
rect 2104 4916 2141 4917
rect 1953 4857 1989 4858
rect 1801 4827 1810 4847
rect 1830 4827 1838 4847
rect 1689 4818 1745 4820
rect 1689 4817 1726 4818
rect 1801 4817 1838 4827
rect 1897 4847 2045 4857
rect 2145 4854 2241 4856
rect 1897 4827 1906 4847
rect 1926 4827 2016 4847
rect 2036 4827 2045 4847
rect 1897 4818 2045 4827
rect 2103 4847 2241 4854
rect 2103 4827 2112 4847
rect 2132 4827 2241 4847
rect 2103 4818 2241 4827
rect 1897 4817 1934 4818
rect 1953 4766 1989 4818
rect 2008 4817 2045 4818
rect 2104 4817 2141 4818
rect 1424 4764 1465 4765
rect 1316 4757 1465 4764
rect 128 4749 165 4751
rect 128 4748 776 4749
rect 127 4742 776 4748
rect 127 4724 137 4742
rect 155 4728 776 4742
rect 1316 4737 1434 4757
rect 1454 4737 1465 4757
rect 1316 4729 1465 4737
rect 1532 4761 1891 4765
rect 1532 4756 1854 4761
rect 1532 4732 1645 4756
rect 1669 4737 1854 4756
rect 1878 4737 1891 4761
rect 1669 4732 1891 4737
rect 1532 4729 1891 4732
rect 1953 4729 1988 4766
rect 2056 4763 2156 4766
rect 2056 4759 2123 4763
rect 2056 4733 2068 4759
rect 2094 4737 2123 4759
rect 2149 4737 2156 4763
rect 2094 4733 2156 4737
rect 2056 4729 2156 4733
rect 155 4724 165 4728
rect 606 4727 776 4728
rect 127 4714 165 4724
rect 127 4636 162 4714
rect 739 4704 776 4727
rect 1532 4708 1563 4729
rect 1953 4708 1989 4729
rect 1375 4707 1412 4708
rect 123 4627 162 4636
rect 123 4609 133 4627
rect 151 4609 162 4627
rect 123 4603 162 4609
rect 318 4679 568 4703
rect 318 4608 355 4679
rect 470 4618 501 4619
rect 123 4599 160 4603
rect 318 4588 327 4608
rect 347 4588 355 4608
rect 318 4578 355 4588
rect 414 4608 501 4618
rect 414 4588 423 4608
rect 443 4588 501 4608
rect 414 4579 501 4588
rect 414 4578 451 4579
rect 126 4528 163 4537
rect 124 4510 135 4528
rect 153 4510 163 4528
rect 470 4526 501 4579
rect 531 4608 568 4679
rect 739 4684 1132 4704
rect 1152 4684 1155 4704
rect 739 4679 1155 4684
rect 1374 4698 1412 4707
rect 739 4678 1080 4679
rect 1374 4678 1383 4698
rect 1403 4678 1412 4698
rect 683 4618 714 4619
rect 531 4588 540 4608
rect 560 4588 568 4608
rect 531 4578 568 4588
rect 627 4611 714 4618
rect 627 4608 688 4611
rect 627 4588 636 4608
rect 656 4591 688 4608
rect 709 4591 714 4611
rect 656 4588 714 4591
rect 627 4581 714 4588
rect 739 4608 776 4678
rect 1042 4677 1079 4678
rect 1374 4670 1412 4678
rect 1478 4702 1563 4708
rect 1588 4707 1625 4708
rect 1478 4682 1486 4702
rect 1506 4682 1563 4702
rect 1478 4674 1563 4682
rect 1587 4698 1625 4707
rect 1587 4678 1596 4698
rect 1616 4678 1625 4698
rect 1478 4673 1514 4674
rect 1587 4670 1625 4678
rect 1691 4702 1776 4708
rect 1796 4707 1833 4708
rect 1691 4682 1699 4702
rect 1719 4701 1776 4702
rect 1719 4682 1748 4701
rect 1691 4681 1748 4682
rect 1769 4681 1776 4701
rect 1691 4674 1776 4681
rect 1795 4698 1833 4707
rect 1795 4678 1804 4698
rect 1824 4678 1833 4698
rect 1691 4673 1727 4674
rect 1795 4670 1833 4678
rect 1899 4702 2043 4708
rect 1899 4682 1907 4702
rect 1927 4701 2015 4702
rect 1927 4682 1960 4701
rect 1983 4682 2015 4701
rect 2035 4682 2043 4702
rect 1899 4674 2043 4682
rect 1899 4673 1935 4674
rect 2007 4673 2043 4674
rect 2109 4707 2146 4708
rect 2109 4706 2147 4707
rect 2109 4698 2173 4706
rect 2109 4678 2118 4698
rect 2138 4684 2173 4698
rect 2193 4684 2196 4704
rect 2138 4679 2196 4684
rect 2138 4678 2173 4679
rect 1375 4641 1412 4670
rect 1376 4639 1412 4641
rect 1588 4639 1625 4670
rect 891 4618 927 4619
rect 739 4588 748 4608
rect 768 4588 776 4608
rect 627 4579 683 4581
rect 627 4578 664 4579
rect 739 4578 776 4588
rect 835 4608 983 4618
rect 1376 4617 1625 4639
rect 1796 4638 1833 4670
rect 2109 4666 2173 4678
rect 2213 4640 2240 4818
rect 2072 4638 2240 4640
rect 1796 4627 2240 4638
rect 2303 4638 2333 5639
rect 2303 4633 2335 4638
rect 1083 4615 1179 4617
rect 835 4588 844 4608
rect 864 4588 954 4608
rect 974 4588 983 4608
rect 835 4579 983 4588
rect 1041 4608 1179 4615
rect 1796 4612 2242 4627
rect 2072 4611 2242 4612
rect 1041 4588 1050 4608
rect 1070 4588 1179 4608
rect 1041 4579 1179 4588
rect 835 4578 872 4579
rect 891 4527 927 4579
rect 946 4578 983 4579
rect 1042 4578 1079 4579
rect 362 4525 403 4526
rect 124 4361 163 4510
rect 254 4518 403 4525
rect 254 4498 372 4518
rect 392 4498 403 4518
rect 254 4490 403 4498
rect 470 4522 829 4526
rect 470 4517 792 4522
rect 470 4493 583 4517
rect 607 4498 792 4517
rect 816 4498 829 4522
rect 607 4493 829 4498
rect 470 4490 829 4493
rect 891 4490 926 4527
rect 994 4524 1094 4527
rect 994 4520 1061 4524
rect 994 4494 1006 4520
rect 1032 4498 1061 4520
rect 1087 4498 1094 4524
rect 1032 4494 1094 4498
rect 994 4490 1094 4494
rect 470 4469 501 4490
rect 891 4469 927 4490
rect 313 4468 350 4469
rect 312 4459 350 4468
rect 312 4439 321 4459
rect 341 4439 350 4459
rect 312 4431 350 4439
rect 416 4463 501 4469
rect 526 4468 563 4469
rect 416 4443 424 4463
rect 444 4443 501 4463
rect 416 4435 501 4443
rect 525 4459 563 4468
rect 525 4439 534 4459
rect 554 4439 563 4459
rect 416 4434 452 4435
rect 525 4431 563 4439
rect 629 4463 714 4469
rect 734 4468 771 4469
rect 629 4443 637 4463
rect 657 4462 714 4463
rect 657 4443 686 4462
rect 629 4442 686 4443
rect 707 4442 714 4462
rect 629 4435 714 4442
rect 733 4459 771 4468
rect 733 4439 742 4459
rect 762 4439 771 4459
rect 629 4434 665 4435
rect 733 4431 771 4439
rect 837 4464 981 4469
rect 837 4463 902 4464
rect 837 4443 845 4463
rect 865 4443 902 4463
rect 924 4463 981 4464
rect 924 4443 953 4463
rect 973 4443 981 4463
rect 837 4435 981 4443
rect 837 4434 873 4435
rect 945 4434 981 4435
rect 1047 4468 1084 4469
rect 1047 4467 1085 4468
rect 1047 4459 1111 4467
rect 1047 4439 1056 4459
rect 1076 4445 1111 4459
rect 1131 4445 1134 4465
rect 1076 4440 1134 4445
rect 1076 4439 1111 4440
rect 313 4402 350 4431
rect 314 4400 350 4402
rect 526 4400 563 4431
rect 314 4378 563 4400
rect 734 4399 771 4431
rect 1047 4427 1111 4439
rect 1151 4401 1178 4579
rect 1010 4399 1178 4401
rect 734 4373 1178 4399
rect 1330 4498 1580 4522
rect 1330 4427 1367 4498
rect 1482 4437 1513 4438
rect 1330 4407 1339 4427
rect 1359 4407 1367 4427
rect 1330 4397 1367 4407
rect 1426 4427 1513 4437
rect 1426 4407 1435 4427
rect 1455 4407 1513 4427
rect 1426 4398 1513 4407
rect 1426 4397 1463 4398
rect 734 4363 756 4373
rect 1010 4372 1178 4373
rect 694 4361 756 4363
rect 124 4354 756 4361
rect 123 4345 756 4354
rect 1482 4345 1513 4398
rect 1543 4427 1580 4498
rect 1751 4503 2144 4523
rect 2164 4503 2167 4523
rect 1751 4498 2167 4503
rect 1751 4497 2092 4498
rect 1695 4437 1726 4438
rect 1543 4407 1552 4427
rect 1572 4407 1580 4427
rect 1543 4397 1580 4407
rect 1639 4430 1726 4437
rect 1639 4427 1700 4430
rect 1639 4407 1648 4427
rect 1668 4410 1700 4427
rect 1721 4410 1726 4430
rect 1668 4407 1726 4410
rect 1639 4400 1726 4407
rect 1751 4427 1788 4497
rect 2054 4496 2091 4497
rect 1903 4437 1939 4438
rect 1751 4407 1760 4427
rect 1780 4407 1788 4427
rect 1639 4398 1695 4400
rect 1639 4397 1676 4398
rect 1751 4397 1788 4407
rect 1847 4427 1995 4437
rect 2095 4434 2191 4436
rect 1847 4407 1856 4427
rect 1876 4407 1966 4427
rect 1986 4407 1995 4427
rect 1847 4398 1995 4407
rect 2053 4427 2191 4434
rect 2053 4407 2062 4427
rect 2082 4407 2191 4427
rect 2053 4398 2191 4407
rect 1847 4397 1884 4398
rect 1903 4346 1939 4398
rect 1958 4397 1995 4398
rect 2054 4397 2091 4398
rect 123 4327 133 4345
rect 151 4344 756 4345
rect 1374 4344 1415 4345
rect 151 4339 172 4344
rect 151 4327 163 4339
rect 1266 4337 1415 4344
rect 123 4319 163 4327
rect 206 4326 232 4327
rect 123 4317 160 4319
rect 206 4308 760 4326
rect 1266 4317 1384 4337
rect 1404 4317 1415 4337
rect 1266 4309 1415 4317
rect 1482 4341 1841 4345
rect 1482 4336 1804 4341
rect 1482 4312 1595 4336
rect 1619 4317 1804 4336
rect 1828 4317 1841 4341
rect 1619 4312 1841 4317
rect 1482 4309 1841 4312
rect 1903 4309 1938 4346
rect 2006 4343 2106 4346
rect 2006 4339 2073 4343
rect 2006 4313 2018 4339
rect 2044 4317 2073 4339
rect 2099 4317 2106 4343
rect 2044 4313 2106 4317
rect 2006 4309 2106 4313
rect 126 4249 163 4255
rect 206 4249 232 4308
rect 739 4289 760 4308
rect 126 4246 232 4249
rect 126 4228 135 4246
rect 153 4232 232 4246
rect 317 4264 567 4288
rect 153 4230 229 4232
rect 153 4228 163 4230
rect 126 4218 163 4228
rect 131 4153 162 4218
rect 317 4193 354 4264
rect 469 4203 500 4204
rect 317 4173 326 4193
rect 346 4173 354 4193
rect 317 4163 354 4173
rect 413 4193 500 4203
rect 413 4173 422 4193
rect 442 4173 500 4193
rect 413 4164 500 4173
rect 413 4163 450 4164
rect 130 4144 167 4153
rect 130 4126 140 4144
rect 158 4126 167 4144
rect 130 4116 167 4126
rect 469 4111 500 4164
rect 530 4193 567 4264
rect 738 4269 1131 4289
rect 1151 4269 1154 4289
rect 1482 4288 1513 4309
rect 1903 4288 1939 4309
rect 1325 4287 1362 4288
rect 738 4264 1154 4269
rect 1324 4278 1362 4287
rect 738 4263 1079 4264
rect 682 4203 713 4204
rect 530 4173 539 4193
rect 559 4173 567 4193
rect 530 4163 567 4173
rect 626 4196 713 4203
rect 626 4193 687 4196
rect 626 4173 635 4193
rect 655 4176 687 4193
rect 708 4176 713 4196
rect 655 4173 713 4176
rect 626 4166 713 4173
rect 738 4193 775 4263
rect 1041 4262 1078 4263
rect 1324 4258 1333 4278
rect 1353 4258 1362 4278
rect 1324 4250 1362 4258
rect 1428 4282 1513 4288
rect 1538 4287 1575 4288
rect 1428 4262 1436 4282
rect 1456 4262 1513 4282
rect 1428 4254 1513 4262
rect 1537 4278 1575 4287
rect 1537 4258 1546 4278
rect 1566 4258 1575 4278
rect 1428 4253 1464 4254
rect 1537 4250 1575 4258
rect 1641 4282 1726 4288
rect 1746 4287 1783 4288
rect 1641 4262 1649 4282
rect 1669 4281 1726 4282
rect 1669 4262 1698 4281
rect 1641 4261 1698 4262
rect 1719 4261 1726 4281
rect 1641 4254 1726 4261
rect 1745 4278 1783 4287
rect 1745 4258 1754 4278
rect 1774 4258 1783 4278
rect 1641 4253 1677 4254
rect 1745 4250 1783 4258
rect 1849 4283 1993 4288
rect 1849 4282 1908 4283
rect 1849 4262 1857 4282
rect 1877 4263 1908 4282
rect 1932 4282 1993 4283
rect 1932 4263 1965 4282
rect 1877 4262 1965 4263
rect 1985 4262 1993 4282
rect 1849 4254 1993 4262
rect 1849 4253 1885 4254
rect 1957 4253 1993 4254
rect 2059 4287 2096 4288
rect 2059 4286 2097 4287
rect 2059 4278 2123 4286
rect 2059 4258 2068 4278
rect 2088 4264 2123 4278
rect 2143 4264 2146 4284
rect 2088 4259 2146 4264
rect 2088 4258 2123 4259
rect 1325 4221 1362 4250
rect 1326 4219 1362 4221
rect 1538 4219 1575 4250
rect 890 4203 926 4204
rect 738 4173 747 4193
rect 767 4173 775 4193
rect 626 4164 682 4166
rect 626 4163 663 4164
rect 738 4163 775 4173
rect 834 4193 982 4203
rect 1082 4200 1178 4202
rect 834 4173 843 4193
rect 863 4173 953 4193
rect 973 4173 982 4193
rect 834 4164 982 4173
rect 1040 4193 1178 4200
rect 1326 4197 1575 4219
rect 1746 4218 1783 4250
rect 2059 4246 2123 4258
rect 2163 4220 2190 4398
rect 2022 4218 2190 4220
rect 1746 4214 2190 4218
rect 1040 4173 1049 4193
rect 1069 4173 1178 4193
rect 1746 4195 1795 4214
rect 1815 4195 2190 4214
rect 1746 4192 2190 4195
rect 2022 4191 2190 4192
rect 2211 4217 2242 4611
rect 2303 4615 2308 4633
rect 2328 4615 2335 4633
rect 2303 4610 2335 4615
rect 2306 4608 2335 4610
rect 2211 4191 2216 4217
rect 2235 4191 2242 4217
rect 2749 4192 2787 6023
rect 2815 5910 2842 6088
rect 2882 6050 2946 6062
rect 3222 6058 3259 6090
rect 3430 6089 3679 6111
rect 4134 6097 4171 6098
rect 4437 6097 4474 6167
rect 4499 6187 4586 6194
rect 4499 6184 4557 6187
rect 4499 6164 4504 6184
rect 4525 6167 4557 6184
rect 4577 6167 4586 6187
rect 4525 6164 4586 6167
rect 4499 6157 4586 6164
rect 4645 6187 4682 6197
rect 4645 6167 4653 6187
rect 4673 6167 4682 6187
rect 4499 6156 4530 6157
rect 4133 6096 4474 6097
rect 3430 6058 3467 6089
rect 3643 6087 3679 6089
rect 4058 6091 4474 6096
rect 3643 6058 3680 6087
rect 4058 6071 4061 6091
rect 4081 6071 4474 6091
rect 4645 6096 4682 6167
rect 4712 6196 4743 6249
rect 5050 6247 5060 6265
rect 5078 6247 5089 6265
rect 5050 6238 5087 6247
rect 4762 6196 4799 6197
rect 4712 6187 4799 6196
rect 4712 6167 4770 6187
rect 4790 6167 4799 6187
rect 4712 6157 4799 6167
rect 4858 6187 4895 6197
rect 4858 6167 4866 6187
rect 4886 6167 4895 6187
rect 5053 6172 5090 6176
rect 4712 6156 4743 6157
rect 4858 6096 4895 6167
rect 4645 6072 4895 6096
rect 5051 6166 5090 6172
rect 5051 6148 5062 6166
rect 5080 6148 5090 6166
rect 5051 6139 5090 6148
rect 2882 6049 2917 6050
rect 2859 6044 2917 6049
rect 2859 6024 2862 6044
rect 2882 6030 2917 6044
rect 2937 6030 2946 6050
rect 2882 6022 2946 6030
rect 2908 6021 2946 6022
rect 2909 6020 2946 6021
rect 3012 6054 3048 6055
rect 3120 6054 3156 6055
rect 3012 6046 3156 6054
rect 3012 6026 3020 6046
rect 3040 6045 3128 6046
rect 3040 6026 3069 6045
rect 3092 6026 3128 6045
rect 3148 6026 3156 6046
rect 3012 6020 3156 6026
rect 3222 6050 3260 6058
rect 3328 6054 3364 6055
rect 3222 6030 3231 6050
rect 3251 6030 3260 6050
rect 3222 6021 3260 6030
rect 3279 6047 3364 6054
rect 3279 6027 3286 6047
rect 3307 6046 3364 6047
rect 3307 6027 3336 6046
rect 3279 6026 3336 6027
rect 3356 6026 3364 6046
rect 3222 6020 3259 6021
rect 3279 6020 3364 6026
rect 3430 6050 3468 6058
rect 3541 6054 3577 6055
rect 3430 6030 3439 6050
rect 3459 6030 3468 6050
rect 3430 6021 3468 6030
rect 3492 6046 3577 6054
rect 3492 6026 3549 6046
rect 3569 6026 3577 6046
rect 3430 6020 3467 6021
rect 3492 6020 3577 6026
rect 3643 6050 3681 6058
rect 3643 6030 3652 6050
rect 3672 6030 3681 6050
rect 3643 6021 3681 6030
rect 4437 6048 4474 6071
rect 5051 6061 5086 6139
rect 5048 6051 5086 6061
rect 4437 6047 4607 6048
rect 5048 6047 5058 6051
rect 4437 6033 5058 6047
rect 5076 6033 5086 6051
rect 4437 6027 5086 6033
rect 4437 6026 5085 6027
rect 5048 6024 5085 6026
rect 3643 6020 3680 6021
rect 3066 5999 3102 6020
rect 3492 5999 3523 6020
rect 2899 5995 2999 5999
rect 2899 5991 2961 5995
rect 2899 5965 2906 5991
rect 2932 5969 2961 5991
rect 2987 5969 2999 5995
rect 2932 5965 2999 5969
rect 2899 5962 2999 5965
rect 3067 5962 3102 5999
rect 3164 5996 3523 5999
rect 3164 5991 3386 5996
rect 3164 5967 3177 5991
rect 3201 5972 3386 5991
rect 3410 5972 3523 5996
rect 3201 5967 3523 5972
rect 3164 5963 3523 5967
rect 3590 5991 3739 5999
rect 3590 5971 3601 5991
rect 3621 5971 3739 5991
rect 3590 5964 3739 5971
rect 3590 5963 3631 5964
rect 2914 5910 2951 5911
rect 3010 5910 3047 5911
rect 3066 5910 3102 5962
rect 3121 5910 3158 5911
rect 2814 5901 2952 5910
rect 2814 5881 2923 5901
rect 2943 5881 2952 5901
rect 2814 5874 2952 5881
rect 3010 5901 3158 5910
rect 3010 5881 3019 5901
rect 3039 5881 3129 5901
rect 3149 5881 3158 5901
rect 2814 5872 2910 5874
rect 3010 5871 3158 5881
rect 3217 5901 3254 5911
rect 3329 5910 3366 5911
rect 3310 5908 3366 5910
rect 3217 5881 3225 5901
rect 3245 5881 3254 5901
rect 3066 5870 3102 5871
rect 2914 5811 2951 5812
rect 3217 5811 3254 5881
rect 3279 5901 3366 5908
rect 3279 5898 3337 5901
rect 3279 5878 3284 5898
rect 3305 5881 3337 5898
rect 3357 5881 3366 5901
rect 3305 5878 3366 5881
rect 3279 5871 3366 5878
rect 3425 5901 3462 5911
rect 3425 5881 3433 5901
rect 3453 5881 3462 5901
rect 3279 5870 3310 5871
rect 2913 5810 3254 5811
rect 2838 5805 3254 5810
rect 2838 5785 2841 5805
rect 2861 5785 3254 5805
rect 3425 5810 3462 5881
rect 3492 5910 3523 5963
rect 5051 5952 5088 5962
rect 5051 5934 5060 5952
rect 5078 5934 5088 5952
rect 5051 5925 5088 5934
rect 3542 5910 3579 5911
rect 3492 5901 3579 5910
rect 3492 5881 3550 5901
rect 3570 5881 3579 5901
rect 3492 5871 3579 5881
rect 3638 5901 3675 5911
rect 3638 5881 3646 5901
rect 3666 5881 3675 5901
rect 3492 5870 3523 5871
rect 3638 5810 3675 5881
rect 5051 5879 5086 5925
rect 5050 5873 5088 5879
rect 4461 5855 5088 5873
rect 3425 5786 3675 5810
rect 4043 5838 4211 5839
rect 4462 5838 4486 5855
rect 4043 5812 4487 5838
rect 4043 5810 4211 5812
rect 4043 5632 4070 5810
rect 4110 5772 4174 5784
rect 4450 5780 4487 5812
rect 4658 5811 4907 5833
rect 4658 5780 4695 5811
rect 4871 5809 4907 5811
rect 5050 5814 5088 5855
rect 4871 5780 4908 5809
rect 4110 5771 4145 5772
rect 4087 5766 4145 5771
rect 4087 5746 4090 5766
rect 4110 5752 4145 5766
rect 4165 5752 4174 5772
rect 4110 5744 4174 5752
rect 4136 5743 4174 5744
rect 4137 5742 4174 5743
rect 4240 5776 4276 5777
rect 4348 5776 4384 5777
rect 4240 5770 4384 5776
rect 4240 5768 4306 5770
rect 4240 5748 4248 5768
rect 4268 5749 4306 5768
rect 4328 5768 4384 5770
rect 4328 5749 4356 5768
rect 4268 5748 4356 5749
rect 4376 5748 4384 5768
rect 4240 5742 4384 5748
rect 4450 5772 4488 5780
rect 4556 5776 4592 5777
rect 4450 5752 4459 5772
rect 4479 5752 4488 5772
rect 4450 5743 4488 5752
rect 4507 5769 4592 5776
rect 4507 5749 4514 5769
rect 4535 5768 4592 5769
rect 4535 5749 4564 5768
rect 4507 5748 4564 5749
rect 4584 5748 4592 5768
rect 4450 5742 4487 5743
rect 4507 5742 4592 5748
rect 4658 5772 4696 5780
rect 4769 5776 4805 5777
rect 4658 5752 4667 5772
rect 4687 5752 4696 5772
rect 4658 5743 4696 5752
rect 4720 5768 4805 5776
rect 4720 5748 4777 5768
rect 4797 5748 4805 5768
rect 4658 5742 4695 5743
rect 4720 5742 4805 5748
rect 4871 5772 4909 5780
rect 4871 5752 4880 5772
rect 4900 5752 4909 5772
rect 4871 5743 4909 5752
rect 5050 5779 5086 5814
rect 5050 5769 5087 5779
rect 5050 5751 5060 5769
rect 5078 5751 5087 5769
rect 4871 5742 4908 5743
rect 5050 5742 5087 5751
rect 4294 5721 4330 5742
rect 4720 5721 4751 5742
rect 4127 5717 4227 5721
rect 4127 5713 4189 5717
rect 4127 5687 4134 5713
rect 4160 5691 4189 5713
rect 4215 5691 4227 5717
rect 4160 5687 4227 5691
rect 4127 5684 4227 5687
rect 4295 5684 4330 5721
rect 4392 5718 4751 5721
rect 4392 5713 4614 5718
rect 4392 5689 4405 5713
rect 4429 5694 4614 5713
rect 4638 5694 4751 5718
rect 4429 5689 4751 5694
rect 4392 5685 4751 5689
rect 4818 5713 4967 5721
rect 4818 5693 4829 5713
rect 4849 5693 4967 5713
rect 4818 5686 4967 5693
rect 4818 5685 4859 5686
rect 4142 5632 4179 5633
rect 4238 5632 4275 5633
rect 4294 5632 4330 5684
rect 4349 5632 4386 5633
rect 4042 5623 4180 5632
rect 2978 5605 3009 5608
rect 2978 5579 2985 5605
rect 3004 5579 3009 5605
rect 2978 5185 3009 5579
rect 3030 5604 3198 5605
rect 3030 5601 3474 5604
rect 3030 5582 3405 5601
rect 3425 5582 3474 5601
rect 4042 5603 4151 5623
rect 4171 5603 4180 5623
rect 3030 5578 3474 5582
rect 3030 5576 3198 5578
rect 3030 5398 3057 5576
rect 3097 5538 3161 5550
rect 3437 5546 3474 5578
rect 3645 5577 3894 5599
rect 4042 5596 4180 5603
rect 4238 5623 4386 5632
rect 4238 5603 4247 5623
rect 4267 5603 4357 5623
rect 4377 5603 4386 5623
rect 4042 5594 4138 5596
rect 4238 5593 4386 5603
rect 4445 5623 4482 5633
rect 4557 5632 4594 5633
rect 4538 5630 4594 5632
rect 4445 5603 4453 5623
rect 4473 5603 4482 5623
rect 4294 5592 4330 5593
rect 3645 5546 3682 5577
rect 3858 5575 3894 5577
rect 3858 5546 3895 5575
rect 3097 5537 3132 5538
rect 3074 5532 3132 5537
rect 3074 5512 3077 5532
rect 3097 5518 3132 5532
rect 3152 5518 3161 5538
rect 3097 5510 3161 5518
rect 3123 5509 3161 5510
rect 3124 5508 3161 5509
rect 3227 5542 3263 5543
rect 3335 5542 3371 5543
rect 3227 5534 3371 5542
rect 3227 5514 3235 5534
rect 3255 5533 3343 5534
rect 3255 5514 3288 5533
rect 3227 5513 3288 5514
rect 3312 5514 3343 5533
rect 3363 5514 3371 5534
rect 3312 5513 3371 5514
rect 3227 5508 3371 5513
rect 3437 5538 3475 5546
rect 3543 5542 3579 5543
rect 3437 5518 3446 5538
rect 3466 5518 3475 5538
rect 3437 5509 3475 5518
rect 3494 5535 3579 5542
rect 3494 5515 3501 5535
rect 3522 5534 3579 5535
rect 3522 5515 3551 5534
rect 3494 5514 3551 5515
rect 3571 5514 3579 5534
rect 3437 5508 3474 5509
rect 3494 5508 3579 5514
rect 3645 5538 3683 5546
rect 3756 5542 3792 5543
rect 3645 5518 3654 5538
rect 3674 5518 3683 5538
rect 3645 5509 3683 5518
rect 3707 5534 3792 5542
rect 3707 5514 3764 5534
rect 3784 5514 3792 5534
rect 3645 5508 3682 5509
rect 3707 5508 3792 5514
rect 3858 5538 3896 5546
rect 3858 5518 3867 5538
rect 3887 5518 3896 5538
rect 4142 5533 4179 5534
rect 4445 5533 4482 5603
rect 4507 5623 4594 5630
rect 4507 5620 4565 5623
rect 4507 5600 4512 5620
rect 4533 5603 4565 5620
rect 4585 5603 4594 5623
rect 4533 5600 4594 5603
rect 4507 5593 4594 5600
rect 4653 5623 4690 5633
rect 4653 5603 4661 5623
rect 4681 5603 4690 5623
rect 4507 5592 4538 5593
rect 4141 5532 4482 5533
rect 3858 5509 3896 5518
rect 4066 5527 4482 5532
rect 3858 5508 3895 5509
rect 3281 5487 3317 5508
rect 3707 5487 3738 5508
rect 4066 5507 4069 5527
rect 4089 5507 4482 5527
rect 4653 5532 4690 5603
rect 4720 5632 4751 5685
rect 5053 5670 5090 5680
rect 5053 5652 5062 5670
rect 5080 5652 5090 5670
rect 5053 5643 5090 5652
rect 4770 5632 4807 5633
rect 4720 5623 4807 5632
rect 4720 5603 4778 5623
rect 4798 5603 4807 5623
rect 4720 5593 4807 5603
rect 4866 5623 4903 5633
rect 4866 5603 4874 5623
rect 4894 5603 4903 5623
rect 4720 5592 4751 5593
rect 4866 5532 4903 5603
rect 5058 5578 5089 5643
rect 5057 5568 5094 5578
rect 5057 5566 5067 5568
rect 4991 5564 5067 5566
rect 4653 5508 4903 5532
rect 4988 5550 5067 5564
rect 5085 5550 5094 5568
rect 4988 5547 5094 5550
rect 4460 5488 4481 5507
rect 4988 5488 5014 5547
rect 5057 5541 5094 5547
rect 3114 5483 3214 5487
rect 3114 5479 3176 5483
rect 3114 5453 3121 5479
rect 3147 5457 3176 5479
rect 3202 5457 3214 5483
rect 3147 5453 3214 5457
rect 3114 5450 3214 5453
rect 3282 5450 3317 5487
rect 3379 5484 3738 5487
rect 3379 5479 3601 5484
rect 3379 5455 3392 5479
rect 3416 5460 3601 5479
rect 3625 5460 3738 5484
rect 3416 5455 3738 5460
rect 3379 5451 3738 5455
rect 3805 5479 3954 5487
rect 3805 5459 3816 5479
rect 3836 5459 3954 5479
rect 4460 5470 5014 5488
rect 5060 5477 5097 5479
rect 4988 5469 5014 5470
rect 5057 5469 5097 5477
rect 3805 5452 3954 5459
rect 5057 5457 5069 5469
rect 5048 5452 5069 5457
rect 3805 5451 3846 5452
rect 4464 5451 5069 5452
rect 5087 5451 5097 5469
rect 3129 5398 3166 5399
rect 3225 5398 3262 5399
rect 3281 5398 3317 5450
rect 3336 5398 3373 5399
rect 3029 5389 3167 5398
rect 3029 5369 3138 5389
rect 3158 5369 3167 5389
rect 3029 5362 3167 5369
rect 3225 5389 3373 5398
rect 3225 5369 3234 5389
rect 3254 5369 3344 5389
rect 3364 5369 3373 5389
rect 3029 5360 3125 5362
rect 3225 5359 3373 5369
rect 3432 5389 3469 5399
rect 3544 5398 3581 5399
rect 3525 5396 3581 5398
rect 3432 5369 3440 5389
rect 3460 5369 3469 5389
rect 3281 5358 3317 5359
rect 3129 5299 3166 5300
rect 3432 5299 3469 5369
rect 3494 5389 3581 5396
rect 3494 5386 3552 5389
rect 3494 5366 3499 5386
rect 3520 5369 3552 5386
rect 3572 5369 3581 5389
rect 3520 5366 3581 5369
rect 3494 5359 3581 5366
rect 3640 5389 3677 5399
rect 3640 5369 3648 5389
rect 3668 5369 3677 5389
rect 3494 5358 3525 5359
rect 3128 5298 3469 5299
rect 3053 5293 3469 5298
rect 3053 5273 3056 5293
rect 3076 5273 3469 5293
rect 3640 5298 3677 5369
rect 3707 5398 3738 5451
rect 4464 5442 5097 5451
rect 4464 5435 5096 5442
rect 4464 5433 4526 5435
rect 4042 5423 4210 5424
rect 4464 5423 4486 5433
rect 3757 5398 3794 5399
rect 3707 5389 3794 5398
rect 3707 5369 3765 5389
rect 3785 5369 3794 5389
rect 3707 5359 3794 5369
rect 3853 5389 3890 5399
rect 3853 5369 3861 5389
rect 3881 5369 3890 5389
rect 3707 5358 3738 5359
rect 3853 5298 3890 5369
rect 3640 5274 3890 5298
rect 4042 5397 4486 5423
rect 4042 5395 4210 5397
rect 4042 5217 4069 5395
rect 4109 5357 4173 5369
rect 4449 5365 4486 5397
rect 4657 5396 4906 5418
rect 4657 5365 4694 5396
rect 4870 5394 4906 5396
rect 4870 5365 4907 5394
rect 4109 5356 4144 5357
rect 4086 5351 4144 5356
rect 4086 5331 4089 5351
rect 4109 5337 4144 5351
rect 4164 5337 4173 5357
rect 4109 5329 4173 5337
rect 4135 5328 4173 5329
rect 4136 5327 4173 5328
rect 4239 5361 4275 5362
rect 4347 5361 4383 5362
rect 4239 5353 4383 5361
rect 4239 5333 4247 5353
rect 4267 5333 4296 5353
rect 4239 5332 4296 5333
rect 4318 5333 4355 5353
rect 4375 5333 4383 5353
rect 4318 5332 4383 5333
rect 4239 5327 4383 5332
rect 4449 5357 4487 5365
rect 4555 5361 4591 5362
rect 4449 5337 4458 5357
rect 4478 5337 4487 5357
rect 4449 5328 4487 5337
rect 4506 5354 4591 5361
rect 4506 5334 4513 5354
rect 4534 5353 4591 5354
rect 4534 5334 4563 5353
rect 4506 5333 4563 5334
rect 4583 5333 4591 5353
rect 4449 5327 4486 5328
rect 4506 5327 4591 5333
rect 4657 5357 4695 5365
rect 4768 5361 4804 5362
rect 4657 5337 4666 5357
rect 4686 5337 4695 5357
rect 4657 5328 4695 5337
rect 4719 5353 4804 5361
rect 4719 5333 4776 5353
rect 4796 5333 4804 5353
rect 4657 5327 4694 5328
rect 4719 5327 4804 5333
rect 4870 5357 4908 5365
rect 4870 5337 4879 5357
rect 4899 5337 4908 5357
rect 4870 5328 4908 5337
rect 4870 5327 4907 5328
rect 4293 5306 4329 5327
rect 4719 5306 4750 5327
rect 4126 5302 4226 5306
rect 4126 5298 4188 5302
rect 4126 5272 4133 5298
rect 4159 5276 4188 5298
rect 4214 5276 4226 5302
rect 4159 5272 4226 5276
rect 4126 5269 4226 5272
rect 4294 5269 4329 5306
rect 4391 5303 4750 5306
rect 4391 5298 4613 5303
rect 4391 5274 4404 5298
rect 4428 5279 4613 5298
rect 4637 5279 4750 5303
rect 4428 5274 4750 5279
rect 4391 5270 4750 5274
rect 4817 5298 4966 5306
rect 4817 5278 4828 5298
rect 4848 5278 4966 5298
rect 4817 5271 4966 5278
rect 5057 5286 5096 5435
rect 4817 5270 4858 5271
rect 4141 5217 4178 5218
rect 4237 5217 4274 5218
rect 4293 5217 4329 5269
rect 4348 5217 4385 5218
rect 4041 5208 4179 5217
rect 4041 5188 4150 5208
rect 4170 5188 4179 5208
rect 2978 5184 3148 5185
rect 2978 5169 3424 5184
rect 4041 5181 4179 5188
rect 4237 5208 4385 5217
rect 4237 5188 4246 5208
rect 4266 5188 4356 5208
rect 4376 5188 4385 5208
rect 4041 5179 4137 5181
rect 2980 5158 3424 5169
rect 2980 5156 3148 5158
rect 2980 4978 3007 5156
rect 3047 5118 3111 5130
rect 3387 5126 3424 5158
rect 3595 5157 3844 5179
rect 4237 5178 4385 5188
rect 4444 5208 4481 5218
rect 4556 5217 4593 5218
rect 4537 5215 4593 5217
rect 4444 5188 4452 5208
rect 4472 5188 4481 5208
rect 4293 5177 4329 5178
rect 3595 5126 3632 5157
rect 3808 5155 3844 5157
rect 3808 5126 3845 5155
rect 3047 5117 3082 5118
rect 3024 5112 3082 5117
rect 3024 5092 3027 5112
rect 3047 5098 3082 5112
rect 3102 5098 3111 5118
rect 3047 5090 3111 5098
rect 3073 5089 3111 5090
rect 3074 5088 3111 5089
rect 3177 5122 3213 5123
rect 3285 5122 3321 5123
rect 3177 5114 3321 5122
rect 3177 5094 3185 5114
rect 3205 5113 3293 5114
rect 3205 5096 3233 5113
rect 3257 5096 3293 5113
rect 3205 5094 3293 5096
rect 3313 5094 3321 5114
rect 3177 5088 3321 5094
rect 3387 5118 3425 5126
rect 3493 5122 3529 5123
rect 3387 5098 3396 5118
rect 3416 5098 3425 5118
rect 3387 5089 3425 5098
rect 3444 5115 3529 5122
rect 3444 5095 3451 5115
rect 3472 5114 3529 5115
rect 3472 5095 3501 5114
rect 3444 5094 3501 5095
rect 3521 5094 3529 5114
rect 3387 5088 3424 5089
rect 3444 5088 3529 5094
rect 3595 5118 3633 5126
rect 3706 5122 3742 5123
rect 3595 5098 3604 5118
rect 3624 5098 3633 5118
rect 3595 5089 3633 5098
rect 3657 5114 3742 5122
rect 3657 5094 3714 5114
rect 3734 5094 3742 5114
rect 3595 5088 3632 5089
rect 3657 5088 3742 5094
rect 3808 5118 3846 5126
rect 4141 5118 4178 5119
rect 4444 5118 4481 5188
rect 4506 5208 4593 5215
rect 4506 5205 4564 5208
rect 4506 5185 4511 5205
rect 4532 5188 4564 5205
rect 4584 5188 4593 5208
rect 4532 5185 4593 5188
rect 4506 5178 4593 5185
rect 4652 5208 4689 5218
rect 4652 5188 4660 5208
rect 4680 5188 4689 5208
rect 4506 5177 4537 5178
rect 3808 5098 3817 5118
rect 3837 5098 3846 5118
rect 4140 5117 4481 5118
rect 3808 5089 3846 5098
rect 4065 5112 4481 5117
rect 4065 5092 4068 5112
rect 4088 5092 4481 5112
rect 4652 5117 4689 5188
rect 4719 5217 4750 5270
rect 5057 5268 5067 5286
rect 5085 5268 5096 5286
rect 5057 5259 5094 5268
rect 4769 5217 4806 5218
rect 4719 5208 4806 5217
rect 4719 5188 4777 5208
rect 4797 5188 4806 5208
rect 4719 5178 4806 5188
rect 4865 5208 4902 5218
rect 4865 5188 4873 5208
rect 4893 5188 4902 5208
rect 5060 5193 5097 5197
rect 4719 5177 4750 5178
rect 4865 5117 4902 5188
rect 4652 5093 4902 5117
rect 5058 5187 5097 5193
rect 5058 5169 5069 5187
rect 5087 5169 5097 5187
rect 5058 5160 5097 5169
rect 3808 5088 3845 5089
rect 3231 5067 3267 5088
rect 3657 5067 3688 5088
rect 4444 5069 4481 5092
rect 5058 5082 5093 5160
rect 5055 5072 5093 5082
rect 4444 5068 4614 5069
rect 5055 5068 5065 5072
rect 3064 5063 3164 5067
rect 3064 5059 3126 5063
rect 3064 5033 3071 5059
rect 3097 5037 3126 5059
rect 3152 5037 3164 5063
rect 3097 5033 3164 5037
rect 3064 5030 3164 5033
rect 3232 5030 3267 5067
rect 3329 5064 3688 5067
rect 3329 5059 3551 5064
rect 3329 5035 3342 5059
rect 3366 5040 3551 5059
rect 3575 5040 3688 5064
rect 3366 5035 3688 5040
rect 3329 5031 3688 5035
rect 3755 5059 3904 5067
rect 3755 5039 3766 5059
rect 3786 5039 3904 5059
rect 4444 5054 5065 5068
rect 5083 5054 5093 5072
rect 4444 5048 5093 5054
rect 4444 5047 5092 5048
rect 5055 5045 5092 5047
rect 3755 5032 3904 5039
rect 3755 5031 3796 5032
rect 3079 4978 3116 4979
rect 3175 4978 3212 4979
rect 3231 4978 3267 5030
rect 3286 4978 3323 4979
rect 2979 4969 3117 4978
rect 2979 4949 3088 4969
rect 3108 4949 3117 4969
rect 2979 4942 3117 4949
rect 3175 4969 3323 4978
rect 3175 4949 3184 4969
rect 3204 4949 3294 4969
rect 3314 4949 3323 4969
rect 2979 4940 3075 4942
rect 3175 4939 3323 4949
rect 3382 4969 3419 4979
rect 3494 4978 3531 4979
rect 3475 4976 3531 4978
rect 3382 4949 3390 4969
rect 3410 4949 3419 4969
rect 3231 4938 3267 4939
rect 3079 4879 3116 4880
rect 3382 4879 3419 4949
rect 3444 4969 3531 4976
rect 3444 4966 3502 4969
rect 3444 4946 3449 4966
rect 3470 4949 3502 4966
rect 3522 4949 3531 4969
rect 3470 4946 3531 4949
rect 3444 4939 3531 4946
rect 3590 4969 3627 4979
rect 3590 4949 3598 4969
rect 3618 4949 3627 4969
rect 3444 4938 3475 4939
rect 3078 4878 3419 4879
rect 3003 4873 3419 4878
rect 3003 4853 3006 4873
rect 3026 4853 3419 4873
rect 3590 4878 3627 4949
rect 3657 4978 3688 5031
rect 3707 4978 3744 4979
rect 3657 4969 3744 4978
rect 3657 4949 3715 4969
rect 3735 4949 3744 4969
rect 3657 4939 3744 4949
rect 3803 4969 3840 4979
rect 3803 4949 3811 4969
rect 3831 4949 3840 4969
rect 3657 4938 3688 4939
rect 3803 4878 3840 4949
rect 5058 4973 5095 4983
rect 5058 4955 5067 4973
rect 5085 4955 5095 4973
rect 5058 4946 5095 4955
rect 5058 4922 5093 4946
rect 5056 4898 5093 4922
rect 5055 4892 5093 4898
rect 3590 4854 3840 4878
rect 4466 4874 5093 4892
rect 4048 4857 4216 4858
rect 4467 4857 4491 4874
rect 4048 4831 4492 4857
rect 4048 4829 4216 4831
rect 4048 4651 4075 4829
rect 4115 4791 4179 4803
rect 4455 4799 4492 4831
rect 4663 4830 4912 4852
rect 4663 4799 4700 4830
rect 4876 4828 4912 4830
rect 5055 4833 5093 4874
rect 4876 4799 4913 4828
rect 4115 4790 4150 4791
rect 4092 4785 4150 4790
rect 4092 4765 4095 4785
rect 4115 4771 4150 4785
rect 4170 4771 4179 4791
rect 4115 4763 4179 4771
rect 4141 4762 4179 4763
rect 4142 4761 4179 4762
rect 4245 4795 4281 4796
rect 4353 4795 4389 4796
rect 4245 4789 4389 4795
rect 4245 4787 4311 4789
rect 4245 4767 4253 4787
rect 4273 4768 4311 4787
rect 4333 4787 4389 4789
rect 4333 4768 4361 4787
rect 4273 4767 4361 4768
rect 4381 4767 4389 4787
rect 4245 4761 4389 4767
rect 4455 4791 4493 4799
rect 4561 4795 4597 4796
rect 4455 4771 4464 4791
rect 4484 4771 4493 4791
rect 4455 4762 4493 4771
rect 4512 4788 4597 4795
rect 4512 4768 4519 4788
rect 4540 4787 4597 4788
rect 4540 4768 4569 4787
rect 4512 4767 4569 4768
rect 4589 4767 4597 4787
rect 4455 4761 4492 4762
rect 4512 4761 4597 4767
rect 4663 4791 4701 4799
rect 4774 4795 4810 4796
rect 4663 4771 4672 4791
rect 4692 4771 4701 4791
rect 4663 4762 4701 4771
rect 4725 4787 4810 4795
rect 4725 4767 4782 4787
rect 4802 4767 4810 4787
rect 4663 4761 4700 4762
rect 4725 4761 4810 4767
rect 4876 4791 4914 4799
rect 4876 4771 4885 4791
rect 4905 4771 4914 4791
rect 4876 4762 4914 4771
rect 5055 4798 5091 4833
rect 5055 4788 5092 4798
rect 5055 4770 5065 4788
rect 5083 4770 5092 4788
rect 4876 4761 4913 4762
rect 5055 4761 5092 4770
rect 4299 4740 4335 4761
rect 4725 4740 4756 4761
rect 4132 4736 4232 4740
rect 4132 4732 4194 4736
rect 4132 4706 4139 4732
rect 4165 4710 4194 4732
rect 4220 4710 4232 4736
rect 4165 4706 4232 4710
rect 4132 4703 4232 4706
rect 4300 4703 4335 4740
rect 4397 4737 4756 4740
rect 4397 4732 4619 4737
rect 4397 4708 4410 4732
rect 4434 4713 4619 4732
rect 4643 4713 4756 4737
rect 4434 4708 4756 4713
rect 4397 4704 4756 4708
rect 4823 4732 4972 4740
rect 4823 4712 4834 4732
rect 4854 4712 4972 4732
rect 4823 4705 4972 4712
rect 4823 4704 4864 4705
rect 4147 4651 4184 4652
rect 4243 4651 4280 4652
rect 4299 4651 4335 4703
rect 4354 4651 4391 4652
rect 4047 4642 4185 4651
rect 3035 4623 3203 4624
rect 3035 4620 3479 4623
rect 3035 4601 3410 4620
rect 3430 4601 3479 4620
rect 4047 4622 4156 4642
rect 4176 4622 4185 4642
rect 3035 4597 3479 4601
rect 3035 4595 3203 4597
rect 3035 4417 3062 4595
rect 3102 4557 3166 4569
rect 3442 4565 3479 4597
rect 3650 4596 3899 4618
rect 4047 4615 4185 4622
rect 4243 4642 4391 4651
rect 4243 4622 4252 4642
rect 4272 4622 4362 4642
rect 4382 4622 4391 4642
rect 4047 4613 4143 4615
rect 4243 4612 4391 4622
rect 4450 4642 4487 4652
rect 4562 4651 4599 4652
rect 4543 4649 4599 4651
rect 4450 4622 4458 4642
rect 4478 4622 4487 4642
rect 4299 4611 4335 4612
rect 3650 4565 3687 4596
rect 3863 4594 3899 4596
rect 3863 4565 3900 4594
rect 3102 4556 3137 4557
rect 3079 4551 3137 4556
rect 3079 4531 3082 4551
rect 3102 4537 3137 4551
rect 3157 4537 3166 4557
rect 3102 4529 3166 4537
rect 3128 4528 3166 4529
rect 3129 4527 3166 4528
rect 3232 4561 3268 4562
rect 3340 4561 3376 4562
rect 3232 4553 3376 4561
rect 3232 4533 3240 4553
rect 3260 4533 3292 4553
rect 3316 4533 3348 4553
rect 3368 4533 3376 4553
rect 3232 4527 3376 4533
rect 3442 4557 3480 4565
rect 3548 4561 3584 4562
rect 3442 4537 3451 4557
rect 3471 4537 3480 4557
rect 3442 4528 3480 4537
rect 3499 4554 3584 4561
rect 3499 4534 3506 4554
rect 3527 4553 3584 4554
rect 3527 4534 3556 4553
rect 3499 4533 3556 4534
rect 3576 4533 3584 4553
rect 3442 4527 3479 4528
rect 3499 4527 3584 4533
rect 3650 4557 3688 4565
rect 3761 4561 3797 4562
rect 3650 4537 3659 4557
rect 3679 4537 3688 4557
rect 3650 4528 3688 4537
rect 3712 4553 3797 4561
rect 3712 4533 3769 4553
rect 3789 4533 3797 4553
rect 3650 4527 3687 4528
rect 3712 4527 3797 4533
rect 3863 4557 3901 4565
rect 3863 4537 3872 4557
rect 3892 4537 3901 4557
rect 4147 4552 4184 4553
rect 4450 4552 4487 4622
rect 4512 4642 4599 4649
rect 4512 4639 4570 4642
rect 4512 4619 4517 4639
rect 4538 4622 4570 4639
rect 4590 4622 4599 4642
rect 4538 4619 4599 4622
rect 4512 4612 4599 4619
rect 4658 4642 4695 4652
rect 4658 4622 4666 4642
rect 4686 4622 4695 4642
rect 4512 4611 4543 4612
rect 4146 4551 4487 4552
rect 3863 4528 3901 4537
rect 4071 4546 4487 4551
rect 3863 4527 3900 4528
rect 3286 4506 3322 4527
rect 3712 4506 3743 4527
rect 4071 4526 4074 4546
rect 4094 4526 4487 4546
rect 4658 4551 4695 4622
rect 4725 4651 4756 4704
rect 5058 4689 5095 4699
rect 5058 4671 5067 4689
rect 5085 4671 5095 4689
rect 5058 4662 5095 4671
rect 4775 4651 4812 4652
rect 4725 4642 4812 4651
rect 4725 4622 4783 4642
rect 4803 4622 4812 4642
rect 4725 4612 4812 4622
rect 4871 4642 4908 4652
rect 4871 4622 4879 4642
rect 4899 4622 4908 4642
rect 4725 4611 4756 4612
rect 4871 4551 4908 4622
rect 5063 4597 5094 4662
rect 5062 4587 5099 4597
rect 5062 4585 5072 4587
rect 4996 4583 5072 4585
rect 4658 4527 4908 4551
rect 4993 4569 5072 4583
rect 5090 4569 5099 4587
rect 4993 4566 5099 4569
rect 4465 4507 4486 4526
rect 4993 4507 5019 4566
rect 5062 4560 5099 4566
rect 3119 4502 3219 4506
rect 3119 4498 3181 4502
rect 3119 4472 3126 4498
rect 3152 4476 3181 4498
rect 3207 4476 3219 4502
rect 3152 4472 3219 4476
rect 3119 4469 3219 4472
rect 3287 4469 3322 4506
rect 3384 4503 3743 4506
rect 3384 4498 3606 4503
rect 3384 4474 3397 4498
rect 3421 4479 3606 4498
rect 3630 4479 3743 4503
rect 3421 4474 3743 4479
rect 3384 4470 3743 4474
rect 3810 4498 3959 4506
rect 3810 4478 3821 4498
rect 3841 4478 3959 4498
rect 4465 4489 5019 4507
rect 5065 4496 5102 4498
rect 4993 4488 5019 4489
rect 5062 4488 5102 4496
rect 3810 4471 3959 4478
rect 5062 4476 5074 4488
rect 5053 4471 5074 4476
rect 3810 4470 3851 4471
rect 4469 4470 5074 4471
rect 5092 4470 5102 4488
rect 3134 4417 3171 4418
rect 3230 4417 3267 4418
rect 3286 4417 3322 4469
rect 3341 4417 3378 4418
rect 3034 4408 3172 4417
rect 3034 4388 3143 4408
rect 3163 4388 3172 4408
rect 3034 4381 3172 4388
rect 3230 4408 3378 4417
rect 3230 4388 3239 4408
rect 3259 4388 3349 4408
rect 3369 4388 3378 4408
rect 3034 4379 3130 4381
rect 3230 4378 3378 4388
rect 3437 4408 3474 4418
rect 3549 4417 3586 4418
rect 3530 4415 3586 4417
rect 3437 4388 3445 4408
rect 3465 4388 3474 4408
rect 3286 4377 3322 4378
rect 3134 4318 3171 4319
rect 3437 4318 3474 4388
rect 3499 4408 3586 4415
rect 3499 4405 3557 4408
rect 3499 4385 3504 4405
rect 3525 4388 3557 4405
rect 3577 4388 3586 4408
rect 3525 4385 3586 4388
rect 3499 4378 3586 4385
rect 3645 4408 3682 4418
rect 3645 4388 3653 4408
rect 3673 4388 3682 4408
rect 3499 4377 3530 4378
rect 3133 4317 3474 4318
rect 3058 4312 3474 4317
rect 3058 4292 3061 4312
rect 3081 4292 3474 4312
rect 3645 4317 3682 4388
rect 3712 4417 3743 4470
rect 4469 4461 5102 4470
rect 4469 4454 5101 4461
rect 4469 4452 4531 4454
rect 4047 4442 4215 4443
rect 4469 4442 4491 4452
rect 3762 4417 3799 4418
rect 3712 4408 3799 4417
rect 3712 4388 3770 4408
rect 3790 4388 3799 4408
rect 3712 4378 3799 4388
rect 3858 4408 3895 4418
rect 3858 4388 3866 4408
rect 3886 4388 3895 4408
rect 3712 4377 3743 4378
rect 3858 4317 3895 4388
rect 3645 4293 3895 4317
rect 4047 4416 4491 4442
rect 4047 4414 4215 4416
rect 4047 4236 4074 4414
rect 4114 4376 4178 4388
rect 4454 4384 4491 4416
rect 4662 4415 4911 4437
rect 4662 4384 4699 4415
rect 4875 4413 4911 4415
rect 4875 4384 4912 4413
rect 4114 4375 4149 4376
rect 4091 4370 4149 4375
rect 4091 4350 4094 4370
rect 4114 4356 4149 4370
rect 4169 4356 4178 4376
rect 4114 4348 4178 4356
rect 4140 4347 4178 4348
rect 4141 4346 4178 4347
rect 4244 4380 4280 4381
rect 4352 4380 4388 4381
rect 4244 4372 4388 4380
rect 4244 4352 4252 4372
rect 4272 4352 4301 4372
rect 4244 4351 4301 4352
rect 4323 4352 4360 4372
rect 4380 4352 4388 4372
rect 4323 4351 4388 4352
rect 4244 4346 4388 4351
rect 4454 4376 4492 4384
rect 4560 4380 4596 4381
rect 4454 4356 4463 4376
rect 4483 4356 4492 4376
rect 4454 4347 4492 4356
rect 4511 4373 4596 4380
rect 4511 4353 4518 4373
rect 4539 4372 4596 4373
rect 4539 4353 4568 4372
rect 4511 4352 4568 4353
rect 4588 4352 4596 4372
rect 4454 4346 4491 4347
rect 4511 4346 4596 4352
rect 4662 4376 4700 4384
rect 4773 4380 4809 4381
rect 4662 4356 4671 4376
rect 4691 4356 4700 4376
rect 4662 4347 4700 4356
rect 4724 4372 4809 4380
rect 4724 4352 4781 4372
rect 4801 4352 4809 4372
rect 4662 4346 4699 4347
rect 4724 4346 4809 4352
rect 4875 4376 4913 4384
rect 4875 4356 4884 4376
rect 4904 4356 4913 4376
rect 4875 4347 4913 4356
rect 4875 4346 4912 4347
rect 4298 4325 4334 4346
rect 4724 4325 4755 4346
rect 4131 4321 4231 4325
rect 4131 4317 4193 4321
rect 4131 4291 4138 4317
rect 4164 4295 4193 4317
rect 4219 4295 4231 4321
rect 4164 4291 4231 4295
rect 4131 4288 4231 4291
rect 4299 4288 4334 4325
rect 4396 4322 4755 4325
rect 4396 4317 4618 4322
rect 4396 4293 4409 4317
rect 4433 4298 4618 4317
rect 4642 4298 4755 4322
rect 4433 4293 4755 4298
rect 4396 4289 4755 4293
rect 4822 4317 4971 4325
rect 4822 4297 4833 4317
rect 4853 4297 4971 4317
rect 4822 4290 4971 4297
rect 5062 4305 5101 4454
rect 4822 4289 4863 4290
rect 4146 4236 4183 4237
rect 4242 4236 4279 4237
rect 4298 4236 4334 4288
rect 4353 4236 4390 4237
rect 4046 4227 4184 4236
rect 4046 4207 4155 4227
rect 4175 4207 4184 4227
rect 4046 4200 4184 4207
rect 4242 4227 4390 4236
rect 4242 4207 4251 4227
rect 4271 4207 4361 4227
rect 4381 4207 4390 4227
rect 4046 4198 4142 4200
rect 4242 4197 4390 4207
rect 4449 4227 4486 4237
rect 4561 4236 4598 4237
rect 4542 4234 4598 4236
rect 4449 4207 4457 4227
rect 4477 4207 4486 4227
rect 4298 4196 4334 4197
rect 2211 4188 2242 4191
rect 2740 4191 2908 4192
rect 1040 4164 1178 4173
rect 2740 4165 3184 4191
rect 834 4163 871 4164
rect 890 4112 926 4164
rect 945 4163 982 4164
rect 1041 4163 1078 4164
rect 361 4110 402 4111
rect 253 4103 402 4110
rect 253 4083 371 4103
rect 391 4083 402 4103
rect 253 4075 402 4083
rect 469 4107 828 4111
rect 469 4102 791 4107
rect 469 4078 582 4102
rect 606 4083 791 4102
rect 815 4083 828 4107
rect 606 4078 828 4083
rect 469 4075 828 4078
rect 890 4075 925 4112
rect 993 4109 1093 4112
rect 993 4105 1060 4109
rect 993 4079 1005 4105
rect 1031 4083 1060 4105
rect 1086 4083 1093 4109
rect 1031 4079 1093 4083
rect 993 4075 1093 4079
rect 469 4054 500 4075
rect 890 4054 926 4075
rect 133 4045 170 4054
rect 312 4053 349 4054
rect 133 4027 142 4045
rect 160 4027 170 4045
rect 133 4017 170 4027
rect 134 3982 170 4017
rect 311 4044 349 4053
rect 311 4024 320 4044
rect 340 4024 349 4044
rect 311 4016 349 4024
rect 415 4048 500 4054
rect 525 4053 562 4054
rect 415 4028 423 4048
rect 443 4028 500 4048
rect 415 4020 500 4028
rect 524 4044 562 4053
rect 524 4024 533 4044
rect 553 4024 562 4044
rect 415 4019 451 4020
rect 524 4016 562 4024
rect 628 4048 713 4054
rect 733 4053 770 4054
rect 628 4028 636 4048
rect 656 4047 713 4048
rect 656 4028 685 4047
rect 628 4027 685 4028
rect 706 4027 713 4047
rect 628 4020 713 4027
rect 732 4044 770 4053
rect 732 4024 741 4044
rect 761 4024 770 4044
rect 628 4019 664 4020
rect 732 4016 770 4024
rect 836 4048 980 4054
rect 836 4028 844 4048
rect 864 4047 952 4048
rect 864 4028 892 4047
rect 836 4026 892 4028
rect 914 4028 952 4047
rect 972 4028 980 4048
rect 914 4026 980 4028
rect 836 4020 980 4026
rect 836 4019 872 4020
rect 944 4019 980 4020
rect 1046 4053 1083 4054
rect 1046 4052 1084 4053
rect 1046 4044 1110 4052
rect 1046 4024 1055 4044
rect 1075 4030 1110 4044
rect 1130 4030 1133 4050
rect 1075 4025 1133 4030
rect 1075 4024 1110 4025
rect 312 3987 349 4016
rect 132 3941 170 3982
rect 313 3985 349 3987
rect 525 3985 562 4016
rect 313 3963 562 3985
rect 733 3984 770 4016
rect 1046 4012 1110 4024
rect 1150 3986 1177 4164
rect 1009 3984 1177 3986
rect 2740 4163 2908 4165
rect 2740 4160 2787 4163
rect 2740 3985 2767 4160
rect 2807 4125 2871 4137
rect 3147 4133 3184 4165
rect 3355 4164 3604 4186
rect 3355 4133 3392 4164
rect 3568 4162 3604 4164
rect 3568 4133 3605 4162
rect 4146 4137 4183 4138
rect 4449 4137 4486 4207
rect 4511 4227 4598 4234
rect 4511 4224 4569 4227
rect 4511 4204 4516 4224
rect 4537 4207 4569 4224
rect 4589 4207 4598 4227
rect 4537 4204 4598 4207
rect 4511 4197 4598 4204
rect 4657 4227 4694 4237
rect 4657 4207 4665 4227
rect 4685 4207 4694 4227
rect 4511 4196 4542 4197
rect 4145 4136 4486 4137
rect 2807 4124 2842 4125
rect 2784 4119 2842 4124
rect 2784 4099 2787 4119
rect 2807 4105 2842 4119
rect 2862 4105 2871 4125
rect 2807 4097 2871 4105
rect 2833 4096 2871 4097
rect 2834 4095 2871 4096
rect 2937 4129 2973 4130
rect 3045 4129 3081 4130
rect 2937 4121 3081 4129
rect 2937 4101 2945 4121
rect 2965 4119 3053 4121
rect 2965 4101 2991 4119
rect 2937 4100 2991 4101
rect 3017 4101 3053 4119
rect 3073 4101 3081 4121
rect 3017 4100 3081 4101
rect 2937 4095 3081 4100
rect 3147 4125 3185 4133
rect 3253 4129 3289 4130
rect 3147 4105 3156 4125
rect 3176 4105 3185 4125
rect 3147 4096 3185 4105
rect 3204 4122 3289 4129
rect 3204 4102 3211 4122
rect 3232 4121 3289 4122
rect 3232 4102 3261 4121
rect 3204 4101 3261 4102
rect 3281 4101 3289 4121
rect 3147 4095 3184 4096
rect 3204 4095 3289 4101
rect 3355 4125 3393 4133
rect 3466 4129 3502 4130
rect 3355 4105 3364 4125
rect 3384 4105 3393 4125
rect 3355 4096 3393 4105
rect 3417 4121 3502 4129
rect 3417 4101 3474 4121
rect 3494 4101 3502 4121
rect 3355 4095 3392 4096
rect 3417 4095 3502 4101
rect 3568 4125 3606 4133
rect 3568 4105 3577 4125
rect 3597 4105 3606 4125
rect 4070 4131 4486 4136
rect 4070 4111 4073 4131
rect 4093 4111 4486 4131
rect 4657 4136 4694 4207
rect 4724 4236 4755 4289
rect 5062 4287 5072 4305
rect 5090 4287 5101 4305
rect 5062 4278 5099 4287
rect 4774 4236 4811 4237
rect 4724 4227 4811 4236
rect 4724 4207 4782 4227
rect 4802 4207 4811 4227
rect 4724 4197 4811 4207
rect 4870 4227 4907 4237
rect 4870 4207 4878 4227
rect 4898 4207 4907 4227
rect 5065 4212 5102 4216
rect 4724 4196 4755 4197
rect 4870 4136 4907 4207
rect 4657 4112 4907 4136
rect 5063 4206 5102 4212
rect 5063 4188 5074 4206
rect 5092 4188 5102 4206
rect 5063 4179 5102 4188
rect 3568 4096 3606 4105
rect 3568 4095 3605 4096
rect 2991 4074 3027 4095
rect 3417 4074 3448 4095
rect 4449 4088 4486 4111
rect 5063 4101 5098 4179
rect 5060 4091 5098 4101
rect 4449 4087 4619 4088
rect 5060 4087 5070 4091
rect 2824 4070 2924 4074
rect 2824 4066 2886 4070
rect 2824 4040 2831 4066
rect 2857 4044 2886 4066
rect 2912 4044 2924 4070
rect 2857 4040 2924 4044
rect 2824 4037 2924 4040
rect 2992 4037 3027 4074
rect 3089 4071 3448 4074
rect 3089 4066 3311 4071
rect 3089 4042 3102 4066
rect 3126 4047 3311 4066
rect 3335 4047 3448 4071
rect 3126 4042 3448 4047
rect 3089 4038 3448 4042
rect 3515 4066 3664 4074
rect 4449 4073 5070 4087
rect 5088 4073 5098 4091
rect 4449 4067 5098 4073
rect 4449 4066 5097 4067
rect 3515 4046 3526 4066
rect 3546 4046 3664 4066
rect 5060 4064 5097 4066
rect 3515 4039 3664 4046
rect 3515 4038 3556 4039
rect 2839 3985 2876 3986
rect 2935 3985 2972 3986
rect 2991 3985 3027 4037
rect 3046 3985 3083 3986
rect 733 3958 1177 3984
rect 734 3941 758 3958
rect 1009 3957 1177 3958
rect 1628 3954 1878 3978
rect 132 3923 759 3941
rect 132 3922 170 3923
rect 130 3917 170 3922
rect 130 3874 165 3917
rect 128 3865 165 3874
rect 128 3847 138 3865
rect 156 3847 165 3865
rect 1628 3883 1665 3954
rect 1780 3893 1811 3894
rect 1628 3863 1637 3883
rect 1657 3863 1665 3883
rect 1628 3853 1665 3863
rect 1724 3883 1811 3893
rect 1724 3863 1733 3883
rect 1753 3863 1811 3883
rect 1724 3854 1811 3863
rect 1724 3853 1761 3854
rect 128 3837 165 3847
rect 1780 3801 1811 3854
rect 1841 3883 1878 3954
rect 2049 3959 2442 3979
rect 2462 3959 2465 3979
rect 2049 3954 2465 3959
rect 2739 3976 2877 3985
rect 2739 3956 2848 3976
rect 2868 3956 2877 3976
rect 2049 3953 2390 3954
rect 1993 3893 2024 3894
rect 1841 3863 1850 3883
rect 1870 3863 1878 3883
rect 1841 3853 1878 3863
rect 1937 3886 2024 3893
rect 1937 3883 1998 3886
rect 1937 3863 1946 3883
rect 1966 3866 1998 3883
rect 2019 3866 2024 3886
rect 1966 3863 2024 3866
rect 1937 3856 2024 3863
rect 2049 3883 2086 3953
rect 2352 3952 2389 3953
rect 2739 3949 2877 3956
rect 2935 3976 3083 3985
rect 2935 3956 2944 3976
rect 2964 3956 3054 3976
rect 3074 3956 3083 3976
rect 2739 3947 2835 3949
rect 2935 3946 3083 3956
rect 3142 3976 3179 3986
rect 3254 3985 3291 3986
rect 3235 3983 3291 3985
rect 3142 3956 3150 3976
rect 3170 3956 3179 3976
rect 2991 3945 3027 3946
rect 2201 3893 2237 3894
rect 2049 3863 2058 3883
rect 2078 3863 2086 3883
rect 1937 3854 1993 3856
rect 1937 3853 1974 3854
rect 2049 3853 2086 3863
rect 2145 3883 2293 3893
rect 2393 3890 2489 3892
rect 2145 3863 2154 3883
rect 2174 3863 2264 3883
rect 2284 3863 2293 3883
rect 2145 3854 2293 3863
rect 2351 3883 2489 3890
rect 2839 3886 2876 3887
rect 3142 3886 3179 3956
rect 3204 3976 3291 3983
rect 3204 3973 3262 3976
rect 3204 3953 3209 3973
rect 3230 3956 3262 3973
rect 3282 3956 3291 3976
rect 3230 3953 3291 3956
rect 3204 3946 3291 3953
rect 3350 3976 3387 3986
rect 3350 3956 3358 3976
rect 3378 3956 3387 3976
rect 3204 3945 3235 3946
rect 2838 3885 3179 3886
rect 2351 3863 2360 3883
rect 2380 3863 2489 3883
rect 2351 3854 2489 3863
rect 2763 3880 3179 3885
rect 2763 3860 2766 3880
rect 2786 3860 3179 3880
rect 3350 3885 3387 3956
rect 3417 3985 3448 4038
rect 5063 3992 5100 4002
rect 3467 3985 3504 3986
rect 3417 3976 3504 3985
rect 3417 3956 3475 3976
rect 3495 3956 3504 3976
rect 3417 3946 3504 3956
rect 3563 3976 3600 3986
rect 3563 3956 3571 3976
rect 3591 3956 3600 3976
rect 3417 3945 3448 3946
rect 3563 3885 3600 3956
rect 5063 3974 5072 3992
rect 5090 3974 5100 3992
rect 5063 3965 5100 3974
rect 5063 3922 5098 3965
rect 5058 3917 5098 3922
rect 5058 3916 5096 3917
rect 4469 3898 5096 3916
rect 3350 3861 3600 3885
rect 4051 3881 4219 3882
rect 4470 3881 4494 3898
rect 4051 3855 4495 3881
rect 2145 3853 2182 3854
rect 2201 3802 2237 3854
rect 2256 3853 2293 3854
rect 2352 3853 2389 3854
rect 1672 3800 1713 3801
rect 1564 3793 1713 3800
rect 131 3773 168 3775
rect 1564 3773 1682 3793
rect 1702 3773 1713 3793
rect 131 3772 779 3773
rect 130 3766 779 3772
rect 130 3748 140 3766
rect 158 3752 779 3766
rect 1564 3765 1713 3773
rect 1780 3797 2139 3801
rect 1780 3792 2102 3797
rect 1780 3768 1893 3792
rect 1917 3773 2102 3792
rect 2126 3773 2139 3797
rect 1917 3768 2139 3773
rect 1780 3765 2139 3768
rect 2201 3765 2236 3802
rect 2304 3799 2404 3802
rect 2304 3795 2371 3799
rect 2304 3769 2316 3795
rect 2342 3773 2371 3795
rect 2397 3773 2404 3799
rect 2342 3769 2404 3773
rect 2304 3765 2404 3769
rect 158 3748 168 3752
rect 609 3751 779 3752
rect 130 3738 168 3748
rect 130 3660 165 3738
rect 742 3728 779 3751
rect 1780 3744 1811 3765
rect 2201 3744 2237 3765
rect 1623 3743 1660 3744
rect 1622 3734 1660 3743
rect 126 3651 165 3660
rect 126 3633 136 3651
rect 154 3633 165 3651
rect 126 3627 165 3633
rect 321 3703 571 3727
rect 321 3632 358 3703
rect 473 3642 504 3643
rect 126 3623 163 3627
rect 321 3612 330 3632
rect 350 3612 358 3632
rect 321 3602 358 3612
rect 417 3632 504 3642
rect 417 3612 426 3632
rect 446 3612 504 3632
rect 417 3603 504 3612
rect 417 3602 454 3603
rect 129 3552 166 3561
rect 127 3534 138 3552
rect 156 3534 166 3552
rect 473 3550 504 3603
rect 534 3632 571 3703
rect 742 3708 1135 3728
rect 1155 3708 1158 3728
rect 742 3703 1158 3708
rect 1622 3714 1631 3734
rect 1651 3714 1660 3734
rect 1622 3706 1660 3714
rect 1726 3738 1811 3744
rect 1836 3743 1873 3744
rect 1726 3718 1734 3738
rect 1754 3718 1811 3738
rect 1726 3710 1811 3718
rect 1835 3734 1873 3743
rect 1835 3714 1844 3734
rect 1864 3714 1873 3734
rect 1726 3709 1762 3710
rect 1835 3706 1873 3714
rect 1939 3738 2024 3744
rect 2044 3743 2081 3744
rect 1939 3718 1947 3738
rect 1967 3737 2024 3738
rect 1967 3718 1996 3737
rect 1939 3717 1996 3718
rect 2017 3717 2024 3737
rect 1939 3710 2024 3717
rect 2043 3734 2081 3743
rect 2043 3714 2052 3734
rect 2072 3714 2081 3734
rect 1939 3709 1975 3710
rect 2043 3706 2081 3714
rect 2147 3739 2291 3744
rect 2147 3738 2211 3739
rect 2147 3718 2155 3738
rect 2175 3720 2211 3738
rect 2237 3738 2291 3739
rect 2237 3720 2263 3738
rect 2175 3718 2263 3720
rect 2283 3718 2291 3738
rect 2147 3710 2291 3718
rect 2147 3709 2183 3710
rect 2255 3709 2291 3710
rect 2357 3743 2394 3744
rect 2357 3742 2395 3743
rect 2357 3734 2421 3742
rect 2357 3714 2366 3734
rect 2386 3720 2421 3734
rect 2441 3720 2444 3740
rect 2386 3715 2444 3720
rect 2386 3714 2421 3715
rect 742 3702 1083 3703
rect 686 3642 717 3643
rect 534 3612 543 3632
rect 563 3612 571 3632
rect 534 3602 571 3612
rect 630 3635 717 3642
rect 630 3632 691 3635
rect 630 3612 639 3632
rect 659 3615 691 3632
rect 712 3615 717 3635
rect 659 3612 717 3615
rect 630 3605 717 3612
rect 742 3632 779 3702
rect 1045 3701 1082 3702
rect 1623 3677 1660 3706
rect 1624 3675 1660 3677
rect 1836 3675 1873 3706
rect 1624 3653 1873 3675
rect 2044 3674 2081 3706
rect 2357 3702 2421 3714
rect 2461 3679 2488 3854
rect 2441 3676 2488 3679
rect 2320 3674 2488 3676
rect 4051 3853 4219 3855
rect 4051 3675 4078 3853
rect 4118 3815 4182 3827
rect 4458 3823 4495 3855
rect 4666 3854 4915 3876
rect 4666 3823 4703 3854
rect 4879 3852 4915 3854
rect 5058 3857 5096 3898
rect 4879 3823 4916 3852
rect 4118 3814 4153 3815
rect 4095 3809 4153 3814
rect 4095 3789 4098 3809
rect 4118 3795 4153 3809
rect 4173 3795 4182 3815
rect 4118 3787 4182 3795
rect 4144 3786 4182 3787
rect 4145 3785 4182 3786
rect 4248 3819 4284 3820
rect 4356 3819 4392 3820
rect 4248 3813 4392 3819
rect 4248 3811 4314 3813
rect 4248 3791 4256 3811
rect 4276 3792 4314 3811
rect 4336 3811 4392 3813
rect 4336 3792 4364 3811
rect 4276 3791 4364 3792
rect 4384 3791 4392 3811
rect 4248 3785 4392 3791
rect 4458 3815 4496 3823
rect 4564 3819 4600 3820
rect 4458 3795 4467 3815
rect 4487 3795 4496 3815
rect 4458 3786 4496 3795
rect 4515 3812 4600 3819
rect 4515 3792 4522 3812
rect 4543 3811 4600 3812
rect 4543 3792 4572 3811
rect 4515 3791 4572 3792
rect 4592 3791 4600 3811
rect 4458 3785 4495 3786
rect 4515 3785 4600 3791
rect 4666 3815 4704 3823
rect 4777 3819 4813 3820
rect 4666 3795 4675 3815
rect 4695 3795 4704 3815
rect 4666 3786 4704 3795
rect 4728 3811 4813 3819
rect 4728 3791 4785 3811
rect 4805 3791 4813 3811
rect 4666 3785 4703 3786
rect 4728 3785 4813 3791
rect 4879 3815 4917 3823
rect 4879 3795 4888 3815
rect 4908 3795 4917 3815
rect 4879 3786 4917 3795
rect 5058 3822 5094 3857
rect 5058 3812 5095 3822
rect 5058 3794 5068 3812
rect 5086 3794 5095 3812
rect 4879 3785 4916 3786
rect 5058 3785 5095 3794
rect 4302 3764 4338 3785
rect 4728 3764 4759 3785
rect 4135 3760 4235 3764
rect 4135 3756 4197 3760
rect 4135 3730 4142 3756
rect 4168 3734 4197 3756
rect 4223 3734 4235 3760
rect 4168 3730 4235 3734
rect 4135 3727 4235 3730
rect 4303 3727 4338 3764
rect 4400 3761 4759 3764
rect 4400 3756 4622 3761
rect 4400 3732 4413 3756
rect 4437 3737 4622 3756
rect 4646 3737 4759 3761
rect 4437 3732 4759 3737
rect 4400 3728 4759 3732
rect 4826 3756 4975 3764
rect 4826 3736 4837 3756
rect 4857 3736 4975 3756
rect 4826 3729 4975 3736
rect 4826 3728 4867 3729
rect 4150 3675 4187 3676
rect 4246 3675 4283 3676
rect 4302 3675 4338 3727
rect 4357 3675 4394 3676
rect 2044 3648 2488 3674
rect 4050 3666 4188 3675
rect 2320 3647 2488 3648
rect 2986 3648 3017 3651
rect 894 3642 930 3643
rect 742 3612 751 3632
rect 771 3612 779 3632
rect 630 3603 686 3605
rect 630 3602 667 3603
rect 742 3602 779 3612
rect 838 3632 986 3642
rect 1086 3639 1182 3641
rect 838 3612 847 3632
rect 867 3612 957 3632
rect 977 3612 986 3632
rect 838 3603 986 3612
rect 1044 3632 1182 3639
rect 1044 3612 1053 3632
rect 1073 3612 1182 3632
rect 1044 3603 1182 3612
rect 838 3602 875 3603
rect 894 3551 930 3603
rect 949 3602 986 3603
rect 1045 3602 1082 3603
rect 365 3549 406 3550
rect 127 3385 166 3534
rect 257 3542 406 3549
rect 257 3522 375 3542
rect 395 3522 406 3542
rect 257 3514 406 3522
rect 473 3546 832 3550
rect 473 3541 795 3546
rect 473 3517 586 3541
rect 610 3522 795 3541
rect 819 3522 832 3546
rect 610 3517 832 3522
rect 473 3514 832 3517
rect 894 3514 929 3551
rect 997 3548 1097 3551
rect 997 3544 1064 3548
rect 997 3518 1009 3544
rect 1035 3522 1064 3544
rect 1090 3522 1097 3548
rect 1035 3518 1097 3522
rect 997 3514 1097 3518
rect 473 3493 504 3514
rect 894 3493 930 3514
rect 316 3492 353 3493
rect 315 3483 353 3492
rect 315 3463 324 3483
rect 344 3463 353 3483
rect 315 3455 353 3463
rect 419 3487 504 3493
rect 529 3492 566 3493
rect 419 3467 427 3487
rect 447 3467 504 3487
rect 419 3459 504 3467
rect 528 3483 566 3492
rect 528 3463 537 3483
rect 557 3463 566 3483
rect 419 3458 455 3459
rect 528 3455 566 3463
rect 632 3487 717 3493
rect 737 3492 774 3493
rect 632 3467 640 3487
rect 660 3486 717 3487
rect 660 3467 689 3486
rect 632 3466 689 3467
rect 710 3466 717 3486
rect 632 3459 717 3466
rect 736 3483 774 3492
rect 736 3463 745 3483
rect 765 3463 774 3483
rect 632 3458 668 3459
rect 736 3455 774 3463
rect 840 3488 984 3493
rect 840 3487 905 3488
rect 840 3467 848 3487
rect 868 3467 905 3487
rect 927 3487 984 3488
rect 927 3467 956 3487
rect 976 3467 984 3487
rect 840 3459 984 3467
rect 840 3458 876 3459
rect 948 3458 984 3459
rect 1050 3492 1087 3493
rect 1050 3491 1088 3492
rect 1050 3483 1114 3491
rect 1050 3463 1059 3483
rect 1079 3469 1114 3483
rect 1134 3469 1137 3489
rect 1079 3464 1137 3469
rect 1079 3463 1114 3464
rect 316 3426 353 3455
rect 317 3424 353 3426
rect 529 3424 566 3455
rect 317 3402 566 3424
rect 737 3423 774 3455
rect 1050 3451 1114 3463
rect 1154 3425 1181 3603
rect 1013 3423 1181 3425
rect 737 3397 1181 3423
rect 1333 3522 1583 3546
rect 1333 3451 1370 3522
rect 1485 3461 1516 3462
rect 1333 3431 1342 3451
rect 1362 3431 1370 3451
rect 1333 3421 1370 3431
rect 1429 3451 1516 3461
rect 1429 3431 1438 3451
rect 1458 3431 1516 3451
rect 1429 3422 1516 3431
rect 1429 3421 1466 3422
rect 737 3387 759 3397
rect 1013 3396 1181 3397
rect 697 3385 759 3387
rect 127 3378 759 3385
rect 126 3369 759 3378
rect 1485 3369 1516 3422
rect 1546 3451 1583 3522
rect 1754 3527 2147 3547
rect 2167 3527 2170 3547
rect 1754 3522 2170 3527
rect 1754 3521 2095 3522
rect 1698 3461 1729 3462
rect 1546 3431 1555 3451
rect 1575 3431 1583 3451
rect 1546 3421 1583 3431
rect 1642 3454 1729 3461
rect 1642 3451 1703 3454
rect 1642 3431 1651 3451
rect 1671 3434 1703 3451
rect 1724 3434 1729 3454
rect 1671 3431 1729 3434
rect 1642 3424 1729 3431
rect 1754 3451 1791 3521
rect 2057 3520 2094 3521
rect 1906 3461 1942 3462
rect 1754 3431 1763 3451
rect 1783 3431 1791 3451
rect 1642 3422 1698 3424
rect 1642 3421 1679 3422
rect 1754 3421 1791 3431
rect 1850 3451 1998 3461
rect 2098 3458 2194 3460
rect 1850 3431 1859 3451
rect 1879 3431 1969 3451
rect 1989 3431 1998 3451
rect 1850 3422 1998 3431
rect 2056 3451 2194 3458
rect 2056 3431 2065 3451
rect 2085 3431 2194 3451
rect 2056 3422 2194 3431
rect 1850 3421 1887 3422
rect 1906 3370 1942 3422
rect 1961 3421 1998 3422
rect 2057 3421 2094 3422
rect 126 3351 136 3369
rect 154 3368 759 3369
rect 1377 3368 1418 3369
rect 154 3363 175 3368
rect 154 3351 166 3363
rect 1269 3361 1418 3368
rect 126 3343 166 3351
rect 209 3350 235 3351
rect 126 3341 163 3343
rect 209 3332 763 3350
rect 1269 3341 1387 3361
rect 1407 3341 1418 3361
rect 1269 3333 1418 3341
rect 1485 3365 1844 3369
rect 1485 3360 1807 3365
rect 1485 3336 1598 3360
rect 1622 3341 1807 3360
rect 1831 3341 1844 3365
rect 1622 3336 1844 3341
rect 1485 3333 1844 3336
rect 1906 3333 1941 3370
rect 2009 3367 2109 3370
rect 2009 3363 2076 3367
rect 2009 3337 2021 3363
rect 2047 3341 2076 3363
rect 2102 3341 2109 3367
rect 2047 3337 2109 3341
rect 2009 3333 2109 3337
rect 129 3273 166 3279
rect 209 3273 235 3332
rect 742 3313 763 3332
rect 129 3270 235 3273
rect 129 3252 138 3270
rect 156 3256 235 3270
rect 320 3288 570 3312
rect 156 3254 232 3256
rect 156 3252 166 3254
rect 129 3242 166 3252
rect 134 3177 165 3242
rect 320 3217 357 3288
rect 472 3227 503 3228
rect 320 3197 329 3217
rect 349 3197 357 3217
rect 320 3187 357 3197
rect 416 3217 503 3227
rect 416 3197 425 3217
rect 445 3197 503 3217
rect 416 3188 503 3197
rect 416 3187 453 3188
rect 133 3168 170 3177
rect 133 3150 143 3168
rect 161 3150 170 3168
rect 133 3140 170 3150
rect 472 3135 503 3188
rect 533 3217 570 3288
rect 741 3293 1134 3313
rect 1154 3293 1157 3313
rect 1485 3312 1516 3333
rect 1906 3312 1942 3333
rect 1328 3311 1365 3312
rect 741 3288 1157 3293
rect 1327 3302 1365 3311
rect 741 3287 1082 3288
rect 685 3227 716 3228
rect 533 3197 542 3217
rect 562 3197 570 3217
rect 533 3187 570 3197
rect 629 3220 716 3227
rect 629 3217 690 3220
rect 629 3197 638 3217
rect 658 3200 690 3217
rect 711 3200 716 3220
rect 658 3197 716 3200
rect 629 3190 716 3197
rect 741 3217 778 3287
rect 1044 3286 1081 3287
rect 1327 3282 1336 3302
rect 1356 3282 1365 3302
rect 1327 3274 1365 3282
rect 1431 3306 1516 3312
rect 1541 3311 1578 3312
rect 1431 3286 1439 3306
rect 1459 3286 1516 3306
rect 1431 3278 1516 3286
rect 1540 3302 1578 3311
rect 1540 3282 1549 3302
rect 1569 3282 1578 3302
rect 1431 3277 1467 3278
rect 1540 3274 1578 3282
rect 1644 3306 1729 3312
rect 1749 3311 1786 3312
rect 1644 3286 1652 3306
rect 1672 3305 1729 3306
rect 1672 3286 1701 3305
rect 1644 3285 1701 3286
rect 1722 3285 1729 3305
rect 1644 3278 1729 3285
rect 1748 3302 1786 3311
rect 1748 3282 1757 3302
rect 1777 3282 1786 3302
rect 1644 3277 1680 3278
rect 1748 3274 1786 3282
rect 1852 3306 1996 3312
rect 1852 3286 1860 3306
rect 1880 3286 1912 3306
rect 1936 3286 1968 3306
rect 1988 3286 1996 3306
rect 1852 3278 1996 3286
rect 1852 3277 1888 3278
rect 1960 3277 1996 3278
rect 2062 3311 2099 3312
rect 2062 3310 2100 3311
rect 2062 3302 2126 3310
rect 2062 3282 2071 3302
rect 2091 3288 2126 3302
rect 2146 3288 2149 3308
rect 2091 3283 2149 3288
rect 2091 3282 2126 3283
rect 1328 3245 1365 3274
rect 1329 3243 1365 3245
rect 1541 3243 1578 3274
rect 893 3227 929 3228
rect 741 3197 750 3217
rect 770 3197 778 3217
rect 629 3188 685 3190
rect 629 3187 666 3188
rect 741 3187 778 3197
rect 837 3217 985 3227
rect 1085 3224 1181 3226
rect 837 3197 846 3217
rect 866 3197 956 3217
rect 976 3197 985 3217
rect 837 3188 985 3197
rect 1043 3217 1181 3224
rect 1329 3221 1578 3243
rect 1749 3242 1786 3274
rect 2062 3270 2126 3282
rect 2166 3244 2193 3422
rect 2025 3242 2193 3244
rect 1749 3238 2193 3242
rect 1043 3197 1052 3217
rect 1072 3197 1181 3217
rect 1749 3219 1798 3238
rect 1818 3219 2193 3238
rect 1749 3216 2193 3219
rect 2025 3215 2193 3216
rect 1043 3188 1181 3197
rect 837 3187 874 3188
rect 893 3136 929 3188
rect 948 3187 985 3188
rect 1044 3187 1081 3188
rect 364 3134 405 3135
rect 256 3127 405 3134
rect 256 3107 374 3127
rect 394 3107 405 3127
rect 256 3099 405 3107
rect 472 3131 831 3135
rect 472 3126 794 3131
rect 472 3102 585 3126
rect 609 3107 794 3126
rect 818 3107 831 3131
rect 609 3102 831 3107
rect 472 3099 831 3102
rect 893 3099 928 3136
rect 996 3133 1096 3136
rect 996 3129 1063 3133
rect 996 3103 1008 3129
rect 1034 3107 1063 3129
rect 1089 3107 1096 3133
rect 1034 3103 1096 3107
rect 996 3099 1096 3103
rect 472 3078 503 3099
rect 893 3078 929 3099
rect 136 3069 173 3078
rect 315 3077 352 3078
rect 136 3051 145 3069
rect 163 3051 173 3069
rect 136 3041 173 3051
rect 137 3006 173 3041
rect 314 3068 352 3077
rect 314 3048 323 3068
rect 343 3048 352 3068
rect 314 3040 352 3048
rect 418 3072 503 3078
rect 528 3077 565 3078
rect 418 3052 426 3072
rect 446 3052 503 3072
rect 418 3044 503 3052
rect 527 3068 565 3077
rect 527 3048 536 3068
rect 556 3048 565 3068
rect 418 3043 454 3044
rect 527 3040 565 3048
rect 631 3072 716 3078
rect 736 3077 773 3078
rect 631 3052 639 3072
rect 659 3071 716 3072
rect 659 3052 688 3071
rect 631 3051 688 3052
rect 709 3051 716 3071
rect 631 3044 716 3051
rect 735 3068 773 3077
rect 735 3048 744 3068
rect 764 3048 773 3068
rect 631 3043 667 3044
rect 735 3040 773 3048
rect 839 3072 983 3078
rect 839 3052 847 3072
rect 867 3071 955 3072
rect 867 3052 895 3071
rect 839 3050 895 3052
rect 917 3052 955 3071
rect 975 3052 983 3072
rect 917 3050 983 3052
rect 839 3044 983 3050
rect 839 3043 875 3044
rect 947 3043 983 3044
rect 1049 3077 1086 3078
rect 1049 3076 1087 3077
rect 1049 3068 1113 3076
rect 1049 3048 1058 3068
rect 1078 3054 1113 3068
rect 1133 3054 1136 3074
rect 1078 3049 1136 3054
rect 1078 3048 1113 3049
rect 315 3011 352 3040
rect 135 2965 173 3006
rect 316 3009 352 3011
rect 528 3009 565 3040
rect 316 2987 565 3009
rect 736 3008 773 3040
rect 1049 3036 1113 3048
rect 1153 3010 1180 3188
rect 1012 3008 1180 3010
rect 736 2982 1180 3008
rect 737 2965 761 2982
rect 1012 2981 1180 2982
rect 135 2947 762 2965
rect 1388 2961 1638 2985
rect 135 2941 173 2947
rect 135 2917 172 2941
rect 135 2893 170 2917
rect 133 2884 170 2893
rect 133 2866 143 2884
rect 161 2866 170 2884
rect 133 2856 170 2866
rect 1388 2890 1425 2961
rect 1540 2900 1571 2901
rect 1388 2870 1397 2890
rect 1417 2870 1425 2890
rect 1388 2860 1425 2870
rect 1484 2890 1571 2900
rect 1484 2870 1493 2890
rect 1513 2870 1571 2890
rect 1484 2861 1571 2870
rect 1484 2860 1521 2861
rect 1540 2808 1571 2861
rect 1601 2890 1638 2961
rect 1809 2966 2202 2986
rect 2222 2966 2225 2986
rect 1809 2961 2225 2966
rect 1809 2960 2150 2961
rect 1753 2900 1784 2901
rect 1601 2870 1610 2890
rect 1630 2870 1638 2890
rect 1601 2860 1638 2870
rect 1697 2893 1784 2900
rect 1697 2890 1758 2893
rect 1697 2870 1706 2890
rect 1726 2873 1758 2890
rect 1779 2873 1784 2893
rect 1726 2870 1784 2873
rect 1697 2863 1784 2870
rect 1809 2890 1846 2960
rect 2112 2959 2149 2960
rect 1961 2900 1997 2901
rect 1809 2870 1818 2890
rect 1838 2870 1846 2890
rect 1697 2861 1753 2863
rect 1697 2860 1734 2861
rect 1809 2860 1846 2870
rect 1905 2890 2053 2900
rect 2153 2897 2249 2899
rect 1905 2870 1914 2890
rect 1934 2870 2024 2890
rect 2044 2870 2053 2890
rect 1905 2861 2053 2870
rect 2111 2890 2249 2897
rect 2111 2870 2120 2890
rect 2140 2870 2249 2890
rect 2111 2861 2249 2870
rect 1905 2860 1942 2861
rect 1961 2809 1997 2861
rect 2016 2860 2053 2861
rect 2112 2860 2149 2861
rect 1432 2807 1473 2808
rect 1324 2800 1473 2807
rect 136 2792 173 2794
rect 136 2791 784 2792
rect 135 2785 784 2791
rect 135 2767 145 2785
rect 163 2771 784 2785
rect 1324 2780 1442 2800
rect 1462 2780 1473 2800
rect 1324 2772 1473 2780
rect 1540 2804 1899 2808
rect 1540 2799 1862 2804
rect 1540 2775 1653 2799
rect 1677 2780 1862 2799
rect 1886 2780 1899 2804
rect 1677 2775 1899 2780
rect 1540 2772 1899 2775
rect 1961 2772 1996 2809
rect 2064 2806 2164 2809
rect 2064 2802 2131 2806
rect 2064 2776 2076 2802
rect 2102 2780 2131 2802
rect 2157 2780 2164 2806
rect 2102 2776 2164 2780
rect 2064 2772 2164 2776
rect 163 2767 173 2771
rect 614 2770 784 2771
rect 135 2757 173 2767
rect 135 2679 170 2757
rect 747 2747 784 2770
rect 1540 2751 1571 2772
rect 1961 2751 1997 2772
rect 1383 2750 1420 2751
rect 131 2670 170 2679
rect 131 2652 141 2670
rect 159 2652 170 2670
rect 131 2646 170 2652
rect 326 2722 576 2746
rect 326 2651 363 2722
rect 478 2661 509 2662
rect 131 2642 168 2646
rect 326 2631 335 2651
rect 355 2631 363 2651
rect 326 2621 363 2631
rect 422 2651 509 2661
rect 422 2631 431 2651
rect 451 2631 509 2651
rect 422 2622 509 2631
rect 422 2621 459 2622
rect 134 2571 171 2580
rect 132 2553 143 2571
rect 161 2553 171 2571
rect 478 2569 509 2622
rect 539 2651 576 2722
rect 747 2727 1140 2747
rect 1160 2727 1163 2747
rect 747 2722 1163 2727
rect 1382 2741 1420 2750
rect 747 2721 1088 2722
rect 1382 2721 1391 2741
rect 1411 2721 1420 2741
rect 691 2661 722 2662
rect 539 2631 548 2651
rect 568 2631 576 2651
rect 539 2621 576 2631
rect 635 2654 722 2661
rect 635 2651 696 2654
rect 635 2631 644 2651
rect 664 2634 696 2651
rect 717 2634 722 2654
rect 664 2631 722 2634
rect 635 2624 722 2631
rect 747 2651 784 2721
rect 1050 2720 1087 2721
rect 1382 2713 1420 2721
rect 1486 2745 1571 2751
rect 1596 2750 1633 2751
rect 1486 2725 1494 2745
rect 1514 2725 1571 2745
rect 1486 2717 1571 2725
rect 1595 2741 1633 2750
rect 1595 2721 1604 2741
rect 1624 2721 1633 2741
rect 1486 2716 1522 2717
rect 1595 2713 1633 2721
rect 1699 2745 1784 2751
rect 1804 2750 1841 2751
rect 1699 2725 1707 2745
rect 1727 2744 1784 2745
rect 1727 2725 1756 2744
rect 1699 2724 1756 2725
rect 1777 2724 1784 2744
rect 1699 2717 1784 2724
rect 1803 2741 1841 2750
rect 1803 2721 1812 2741
rect 1832 2721 1841 2741
rect 1699 2716 1735 2717
rect 1803 2713 1841 2721
rect 1907 2745 2051 2751
rect 1907 2725 1915 2745
rect 1935 2743 2023 2745
rect 1935 2726 1971 2743
rect 1995 2726 2023 2743
rect 1935 2725 2023 2726
rect 2043 2725 2051 2745
rect 1907 2717 2051 2725
rect 1907 2716 1943 2717
rect 2015 2716 2051 2717
rect 2117 2750 2154 2751
rect 2117 2749 2155 2750
rect 2117 2741 2181 2749
rect 2117 2721 2126 2741
rect 2146 2727 2181 2741
rect 2201 2727 2204 2747
rect 2146 2722 2204 2727
rect 2146 2721 2181 2722
rect 1383 2684 1420 2713
rect 1384 2682 1420 2684
rect 1596 2682 1633 2713
rect 899 2661 935 2662
rect 747 2631 756 2651
rect 776 2631 784 2651
rect 635 2622 691 2624
rect 635 2621 672 2622
rect 747 2621 784 2631
rect 843 2651 991 2661
rect 1384 2660 1633 2682
rect 1804 2681 1841 2713
rect 2117 2709 2181 2721
rect 2221 2683 2248 2861
rect 2080 2681 2248 2683
rect 1804 2670 2248 2681
rect 1091 2658 1187 2660
rect 843 2631 852 2651
rect 872 2631 962 2651
rect 982 2631 991 2651
rect 843 2622 991 2631
rect 1049 2651 1187 2658
rect 1804 2655 2250 2670
rect 2080 2654 2250 2655
rect 1049 2631 1058 2651
rect 1078 2631 1187 2651
rect 1049 2622 1187 2631
rect 843 2621 880 2622
rect 899 2570 935 2622
rect 954 2621 991 2622
rect 1050 2621 1087 2622
rect 370 2568 411 2569
rect 132 2404 171 2553
rect 262 2561 411 2568
rect 262 2541 380 2561
rect 400 2541 411 2561
rect 262 2533 411 2541
rect 478 2565 837 2569
rect 478 2560 800 2565
rect 478 2536 591 2560
rect 615 2541 800 2560
rect 824 2541 837 2565
rect 615 2536 837 2541
rect 478 2533 837 2536
rect 899 2533 934 2570
rect 1002 2567 1102 2570
rect 1002 2563 1069 2567
rect 1002 2537 1014 2563
rect 1040 2541 1069 2563
rect 1095 2541 1102 2567
rect 1040 2537 1102 2541
rect 1002 2533 1102 2537
rect 478 2512 509 2533
rect 899 2512 935 2533
rect 321 2511 358 2512
rect 320 2502 358 2511
rect 320 2482 329 2502
rect 349 2482 358 2502
rect 320 2474 358 2482
rect 424 2506 509 2512
rect 534 2511 571 2512
rect 424 2486 432 2506
rect 452 2486 509 2506
rect 424 2478 509 2486
rect 533 2502 571 2511
rect 533 2482 542 2502
rect 562 2482 571 2502
rect 424 2477 460 2478
rect 533 2474 571 2482
rect 637 2506 722 2512
rect 742 2511 779 2512
rect 637 2486 645 2506
rect 665 2505 722 2506
rect 665 2486 694 2505
rect 637 2485 694 2486
rect 715 2485 722 2505
rect 637 2478 722 2485
rect 741 2502 779 2511
rect 741 2482 750 2502
rect 770 2482 779 2502
rect 637 2477 673 2478
rect 741 2474 779 2482
rect 845 2507 989 2512
rect 845 2506 910 2507
rect 845 2486 853 2506
rect 873 2486 910 2506
rect 932 2506 989 2507
rect 932 2486 961 2506
rect 981 2486 989 2506
rect 845 2478 989 2486
rect 845 2477 881 2478
rect 953 2477 989 2478
rect 1055 2511 1092 2512
rect 1055 2510 1093 2511
rect 1055 2502 1119 2510
rect 1055 2482 1064 2502
rect 1084 2488 1119 2502
rect 1139 2488 1142 2508
rect 1084 2483 1142 2488
rect 1084 2482 1119 2483
rect 321 2445 358 2474
rect 322 2443 358 2445
rect 534 2443 571 2474
rect 322 2421 571 2443
rect 742 2442 779 2474
rect 1055 2470 1119 2482
rect 1159 2444 1186 2622
rect 1018 2442 1186 2444
rect 742 2416 1186 2442
rect 1338 2541 1588 2565
rect 1338 2470 1375 2541
rect 1490 2480 1521 2481
rect 1338 2450 1347 2470
rect 1367 2450 1375 2470
rect 1338 2440 1375 2450
rect 1434 2470 1521 2480
rect 1434 2450 1443 2470
rect 1463 2450 1521 2470
rect 1434 2441 1521 2450
rect 1434 2440 1471 2441
rect 742 2406 764 2416
rect 1018 2415 1186 2416
rect 702 2404 764 2406
rect 132 2397 764 2404
rect 131 2388 764 2397
rect 1490 2388 1521 2441
rect 1551 2470 1588 2541
rect 1759 2546 2152 2566
rect 2172 2546 2175 2566
rect 1759 2541 2175 2546
rect 1759 2540 2100 2541
rect 1703 2480 1734 2481
rect 1551 2450 1560 2470
rect 1580 2450 1588 2470
rect 1551 2440 1588 2450
rect 1647 2473 1734 2480
rect 1647 2470 1708 2473
rect 1647 2450 1656 2470
rect 1676 2453 1708 2470
rect 1729 2453 1734 2473
rect 1676 2450 1734 2453
rect 1647 2443 1734 2450
rect 1759 2470 1796 2540
rect 2062 2539 2099 2540
rect 1911 2480 1947 2481
rect 1759 2450 1768 2470
rect 1788 2450 1796 2470
rect 1647 2441 1703 2443
rect 1647 2440 1684 2441
rect 1759 2440 1796 2450
rect 1855 2470 2003 2480
rect 2103 2477 2199 2479
rect 1855 2450 1864 2470
rect 1884 2450 1974 2470
rect 1994 2450 2003 2470
rect 1855 2441 2003 2450
rect 2061 2470 2199 2477
rect 2061 2450 2070 2470
rect 2090 2450 2199 2470
rect 2061 2441 2199 2450
rect 1855 2440 1892 2441
rect 1911 2389 1947 2441
rect 1966 2440 2003 2441
rect 2062 2440 2099 2441
rect 131 2370 141 2388
rect 159 2387 764 2388
rect 1382 2387 1423 2388
rect 159 2382 180 2387
rect 159 2370 171 2382
rect 1274 2380 1423 2387
rect 131 2362 171 2370
rect 214 2369 240 2370
rect 131 2360 168 2362
rect 214 2351 768 2369
rect 1274 2360 1392 2380
rect 1412 2360 1423 2380
rect 1274 2352 1423 2360
rect 1490 2384 1849 2388
rect 1490 2379 1812 2384
rect 1490 2355 1603 2379
rect 1627 2360 1812 2379
rect 1836 2360 1849 2384
rect 1627 2355 1849 2360
rect 1490 2352 1849 2355
rect 1911 2352 1946 2389
rect 2014 2386 2114 2389
rect 2014 2382 2081 2386
rect 2014 2356 2026 2382
rect 2052 2360 2081 2382
rect 2107 2360 2114 2386
rect 2052 2356 2114 2360
rect 2014 2352 2114 2356
rect 134 2292 171 2298
rect 214 2292 240 2351
rect 747 2332 768 2351
rect 134 2289 240 2292
rect 134 2271 143 2289
rect 161 2275 240 2289
rect 325 2307 575 2331
rect 161 2273 237 2275
rect 161 2271 171 2273
rect 134 2261 171 2271
rect 139 2196 170 2261
rect 325 2236 362 2307
rect 477 2246 508 2247
rect 325 2216 334 2236
rect 354 2216 362 2236
rect 325 2206 362 2216
rect 421 2236 508 2246
rect 421 2216 430 2236
rect 450 2216 508 2236
rect 421 2207 508 2216
rect 421 2206 458 2207
rect 138 2187 175 2196
rect 138 2169 148 2187
rect 166 2169 175 2187
rect 138 2159 175 2169
rect 477 2154 508 2207
rect 538 2236 575 2307
rect 746 2312 1139 2332
rect 1159 2312 1162 2332
rect 1490 2331 1521 2352
rect 1911 2331 1947 2352
rect 1333 2330 1370 2331
rect 746 2307 1162 2312
rect 1332 2321 1370 2330
rect 746 2306 1087 2307
rect 690 2246 721 2247
rect 538 2216 547 2236
rect 567 2216 575 2236
rect 538 2206 575 2216
rect 634 2239 721 2246
rect 634 2236 695 2239
rect 634 2216 643 2236
rect 663 2219 695 2236
rect 716 2219 721 2239
rect 663 2216 721 2219
rect 634 2209 721 2216
rect 746 2236 783 2306
rect 1049 2305 1086 2306
rect 1332 2301 1341 2321
rect 1361 2301 1370 2321
rect 1332 2293 1370 2301
rect 1436 2325 1521 2331
rect 1546 2330 1583 2331
rect 1436 2305 1444 2325
rect 1464 2305 1521 2325
rect 1436 2297 1521 2305
rect 1545 2321 1583 2330
rect 1545 2301 1554 2321
rect 1574 2301 1583 2321
rect 1436 2296 1472 2297
rect 1545 2293 1583 2301
rect 1649 2325 1734 2331
rect 1754 2330 1791 2331
rect 1649 2305 1657 2325
rect 1677 2324 1734 2325
rect 1677 2305 1706 2324
rect 1649 2304 1706 2305
rect 1727 2304 1734 2324
rect 1649 2297 1734 2304
rect 1753 2321 1791 2330
rect 1753 2301 1762 2321
rect 1782 2301 1791 2321
rect 1649 2296 1685 2297
rect 1753 2293 1791 2301
rect 1857 2326 2001 2331
rect 1857 2325 1916 2326
rect 1857 2305 1865 2325
rect 1885 2306 1916 2325
rect 1940 2325 2001 2326
rect 1940 2306 1973 2325
rect 1885 2305 1973 2306
rect 1993 2305 2001 2325
rect 1857 2297 2001 2305
rect 1857 2296 1893 2297
rect 1965 2296 2001 2297
rect 2067 2330 2104 2331
rect 2067 2329 2105 2330
rect 2067 2321 2131 2329
rect 2067 2301 2076 2321
rect 2096 2307 2131 2321
rect 2151 2307 2154 2327
rect 2096 2302 2154 2307
rect 2096 2301 2131 2302
rect 1333 2264 1370 2293
rect 1334 2262 1370 2264
rect 1546 2262 1583 2293
rect 898 2246 934 2247
rect 746 2216 755 2236
rect 775 2216 783 2236
rect 634 2207 690 2209
rect 634 2206 671 2207
rect 746 2206 783 2216
rect 842 2236 990 2246
rect 1090 2243 1186 2245
rect 842 2216 851 2236
rect 871 2216 961 2236
rect 981 2216 990 2236
rect 842 2207 990 2216
rect 1048 2236 1186 2243
rect 1334 2240 1583 2262
rect 1754 2261 1791 2293
rect 2067 2289 2131 2301
rect 2171 2263 2198 2441
rect 2030 2261 2198 2263
rect 1754 2257 2198 2261
rect 1048 2216 1057 2236
rect 1077 2216 1186 2236
rect 1754 2238 1803 2257
rect 1823 2238 2198 2257
rect 1754 2235 2198 2238
rect 2030 2234 2198 2235
rect 2219 2260 2250 2654
rect 2219 2234 2224 2260
rect 2243 2234 2250 2260
rect 2219 2231 2250 2234
rect 1048 2207 1186 2216
rect 842 2206 879 2207
rect 898 2155 934 2207
rect 953 2206 990 2207
rect 1049 2206 1086 2207
rect 369 2153 410 2154
rect 261 2146 410 2153
rect 261 2126 379 2146
rect 399 2126 410 2146
rect 261 2118 410 2126
rect 477 2150 836 2154
rect 477 2145 799 2150
rect 477 2121 590 2145
rect 614 2126 799 2145
rect 823 2126 836 2150
rect 614 2121 836 2126
rect 477 2118 836 2121
rect 898 2118 933 2155
rect 1001 2152 1101 2155
rect 1001 2148 1068 2152
rect 1001 2122 1013 2148
rect 1039 2126 1068 2148
rect 1094 2126 1101 2152
rect 1039 2122 1101 2126
rect 1001 2118 1101 2122
rect 477 2097 508 2118
rect 898 2097 934 2118
rect 141 2088 178 2097
rect 320 2096 357 2097
rect 141 2070 150 2088
rect 168 2070 178 2088
rect 141 2060 178 2070
rect 142 2025 178 2060
rect 319 2087 357 2096
rect 319 2067 328 2087
rect 348 2067 357 2087
rect 319 2059 357 2067
rect 423 2091 508 2097
rect 533 2096 570 2097
rect 423 2071 431 2091
rect 451 2071 508 2091
rect 423 2063 508 2071
rect 532 2087 570 2096
rect 532 2067 541 2087
rect 561 2067 570 2087
rect 423 2062 459 2063
rect 532 2059 570 2067
rect 636 2091 721 2097
rect 741 2096 778 2097
rect 636 2071 644 2091
rect 664 2090 721 2091
rect 664 2071 693 2090
rect 636 2070 693 2071
rect 714 2070 721 2090
rect 636 2063 721 2070
rect 740 2087 778 2096
rect 740 2067 749 2087
rect 769 2067 778 2087
rect 636 2062 672 2063
rect 740 2059 778 2067
rect 844 2091 988 2097
rect 844 2071 852 2091
rect 872 2090 960 2091
rect 872 2071 900 2090
rect 844 2069 900 2071
rect 922 2071 960 2090
rect 980 2071 988 2091
rect 922 2069 988 2071
rect 844 2063 988 2069
rect 844 2062 880 2063
rect 952 2062 988 2063
rect 1054 2096 1091 2097
rect 1054 2095 1092 2096
rect 1054 2087 1118 2095
rect 1054 2067 1063 2087
rect 1083 2073 1118 2087
rect 1138 2073 1141 2093
rect 1083 2068 1141 2073
rect 1083 2067 1118 2068
rect 320 2030 357 2059
rect 140 1984 178 2025
rect 321 2028 357 2030
rect 533 2028 570 2059
rect 321 2006 570 2028
rect 741 2027 778 2059
rect 1054 2055 1118 2067
rect 1158 2029 1185 2207
rect 1017 2027 1185 2029
rect 741 2001 1185 2027
rect 742 1984 766 2001
rect 1017 2000 1185 2001
rect 1553 2029 1803 2053
rect 140 1966 767 1984
rect 140 1960 178 1966
rect 142 1914 177 1960
rect 1553 1958 1590 2029
rect 1705 1968 1736 1969
rect 1553 1938 1562 1958
rect 1582 1938 1590 1958
rect 1553 1928 1590 1938
rect 1649 1958 1736 1968
rect 1649 1938 1658 1958
rect 1678 1938 1736 1958
rect 1649 1929 1736 1938
rect 1649 1928 1686 1929
rect 140 1905 177 1914
rect 140 1887 150 1905
rect 168 1887 177 1905
rect 140 1877 177 1887
rect 1705 1876 1736 1929
rect 1766 1958 1803 2029
rect 1974 2034 2367 2054
rect 2387 2034 2390 2054
rect 1974 2029 2390 2034
rect 1974 2028 2315 2029
rect 1918 1968 1949 1969
rect 1766 1938 1775 1958
rect 1795 1938 1803 1958
rect 1766 1928 1803 1938
rect 1862 1961 1949 1968
rect 1862 1958 1923 1961
rect 1862 1938 1871 1958
rect 1891 1941 1923 1958
rect 1944 1941 1949 1961
rect 1891 1938 1949 1941
rect 1862 1931 1949 1938
rect 1974 1958 2011 2028
rect 2277 2027 2314 2028
rect 2126 1968 2162 1969
rect 1974 1938 1983 1958
rect 2003 1938 2011 1958
rect 1862 1929 1918 1931
rect 1862 1928 1899 1929
rect 1974 1928 2011 1938
rect 2070 1958 2218 1968
rect 2318 1965 2414 1967
rect 2070 1938 2079 1958
rect 2099 1938 2189 1958
rect 2209 1938 2218 1958
rect 2070 1929 2218 1938
rect 2276 1958 2414 1965
rect 2276 1938 2285 1958
rect 2305 1938 2414 1958
rect 2276 1929 2414 1938
rect 2070 1928 2107 1929
rect 2126 1877 2162 1929
rect 2181 1928 2218 1929
rect 2277 1928 2314 1929
rect 1597 1875 1638 1876
rect 1489 1868 1638 1875
rect 1489 1848 1607 1868
rect 1627 1848 1638 1868
rect 1489 1840 1638 1848
rect 1705 1872 2064 1876
rect 1705 1867 2027 1872
rect 1705 1843 1818 1867
rect 1842 1848 2027 1867
rect 2051 1848 2064 1872
rect 1842 1843 2064 1848
rect 1705 1840 2064 1843
rect 2126 1840 2161 1877
rect 2229 1874 2329 1877
rect 2229 1870 2296 1874
rect 2229 1844 2241 1870
rect 2267 1848 2296 1870
rect 2322 1848 2329 1874
rect 2267 1844 2329 1848
rect 2229 1840 2329 1844
rect 1705 1819 1736 1840
rect 2126 1819 2162 1840
rect 1548 1818 1585 1819
rect 143 1813 180 1815
rect 143 1812 791 1813
rect 142 1806 791 1812
rect 142 1788 152 1806
rect 170 1792 791 1806
rect 170 1788 180 1792
rect 621 1791 791 1792
rect 142 1778 180 1788
rect 142 1700 177 1778
rect 754 1768 791 1791
rect 1547 1809 1585 1818
rect 1547 1789 1556 1809
rect 1576 1789 1585 1809
rect 1547 1781 1585 1789
rect 1651 1813 1736 1819
rect 1761 1818 1798 1819
rect 1651 1793 1659 1813
rect 1679 1793 1736 1813
rect 1651 1785 1736 1793
rect 1760 1809 1798 1818
rect 1760 1789 1769 1809
rect 1789 1789 1798 1809
rect 1651 1784 1687 1785
rect 1760 1781 1798 1789
rect 1864 1813 1949 1819
rect 1969 1818 2006 1819
rect 1864 1793 1872 1813
rect 1892 1812 1949 1813
rect 1892 1793 1921 1812
rect 1864 1792 1921 1793
rect 1942 1792 1949 1812
rect 1864 1785 1949 1792
rect 1968 1809 2006 1818
rect 1968 1789 1977 1809
rect 1997 1789 2006 1809
rect 1864 1784 1900 1785
rect 1968 1781 2006 1789
rect 2072 1813 2216 1819
rect 2072 1793 2080 1813
rect 2100 1794 2136 1813
rect 2159 1794 2188 1813
rect 2100 1793 2188 1794
rect 2208 1793 2216 1813
rect 2072 1785 2216 1793
rect 2072 1784 2108 1785
rect 2180 1784 2216 1785
rect 2282 1818 2319 1819
rect 2282 1817 2320 1818
rect 2282 1809 2346 1817
rect 2282 1789 2291 1809
rect 2311 1795 2346 1809
rect 2366 1795 2369 1815
rect 2311 1790 2369 1795
rect 2311 1789 2346 1790
rect 138 1691 177 1700
rect 138 1673 148 1691
rect 166 1673 177 1691
rect 138 1667 177 1673
rect 333 1743 583 1767
rect 333 1672 370 1743
rect 485 1682 516 1683
rect 138 1663 175 1667
rect 333 1652 342 1672
rect 362 1652 370 1672
rect 333 1642 370 1652
rect 429 1672 516 1682
rect 429 1652 438 1672
rect 458 1652 516 1672
rect 429 1643 516 1652
rect 429 1642 466 1643
rect 141 1592 178 1601
rect 139 1574 150 1592
rect 168 1574 178 1592
rect 485 1590 516 1643
rect 546 1672 583 1743
rect 754 1748 1147 1768
rect 1167 1748 1170 1768
rect 1548 1752 1585 1781
rect 754 1743 1170 1748
rect 1549 1750 1585 1752
rect 1761 1750 1798 1781
rect 754 1742 1095 1743
rect 698 1682 729 1683
rect 546 1652 555 1672
rect 575 1652 583 1672
rect 546 1642 583 1652
rect 642 1675 729 1682
rect 642 1672 703 1675
rect 642 1652 651 1672
rect 671 1655 703 1672
rect 724 1655 729 1675
rect 671 1652 729 1655
rect 642 1645 729 1652
rect 754 1672 791 1742
rect 1057 1741 1094 1742
rect 1549 1728 1798 1750
rect 1969 1749 2006 1781
rect 2282 1777 2346 1789
rect 2386 1751 2413 1929
rect 2441 1816 2479 3647
rect 2986 3622 2993 3648
rect 3012 3622 3017 3648
rect 2893 3229 2922 3231
rect 2893 3224 2925 3229
rect 2893 3206 2900 3224
rect 2920 3206 2925 3224
rect 2986 3228 3017 3622
rect 3038 3647 3206 3648
rect 3038 3644 3482 3647
rect 3038 3625 3413 3644
rect 3433 3625 3482 3644
rect 4050 3646 4159 3666
rect 4179 3646 4188 3666
rect 3038 3621 3482 3625
rect 3038 3619 3206 3621
rect 3038 3441 3065 3619
rect 3105 3581 3169 3593
rect 3445 3589 3482 3621
rect 3653 3620 3902 3642
rect 4050 3639 4188 3646
rect 4246 3666 4394 3675
rect 4246 3646 4255 3666
rect 4275 3646 4365 3666
rect 4385 3646 4394 3666
rect 4050 3637 4146 3639
rect 4246 3636 4394 3646
rect 4453 3666 4490 3676
rect 4565 3675 4602 3676
rect 4546 3673 4602 3675
rect 4453 3646 4461 3666
rect 4481 3646 4490 3666
rect 4302 3635 4338 3636
rect 3653 3589 3690 3620
rect 3866 3618 3902 3620
rect 3866 3589 3903 3618
rect 3105 3580 3140 3581
rect 3082 3575 3140 3580
rect 3082 3555 3085 3575
rect 3105 3561 3140 3575
rect 3160 3561 3169 3581
rect 3105 3553 3169 3561
rect 3131 3552 3169 3553
rect 3132 3551 3169 3552
rect 3235 3585 3271 3586
rect 3343 3585 3379 3586
rect 3235 3577 3379 3585
rect 3235 3557 3243 3577
rect 3263 3576 3351 3577
rect 3263 3557 3296 3576
rect 3235 3556 3296 3557
rect 3320 3557 3351 3576
rect 3371 3557 3379 3577
rect 3320 3556 3379 3557
rect 3235 3551 3379 3556
rect 3445 3581 3483 3589
rect 3551 3585 3587 3586
rect 3445 3561 3454 3581
rect 3474 3561 3483 3581
rect 3445 3552 3483 3561
rect 3502 3578 3587 3585
rect 3502 3558 3509 3578
rect 3530 3577 3587 3578
rect 3530 3558 3559 3577
rect 3502 3557 3559 3558
rect 3579 3557 3587 3577
rect 3445 3551 3482 3552
rect 3502 3551 3587 3557
rect 3653 3581 3691 3589
rect 3764 3585 3800 3586
rect 3653 3561 3662 3581
rect 3682 3561 3691 3581
rect 3653 3552 3691 3561
rect 3715 3577 3800 3585
rect 3715 3557 3772 3577
rect 3792 3557 3800 3577
rect 3653 3551 3690 3552
rect 3715 3551 3800 3557
rect 3866 3581 3904 3589
rect 3866 3561 3875 3581
rect 3895 3561 3904 3581
rect 4150 3576 4187 3577
rect 4453 3576 4490 3646
rect 4515 3666 4602 3673
rect 4515 3663 4573 3666
rect 4515 3643 4520 3663
rect 4541 3646 4573 3663
rect 4593 3646 4602 3666
rect 4541 3643 4602 3646
rect 4515 3636 4602 3643
rect 4661 3666 4698 3676
rect 4661 3646 4669 3666
rect 4689 3646 4698 3666
rect 4515 3635 4546 3636
rect 4149 3575 4490 3576
rect 3866 3552 3904 3561
rect 4074 3570 4490 3575
rect 3866 3551 3903 3552
rect 3289 3530 3325 3551
rect 3715 3530 3746 3551
rect 4074 3550 4077 3570
rect 4097 3550 4490 3570
rect 4661 3575 4698 3646
rect 4728 3675 4759 3728
rect 5061 3713 5098 3723
rect 5061 3695 5070 3713
rect 5088 3695 5098 3713
rect 5061 3686 5098 3695
rect 4778 3675 4815 3676
rect 4728 3666 4815 3675
rect 4728 3646 4786 3666
rect 4806 3646 4815 3666
rect 4728 3636 4815 3646
rect 4874 3666 4911 3676
rect 4874 3646 4882 3666
rect 4902 3646 4911 3666
rect 4728 3635 4759 3636
rect 4874 3575 4911 3646
rect 5066 3621 5097 3686
rect 5065 3611 5102 3621
rect 5065 3609 5075 3611
rect 4999 3607 5075 3609
rect 4661 3551 4911 3575
rect 4996 3593 5075 3607
rect 5093 3593 5102 3611
rect 4996 3590 5102 3593
rect 4468 3531 4489 3550
rect 4996 3531 5022 3590
rect 5065 3584 5102 3590
rect 3122 3526 3222 3530
rect 3122 3522 3184 3526
rect 3122 3496 3129 3522
rect 3155 3500 3184 3522
rect 3210 3500 3222 3526
rect 3155 3496 3222 3500
rect 3122 3493 3222 3496
rect 3290 3493 3325 3530
rect 3387 3527 3746 3530
rect 3387 3522 3609 3527
rect 3387 3498 3400 3522
rect 3424 3503 3609 3522
rect 3633 3503 3746 3527
rect 3424 3498 3746 3503
rect 3387 3494 3746 3498
rect 3813 3522 3962 3530
rect 3813 3502 3824 3522
rect 3844 3502 3962 3522
rect 4468 3513 5022 3531
rect 5068 3520 5105 3522
rect 4996 3512 5022 3513
rect 5065 3512 5105 3520
rect 3813 3495 3962 3502
rect 5065 3500 5077 3512
rect 5056 3495 5077 3500
rect 3813 3494 3854 3495
rect 4472 3494 5077 3495
rect 5095 3494 5105 3512
rect 3137 3441 3174 3442
rect 3233 3441 3270 3442
rect 3289 3441 3325 3493
rect 3344 3441 3381 3442
rect 3037 3432 3175 3441
rect 3037 3412 3146 3432
rect 3166 3412 3175 3432
rect 3037 3405 3175 3412
rect 3233 3432 3381 3441
rect 3233 3412 3242 3432
rect 3262 3412 3352 3432
rect 3372 3412 3381 3432
rect 3037 3403 3133 3405
rect 3233 3402 3381 3412
rect 3440 3432 3477 3442
rect 3552 3441 3589 3442
rect 3533 3439 3589 3441
rect 3440 3412 3448 3432
rect 3468 3412 3477 3432
rect 3289 3401 3325 3402
rect 3137 3342 3174 3343
rect 3440 3342 3477 3412
rect 3502 3432 3589 3439
rect 3502 3429 3560 3432
rect 3502 3409 3507 3429
rect 3528 3412 3560 3429
rect 3580 3412 3589 3432
rect 3528 3409 3589 3412
rect 3502 3402 3589 3409
rect 3648 3432 3685 3442
rect 3648 3412 3656 3432
rect 3676 3412 3685 3432
rect 3502 3401 3533 3402
rect 3136 3341 3477 3342
rect 3061 3336 3477 3341
rect 3061 3316 3064 3336
rect 3084 3316 3477 3336
rect 3648 3341 3685 3412
rect 3715 3441 3746 3494
rect 4472 3485 5105 3494
rect 4472 3478 5104 3485
rect 4472 3476 4534 3478
rect 4050 3466 4218 3467
rect 4472 3466 4494 3476
rect 3765 3441 3802 3442
rect 3715 3432 3802 3441
rect 3715 3412 3773 3432
rect 3793 3412 3802 3432
rect 3715 3402 3802 3412
rect 3861 3432 3898 3442
rect 3861 3412 3869 3432
rect 3889 3412 3898 3432
rect 3715 3401 3746 3402
rect 3861 3341 3898 3412
rect 3648 3317 3898 3341
rect 4050 3440 4494 3466
rect 4050 3438 4218 3440
rect 4050 3260 4077 3438
rect 4117 3400 4181 3412
rect 4457 3408 4494 3440
rect 4665 3439 4914 3461
rect 4665 3408 4702 3439
rect 4878 3437 4914 3439
rect 4878 3408 4915 3437
rect 4117 3399 4152 3400
rect 4094 3394 4152 3399
rect 4094 3374 4097 3394
rect 4117 3380 4152 3394
rect 4172 3380 4181 3400
rect 4117 3372 4181 3380
rect 4143 3371 4181 3372
rect 4144 3370 4181 3371
rect 4247 3404 4283 3405
rect 4355 3404 4391 3405
rect 4247 3396 4391 3404
rect 4247 3376 4255 3396
rect 4275 3376 4304 3396
rect 4247 3375 4304 3376
rect 4326 3376 4363 3396
rect 4383 3376 4391 3396
rect 4326 3375 4391 3376
rect 4247 3370 4391 3375
rect 4457 3400 4495 3408
rect 4563 3404 4599 3405
rect 4457 3380 4466 3400
rect 4486 3380 4495 3400
rect 4457 3371 4495 3380
rect 4514 3397 4599 3404
rect 4514 3377 4521 3397
rect 4542 3396 4599 3397
rect 4542 3377 4571 3396
rect 4514 3376 4571 3377
rect 4591 3376 4599 3396
rect 4457 3370 4494 3371
rect 4514 3370 4599 3376
rect 4665 3400 4703 3408
rect 4776 3404 4812 3405
rect 4665 3380 4674 3400
rect 4694 3380 4703 3400
rect 4665 3371 4703 3380
rect 4727 3396 4812 3404
rect 4727 3376 4784 3396
rect 4804 3376 4812 3396
rect 4665 3370 4702 3371
rect 4727 3370 4812 3376
rect 4878 3400 4916 3408
rect 4878 3380 4887 3400
rect 4907 3380 4916 3400
rect 4878 3371 4916 3380
rect 4878 3370 4915 3371
rect 4301 3349 4337 3370
rect 4727 3349 4758 3370
rect 4134 3345 4234 3349
rect 4134 3341 4196 3345
rect 4134 3315 4141 3341
rect 4167 3319 4196 3341
rect 4222 3319 4234 3345
rect 4167 3315 4234 3319
rect 4134 3312 4234 3315
rect 4302 3312 4337 3349
rect 4399 3346 4758 3349
rect 4399 3341 4621 3346
rect 4399 3317 4412 3341
rect 4436 3322 4621 3341
rect 4645 3322 4758 3346
rect 4436 3317 4758 3322
rect 4399 3313 4758 3317
rect 4825 3341 4974 3349
rect 4825 3321 4836 3341
rect 4856 3321 4974 3341
rect 4825 3314 4974 3321
rect 5065 3329 5104 3478
rect 4825 3313 4866 3314
rect 4149 3260 4186 3261
rect 4245 3260 4282 3261
rect 4301 3260 4337 3312
rect 4356 3260 4393 3261
rect 4049 3251 4187 3260
rect 4049 3231 4158 3251
rect 4178 3231 4187 3251
rect 2986 3227 3156 3228
rect 2986 3212 3432 3227
rect 4049 3224 4187 3231
rect 4245 3251 4393 3260
rect 4245 3231 4254 3251
rect 4274 3231 4364 3251
rect 4384 3231 4393 3251
rect 4049 3222 4145 3224
rect 2893 3201 2925 3206
rect 2895 2200 2925 3201
rect 2988 3201 3432 3212
rect 2988 3199 3156 3201
rect 2988 3021 3015 3199
rect 3055 3161 3119 3173
rect 3395 3169 3432 3201
rect 3603 3200 3852 3222
rect 4245 3221 4393 3231
rect 4452 3251 4489 3261
rect 4564 3260 4601 3261
rect 4545 3258 4601 3260
rect 4452 3231 4460 3251
rect 4480 3231 4489 3251
rect 4301 3220 4337 3221
rect 3603 3169 3640 3200
rect 3816 3198 3852 3200
rect 3816 3169 3853 3198
rect 3055 3160 3090 3161
rect 3032 3155 3090 3160
rect 3032 3135 3035 3155
rect 3055 3141 3090 3155
rect 3110 3141 3119 3161
rect 3055 3133 3119 3141
rect 3081 3132 3119 3133
rect 3082 3131 3119 3132
rect 3185 3165 3221 3166
rect 3293 3165 3329 3166
rect 3185 3157 3329 3165
rect 3185 3137 3193 3157
rect 3213 3138 3245 3157
rect 3268 3138 3301 3157
rect 3213 3137 3301 3138
rect 3321 3137 3329 3157
rect 3185 3131 3329 3137
rect 3395 3161 3433 3169
rect 3501 3165 3537 3166
rect 3395 3141 3404 3161
rect 3424 3141 3433 3161
rect 3395 3132 3433 3141
rect 3452 3158 3537 3165
rect 3452 3138 3459 3158
rect 3480 3157 3537 3158
rect 3480 3138 3509 3157
rect 3452 3137 3509 3138
rect 3529 3137 3537 3157
rect 3395 3131 3432 3132
rect 3452 3131 3537 3137
rect 3603 3161 3641 3169
rect 3714 3165 3750 3166
rect 3603 3141 3612 3161
rect 3632 3141 3641 3161
rect 3603 3132 3641 3141
rect 3665 3157 3750 3165
rect 3665 3137 3722 3157
rect 3742 3137 3750 3157
rect 3603 3131 3640 3132
rect 3665 3131 3750 3137
rect 3816 3161 3854 3169
rect 4149 3161 4186 3162
rect 4452 3161 4489 3231
rect 4514 3251 4601 3258
rect 4514 3248 4572 3251
rect 4514 3228 4519 3248
rect 4540 3231 4572 3248
rect 4592 3231 4601 3251
rect 4540 3228 4601 3231
rect 4514 3221 4601 3228
rect 4660 3251 4697 3261
rect 4660 3231 4668 3251
rect 4688 3231 4697 3251
rect 4514 3220 4545 3221
rect 3816 3141 3825 3161
rect 3845 3141 3854 3161
rect 4148 3160 4489 3161
rect 3816 3132 3854 3141
rect 4073 3155 4489 3160
rect 4073 3135 4076 3155
rect 4096 3135 4489 3155
rect 4660 3160 4697 3231
rect 4727 3260 4758 3313
rect 5065 3311 5075 3329
rect 5093 3311 5104 3329
rect 5065 3302 5102 3311
rect 4777 3260 4814 3261
rect 4727 3251 4814 3260
rect 4727 3231 4785 3251
rect 4805 3231 4814 3251
rect 4727 3221 4814 3231
rect 4873 3251 4910 3261
rect 4873 3231 4881 3251
rect 4901 3231 4910 3251
rect 5068 3236 5105 3240
rect 4727 3220 4758 3221
rect 4873 3160 4910 3231
rect 4660 3136 4910 3160
rect 5066 3230 5105 3236
rect 5066 3212 5077 3230
rect 5095 3212 5105 3230
rect 5066 3203 5105 3212
rect 3816 3131 3853 3132
rect 3239 3110 3275 3131
rect 3665 3110 3696 3131
rect 4452 3112 4489 3135
rect 5066 3125 5101 3203
rect 5063 3115 5101 3125
rect 4452 3111 4622 3112
rect 5063 3111 5073 3115
rect 3072 3106 3172 3110
rect 3072 3102 3134 3106
rect 3072 3076 3079 3102
rect 3105 3080 3134 3102
rect 3160 3080 3172 3106
rect 3105 3076 3172 3080
rect 3072 3073 3172 3076
rect 3240 3073 3275 3110
rect 3337 3107 3696 3110
rect 3337 3102 3559 3107
rect 3337 3078 3350 3102
rect 3374 3083 3559 3102
rect 3583 3083 3696 3107
rect 3374 3078 3696 3083
rect 3337 3074 3696 3078
rect 3763 3102 3912 3110
rect 3763 3082 3774 3102
rect 3794 3082 3912 3102
rect 4452 3097 5073 3111
rect 5091 3097 5101 3115
rect 4452 3091 5101 3097
rect 4452 3090 5100 3091
rect 5063 3088 5100 3090
rect 3763 3075 3912 3082
rect 3763 3074 3804 3075
rect 3087 3021 3124 3022
rect 3183 3021 3220 3022
rect 3239 3021 3275 3073
rect 3294 3021 3331 3022
rect 2987 3012 3125 3021
rect 2987 2992 3096 3012
rect 3116 2992 3125 3012
rect 2987 2985 3125 2992
rect 3183 3012 3331 3021
rect 3183 2992 3192 3012
rect 3212 2992 3302 3012
rect 3322 2992 3331 3012
rect 2987 2983 3083 2985
rect 3183 2982 3331 2992
rect 3390 3012 3427 3022
rect 3502 3021 3539 3022
rect 3483 3019 3539 3021
rect 3390 2992 3398 3012
rect 3418 2992 3427 3012
rect 3239 2981 3275 2982
rect 3087 2922 3124 2923
rect 3390 2922 3427 2992
rect 3452 3012 3539 3019
rect 3452 3009 3510 3012
rect 3452 2989 3457 3009
rect 3478 2992 3510 3009
rect 3530 2992 3539 3012
rect 3478 2989 3539 2992
rect 3452 2982 3539 2989
rect 3598 3012 3635 3022
rect 3598 2992 3606 3012
rect 3626 2992 3635 3012
rect 3452 2981 3483 2982
rect 3086 2921 3427 2922
rect 3011 2916 3427 2921
rect 3011 2896 3014 2916
rect 3034 2896 3427 2916
rect 3598 2921 3635 2992
rect 3665 3021 3696 3074
rect 3715 3021 3752 3022
rect 3665 3012 3752 3021
rect 3665 2992 3723 3012
rect 3743 2992 3752 3012
rect 3665 2982 3752 2992
rect 3811 3012 3848 3022
rect 3811 2992 3819 3012
rect 3839 2992 3848 3012
rect 3665 2981 3696 2982
rect 3811 2921 3848 2992
rect 5066 3016 5103 3026
rect 5066 2998 5075 3016
rect 5093 2998 5103 3016
rect 5066 2989 5103 2998
rect 5066 2965 5101 2989
rect 5064 2941 5101 2965
rect 5063 2935 5101 2941
rect 3598 2897 3848 2921
rect 4474 2917 5101 2935
rect 4056 2900 4224 2901
rect 4475 2900 4499 2917
rect 4056 2874 4500 2900
rect 4056 2872 4224 2874
rect 4056 2694 4083 2872
rect 4123 2834 4187 2846
rect 4463 2842 4500 2874
rect 4671 2873 4920 2895
rect 4671 2842 4708 2873
rect 4884 2871 4920 2873
rect 5063 2876 5101 2917
rect 4884 2842 4921 2871
rect 4123 2833 4158 2834
rect 4100 2828 4158 2833
rect 4100 2808 4103 2828
rect 4123 2814 4158 2828
rect 4178 2814 4187 2834
rect 4123 2806 4187 2814
rect 4149 2805 4187 2806
rect 4150 2804 4187 2805
rect 4253 2838 4289 2839
rect 4361 2838 4397 2839
rect 4253 2832 4397 2838
rect 4253 2830 4319 2832
rect 4253 2810 4261 2830
rect 4281 2811 4319 2830
rect 4341 2830 4397 2832
rect 4341 2811 4369 2830
rect 4281 2810 4369 2811
rect 4389 2810 4397 2830
rect 4253 2804 4397 2810
rect 4463 2834 4501 2842
rect 4569 2838 4605 2839
rect 4463 2814 4472 2834
rect 4492 2814 4501 2834
rect 4463 2805 4501 2814
rect 4520 2831 4605 2838
rect 4520 2811 4527 2831
rect 4548 2830 4605 2831
rect 4548 2811 4577 2830
rect 4520 2810 4577 2811
rect 4597 2810 4605 2830
rect 4463 2804 4500 2805
rect 4520 2804 4605 2810
rect 4671 2834 4709 2842
rect 4782 2838 4818 2839
rect 4671 2814 4680 2834
rect 4700 2814 4709 2834
rect 4671 2805 4709 2814
rect 4733 2830 4818 2838
rect 4733 2810 4790 2830
rect 4810 2810 4818 2830
rect 4671 2804 4708 2805
rect 4733 2804 4818 2810
rect 4884 2834 4922 2842
rect 4884 2814 4893 2834
rect 4913 2814 4922 2834
rect 4884 2805 4922 2814
rect 5063 2841 5099 2876
rect 5063 2831 5100 2841
rect 5063 2813 5073 2831
rect 5091 2813 5100 2831
rect 4884 2804 4921 2805
rect 5063 2804 5100 2813
rect 4307 2783 4343 2804
rect 4733 2783 4764 2804
rect 4140 2779 4240 2783
rect 4140 2775 4202 2779
rect 4140 2749 4147 2775
rect 4173 2753 4202 2775
rect 4228 2753 4240 2779
rect 4173 2749 4240 2753
rect 4140 2746 4240 2749
rect 4308 2746 4343 2783
rect 4405 2780 4764 2783
rect 4405 2775 4627 2780
rect 4405 2751 4418 2775
rect 4442 2756 4627 2775
rect 4651 2756 4764 2780
rect 4442 2751 4764 2756
rect 4405 2747 4764 2751
rect 4831 2775 4980 2783
rect 4831 2755 4842 2775
rect 4862 2755 4980 2775
rect 4831 2748 4980 2755
rect 4831 2747 4872 2748
rect 4155 2694 4192 2695
rect 4251 2694 4288 2695
rect 4307 2694 4343 2746
rect 4362 2694 4399 2695
rect 4055 2685 4193 2694
rect 3043 2666 3211 2667
rect 3043 2663 3487 2666
rect 3043 2644 3418 2663
rect 3438 2644 3487 2663
rect 4055 2665 4164 2685
rect 4184 2665 4193 2685
rect 3043 2640 3487 2644
rect 3043 2638 3211 2640
rect 3043 2460 3070 2638
rect 3110 2600 3174 2612
rect 3450 2608 3487 2640
rect 3658 2639 3907 2661
rect 4055 2658 4193 2665
rect 4251 2685 4399 2694
rect 4251 2665 4260 2685
rect 4280 2665 4370 2685
rect 4390 2665 4399 2685
rect 4055 2656 4151 2658
rect 4251 2655 4399 2665
rect 4458 2685 4495 2695
rect 4570 2694 4607 2695
rect 4551 2692 4607 2694
rect 4458 2665 4466 2685
rect 4486 2665 4495 2685
rect 4307 2654 4343 2655
rect 3658 2608 3695 2639
rect 3871 2637 3907 2639
rect 3871 2608 3908 2637
rect 3110 2599 3145 2600
rect 3087 2594 3145 2599
rect 3087 2574 3090 2594
rect 3110 2580 3145 2594
rect 3165 2580 3174 2600
rect 3110 2572 3174 2580
rect 3136 2571 3174 2572
rect 3137 2570 3174 2571
rect 3240 2604 3276 2605
rect 3348 2604 3384 2605
rect 3240 2596 3384 2604
rect 3240 2576 3248 2596
rect 3268 2576 3300 2596
rect 3324 2576 3356 2596
rect 3376 2576 3384 2596
rect 3240 2570 3384 2576
rect 3450 2600 3488 2608
rect 3556 2604 3592 2605
rect 3450 2580 3459 2600
rect 3479 2580 3488 2600
rect 3450 2571 3488 2580
rect 3507 2597 3592 2604
rect 3507 2577 3514 2597
rect 3535 2596 3592 2597
rect 3535 2577 3564 2596
rect 3507 2576 3564 2577
rect 3584 2576 3592 2596
rect 3450 2570 3487 2571
rect 3507 2570 3592 2576
rect 3658 2600 3696 2608
rect 3769 2604 3805 2605
rect 3658 2580 3667 2600
rect 3687 2580 3696 2600
rect 3658 2571 3696 2580
rect 3720 2596 3805 2604
rect 3720 2576 3777 2596
rect 3797 2576 3805 2596
rect 3658 2570 3695 2571
rect 3720 2570 3805 2576
rect 3871 2600 3909 2608
rect 3871 2580 3880 2600
rect 3900 2580 3909 2600
rect 4155 2595 4192 2596
rect 4458 2595 4495 2665
rect 4520 2685 4607 2692
rect 4520 2682 4578 2685
rect 4520 2662 4525 2682
rect 4546 2665 4578 2682
rect 4598 2665 4607 2685
rect 4546 2662 4607 2665
rect 4520 2655 4607 2662
rect 4666 2685 4703 2695
rect 4666 2665 4674 2685
rect 4694 2665 4703 2685
rect 4520 2654 4551 2655
rect 4154 2594 4495 2595
rect 3871 2571 3909 2580
rect 4079 2589 4495 2594
rect 3871 2570 3908 2571
rect 3294 2549 3330 2570
rect 3720 2549 3751 2570
rect 4079 2569 4082 2589
rect 4102 2569 4495 2589
rect 4666 2594 4703 2665
rect 4733 2694 4764 2747
rect 5066 2732 5103 2742
rect 5066 2714 5075 2732
rect 5093 2714 5103 2732
rect 5066 2705 5103 2714
rect 4783 2694 4820 2695
rect 4733 2685 4820 2694
rect 4733 2665 4791 2685
rect 4811 2665 4820 2685
rect 4733 2655 4820 2665
rect 4879 2685 4916 2695
rect 4879 2665 4887 2685
rect 4907 2665 4916 2685
rect 4733 2654 4764 2655
rect 4879 2594 4916 2665
rect 5071 2640 5102 2705
rect 5070 2630 5107 2640
rect 5070 2628 5080 2630
rect 5004 2626 5080 2628
rect 4666 2570 4916 2594
rect 5001 2612 5080 2626
rect 5098 2612 5107 2630
rect 5001 2609 5107 2612
rect 4473 2550 4494 2569
rect 5001 2550 5027 2609
rect 5070 2603 5107 2609
rect 3127 2545 3227 2549
rect 3127 2541 3189 2545
rect 3127 2515 3134 2541
rect 3160 2519 3189 2541
rect 3215 2519 3227 2545
rect 3160 2515 3227 2519
rect 3127 2512 3227 2515
rect 3295 2512 3330 2549
rect 3392 2546 3751 2549
rect 3392 2541 3614 2546
rect 3392 2517 3405 2541
rect 3429 2522 3614 2541
rect 3638 2522 3751 2546
rect 3429 2517 3751 2522
rect 3392 2513 3751 2517
rect 3818 2541 3967 2549
rect 3818 2521 3829 2541
rect 3849 2521 3967 2541
rect 4473 2532 5027 2550
rect 5073 2539 5110 2541
rect 5001 2531 5027 2532
rect 5070 2531 5110 2539
rect 3818 2514 3967 2521
rect 5070 2519 5082 2531
rect 5061 2514 5082 2519
rect 3818 2513 3859 2514
rect 4477 2513 5082 2514
rect 5100 2513 5110 2531
rect 3142 2460 3179 2461
rect 3238 2460 3275 2461
rect 3294 2460 3330 2512
rect 3349 2460 3386 2461
rect 3042 2451 3180 2460
rect 3042 2431 3151 2451
rect 3171 2431 3180 2451
rect 3042 2424 3180 2431
rect 3238 2451 3386 2460
rect 3238 2431 3247 2451
rect 3267 2431 3357 2451
rect 3377 2431 3386 2451
rect 3042 2422 3138 2424
rect 3238 2421 3386 2431
rect 3445 2451 3482 2461
rect 3557 2460 3594 2461
rect 3538 2458 3594 2460
rect 3445 2431 3453 2451
rect 3473 2431 3482 2451
rect 3294 2420 3330 2421
rect 3142 2361 3179 2362
rect 3445 2361 3482 2431
rect 3507 2451 3594 2458
rect 3507 2448 3565 2451
rect 3507 2428 3512 2448
rect 3533 2431 3565 2448
rect 3585 2431 3594 2451
rect 3533 2428 3594 2431
rect 3507 2421 3594 2428
rect 3653 2451 3690 2461
rect 3653 2431 3661 2451
rect 3681 2431 3690 2451
rect 3507 2420 3538 2421
rect 3141 2360 3482 2361
rect 3066 2355 3482 2360
rect 3066 2335 3069 2355
rect 3089 2335 3482 2355
rect 3653 2360 3690 2431
rect 3720 2460 3751 2513
rect 4477 2504 5110 2513
rect 4477 2497 5109 2504
rect 4477 2495 4539 2497
rect 4055 2485 4223 2486
rect 4477 2485 4499 2495
rect 3770 2460 3807 2461
rect 3720 2451 3807 2460
rect 3720 2431 3778 2451
rect 3798 2431 3807 2451
rect 3720 2421 3807 2431
rect 3866 2451 3903 2461
rect 3866 2431 3874 2451
rect 3894 2431 3903 2451
rect 3720 2420 3751 2421
rect 3866 2360 3903 2431
rect 3653 2336 3903 2360
rect 4055 2459 4499 2485
rect 4055 2457 4223 2459
rect 4055 2279 4082 2457
rect 4122 2419 4186 2431
rect 4462 2427 4499 2459
rect 4670 2458 4919 2480
rect 4670 2427 4707 2458
rect 4883 2456 4919 2458
rect 4883 2427 4920 2456
rect 4122 2418 4157 2419
rect 4099 2413 4157 2418
rect 4099 2393 4102 2413
rect 4122 2399 4157 2413
rect 4177 2399 4186 2419
rect 4122 2391 4186 2399
rect 4148 2390 4186 2391
rect 4149 2389 4186 2390
rect 4252 2423 4288 2424
rect 4360 2423 4396 2424
rect 4252 2415 4396 2423
rect 4252 2395 4260 2415
rect 4280 2395 4309 2415
rect 4252 2394 4309 2395
rect 4331 2395 4368 2415
rect 4388 2395 4396 2415
rect 4331 2394 4396 2395
rect 4252 2389 4396 2394
rect 4462 2419 4500 2427
rect 4568 2423 4604 2424
rect 4462 2399 4471 2419
rect 4491 2399 4500 2419
rect 4462 2390 4500 2399
rect 4519 2416 4604 2423
rect 4519 2396 4526 2416
rect 4547 2415 4604 2416
rect 4547 2396 4576 2415
rect 4519 2395 4576 2396
rect 4596 2395 4604 2415
rect 4462 2389 4499 2390
rect 4519 2389 4604 2395
rect 4670 2419 4708 2427
rect 4781 2423 4817 2424
rect 4670 2399 4679 2419
rect 4699 2399 4708 2419
rect 4670 2390 4708 2399
rect 4732 2415 4817 2423
rect 4732 2395 4789 2415
rect 4809 2395 4817 2415
rect 4670 2389 4707 2390
rect 4732 2389 4817 2395
rect 4883 2419 4921 2427
rect 4883 2399 4892 2419
rect 4912 2399 4921 2419
rect 4883 2390 4921 2399
rect 4883 2389 4920 2390
rect 4306 2368 4342 2389
rect 4732 2368 4763 2389
rect 4139 2364 4239 2368
rect 4139 2360 4201 2364
rect 4139 2334 4146 2360
rect 4172 2338 4201 2360
rect 4227 2338 4239 2364
rect 4172 2334 4239 2338
rect 4139 2331 4239 2334
rect 4307 2331 4342 2368
rect 4404 2365 4763 2368
rect 4404 2360 4626 2365
rect 4404 2336 4417 2360
rect 4441 2341 4626 2360
rect 4650 2341 4763 2365
rect 4441 2336 4763 2341
rect 4404 2332 4763 2336
rect 4830 2360 4979 2368
rect 4830 2340 4841 2360
rect 4861 2340 4979 2360
rect 4830 2333 4979 2340
rect 5070 2348 5109 2497
rect 4830 2332 4871 2333
rect 4154 2279 4191 2280
rect 4250 2279 4287 2280
rect 4306 2279 4342 2331
rect 4361 2279 4398 2280
rect 4054 2270 4192 2279
rect 4054 2250 4163 2270
rect 4183 2250 4192 2270
rect 4054 2243 4192 2250
rect 4250 2270 4398 2279
rect 4250 2250 4259 2270
rect 4279 2250 4369 2270
rect 4389 2250 4398 2270
rect 4054 2241 4150 2243
rect 4250 2240 4398 2250
rect 4457 2270 4494 2280
rect 4569 2279 4606 2280
rect 4550 2277 4606 2279
rect 4457 2250 4465 2270
rect 4485 2250 4494 2270
rect 4306 2239 4342 2240
rect 2835 2199 3003 2200
rect 2835 2173 3279 2199
rect 2835 2171 3003 2173
rect 2835 1993 2862 2171
rect 2902 2133 2966 2145
rect 3242 2141 3279 2173
rect 3450 2172 3699 2194
rect 4154 2180 4191 2181
rect 4457 2180 4494 2250
rect 4519 2270 4606 2277
rect 4519 2267 4577 2270
rect 4519 2247 4524 2267
rect 4545 2250 4577 2267
rect 4597 2250 4606 2270
rect 4545 2247 4606 2250
rect 4519 2240 4606 2247
rect 4665 2270 4702 2280
rect 4665 2250 4673 2270
rect 4693 2250 4702 2270
rect 4519 2239 4550 2240
rect 4153 2179 4494 2180
rect 3450 2141 3487 2172
rect 3663 2170 3699 2172
rect 4078 2174 4494 2179
rect 3663 2141 3700 2170
rect 4078 2154 4081 2174
rect 4101 2154 4494 2174
rect 4665 2179 4702 2250
rect 4732 2279 4763 2332
rect 5070 2330 5080 2348
rect 5098 2330 5109 2348
rect 5070 2321 5107 2330
rect 4782 2279 4819 2280
rect 4732 2270 4819 2279
rect 4732 2250 4790 2270
rect 4810 2250 4819 2270
rect 4732 2240 4819 2250
rect 4878 2270 4915 2280
rect 4878 2250 4886 2270
rect 4906 2250 4915 2270
rect 5073 2255 5110 2259
rect 4732 2239 4763 2240
rect 4878 2179 4915 2250
rect 4665 2155 4915 2179
rect 5071 2249 5110 2255
rect 5071 2231 5082 2249
rect 5100 2231 5110 2249
rect 5071 2222 5110 2231
rect 2902 2132 2937 2133
rect 2879 2127 2937 2132
rect 2879 2107 2882 2127
rect 2902 2113 2937 2127
rect 2957 2113 2966 2133
rect 2902 2105 2966 2113
rect 2928 2104 2966 2105
rect 2929 2103 2966 2104
rect 3032 2137 3068 2138
rect 3140 2137 3176 2138
rect 3032 2131 3176 2137
rect 3032 2129 3093 2131
rect 3032 2109 3040 2129
rect 3060 2109 3093 2129
rect 3032 2105 3093 2109
rect 3118 2129 3176 2131
rect 3118 2109 3148 2129
rect 3168 2109 3176 2129
rect 3118 2105 3176 2109
rect 3032 2103 3176 2105
rect 3242 2133 3280 2141
rect 3348 2137 3384 2138
rect 3242 2113 3251 2133
rect 3271 2113 3280 2133
rect 3242 2104 3280 2113
rect 3299 2130 3384 2137
rect 3299 2110 3306 2130
rect 3327 2129 3384 2130
rect 3327 2110 3356 2129
rect 3299 2109 3356 2110
rect 3376 2109 3384 2129
rect 3242 2103 3279 2104
rect 3299 2103 3384 2109
rect 3450 2133 3488 2141
rect 3561 2137 3597 2138
rect 3450 2113 3459 2133
rect 3479 2113 3488 2133
rect 3450 2104 3488 2113
rect 3512 2129 3597 2137
rect 3512 2109 3569 2129
rect 3589 2109 3597 2129
rect 3450 2103 3487 2104
rect 3512 2103 3597 2109
rect 3663 2133 3701 2141
rect 3663 2113 3672 2133
rect 3692 2113 3701 2133
rect 3663 2104 3701 2113
rect 4457 2131 4494 2154
rect 5071 2144 5106 2222
rect 5068 2134 5106 2144
rect 4457 2130 4627 2131
rect 5068 2130 5078 2134
rect 4457 2116 5078 2130
rect 5096 2116 5106 2134
rect 4457 2110 5106 2116
rect 4457 2109 5105 2110
rect 5068 2107 5105 2109
rect 3663 2103 3700 2104
rect 3086 2082 3122 2103
rect 3512 2082 3543 2103
rect 2919 2078 3019 2082
rect 2919 2074 2981 2078
rect 2919 2048 2926 2074
rect 2952 2052 2981 2074
rect 3007 2052 3019 2078
rect 2952 2048 3019 2052
rect 2919 2045 3019 2048
rect 3087 2045 3122 2082
rect 3184 2079 3543 2082
rect 3184 2074 3406 2079
rect 3184 2050 3197 2074
rect 3221 2055 3406 2074
rect 3430 2055 3543 2079
rect 3221 2050 3543 2055
rect 3184 2046 3543 2050
rect 3610 2074 3759 2082
rect 3610 2054 3621 2074
rect 3641 2054 3759 2074
rect 3610 2047 3759 2054
rect 3610 2046 3651 2047
rect 2934 1993 2971 1994
rect 3030 1993 3067 1994
rect 3086 1993 3122 2045
rect 3141 1993 3178 1994
rect 2834 1984 2972 1993
rect 2834 1964 2943 1984
rect 2963 1964 2972 1984
rect 2834 1957 2972 1964
rect 3030 1984 3178 1993
rect 3030 1964 3039 1984
rect 3059 1964 3149 1984
rect 3169 1964 3178 1984
rect 2834 1955 2930 1957
rect 3030 1954 3178 1964
rect 3237 1984 3274 1994
rect 3349 1993 3386 1994
rect 3330 1991 3386 1993
rect 3237 1964 3245 1984
rect 3265 1964 3274 1984
rect 3086 1953 3122 1954
rect 2934 1894 2971 1895
rect 3237 1894 3274 1964
rect 3299 1984 3386 1991
rect 3299 1981 3357 1984
rect 3299 1961 3304 1981
rect 3325 1964 3357 1981
rect 3377 1964 3386 1984
rect 3325 1961 3386 1964
rect 3299 1954 3386 1961
rect 3445 1984 3482 1994
rect 3445 1964 3453 1984
rect 3473 1964 3482 1984
rect 3299 1953 3330 1954
rect 2933 1893 3274 1894
rect 2858 1888 3274 1893
rect 2858 1868 2861 1888
rect 2881 1868 3274 1888
rect 3445 1893 3482 1964
rect 3512 1993 3543 2046
rect 5071 2035 5108 2045
rect 5071 2017 5080 2035
rect 5098 2017 5108 2035
rect 5071 2008 5108 2017
rect 3562 1993 3599 1994
rect 3512 1984 3599 1993
rect 3512 1964 3570 1984
rect 3590 1964 3599 1984
rect 3512 1954 3599 1964
rect 3658 1984 3695 1994
rect 3658 1964 3666 1984
rect 3686 1964 3695 1984
rect 3512 1953 3543 1954
rect 3658 1893 3695 1964
rect 5071 1962 5106 2008
rect 5070 1956 5108 1962
rect 4481 1938 5108 1956
rect 3445 1869 3695 1893
rect 4063 1921 4231 1922
rect 4482 1921 4506 1938
rect 4063 1895 4507 1921
rect 4063 1893 4231 1895
rect 2443 1756 2476 1816
rect 2245 1749 2413 1751
rect 1969 1723 2413 1749
rect 2245 1722 2413 1723
rect 2442 1745 2479 1756
rect 2442 1726 2448 1745
rect 2471 1726 2479 1745
rect 906 1682 942 1683
rect 754 1652 763 1672
rect 783 1652 791 1672
rect 642 1643 698 1645
rect 642 1642 679 1643
rect 754 1642 791 1652
rect 850 1672 998 1682
rect 1098 1679 1194 1681
rect 850 1652 859 1672
rect 879 1652 969 1672
rect 989 1652 998 1672
rect 850 1643 998 1652
rect 1056 1672 1194 1679
rect 1056 1652 1065 1672
rect 1085 1652 1194 1672
rect 1056 1643 1194 1652
rect 850 1642 887 1643
rect 906 1591 942 1643
rect 961 1642 998 1643
rect 1057 1642 1094 1643
rect 377 1589 418 1590
rect 139 1425 178 1574
rect 269 1582 418 1589
rect 269 1562 387 1582
rect 407 1562 418 1582
rect 269 1554 418 1562
rect 485 1586 844 1590
rect 485 1581 807 1586
rect 485 1557 598 1581
rect 622 1562 807 1581
rect 831 1562 844 1586
rect 622 1557 844 1562
rect 485 1554 844 1557
rect 906 1554 941 1591
rect 1009 1588 1109 1591
rect 1009 1584 1076 1588
rect 1009 1558 1021 1584
rect 1047 1562 1076 1584
rect 1102 1562 1109 1588
rect 1047 1558 1109 1562
rect 1009 1554 1109 1558
rect 485 1533 516 1554
rect 906 1533 942 1554
rect 328 1532 365 1533
rect 327 1523 365 1532
rect 327 1503 336 1523
rect 356 1503 365 1523
rect 327 1495 365 1503
rect 431 1527 516 1533
rect 541 1532 578 1533
rect 431 1507 439 1527
rect 459 1507 516 1527
rect 431 1499 516 1507
rect 540 1523 578 1532
rect 540 1503 549 1523
rect 569 1503 578 1523
rect 431 1498 467 1499
rect 540 1495 578 1503
rect 644 1527 729 1533
rect 749 1532 786 1533
rect 644 1507 652 1527
rect 672 1526 729 1527
rect 672 1507 701 1526
rect 644 1506 701 1507
rect 722 1506 729 1526
rect 644 1499 729 1506
rect 748 1523 786 1532
rect 748 1503 757 1523
rect 777 1503 786 1523
rect 644 1498 680 1499
rect 748 1495 786 1503
rect 852 1528 996 1533
rect 852 1527 917 1528
rect 852 1507 860 1527
rect 880 1507 917 1527
rect 939 1527 996 1528
rect 939 1507 968 1527
rect 988 1507 996 1527
rect 852 1499 996 1507
rect 852 1498 888 1499
rect 960 1498 996 1499
rect 1062 1532 1099 1533
rect 1062 1531 1100 1532
rect 1062 1523 1126 1531
rect 1062 1503 1071 1523
rect 1091 1509 1126 1523
rect 1146 1509 1149 1529
rect 1091 1504 1149 1509
rect 1091 1503 1126 1504
rect 328 1466 365 1495
rect 329 1464 365 1466
rect 541 1464 578 1495
rect 329 1442 578 1464
rect 749 1463 786 1495
rect 1062 1491 1126 1503
rect 1166 1465 1193 1643
rect 1025 1463 1193 1465
rect 749 1437 1193 1463
rect 1345 1562 1595 1586
rect 1345 1491 1382 1562
rect 1497 1501 1528 1502
rect 1345 1471 1354 1491
rect 1374 1471 1382 1491
rect 1345 1461 1382 1471
rect 1441 1491 1528 1501
rect 1441 1471 1450 1491
rect 1470 1471 1528 1491
rect 1441 1462 1528 1471
rect 1441 1461 1478 1462
rect 749 1427 771 1437
rect 1025 1436 1193 1437
rect 709 1425 771 1427
rect 139 1418 771 1425
rect 138 1409 771 1418
rect 1497 1409 1528 1462
rect 1558 1491 1595 1562
rect 1766 1567 2159 1587
rect 2179 1567 2182 1587
rect 1766 1562 2182 1567
rect 1766 1561 2107 1562
rect 1710 1501 1741 1502
rect 1558 1471 1567 1491
rect 1587 1471 1595 1491
rect 1558 1461 1595 1471
rect 1654 1494 1741 1501
rect 1654 1491 1715 1494
rect 1654 1471 1663 1491
rect 1683 1474 1715 1491
rect 1736 1474 1741 1494
rect 1683 1471 1741 1474
rect 1654 1464 1741 1471
rect 1766 1491 1803 1561
rect 2069 1560 2106 1561
rect 1918 1501 1954 1502
rect 1766 1471 1775 1491
rect 1795 1471 1803 1491
rect 1654 1462 1710 1464
rect 1654 1461 1691 1462
rect 1766 1461 1803 1471
rect 1862 1491 2010 1501
rect 2110 1498 2206 1500
rect 1862 1471 1871 1491
rect 1891 1471 1981 1491
rect 2001 1471 2010 1491
rect 1862 1462 2010 1471
rect 2068 1491 2206 1498
rect 2068 1471 2077 1491
rect 2097 1471 2206 1491
rect 2068 1462 2206 1471
rect 1862 1461 1899 1462
rect 1918 1410 1954 1462
rect 1973 1461 2010 1462
rect 2069 1461 2106 1462
rect 138 1391 148 1409
rect 166 1408 771 1409
rect 1389 1408 1430 1409
rect 166 1403 187 1408
rect 166 1391 178 1403
rect 1281 1401 1430 1408
rect 138 1383 178 1391
rect 221 1390 247 1391
rect 138 1381 175 1383
rect 221 1372 775 1390
rect 1281 1381 1399 1401
rect 1419 1381 1430 1401
rect 1281 1373 1430 1381
rect 1497 1405 1856 1409
rect 1497 1400 1819 1405
rect 1497 1376 1610 1400
rect 1634 1381 1819 1400
rect 1843 1381 1856 1405
rect 1634 1376 1856 1381
rect 1497 1373 1856 1376
rect 1918 1373 1953 1410
rect 2021 1407 2121 1410
rect 2021 1403 2088 1407
rect 2021 1377 2033 1403
rect 2059 1381 2088 1403
rect 2114 1381 2121 1407
rect 2059 1377 2121 1381
rect 2021 1373 2121 1377
rect 141 1313 178 1319
rect 221 1313 247 1372
rect 754 1353 775 1372
rect 141 1310 247 1313
rect 141 1292 150 1310
rect 168 1296 247 1310
rect 332 1328 582 1352
rect 168 1294 244 1296
rect 168 1292 178 1294
rect 141 1282 178 1292
rect 146 1217 177 1282
rect 332 1257 369 1328
rect 484 1267 515 1268
rect 332 1237 341 1257
rect 361 1237 369 1257
rect 332 1227 369 1237
rect 428 1257 515 1267
rect 428 1237 437 1257
rect 457 1237 515 1257
rect 428 1228 515 1237
rect 428 1227 465 1228
rect 145 1208 182 1217
rect 145 1190 155 1208
rect 173 1190 182 1208
rect 145 1180 182 1190
rect 484 1175 515 1228
rect 545 1257 582 1328
rect 753 1333 1146 1353
rect 1166 1333 1169 1353
rect 1497 1352 1528 1373
rect 1918 1352 1954 1373
rect 1340 1351 1377 1352
rect 753 1328 1169 1333
rect 1339 1342 1377 1351
rect 753 1327 1094 1328
rect 697 1267 728 1268
rect 545 1237 554 1257
rect 574 1237 582 1257
rect 545 1227 582 1237
rect 641 1260 728 1267
rect 641 1257 702 1260
rect 641 1237 650 1257
rect 670 1240 702 1257
rect 723 1240 728 1260
rect 670 1237 728 1240
rect 641 1230 728 1237
rect 753 1257 790 1327
rect 1056 1326 1093 1327
rect 1339 1322 1348 1342
rect 1368 1322 1377 1342
rect 1339 1314 1377 1322
rect 1443 1346 1528 1352
rect 1553 1351 1590 1352
rect 1443 1326 1451 1346
rect 1471 1326 1528 1346
rect 1443 1318 1528 1326
rect 1552 1342 1590 1351
rect 1552 1322 1561 1342
rect 1581 1322 1590 1342
rect 1443 1317 1479 1318
rect 1552 1314 1590 1322
rect 1656 1346 1741 1352
rect 1761 1351 1798 1352
rect 1656 1326 1664 1346
rect 1684 1345 1741 1346
rect 1684 1326 1713 1345
rect 1656 1325 1713 1326
rect 1734 1325 1741 1345
rect 1656 1318 1741 1325
rect 1760 1342 1798 1351
rect 1760 1322 1769 1342
rect 1789 1322 1798 1342
rect 1656 1317 1692 1318
rect 1760 1314 1798 1322
rect 1864 1346 2008 1352
rect 1864 1326 1872 1346
rect 1892 1326 1924 1346
rect 1948 1326 1980 1346
rect 2000 1326 2008 1346
rect 1864 1318 2008 1326
rect 1864 1317 1900 1318
rect 1972 1317 2008 1318
rect 2074 1351 2111 1352
rect 2074 1350 2112 1351
rect 2074 1342 2138 1350
rect 2074 1322 2083 1342
rect 2103 1328 2138 1342
rect 2158 1328 2161 1348
rect 2103 1323 2161 1328
rect 2103 1322 2138 1323
rect 1340 1285 1377 1314
rect 1341 1283 1377 1285
rect 1553 1283 1590 1314
rect 905 1267 941 1268
rect 753 1237 762 1257
rect 782 1237 790 1257
rect 641 1228 697 1230
rect 641 1227 678 1228
rect 753 1227 790 1237
rect 849 1257 997 1267
rect 1097 1264 1193 1266
rect 849 1237 858 1257
rect 878 1237 968 1257
rect 988 1237 997 1257
rect 849 1228 997 1237
rect 1055 1257 1193 1264
rect 1341 1261 1590 1283
rect 1761 1282 1798 1314
rect 2074 1310 2138 1322
rect 2178 1284 2205 1462
rect 2037 1282 2205 1284
rect 1761 1278 2205 1282
rect 1055 1237 1064 1257
rect 1084 1237 1193 1257
rect 1761 1259 1810 1278
rect 1830 1259 2205 1278
rect 1761 1256 2205 1259
rect 2037 1255 2205 1256
rect 1055 1228 1193 1237
rect 849 1227 886 1228
rect 905 1176 941 1228
rect 960 1227 997 1228
rect 1056 1227 1093 1228
rect 376 1174 417 1175
rect 268 1167 417 1174
rect 268 1147 386 1167
rect 406 1147 417 1167
rect 268 1139 417 1147
rect 484 1171 843 1175
rect 484 1166 806 1171
rect 484 1142 597 1166
rect 621 1147 806 1166
rect 830 1147 843 1171
rect 621 1142 843 1147
rect 484 1139 843 1142
rect 905 1139 940 1176
rect 1008 1173 1108 1176
rect 1008 1169 1075 1173
rect 1008 1143 1020 1169
rect 1046 1147 1075 1169
rect 1101 1147 1108 1173
rect 1046 1143 1108 1147
rect 1008 1139 1108 1143
rect 484 1118 515 1139
rect 905 1118 941 1139
rect 148 1109 185 1118
rect 327 1117 364 1118
rect 148 1091 157 1109
rect 175 1091 185 1109
rect 148 1081 185 1091
rect 149 1046 185 1081
rect 326 1108 364 1117
rect 326 1088 335 1108
rect 355 1088 364 1108
rect 326 1080 364 1088
rect 430 1112 515 1118
rect 540 1117 577 1118
rect 430 1092 438 1112
rect 458 1092 515 1112
rect 430 1084 515 1092
rect 539 1108 577 1117
rect 539 1088 548 1108
rect 568 1088 577 1108
rect 430 1083 466 1084
rect 539 1080 577 1088
rect 643 1112 728 1118
rect 748 1117 785 1118
rect 643 1092 651 1112
rect 671 1111 728 1112
rect 671 1092 700 1111
rect 643 1091 700 1092
rect 721 1091 728 1111
rect 643 1084 728 1091
rect 747 1108 785 1117
rect 747 1088 756 1108
rect 776 1088 785 1108
rect 643 1083 679 1084
rect 747 1080 785 1088
rect 851 1112 995 1118
rect 851 1092 859 1112
rect 879 1111 967 1112
rect 879 1092 907 1111
rect 851 1090 907 1092
rect 929 1092 967 1111
rect 987 1092 995 1112
rect 929 1090 995 1092
rect 851 1084 995 1090
rect 851 1083 887 1084
rect 959 1083 995 1084
rect 1061 1117 1098 1118
rect 1061 1116 1099 1117
rect 1061 1108 1125 1116
rect 1061 1088 1070 1108
rect 1090 1094 1125 1108
rect 1145 1094 1148 1114
rect 1090 1089 1148 1094
rect 1090 1088 1125 1089
rect 327 1051 364 1080
rect 147 1005 185 1046
rect 328 1049 364 1051
rect 540 1049 577 1080
rect 328 1027 577 1049
rect 748 1048 785 1080
rect 1061 1076 1125 1088
rect 1165 1050 1192 1228
rect 1024 1048 1192 1050
rect 748 1022 1192 1048
rect 749 1005 773 1022
rect 1024 1021 1192 1022
rect 147 987 774 1005
rect 1400 1001 1650 1025
rect 147 981 185 987
rect 147 957 184 981
rect 147 933 182 957
rect 145 924 182 933
rect 145 906 155 924
rect 173 906 182 924
rect 145 896 182 906
rect 1400 930 1437 1001
rect 1552 940 1583 941
rect 1400 910 1409 930
rect 1429 910 1437 930
rect 1400 900 1437 910
rect 1496 930 1583 940
rect 1496 910 1505 930
rect 1525 910 1583 930
rect 1496 901 1583 910
rect 1496 900 1533 901
rect 1552 848 1583 901
rect 1613 930 1650 1001
rect 1821 1006 2214 1026
rect 2234 1006 2237 1026
rect 1821 1001 2237 1006
rect 1821 1000 2162 1001
rect 1765 940 1796 941
rect 1613 910 1622 930
rect 1642 910 1650 930
rect 1613 900 1650 910
rect 1709 933 1796 940
rect 1709 930 1770 933
rect 1709 910 1718 930
rect 1738 913 1770 930
rect 1791 913 1796 933
rect 1738 910 1796 913
rect 1709 903 1796 910
rect 1821 930 1858 1000
rect 2124 999 2161 1000
rect 1973 940 2009 941
rect 1821 910 1830 930
rect 1850 910 1858 930
rect 1709 901 1765 903
rect 1709 900 1746 901
rect 1821 900 1858 910
rect 1917 930 2065 940
rect 2165 937 2261 939
rect 1917 910 1926 930
rect 1946 910 2036 930
rect 2056 910 2065 930
rect 1917 901 2065 910
rect 2123 930 2261 937
rect 2123 910 2132 930
rect 2152 910 2261 930
rect 2123 901 2261 910
rect 1917 900 1954 901
rect 1973 849 2009 901
rect 2028 900 2065 901
rect 2124 900 2161 901
rect 1444 847 1485 848
rect 1336 840 1485 847
rect 148 832 185 834
rect 148 831 796 832
rect 147 825 796 831
rect 147 807 157 825
rect 175 811 796 825
rect 1336 820 1454 840
rect 1474 820 1485 840
rect 1336 812 1485 820
rect 1552 844 1911 848
rect 1552 839 1874 844
rect 1552 815 1665 839
rect 1689 820 1874 839
rect 1898 820 1911 844
rect 1689 815 1911 820
rect 1552 812 1911 815
rect 1973 812 2008 849
rect 2076 846 2176 849
rect 2076 842 2143 846
rect 2076 816 2088 842
rect 2114 820 2143 842
rect 2169 820 2176 846
rect 2114 816 2176 820
rect 2076 812 2176 816
rect 175 807 185 811
rect 626 810 796 811
rect 147 797 185 807
rect 147 719 182 797
rect 759 787 796 810
rect 1552 791 1583 812
rect 1973 791 2009 812
rect 1395 790 1432 791
rect 143 710 182 719
rect 143 692 153 710
rect 171 692 182 710
rect 143 686 182 692
rect 338 762 588 786
rect 338 691 375 762
rect 490 701 521 702
rect 143 682 180 686
rect 338 671 347 691
rect 367 671 375 691
rect 338 661 375 671
rect 434 691 521 701
rect 434 671 443 691
rect 463 671 521 691
rect 434 662 521 671
rect 434 661 471 662
rect 146 611 183 620
rect 144 593 155 611
rect 173 593 183 611
rect 490 609 521 662
rect 551 691 588 762
rect 759 767 1152 787
rect 1172 767 1175 787
rect 759 762 1175 767
rect 1394 781 1432 790
rect 759 761 1100 762
rect 1394 761 1403 781
rect 1423 761 1432 781
rect 703 701 734 702
rect 551 671 560 691
rect 580 671 588 691
rect 551 661 588 671
rect 647 694 734 701
rect 647 691 708 694
rect 647 671 656 691
rect 676 674 708 691
rect 729 674 734 694
rect 676 671 734 674
rect 647 664 734 671
rect 759 691 796 761
rect 1062 760 1099 761
rect 1394 753 1432 761
rect 1498 785 1583 791
rect 1608 790 1645 791
rect 1498 765 1506 785
rect 1526 765 1583 785
rect 1498 757 1583 765
rect 1607 781 1645 790
rect 1607 761 1616 781
rect 1636 761 1645 781
rect 1498 756 1534 757
rect 1607 753 1645 761
rect 1711 785 1796 791
rect 1816 790 1853 791
rect 1711 765 1719 785
rect 1739 784 1796 785
rect 1739 765 1768 784
rect 1711 764 1768 765
rect 1789 764 1796 784
rect 1711 757 1796 764
rect 1815 781 1853 790
rect 1815 761 1824 781
rect 1844 761 1853 781
rect 1711 756 1747 757
rect 1815 753 1853 761
rect 1919 785 2063 791
rect 1919 765 1927 785
rect 1947 784 2035 785
rect 1947 765 1980 784
rect 2003 765 2035 784
rect 2055 765 2063 785
rect 1919 757 2063 765
rect 1919 756 1955 757
rect 2027 756 2063 757
rect 2129 790 2166 791
rect 2129 789 2167 790
rect 2129 781 2193 789
rect 2129 761 2138 781
rect 2158 767 2193 781
rect 2213 767 2216 787
rect 2158 762 2216 767
rect 2158 761 2193 762
rect 1395 724 1432 753
rect 1396 722 1432 724
rect 1608 722 1645 753
rect 911 701 947 702
rect 759 671 768 691
rect 788 671 796 691
rect 647 662 703 664
rect 647 661 684 662
rect 759 661 796 671
rect 855 691 1003 701
rect 1396 700 1645 722
rect 1816 721 1853 753
rect 2129 749 2193 761
rect 2233 723 2260 901
rect 2092 721 2260 723
rect 1816 710 2260 721
rect 2323 721 2353 1722
rect 2442 1715 2479 1726
rect 4063 1715 4090 1893
rect 4130 1855 4194 1867
rect 4470 1863 4507 1895
rect 4678 1894 4927 1916
rect 4678 1863 4715 1894
rect 4891 1892 4927 1894
rect 5070 1897 5108 1938
rect 4891 1863 4928 1892
rect 4130 1854 4165 1855
rect 4107 1849 4165 1854
rect 4107 1829 4110 1849
rect 4130 1835 4165 1849
rect 4185 1835 4194 1855
rect 4130 1827 4194 1835
rect 4156 1826 4194 1827
rect 4157 1825 4194 1826
rect 4260 1859 4296 1860
rect 4368 1859 4404 1860
rect 4260 1853 4404 1859
rect 4260 1851 4326 1853
rect 4260 1831 4268 1851
rect 4288 1832 4326 1851
rect 4348 1851 4404 1853
rect 4348 1832 4376 1851
rect 4288 1831 4376 1832
rect 4396 1831 4404 1851
rect 4260 1825 4404 1831
rect 4470 1855 4508 1863
rect 4576 1859 4612 1860
rect 4470 1835 4479 1855
rect 4499 1835 4508 1855
rect 4470 1826 4508 1835
rect 4527 1852 4612 1859
rect 4527 1832 4534 1852
rect 4555 1851 4612 1852
rect 4555 1832 4584 1851
rect 4527 1831 4584 1832
rect 4604 1831 4612 1851
rect 4470 1825 4507 1826
rect 4527 1825 4612 1831
rect 4678 1855 4716 1863
rect 4789 1859 4825 1860
rect 4678 1835 4687 1855
rect 4707 1835 4716 1855
rect 4678 1826 4716 1835
rect 4740 1851 4825 1859
rect 4740 1831 4797 1851
rect 4817 1831 4825 1851
rect 4678 1825 4715 1826
rect 4740 1825 4825 1831
rect 4891 1855 4929 1863
rect 4891 1835 4900 1855
rect 4920 1835 4929 1855
rect 4891 1826 4929 1835
rect 5070 1862 5106 1897
rect 5070 1852 5107 1862
rect 5070 1834 5080 1852
rect 5098 1834 5107 1852
rect 4891 1825 4928 1826
rect 5070 1825 5107 1834
rect 4314 1804 4350 1825
rect 4740 1804 4771 1825
rect 4147 1800 4247 1804
rect 4147 1796 4209 1800
rect 4147 1770 4154 1796
rect 4180 1774 4209 1796
rect 4235 1774 4247 1800
rect 4180 1770 4247 1774
rect 4147 1767 4247 1770
rect 4315 1767 4350 1804
rect 4412 1801 4771 1804
rect 4412 1796 4634 1801
rect 4412 1772 4425 1796
rect 4449 1777 4634 1796
rect 4658 1777 4771 1801
rect 4449 1772 4771 1777
rect 4412 1768 4771 1772
rect 4838 1796 4987 1804
rect 4838 1776 4849 1796
rect 4869 1776 4987 1796
rect 4838 1769 4987 1776
rect 4838 1768 4879 1769
rect 4162 1715 4199 1716
rect 4258 1715 4295 1716
rect 4314 1715 4350 1767
rect 4369 1715 4406 1716
rect 4062 1706 4200 1715
rect 2998 1688 3029 1691
rect 2998 1662 3005 1688
rect 3024 1662 3029 1688
rect 2998 1268 3029 1662
rect 3050 1687 3218 1688
rect 3050 1684 3494 1687
rect 3050 1665 3425 1684
rect 3445 1665 3494 1684
rect 4062 1686 4171 1706
rect 4191 1686 4200 1706
rect 3050 1661 3494 1665
rect 3050 1659 3218 1661
rect 3050 1481 3077 1659
rect 3117 1621 3181 1633
rect 3457 1629 3494 1661
rect 3665 1660 3914 1682
rect 4062 1679 4200 1686
rect 4258 1706 4406 1715
rect 4258 1686 4267 1706
rect 4287 1686 4377 1706
rect 4397 1686 4406 1706
rect 4062 1677 4158 1679
rect 4258 1676 4406 1686
rect 4465 1706 4502 1716
rect 4577 1715 4614 1716
rect 4558 1713 4614 1715
rect 4465 1686 4473 1706
rect 4493 1686 4502 1706
rect 4314 1675 4350 1676
rect 3665 1629 3702 1660
rect 3878 1658 3914 1660
rect 3878 1629 3915 1658
rect 3117 1620 3152 1621
rect 3094 1615 3152 1620
rect 3094 1595 3097 1615
rect 3117 1601 3152 1615
rect 3172 1601 3181 1621
rect 3117 1593 3181 1601
rect 3143 1592 3181 1593
rect 3144 1591 3181 1592
rect 3247 1625 3283 1626
rect 3355 1625 3391 1626
rect 3247 1617 3391 1625
rect 3247 1597 3255 1617
rect 3275 1616 3363 1617
rect 3275 1597 3308 1616
rect 3247 1596 3308 1597
rect 3332 1597 3363 1616
rect 3383 1597 3391 1617
rect 3332 1596 3391 1597
rect 3247 1591 3391 1596
rect 3457 1621 3495 1629
rect 3563 1625 3599 1626
rect 3457 1601 3466 1621
rect 3486 1601 3495 1621
rect 3457 1592 3495 1601
rect 3514 1618 3599 1625
rect 3514 1598 3521 1618
rect 3542 1617 3599 1618
rect 3542 1598 3571 1617
rect 3514 1597 3571 1598
rect 3591 1597 3599 1617
rect 3457 1591 3494 1592
rect 3514 1591 3599 1597
rect 3665 1621 3703 1629
rect 3776 1625 3812 1626
rect 3665 1601 3674 1621
rect 3694 1601 3703 1621
rect 3665 1592 3703 1601
rect 3727 1617 3812 1625
rect 3727 1597 3784 1617
rect 3804 1597 3812 1617
rect 3665 1591 3702 1592
rect 3727 1591 3812 1597
rect 3878 1621 3916 1629
rect 3878 1601 3887 1621
rect 3907 1601 3916 1621
rect 4162 1616 4199 1617
rect 4465 1616 4502 1686
rect 4527 1706 4614 1713
rect 4527 1703 4585 1706
rect 4527 1683 4532 1703
rect 4553 1686 4585 1703
rect 4605 1686 4614 1706
rect 4553 1683 4614 1686
rect 4527 1676 4614 1683
rect 4673 1706 4710 1716
rect 4673 1686 4681 1706
rect 4701 1686 4710 1706
rect 4527 1675 4558 1676
rect 4161 1615 4502 1616
rect 3878 1592 3916 1601
rect 4086 1610 4502 1615
rect 3878 1591 3915 1592
rect 3301 1570 3337 1591
rect 3727 1570 3758 1591
rect 4086 1590 4089 1610
rect 4109 1590 4502 1610
rect 4673 1615 4710 1686
rect 4740 1715 4771 1768
rect 5073 1753 5110 1763
rect 5073 1735 5082 1753
rect 5100 1735 5110 1753
rect 5073 1726 5110 1735
rect 4790 1715 4827 1716
rect 4740 1706 4827 1715
rect 4740 1686 4798 1706
rect 4818 1686 4827 1706
rect 4740 1676 4827 1686
rect 4886 1706 4923 1716
rect 4886 1686 4894 1706
rect 4914 1686 4923 1706
rect 4740 1675 4771 1676
rect 4886 1615 4923 1686
rect 5078 1661 5109 1726
rect 5077 1651 5114 1661
rect 5077 1649 5087 1651
rect 5011 1647 5087 1649
rect 4673 1591 4923 1615
rect 5008 1633 5087 1647
rect 5105 1633 5114 1651
rect 5008 1630 5114 1633
rect 4480 1571 4501 1590
rect 5008 1571 5034 1630
rect 5077 1624 5114 1630
rect 3134 1566 3234 1570
rect 3134 1562 3196 1566
rect 3134 1536 3141 1562
rect 3167 1540 3196 1562
rect 3222 1540 3234 1566
rect 3167 1536 3234 1540
rect 3134 1533 3234 1536
rect 3302 1533 3337 1570
rect 3399 1567 3758 1570
rect 3399 1562 3621 1567
rect 3399 1538 3412 1562
rect 3436 1543 3621 1562
rect 3645 1543 3758 1567
rect 3436 1538 3758 1543
rect 3399 1534 3758 1538
rect 3825 1562 3974 1570
rect 3825 1542 3836 1562
rect 3856 1542 3974 1562
rect 4480 1553 5034 1571
rect 5080 1560 5117 1562
rect 5008 1552 5034 1553
rect 5077 1552 5117 1560
rect 3825 1535 3974 1542
rect 5077 1540 5089 1552
rect 5068 1535 5089 1540
rect 3825 1534 3866 1535
rect 4484 1534 5089 1535
rect 5107 1534 5117 1552
rect 3149 1481 3186 1482
rect 3245 1481 3282 1482
rect 3301 1481 3337 1533
rect 3356 1481 3393 1482
rect 3049 1472 3187 1481
rect 3049 1452 3158 1472
rect 3178 1452 3187 1472
rect 3049 1445 3187 1452
rect 3245 1472 3393 1481
rect 3245 1452 3254 1472
rect 3274 1452 3364 1472
rect 3384 1452 3393 1472
rect 3049 1443 3145 1445
rect 3245 1442 3393 1452
rect 3452 1472 3489 1482
rect 3564 1481 3601 1482
rect 3545 1479 3601 1481
rect 3452 1452 3460 1472
rect 3480 1452 3489 1472
rect 3301 1441 3337 1442
rect 3149 1382 3186 1383
rect 3452 1382 3489 1452
rect 3514 1472 3601 1479
rect 3514 1469 3572 1472
rect 3514 1449 3519 1469
rect 3540 1452 3572 1469
rect 3592 1452 3601 1472
rect 3540 1449 3601 1452
rect 3514 1442 3601 1449
rect 3660 1472 3697 1482
rect 3660 1452 3668 1472
rect 3688 1452 3697 1472
rect 3514 1441 3545 1442
rect 3148 1381 3489 1382
rect 3073 1376 3489 1381
rect 3073 1356 3076 1376
rect 3096 1356 3489 1376
rect 3660 1381 3697 1452
rect 3727 1481 3758 1534
rect 4484 1525 5117 1534
rect 4484 1518 5116 1525
rect 4484 1516 4546 1518
rect 4062 1506 4230 1507
rect 4484 1506 4506 1516
rect 3777 1481 3814 1482
rect 3727 1472 3814 1481
rect 3727 1452 3785 1472
rect 3805 1452 3814 1472
rect 3727 1442 3814 1452
rect 3873 1472 3910 1482
rect 3873 1452 3881 1472
rect 3901 1452 3910 1472
rect 3727 1441 3758 1442
rect 3873 1381 3910 1452
rect 3660 1357 3910 1381
rect 4062 1480 4506 1506
rect 4062 1478 4230 1480
rect 4062 1300 4089 1478
rect 4129 1440 4193 1452
rect 4469 1448 4506 1480
rect 4677 1479 4926 1501
rect 4677 1448 4714 1479
rect 4890 1477 4926 1479
rect 4890 1448 4927 1477
rect 4129 1439 4164 1440
rect 4106 1434 4164 1439
rect 4106 1414 4109 1434
rect 4129 1420 4164 1434
rect 4184 1420 4193 1440
rect 4129 1412 4193 1420
rect 4155 1411 4193 1412
rect 4156 1410 4193 1411
rect 4259 1444 4295 1445
rect 4367 1444 4403 1445
rect 4259 1436 4403 1444
rect 4259 1416 4267 1436
rect 4287 1416 4316 1436
rect 4259 1415 4316 1416
rect 4338 1416 4375 1436
rect 4395 1416 4403 1436
rect 4338 1415 4403 1416
rect 4259 1410 4403 1415
rect 4469 1440 4507 1448
rect 4575 1444 4611 1445
rect 4469 1420 4478 1440
rect 4498 1420 4507 1440
rect 4469 1411 4507 1420
rect 4526 1437 4611 1444
rect 4526 1417 4533 1437
rect 4554 1436 4611 1437
rect 4554 1417 4583 1436
rect 4526 1416 4583 1417
rect 4603 1416 4611 1436
rect 4469 1410 4506 1411
rect 4526 1410 4611 1416
rect 4677 1440 4715 1448
rect 4788 1444 4824 1445
rect 4677 1420 4686 1440
rect 4706 1420 4715 1440
rect 4677 1411 4715 1420
rect 4739 1436 4824 1444
rect 4739 1416 4796 1436
rect 4816 1416 4824 1436
rect 4677 1410 4714 1411
rect 4739 1410 4824 1416
rect 4890 1440 4928 1448
rect 4890 1420 4899 1440
rect 4919 1420 4928 1440
rect 4890 1411 4928 1420
rect 4890 1410 4927 1411
rect 4313 1389 4349 1410
rect 4739 1389 4770 1410
rect 4146 1385 4246 1389
rect 4146 1381 4208 1385
rect 4146 1355 4153 1381
rect 4179 1359 4208 1381
rect 4234 1359 4246 1385
rect 4179 1355 4246 1359
rect 4146 1352 4246 1355
rect 4314 1352 4349 1389
rect 4411 1386 4770 1389
rect 4411 1381 4633 1386
rect 4411 1357 4424 1381
rect 4448 1362 4633 1381
rect 4657 1362 4770 1386
rect 4448 1357 4770 1362
rect 4411 1353 4770 1357
rect 4837 1381 4986 1389
rect 4837 1361 4848 1381
rect 4868 1361 4986 1381
rect 4837 1354 4986 1361
rect 5077 1369 5116 1518
rect 4837 1353 4878 1354
rect 4161 1300 4198 1301
rect 4257 1300 4294 1301
rect 4313 1300 4349 1352
rect 4368 1300 4405 1301
rect 4061 1291 4199 1300
rect 4061 1271 4170 1291
rect 4190 1271 4199 1291
rect 2998 1267 3168 1268
rect 2998 1252 3444 1267
rect 4061 1264 4199 1271
rect 4257 1291 4405 1300
rect 4257 1271 4266 1291
rect 4286 1271 4376 1291
rect 4396 1271 4405 1291
rect 4061 1262 4157 1264
rect 3000 1241 3444 1252
rect 3000 1239 3168 1241
rect 3000 1061 3027 1239
rect 3067 1201 3131 1213
rect 3407 1209 3444 1241
rect 3615 1240 3864 1262
rect 4257 1261 4405 1271
rect 4464 1291 4501 1301
rect 4576 1300 4613 1301
rect 4557 1298 4613 1300
rect 4464 1271 4472 1291
rect 4492 1271 4501 1291
rect 4313 1260 4349 1261
rect 3615 1209 3652 1240
rect 3828 1238 3864 1240
rect 3828 1209 3865 1238
rect 3067 1200 3102 1201
rect 3044 1195 3102 1200
rect 3044 1175 3047 1195
rect 3067 1181 3102 1195
rect 3122 1181 3131 1201
rect 3067 1173 3131 1181
rect 3093 1172 3131 1173
rect 3094 1171 3131 1172
rect 3197 1205 3233 1206
rect 3305 1205 3341 1206
rect 3197 1197 3341 1205
rect 3197 1177 3205 1197
rect 3225 1196 3313 1197
rect 3225 1179 3253 1196
rect 3277 1179 3313 1196
rect 3225 1177 3313 1179
rect 3333 1177 3341 1197
rect 3197 1171 3341 1177
rect 3407 1201 3445 1209
rect 3513 1205 3549 1206
rect 3407 1181 3416 1201
rect 3436 1181 3445 1201
rect 3407 1172 3445 1181
rect 3464 1198 3549 1205
rect 3464 1178 3471 1198
rect 3492 1197 3549 1198
rect 3492 1178 3521 1197
rect 3464 1177 3521 1178
rect 3541 1177 3549 1197
rect 3407 1171 3444 1172
rect 3464 1171 3549 1177
rect 3615 1201 3653 1209
rect 3726 1205 3762 1206
rect 3615 1181 3624 1201
rect 3644 1181 3653 1201
rect 3615 1172 3653 1181
rect 3677 1197 3762 1205
rect 3677 1177 3734 1197
rect 3754 1177 3762 1197
rect 3615 1171 3652 1172
rect 3677 1171 3762 1177
rect 3828 1201 3866 1209
rect 4161 1201 4198 1202
rect 4464 1201 4501 1271
rect 4526 1291 4613 1298
rect 4526 1288 4584 1291
rect 4526 1268 4531 1288
rect 4552 1271 4584 1288
rect 4604 1271 4613 1291
rect 4552 1268 4613 1271
rect 4526 1261 4613 1268
rect 4672 1291 4709 1301
rect 4672 1271 4680 1291
rect 4700 1271 4709 1291
rect 4526 1260 4557 1261
rect 3828 1181 3837 1201
rect 3857 1181 3866 1201
rect 4160 1200 4501 1201
rect 3828 1172 3866 1181
rect 4085 1195 4501 1200
rect 4085 1175 4088 1195
rect 4108 1175 4501 1195
rect 4672 1200 4709 1271
rect 4739 1300 4770 1353
rect 5077 1351 5087 1369
rect 5105 1351 5116 1369
rect 5077 1342 5114 1351
rect 4789 1300 4826 1301
rect 4739 1291 4826 1300
rect 4739 1271 4797 1291
rect 4817 1271 4826 1291
rect 4739 1261 4826 1271
rect 4885 1291 4922 1301
rect 4885 1271 4893 1291
rect 4913 1271 4922 1291
rect 5080 1276 5117 1280
rect 4739 1260 4770 1261
rect 4885 1200 4922 1271
rect 4672 1176 4922 1200
rect 5078 1270 5117 1276
rect 5078 1252 5089 1270
rect 5107 1252 5117 1270
rect 5078 1243 5117 1252
rect 3828 1171 3865 1172
rect 3251 1150 3287 1171
rect 3677 1150 3708 1171
rect 4464 1152 4501 1175
rect 5078 1165 5113 1243
rect 5075 1155 5113 1165
rect 4464 1151 4634 1152
rect 5075 1151 5085 1155
rect 3084 1146 3184 1150
rect 3084 1142 3146 1146
rect 3084 1116 3091 1142
rect 3117 1120 3146 1142
rect 3172 1120 3184 1146
rect 3117 1116 3184 1120
rect 3084 1113 3184 1116
rect 3252 1113 3287 1150
rect 3349 1147 3708 1150
rect 3349 1142 3571 1147
rect 3349 1118 3362 1142
rect 3386 1123 3571 1142
rect 3595 1123 3708 1147
rect 3386 1118 3708 1123
rect 3349 1114 3708 1118
rect 3775 1142 3924 1150
rect 3775 1122 3786 1142
rect 3806 1122 3924 1142
rect 4464 1137 5085 1151
rect 5103 1137 5113 1155
rect 4464 1131 5113 1137
rect 4464 1130 5112 1131
rect 5075 1128 5112 1130
rect 3775 1115 3924 1122
rect 3775 1114 3816 1115
rect 3099 1061 3136 1062
rect 3195 1061 3232 1062
rect 3251 1061 3287 1113
rect 3306 1061 3343 1062
rect 2999 1052 3137 1061
rect 2999 1032 3108 1052
rect 3128 1032 3137 1052
rect 2999 1025 3137 1032
rect 3195 1052 3343 1061
rect 3195 1032 3204 1052
rect 3224 1032 3314 1052
rect 3334 1032 3343 1052
rect 2999 1023 3095 1025
rect 3195 1022 3343 1032
rect 3402 1052 3439 1062
rect 3514 1061 3551 1062
rect 3495 1059 3551 1061
rect 3402 1032 3410 1052
rect 3430 1032 3439 1052
rect 3251 1021 3287 1022
rect 3099 962 3136 963
rect 3402 962 3439 1032
rect 3464 1052 3551 1059
rect 3464 1049 3522 1052
rect 3464 1029 3469 1049
rect 3490 1032 3522 1049
rect 3542 1032 3551 1052
rect 3490 1029 3551 1032
rect 3464 1022 3551 1029
rect 3610 1052 3647 1062
rect 3610 1032 3618 1052
rect 3638 1032 3647 1052
rect 3464 1021 3495 1022
rect 3098 961 3439 962
rect 3023 956 3439 961
rect 3023 936 3026 956
rect 3046 936 3439 956
rect 3610 961 3647 1032
rect 3677 1061 3708 1114
rect 3727 1061 3764 1062
rect 3677 1052 3764 1061
rect 3677 1032 3735 1052
rect 3755 1032 3764 1052
rect 3677 1022 3764 1032
rect 3823 1052 3860 1062
rect 3823 1032 3831 1052
rect 3851 1032 3860 1052
rect 3677 1021 3708 1022
rect 3823 961 3860 1032
rect 5078 1056 5115 1066
rect 5078 1038 5087 1056
rect 5105 1038 5115 1056
rect 5078 1029 5115 1038
rect 5078 1005 5113 1029
rect 5076 981 5113 1005
rect 5075 975 5113 981
rect 3610 937 3860 961
rect 4486 957 5113 975
rect 4068 940 4236 941
rect 4487 940 4511 957
rect 4068 914 4512 940
rect 4068 912 4236 914
rect 4068 734 4095 912
rect 4135 874 4199 886
rect 4475 882 4512 914
rect 4683 913 4932 935
rect 4683 882 4720 913
rect 4896 911 4932 913
rect 5075 916 5113 957
rect 4896 882 4933 911
rect 4135 873 4170 874
rect 4112 868 4170 873
rect 4112 848 4115 868
rect 4135 854 4170 868
rect 4190 854 4199 874
rect 4135 846 4199 854
rect 4161 845 4199 846
rect 4162 844 4199 845
rect 4265 878 4301 879
rect 4373 878 4409 879
rect 4265 872 4409 878
rect 4265 870 4331 872
rect 4265 850 4273 870
rect 4293 851 4331 870
rect 4353 870 4409 872
rect 4353 851 4381 870
rect 4293 850 4381 851
rect 4401 850 4409 870
rect 4265 844 4409 850
rect 4475 874 4513 882
rect 4581 878 4617 879
rect 4475 854 4484 874
rect 4504 854 4513 874
rect 4475 845 4513 854
rect 4532 871 4617 878
rect 4532 851 4539 871
rect 4560 870 4617 871
rect 4560 851 4589 870
rect 4532 850 4589 851
rect 4609 850 4617 870
rect 4475 844 4512 845
rect 4532 844 4617 850
rect 4683 874 4721 882
rect 4794 878 4830 879
rect 4683 854 4692 874
rect 4712 854 4721 874
rect 4683 845 4721 854
rect 4745 870 4830 878
rect 4745 850 4802 870
rect 4822 850 4830 870
rect 4683 844 4720 845
rect 4745 844 4830 850
rect 4896 874 4934 882
rect 4896 854 4905 874
rect 4925 854 4934 874
rect 4896 845 4934 854
rect 5075 881 5111 916
rect 5075 871 5112 881
rect 5075 853 5085 871
rect 5103 853 5112 871
rect 4896 844 4933 845
rect 5075 844 5112 853
rect 4319 823 4355 844
rect 4745 823 4776 844
rect 4152 819 4252 823
rect 4152 815 4214 819
rect 4152 789 4159 815
rect 4185 793 4214 815
rect 4240 793 4252 819
rect 4185 789 4252 793
rect 4152 786 4252 789
rect 4320 786 4355 823
rect 4417 820 4776 823
rect 4417 815 4639 820
rect 4417 791 4430 815
rect 4454 796 4639 815
rect 4663 796 4776 820
rect 4454 791 4776 796
rect 4417 787 4776 791
rect 4843 815 4992 823
rect 4843 795 4854 815
rect 4874 795 4992 815
rect 4843 788 4992 795
rect 4843 787 4884 788
rect 4167 734 4204 735
rect 4263 734 4300 735
rect 4319 734 4355 786
rect 4374 734 4411 735
rect 4067 725 4205 734
rect 2323 716 2355 721
rect 1103 698 1199 700
rect 855 671 864 691
rect 884 671 974 691
rect 994 671 1003 691
rect 855 662 1003 671
rect 1061 691 1199 698
rect 1816 695 2262 710
rect 2092 694 2262 695
rect 1061 671 1070 691
rect 1090 671 1199 691
rect 1061 662 1199 671
rect 855 661 892 662
rect 911 610 947 662
rect 966 661 1003 662
rect 1062 661 1099 662
rect 382 608 423 609
rect 144 444 183 593
rect 274 601 423 608
rect 274 581 392 601
rect 412 581 423 601
rect 274 573 423 581
rect 490 605 849 609
rect 490 600 812 605
rect 490 576 603 600
rect 627 581 812 600
rect 836 581 849 605
rect 627 576 849 581
rect 490 573 849 576
rect 911 573 946 610
rect 1014 607 1114 610
rect 1014 603 1081 607
rect 1014 577 1026 603
rect 1052 581 1081 603
rect 1107 581 1114 607
rect 1052 577 1114 581
rect 1014 573 1114 577
rect 490 552 521 573
rect 911 552 947 573
rect 333 551 370 552
rect 332 542 370 551
rect 332 522 341 542
rect 361 522 370 542
rect 332 514 370 522
rect 436 546 521 552
rect 546 551 583 552
rect 436 526 444 546
rect 464 526 521 546
rect 436 518 521 526
rect 545 542 583 551
rect 545 522 554 542
rect 574 522 583 542
rect 436 517 472 518
rect 545 514 583 522
rect 649 546 734 552
rect 754 551 791 552
rect 649 526 657 546
rect 677 545 734 546
rect 677 526 706 545
rect 649 525 706 526
rect 727 525 734 545
rect 649 518 734 525
rect 753 542 791 551
rect 753 522 762 542
rect 782 522 791 542
rect 649 517 685 518
rect 753 514 791 522
rect 857 547 1001 552
rect 857 546 922 547
rect 857 526 865 546
rect 885 526 922 546
rect 944 546 1001 547
rect 944 526 973 546
rect 993 526 1001 546
rect 857 518 1001 526
rect 857 517 893 518
rect 965 517 1001 518
rect 1067 551 1104 552
rect 1067 550 1105 551
rect 1067 542 1131 550
rect 1067 522 1076 542
rect 1096 528 1131 542
rect 1151 528 1154 548
rect 1096 523 1154 528
rect 1096 522 1131 523
rect 333 485 370 514
rect 334 483 370 485
rect 546 483 583 514
rect 334 461 583 483
rect 754 482 791 514
rect 1067 510 1131 522
rect 1171 484 1198 662
rect 1030 482 1198 484
rect 754 456 1198 482
rect 1350 581 1600 605
rect 1350 510 1387 581
rect 1502 520 1533 521
rect 1350 490 1359 510
rect 1379 490 1387 510
rect 1350 480 1387 490
rect 1446 510 1533 520
rect 1446 490 1455 510
rect 1475 490 1533 510
rect 1446 481 1533 490
rect 1446 480 1483 481
rect 754 446 776 456
rect 1030 455 1198 456
rect 714 444 776 446
rect 144 437 776 444
rect 143 428 776 437
rect 1502 428 1533 481
rect 1563 510 1600 581
rect 1771 586 2164 606
rect 2184 586 2187 606
rect 1771 581 2187 586
rect 1771 580 2112 581
rect 1715 520 1746 521
rect 1563 490 1572 510
rect 1592 490 1600 510
rect 1563 480 1600 490
rect 1659 513 1746 520
rect 1659 510 1720 513
rect 1659 490 1668 510
rect 1688 493 1720 510
rect 1741 493 1746 513
rect 1688 490 1746 493
rect 1659 483 1746 490
rect 1771 510 1808 580
rect 2074 579 2111 580
rect 1923 520 1959 521
rect 1771 490 1780 510
rect 1800 490 1808 510
rect 1659 481 1715 483
rect 1659 480 1696 481
rect 1771 480 1808 490
rect 1867 510 2015 520
rect 2115 517 2211 519
rect 1867 490 1876 510
rect 1896 490 1986 510
rect 2006 490 2015 510
rect 1867 481 2015 490
rect 2073 510 2211 517
rect 2073 490 2082 510
rect 2102 490 2211 510
rect 2073 481 2211 490
rect 1867 480 1904 481
rect 1923 429 1959 481
rect 1978 480 2015 481
rect 2074 480 2111 481
rect 143 410 153 428
rect 171 427 776 428
rect 1394 427 1435 428
rect 171 422 192 427
rect 171 410 183 422
rect 1286 420 1435 427
rect 143 402 183 410
rect 226 409 252 410
rect 143 400 180 402
rect 226 391 780 409
rect 1286 400 1404 420
rect 1424 400 1435 420
rect 1286 392 1435 400
rect 1502 424 1861 428
rect 1502 419 1824 424
rect 1502 395 1615 419
rect 1639 400 1824 419
rect 1848 400 1861 424
rect 1639 395 1861 400
rect 1502 392 1861 395
rect 1923 392 1958 429
rect 2026 426 2126 429
rect 2026 422 2093 426
rect 2026 396 2038 422
rect 2064 400 2093 422
rect 2119 400 2126 426
rect 2064 396 2126 400
rect 2026 392 2126 396
rect 146 332 183 338
rect 226 332 252 391
rect 759 372 780 391
rect 146 329 252 332
rect 146 311 155 329
rect 173 315 252 329
rect 337 347 587 371
rect 173 313 249 315
rect 173 311 183 313
rect 146 301 183 311
rect 151 236 182 301
rect 337 276 374 347
rect 489 286 520 287
rect 337 256 346 276
rect 366 256 374 276
rect 337 246 374 256
rect 433 276 520 286
rect 433 256 442 276
rect 462 256 520 276
rect 433 247 520 256
rect 433 246 470 247
rect 150 227 187 236
rect 150 209 160 227
rect 178 209 187 227
rect 150 199 187 209
rect 489 194 520 247
rect 550 276 587 347
rect 758 352 1151 372
rect 1171 352 1174 372
rect 1502 371 1533 392
rect 1923 371 1959 392
rect 1345 370 1382 371
rect 758 347 1174 352
rect 1344 361 1382 370
rect 758 346 1099 347
rect 702 286 733 287
rect 550 256 559 276
rect 579 256 587 276
rect 550 246 587 256
rect 646 279 733 286
rect 646 276 707 279
rect 646 256 655 276
rect 675 259 707 276
rect 728 259 733 279
rect 675 256 733 259
rect 646 249 733 256
rect 758 276 795 346
rect 1061 345 1098 346
rect 1344 341 1353 361
rect 1373 341 1382 361
rect 1344 333 1382 341
rect 1448 365 1533 371
rect 1558 370 1595 371
rect 1448 345 1456 365
rect 1476 345 1533 365
rect 1448 337 1533 345
rect 1557 361 1595 370
rect 1557 341 1566 361
rect 1586 341 1595 361
rect 1448 336 1484 337
rect 1557 333 1595 341
rect 1661 365 1746 371
rect 1766 370 1803 371
rect 1661 345 1669 365
rect 1689 364 1746 365
rect 1689 345 1718 364
rect 1661 344 1718 345
rect 1739 344 1746 364
rect 1661 337 1746 344
rect 1765 361 1803 370
rect 1765 341 1774 361
rect 1794 341 1803 361
rect 1661 336 1697 337
rect 1765 333 1803 341
rect 1869 366 2013 371
rect 1869 365 1928 366
rect 1869 345 1877 365
rect 1897 346 1928 365
rect 1952 365 2013 366
rect 1952 346 1985 365
rect 1897 345 1985 346
rect 2005 345 2013 365
rect 1869 337 2013 345
rect 1869 336 1905 337
rect 1977 336 2013 337
rect 2079 370 2116 371
rect 2079 369 2117 370
rect 2079 361 2143 369
rect 2079 341 2088 361
rect 2108 347 2143 361
rect 2163 347 2166 367
rect 2108 342 2166 347
rect 2108 341 2143 342
rect 1345 304 1382 333
rect 1346 302 1382 304
rect 1558 302 1595 333
rect 910 286 946 287
rect 758 256 767 276
rect 787 256 795 276
rect 646 247 702 249
rect 646 246 683 247
rect 758 246 795 256
rect 854 276 1002 286
rect 1102 283 1198 285
rect 854 256 863 276
rect 883 256 973 276
rect 993 256 1002 276
rect 854 247 1002 256
rect 1060 276 1198 283
rect 1346 280 1595 302
rect 1766 301 1803 333
rect 2079 329 2143 341
rect 2183 303 2210 481
rect 2042 301 2210 303
rect 1766 297 2210 301
rect 1060 256 1069 276
rect 1089 256 1198 276
rect 1766 278 1815 297
rect 1835 278 2210 297
rect 1766 275 2210 278
rect 2042 274 2210 275
rect 2231 300 2262 694
rect 2323 698 2328 716
rect 2348 698 2355 716
rect 2323 693 2355 698
rect 2326 691 2355 693
rect 3055 706 3223 707
rect 3055 703 3499 706
rect 3055 684 3430 703
rect 3450 684 3499 703
rect 4067 705 4176 725
rect 4196 705 4205 725
rect 3055 680 3499 684
rect 3055 678 3223 680
rect 3055 500 3082 678
rect 3122 640 3186 652
rect 3462 648 3499 680
rect 3670 679 3919 701
rect 4067 698 4205 705
rect 4263 725 4411 734
rect 4263 705 4272 725
rect 4292 705 4382 725
rect 4402 705 4411 725
rect 4067 696 4163 698
rect 4263 695 4411 705
rect 4470 725 4507 735
rect 4582 734 4619 735
rect 4563 732 4619 734
rect 4470 705 4478 725
rect 4498 705 4507 725
rect 4319 694 4355 695
rect 3670 648 3707 679
rect 3883 677 3919 679
rect 3883 648 3920 677
rect 3122 639 3157 640
rect 3099 634 3157 639
rect 3099 614 3102 634
rect 3122 620 3157 634
rect 3177 620 3186 640
rect 3122 612 3186 620
rect 3148 611 3186 612
rect 3149 610 3186 611
rect 3252 644 3288 645
rect 3360 644 3396 645
rect 3252 636 3396 644
rect 3252 616 3260 636
rect 3280 616 3312 636
rect 3336 616 3368 636
rect 3388 616 3396 636
rect 3252 610 3396 616
rect 3462 640 3500 648
rect 3568 644 3604 645
rect 3462 620 3471 640
rect 3491 620 3500 640
rect 3462 611 3500 620
rect 3519 637 3604 644
rect 3519 617 3526 637
rect 3547 636 3604 637
rect 3547 617 3576 636
rect 3519 616 3576 617
rect 3596 616 3604 636
rect 3462 610 3499 611
rect 3519 610 3604 616
rect 3670 640 3708 648
rect 3781 644 3817 645
rect 3670 620 3679 640
rect 3699 620 3708 640
rect 3670 611 3708 620
rect 3732 636 3817 644
rect 3732 616 3789 636
rect 3809 616 3817 636
rect 3670 610 3707 611
rect 3732 610 3817 616
rect 3883 640 3921 648
rect 3883 620 3892 640
rect 3912 620 3921 640
rect 4167 635 4204 636
rect 4470 635 4507 705
rect 4532 725 4619 732
rect 4532 722 4590 725
rect 4532 702 4537 722
rect 4558 705 4590 722
rect 4610 705 4619 725
rect 4558 702 4619 705
rect 4532 695 4619 702
rect 4678 725 4715 735
rect 4678 705 4686 725
rect 4706 705 4715 725
rect 4532 694 4563 695
rect 4166 634 4507 635
rect 3883 611 3921 620
rect 4091 629 4507 634
rect 3883 610 3920 611
rect 3306 589 3342 610
rect 3732 589 3763 610
rect 4091 609 4094 629
rect 4114 609 4507 629
rect 4678 634 4715 705
rect 4745 734 4776 787
rect 5078 772 5115 782
rect 5078 754 5087 772
rect 5105 754 5115 772
rect 5078 745 5115 754
rect 4795 734 4832 735
rect 4745 725 4832 734
rect 4745 705 4803 725
rect 4823 705 4832 725
rect 4745 695 4832 705
rect 4891 725 4928 735
rect 4891 705 4899 725
rect 4919 705 4928 725
rect 4745 694 4776 695
rect 4891 634 4928 705
rect 5083 680 5114 745
rect 5082 670 5119 680
rect 5082 668 5092 670
rect 5016 666 5092 668
rect 4678 610 4928 634
rect 5013 652 5092 666
rect 5110 652 5119 670
rect 5013 649 5119 652
rect 4485 590 4506 609
rect 5013 590 5039 649
rect 5082 643 5119 649
rect 3139 585 3239 589
rect 3139 581 3201 585
rect 3139 555 3146 581
rect 3172 559 3201 581
rect 3227 559 3239 585
rect 3172 555 3239 559
rect 3139 552 3239 555
rect 3307 552 3342 589
rect 3404 586 3763 589
rect 3404 581 3626 586
rect 3404 557 3417 581
rect 3441 562 3626 581
rect 3650 562 3763 586
rect 3441 557 3763 562
rect 3404 553 3763 557
rect 3830 581 3979 589
rect 3830 561 3841 581
rect 3861 561 3979 581
rect 4485 572 5039 590
rect 5085 579 5122 581
rect 5013 571 5039 572
rect 5082 571 5122 579
rect 3830 554 3979 561
rect 5082 559 5094 571
rect 5073 554 5094 559
rect 3830 553 3871 554
rect 4489 553 5094 554
rect 5112 553 5122 571
rect 3154 500 3191 501
rect 3250 500 3287 501
rect 3306 500 3342 552
rect 3361 500 3398 501
rect 3054 491 3192 500
rect 3054 471 3163 491
rect 3183 471 3192 491
rect 3054 464 3192 471
rect 3250 491 3398 500
rect 3250 471 3259 491
rect 3279 471 3369 491
rect 3389 471 3398 491
rect 3054 462 3150 464
rect 3250 461 3398 471
rect 3457 491 3494 501
rect 3569 500 3606 501
rect 3550 498 3606 500
rect 3457 471 3465 491
rect 3485 471 3494 491
rect 3306 460 3342 461
rect 3154 401 3191 402
rect 3457 401 3494 471
rect 3519 491 3606 498
rect 3519 488 3577 491
rect 3519 468 3524 488
rect 3545 471 3577 488
rect 3597 471 3606 491
rect 3545 468 3606 471
rect 3519 461 3606 468
rect 3665 491 3702 501
rect 3665 471 3673 491
rect 3693 471 3702 491
rect 3519 460 3550 461
rect 3153 400 3494 401
rect 3078 395 3494 400
rect 3078 375 3081 395
rect 3101 375 3494 395
rect 3665 400 3702 471
rect 3732 500 3763 553
rect 4489 544 5122 553
rect 4489 537 5121 544
rect 4489 535 4551 537
rect 4067 525 4235 526
rect 4489 525 4511 535
rect 3782 500 3819 501
rect 3732 491 3819 500
rect 3732 471 3790 491
rect 3810 471 3819 491
rect 3732 461 3819 471
rect 3878 491 3915 501
rect 3878 471 3886 491
rect 3906 471 3915 491
rect 3732 460 3763 461
rect 3878 400 3915 471
rect 3665 376 3915 400
rect 4067 499 4511 525
rect 4067 497 4235 499
rect 4067 319 4094 497
rect 4134 459 4198 471
rect 4474 467 4511 499
rect 4682 498 4931 520
rect 4682 467 4719 498
rect 4895 496 4931 498
rect 4895 467 4932 496
rect 4134 458 4169 459
rect 4111 453 4169 458
rect 4111 433 4114 453
rect 4134 439 4169 453
rect 4189 439 4198 459
rect 4134 431 4198 439
rect 4160 430 4198 431
rect 4161 429 4198 430
rect 4264 463 4300 464
rect 4372 463 4408 464
rect 4264 455 4408 463
rect 4264 435 4272 455
rect 4292 435 4321 455
rect 4264 434 4321 435
rect 4343 435 4380 455
rect 4400 435 4408 455
rect 4343 434 4408 435
rect 4264 429 4408 434
rect 4474 459 4512 467
rect 4580 463 4616 464
rect 4474 439 4483 459
rect 4503 439 4512 459
rect 4474 430 4512 439
rect 4531 456 4616 463
rect 4531 436 4538 456
rect 4559 455 4616 456
rect 4559 436 4588 455
rect 4531 435 4588 436
rect 4608 435 4616 455
rect 4474 429 4511 430
rect 4531 429 4616 435
rect 4682 459 4720 467
rect 4793 463 4829 464
rect 4682 439 4691 459
rect 4711 439 4720 459
rect 4682 430 4720 439
rect 4744 455 4829 463
rect 4744 435 4801 455
rect 4821 435 4829 455
rect 4682 429 4719 430
rect 4744 429 4829 435
rect 4895 459 4933 467
rect 4895 439 4904 459
rect 4924 439 4933 459
rect 4895 430 4933 439
rect 4895 429 4932 430
rect 4318 408 4354 429
rect 4744 408 4775 429
rect 4151 404 4251 408
rect 4151 400 4213 404
rect 4151 374 4158 400
rect 4184 378 4213 400
rect 4239 378 4251 404
rect 4184 374 4251 378
rect 4151 371 4251 374
rect 4319 371 4354 408
rect 4416 405 4775 408
rect 4416 400 4638 405
rect 4416 376 4429 400
rect 4453 381 4638 400
rect 4662 381 4775 405
rect 4453 376 4775 381
rect 4416 372 4775 376
rect 4842 400 4991 408
rect 4842 380 4853 400
rect 4873 380 4991 400
rect 4842 373 4991 380
rect 5082 388 5121 537
rect 4842 372 4883 373
rect 4166 319 4203 320
rect 4262 319 4299 320
rect 4318 319 4354 371
rect 4373 319 4410 320
rect 2231 274 2236 300
rect 2255 274 2262 300
rect 4066 310 4204 319
rect 4066 290 4175 310
rect 4195 290 4204 310
rect 4066 283 4204 290
rect 4262 310 4410 319
rect 4262 290 4271 310
rect 4291 290 4381 310
rect 4401 290 4410 310
rect 4066 281 4162 283
rect 4262 280 4410 290
rect 4469 310 4506 320
rect 4581 319 4618 320
rect 4562 317 4618 319
rect 4469 290 4477 310
rect 4497 290 4506 310
rect 4318 279 4354 280
rect 2231 271 2262 274
rect 1060 247 1198 256
rect 854 246 891 247
rect 910 195 946 247
rect 965 246 1002 247
rect 1061 246 1098 247
rect 381 193 422 194
rect 273 186 422 193
rect 273 166 391 186
rect 411 166 422 186
rect 273 158 422 166
rect 489 190 848 194
rect 489 185 811 190
rect 489 161 602 185
rect 626 166 811 185
rect 835 166 848 190
rect 626 161 848 166
rect 489 158 848 161
rect 910 158 945 195
rect 1013 192 1113 195
rect 1013 188 1080 192
rect 1013 162 1025 188
rect 1051 166 1080 188
rect 1106 166 1113 192
rect 1051 162 1113 166
rect 1013 158 1113 162
rect 489 137 520 158
rect 910 137 946 158
rect 153 128 190 137
rect 332 136 369 137
rect 153 110 162 128
rect 180 110 190 128
rect 153 100 190 110
rect 154 65 190 100
rect 331 127 369 136
rect 331 107 340 127
rect 360 107 369 127
rect 331 99 369 107
rect 435 131 520 137
rect 545 136 582 137
rect 435 111 443 131
rect 463 111 520 131
rect 435 103 520 111
rect 544 127 582 136
rect 544 107 553 127
rect 573 107 582 127
rect 435 102 471 103
rect 544 99 582 107
rect 648 131 733 137
rect 753 136 790 137
rect 648 111 656 131
rect 676 130 733 131
rect 676 111 705 130
rect 648 110 705 111
rect 726 110 733 130
rect 648 103 733 110
rect 752 127 790 136
rect 752 107 761 127
rect 781 107 790 127
rect 648 102 684 103
rect 752 99 790 107
rect 856 131 1000 137
rect 856 111 864 131
rect 884 130 972 131
rect 884 111 912 130
rect 856 109 912 111
rect 934 111 972 130
rect 992 111 1000 131
rect 934 109 1000 111
rect 856 103 1000 109
rect 856 102 892 103
rect 964 102 1000 103
rect 1066 136 1103 137
rect 1066 135 1104 136
rect 1066 127 1130 135
rect 1066 107 1075 127
rect 1095 113 1130 127
rect 1150 113 1153 133
rect 1095 108 1153 113
rect 1095 107 1130 108
rect 332 70 369 99
rect 152 0 190 65
rect 333 68 369 70
rect 545 68 582 99
rect 333 46 582 68
rect 753 67 790 99
rect 1066 95 1130 107
rect 1170 69 1197 247
rect 4166 220 4203 221
rect 4469 220 4506 290
rect 4531 310 4618 317
rect 4531 307 4589 310
rect 4531 287 4536 307
rect 4557 290 4589 307
rect 4609 290 4618 310
rect 4557 287 4618 290
rect 4531 280 4618 287
rect 4677 310 4714 320
rect 4677 290 4685 310
rect 4705 290 4714 310
rect 4531 279 4562 280
rect 4165 219 4506 220
rect 4090 214 4506 219
rect 4090 194 4093 214
rect 4113 194 4506 214
rect 4677 219 4714 290
rect 4744 319 4775 372
rect 5082 370 5092 388
rect 5110 370 5121 388
rect 5082 361 5119 370
rect 4794 319 4831 320
rect 4744 310 4831 319
rect 4744 290 4802 310
rect 4822 290 4831 310
rect 4744 280 4831 290
rect 4890 310 4927 320
rect 4890 290 4898 310
rect 4918 290 4927 310
rect 5085 295 5122 299
rect 4744 279 4775 280
rect 4890 219 4927 290
rect 4677 195 4927 219
rect 5083 289 5122 295
rect 5083 271 5094 289
rect 5112 271 5122 289
rect 5083 262 5122 271
rect 4469 171 4506 194
rect 5083 184 5118 262
rect 5080 174 5118 184
rect 4469 170 4639 171
rect 5080 170 5090 174
rect 4469 156 5090 170
rect 5108 156 5118 174
rect 4469 150 5118 156
rect 4469 149 5117 150
rect 5080 147 5117 149
rect 5083 83 5120 85
rect 1029 67 1197 69
rect 753 41 1197 67
rect 754 15 778 41
rect 1029 40 1197 41
rect 5078 75 5120 83
rect 5078 57 5092 75
rect 5110 57 5120 75
rect 5078 48 5120 57
rect 747 7 787 15
rect 747 0 756 7
rect 152 -15 756 0
rect 779 -15 787 7
rect 152 -18 787 -15
rect 152 -24 190 -18
rect 747 -30 787 -18
rect 5078 7 5119 48
rect 5078 -15 5089 7
rect 5112 -15 5119 7
rect 5078 -20 5119 -15
rect 1740 -134 1990 -110
rect 1740 -205 1777 -134
rect 1892 -195 1923 -194
rect 1740 -225 1749 -205
rect 1769 -225 1777 -205
rect 1740 -235 1777 -225
rect 1836 -205 1923 -195
rect 1836 -225 1845 -205
rect 1865 -225 1923 -205
rect 1836 -234 1923 -225
rect 1836 -235 1873 -234
rect 1892 -287 1923 -234
rect 1953 -205 1990 -134
rect 2161 -129 2554 -109
rect 2574 -129 2577 -109
rect 2161 -134 2577 -129
rect 2161 -135 2502 -134
rect 2105 -195 2136 -194
rect 1953 -225 1962 -205
rect 1982 -225 1990 -205
rect 1953 -235 1990 -225
rect 2049 -202 2136 -195
rect 2049 -205 2110 -202
rect 2049 -225 2058 -205
rect 2078 -222 2110 -205
rect 2131 -222 2136 -202
rect 2078 -225 2136 -222
rect 2049 -232 2136 -225
rect 2161 -205 2198 -135
rect 2464 -136 2501 -135
rect 2313 -195 2349 -194
rect 2161 -225 2170 -205
rect 2190 -225 2198 -205
rect 2049 -234 2105 -232
rect 2049 -235 2086 -234
rect 2161 -235 2198 -225
rect 2257 -205 2405 -195
rect 2505 -198 2601 -196
rect 2257 -225 2266 -205
rect 2286 -225 2376 -205
rect 2396 -225 2405 -205
rect 2257 -234 2405 -225
rect 2463 -199 2601 -198
rect 2463 -204 2687 -199
rect 2463 -205 2651 -204
rect 2463 -225 2472 -205
rect 2492 -224 2651 -205
rect 2679 -224 2687 -204
rect 2492 -225 2687 -224
rect 2463 -232 2687 -225
rect 2463 -234 2601 -232
rect 2257 -235 2294 -234
rect 2313 -286 2349 -234
rect 2368 -235 2405 -234
rect 2464 -235 2501 -234
rect 1784 -288 1825 -287
rect 1676 -295 1825 -288
rect 1676 -315 1794 -295
rect 1814 -315 1825 -295
rect 1676 -323 1825 -315
rect 1892 -291 2251 -287
rect 1892 -296 2214 -291
rect 1892 -320 2005 -296
rect 2029 -315 2214 -296
rect 2238 -315 2251 -291
rect 2029 -320 2251 -315
rect 1892 -323 2251 -320
rect 2313 -323 2348 -286
rect 2416 -289 2516 -286
rect 2416 -293 2483 -289
rect 2416 -319 2428 -293
rect 2454 -315 2483 -293
rect 2509 -315 2516 -289
rect 2454 -319 2516 -315
rect 2416 -323 2516 -319
rect 1892 -344 1923 -323
rect 2313 -344 2349 -323
rect 1735 -345 1772 -344
rect 1734 -354 1772 -345
rect 1734 -374 1743 -354
rect 1763 -374 1772 -354
rect 1734 -382 1772 -374
rect 1838 -350 1923 -344
rect 1948 -345 1985 -344
rect 1838 -370 1846 -350
rect 1866 -370 1923 -350
rect 1838 -378 1923 -370
rect 1947 -354 1985 -345
rect 1947 -374 1956 -354
rect 1976 -374 1985 -354
rect 1838 -379 1874 -378
rect 1947 -382 1985 -374
rect 2051 -350 2136 -344
rect 2156 -345 2193 -344
rect 2051 -370 2059 -350
rect 2079 -351 2136 -350
rect 2079 -370 2108 -351
rect 2051 -371 2108 -370
rect 2129 -371 2136 -351
rect 2051 -378 2136 -371
rect 2155 -354 2193 -345
rect 2155 -374 2164 -354
rect 2184 -374 2193 -354
rect 2051 -379 2087 -378
rect 2155 -382 2193 -374
rect 2259 -350 2403 -344
rect 2259 -370 2267 -350
rect 2287 -351 2375 -350
rect 2287 -370 2322 -351
rect 2259 -373 2322 -370
rect 2347 -370 2375 -351
rect 2395 -370 2403 -350
rect 2347 -373 2403 -370
rect 2259 -378 2403 -373
rect 2259 -379 2295 -378
rect 2367 -379 2403 -378
rect 2469 -345 2506 -344
rect 2469 -346 2507 -345
rect 2469 -354 2533 -346
rect 2469 -374 2478 -354
rect 2498 -368 2533 -354
rect 2553 -368 2556 -348
rect 2498 -373 2556 -368
rect 2498 -374 2533 -373
rect 1735 -411 1772 -382
rect 1736 -413 1772 -411
rect 1948 -413 1985 -382
rect 1736 -435 1985 -413
rect 2156 -414 2193 -382
rect 2469 -386 2533 -374
rect 2573 -412 2600 -234
rect 2432 -414 2600 -412
rect 2156 -440 2600 -414
rect 2432 -441 2600 -440
<< viali >>
rect 1115 7625 1135 7645
rect 671 7532 692 7552
rect 4078 7706 4098 7726
rect 4294 7709 4316 7730
rect 4502 7709 4523 7729
rect 4122 7647 4148 7673
rect 2973 7539 2992 7565
rect 1044 7439 1070 7465
rect 669 7383 690 7403
rect 885 7384 907 7405
rect 1094 7386 1114 7406
rect 2127 7444 2147 7464
rect 1683 7351 1704 7371
rect 2056 7258 2082 7284
rect 1114 7210 1134 7230
rect 670 7117 691 7137
rect 1681 7202 1702 7222
rect 1892 7203 1916 7223
rect 2106 7205 2126 7225
rect 1778 7136 1798 7155
rect 2880 7123 2900 7141
rect 3393 7542 3413 7561
rect 3065 7472 3085 7492
rect 3276 7473 3300 7493
rect 3489 7475 3510 7495
rect 4500 7560 4521 7580
rect 4057 7467 4077 7487
rect 3109 7413 3135 7439
rect 3487 7326 3508 7346
rect 3044 7233 3064 7253
rect 4077 7291 4097 7311
rect 4284 7292 4306 7313
rect 4501 7294 4522 7314
rect 4121 7232 4147 7258
rect 1043 7024 1069 7050
rect 668 6968 689 6988
rect 875 6967 897 6988
rect 1093 6971 1113 6991
rect 2182 6883 2202 6903
rect 1738 6790 1759 6810
rect 2111 6697 2137 6723
rect 1120 6644 1140 6664
rect 676 6551 697 6571
rect 1736 6641 1757 6661
rect 1951 6643 1975 6660
rect 2161 6644 2181 6664
rect 1049 6458 1075 6484
rect 674 6402 695 6422
rect 890 6403 912 6424
rect 1099 6405 1119 6425
rect 2132 6463 2152 6483
rect 1688 6370 1709 6390
rect 2061 6277 2087 6303
rect 1119 6229 1139 6249
rect 675 6136 696 6156
rect 1686 6221 1707 6241
rect 1896 6223 1920 6243
rect 2111 6224 2131 6244
rect 1783 6155 1803 6174
rect 2204 6151 2223 6177
rect 1048 6043 1074 6069
rect 673 5987 694 6007
rect 880 5986 902 6007
rect 1098 5990 1118 6010
rect 3015 7052 3035 7072
rect 3225 7055 3248 7074
rect 3439 7055 3460 7075
rect 4499 7145 4520 7165
rect 4056 7052 4076 7072
rect 3059 6993 3085 7019
rect 3437 6906 3458 6926
rect 2994 6813 3014 6833
rect 4083 6725 4103 6745
rect 4299 6728 4321 6749
rect 4507 6728 4528 6748
rect 4127 6666 4153 6692
rect 3398 6561 3418 6580
rect 3070 6491 3090 6511
rect 3280 6493 3304 6513
rect 3494 6494 3515 6514
rect 4505 6579 4526 6599
rect 4062 6486 4082 6506
rect 3114 6432 3140 6458
rect 3492 6345 3513 6365
rect 3049 6252 3069 6272
rect 4082 6310 4102 6330
rect 4289 6311 4311 6332
rect 4506 6313 4527 6333
rect 4126 6251 4152 6277
rect 2757 6094 2780 6113
rect 2347 5951 2367 5971
rect 1903 5858 1924 5878
rect 2276 5765 2302 5791
rect 1901 5709 1922 5729
rect 2110 5708 2135 5734
rect 2326 5712 2346 5732
rect 1127 5665 1147 5685
rect 683 5572 704 5592
rect 1056 5479 1082 5505
rect 681 5423 702 5443
rect 897 5424 919 5445
rect 1106 5426 1126 5446
rect 2139 5484 2159 5504
rect 1695 5391 1716 5411
rect 2068 5298 2094 5324
rect 1126 5250 1146 5270
rect 682 5157 703 5177
rect 1693 5242 1714 5262
rect 1904 5243 1928 5263
rect 2118 5245 2138 5265
rect 1790 5176 1810 5195
rect 1055 5064 1081 5090
rect 680 5008 701 5028
rect 887 5007 909 5028
rect 1105 5011 1125 5031
rect 2194 4923 2214 4943
rect 1750 4830 1771 4850
rect 2123 4737 2149 4763
rect 1132 4684 1152 4704
rect 688 4591 709 4611
rect 1748 4681 1769 4701
rect 1960 4682 1983 4701
rect 2173 4684 2193 4704
rect 1061 4498 1087 4524
rect 686 4442 707 4462
rect 902 4443 924 4464
rect 1111 4445 1131 4465
rect 2144 4503 2164 4523
rect 1700 4410 1721 4430
rect 2073 4317 2099 4343
rect 1131 4269 1151 4289
rect 687 4176 708 4196
rect 1698 4261 1719 4281
rect 1908 4263 1932 4283
rect 2123 4264 2143 4284
rect 1795 4195 1815 4214
rect 2308 4615 2328 4633
rect 2216 4191 2235 4217
rect 4504 6164 4525 6184
rect 4061 6071 4081 6091
rect 2862 6024 2882 6044
rect 3069 6026 3092 6045
rect 3286 6027 3307 6047
rect 2906 5965 2932 5991
rect 3284 5878 3305 5898
rect 2841 5785 2861 5805
rect 4090 5746 4110 5766
rect 4306 5749 4328 5770
rect 4514 5749 4535 5769
rect 4134 5687 4160 5713
rect 2985 5579 3004 5605
rect 3405 5582 3425 5601
rect 3077 5512 3097 5532
rect 3288 5513 3312 5533
rect 3501 5515 3522 5535
rect 4512 5600 4533 5620
rect 4069 5507 4089 5527
rect 3121 5453 3147 5479
rect 3499 5366 3520 5386
rect 3056 5273 3076 5293
rect 4089 5331 4109 5351
rect 4296 5332 4318 5353
rect 4513 5334 4534 5354
rect 4133 5272 4159 5298
rect 3027 5092 3047 5112
rect 3233 5096 3257 5113
rect 3451 5095 3472 5115
rect 4511 5185 4532 5205
rect 4068 5092 4088 5112
rect 3071 5033 3097 5059
rect 3449 4946 3470 4966
rect 3006 4853 3026 4873
rect 4095 4765 4115 4785
rect 4311 4768 4333 4789
rect 4519 4768 4540 4788
rect 4139 4706 4165 4732
rect 3410 4601 3430 4620
rect 3082 4531 3102 4551
rect 3292 4533 3316 4553
rect 3506 4534 3527 4554
rect 4517 4619 4538 4639
rect 4074 4526 4094 4546
rect 3126 4472 3152 4498
rect 3504 4385 3525 4405
rect 3061 4292 3081 4312
rect 4094 4350 4114 4370
rect 4301 4351 4323 4372
rect 4518 4353 4539 4373
rect 4138 4291 4164 4317
rect 1060 4083 1086 4109
rect 685 4027 706 4047
rect 892 4026 914 4047
rect 1110 4030 1130 4050
rect 4516 4204 4537 4224
rect 2787 4099 2807 4119
rect 2991 4100 3017 4119
rect 3211 4102 3232 4122
rect 4073 4111 4093 4131
rect 2831 4040 2857 4066
rect 2442 3959 2462 3979
rect 1998 3866 2019 3886
rect 3209 3953 3230 3973
rect 2766 3860 2786 3880
rect 2371 3773 2397 3799
rect 1135 3708 1155 3728
rect 1996 3717 2017 3737
rect 2211 3720 2237 3739
rect 2421 3720 2441 3740
rect 691 3615 712 3635
rect 4098 3789 4118 3809
rect 4314 3792 4336 3813
rect 4522 3792 4543 3812
rect 4142 3730 4168 3756
rect 1064 3522 1090 3548
rect 689 3466 710 3486
rect 905 3467 927 3488
rect 1114 3469 1134 3489
rect 2147 3527 2167 3547
rect 1703 3434 1724 3454
rect 2076 3341 2102 3367
rect 1134 3293 1154 3313
rect 690 3200 711 3220
rect 1701 3285 1722 3305
rect 1912 3286 1936 3306
rect 2126 3288 2146 3308
rect 1798 3219 1818 3238
rect 1063 3107 1089 3133
rect 688 3051 709 3071
rect 895 3050 917 3071
rect 1113 3054 1133 3074
rect 2202 2966 2222 2986
rect 1758 2873 1779 2893
rect 2131 2780 2157 2806
rect 1140 2727 1160 2747
rect 696 2634 717 2654
rect 1756 2724 1777 2744
rect 1971 2726 1995 2743
rect 2181 2727 2201 2747
rect 1069 2541 1095 2567
rect 694 2485 715 2505
rect 910 2486 932 2507
rect 1119 2488 1139 2508
rect 2152 2546 2172 2566
rect 1708 2453 1729 2473
rect 2081 2360 2107 2386
rect 1139 2312 1159 2332
rect 695 2219 716 2239
rect 1706 2304 1727 2324
rect 1916 2306 1940 2326
rect 2131 2307 2151 2327
rect 1803 2238 1823 2257
rect 2224 2234 2243 2260
rect 1068 2126 1094 2152
rect 693 2070 714 2090
rect 900 2069 922 2090
rect 1118 2073 1138 2093
rect 2367 2034 2387 2054
rect 1923 1941 1944 1961
rect 2296 1848 2322 1874
rect 1921 1792 1942 1812
rect 2136 1794 2159 1813
rect 2346 1795 2366 1815
rect 1147 1748 1167 1768
rect 703 1655 724 1675
rect 2993 3622 3012 3648
rect 2900 3206 2920 3224
rect 3413 3625 3433 3644
rect 3085 3555 3105 3575
rect 3296 3556 3320 3576
rect 3509 3558 3530 3578
rect 4520 3643 4541 3663
rect 4077 3550 4097 3570
rect 3129 3496 3155 3522
rect 3507 3409 3528 3429
rect 3064 3316 3084 3336
rect 4097 3374 4117 3394
rect 4304 3375 4326 3396
rect 4521 3377 4542 3397
rect 4141 3315 4167 3341
rect 3035 3135 3055 3155
rect 3245 3138 3268 3157
rect 3459 3138 3480 3158
rect 4519 3228 4540 3248
rect 4076 3135 4096 3155
rect 3079 3076 3105 3102
rect 3457 2989 3478 3009
rect 3014 2896 3034 2916
rect 4103 2808 4123 2828
rect 4319 2811 4341 2832
rect 4527 2811 4548 2831
rect 4147 2749 4173 2775
rect 3418 2644 3438 2663
rect 3090 2574 3110 2594
rect 3300 2576 3324 2596
rect 3514 2577 3535 2597
rect 4525 2662 4546 2682
rect 4082 2569 4102 2589
rect 3134 2515 3160 2541
rect 3512 2428 3533 2448
rect 3069 2335 3089 2355
rect 4102 2393 4122 2413
rect 4309 2394 4331 2415
rect 4526 2396 4547 2416
rect 4146 2334 4172 2360
rect 4524 2247 4545 2267
rect 4081 2154 4101 2174
rect 2882 2107 2902 2127
rect 3093 2105 3118 2131
rect 3306 2110 3327 2130
rect 2926 2048 2952 2074
rect 3304 1961 3325 1981
rect 2861 1868 2881 1888
rect 2448 1726 2471 1745
rect 1076 1562 1102 1588
rect 701 1506 722 1526
rect 917 1507 939 1528
rect 1126 1509 1146 1529
rect 2159 1567 2179 1587
rect 1715 1474 1736 1494
rect 2088 1381 2114 1407
rect 1146 1333 1166 1353
rect 702 1240 723 1260
rect 1713 1325 1734 1345
rect 1924 1326 1948 1346
rect 2138 1328 2158 1348
rect 1810 1259 1830 1278
rect 1075 1147 1101 1173
rect 700 1091 721 1111
rect 907 1090 929 1111
rect 1125 1094 1145 1114
rect 2214 1006 2234 1026
rect 1770 913 1791 933
rect 2143 820 2169 846
rect 1152 767 1172 787
rect 708 674 729 694
rect 1768 764 1789 784
rect 1980 765 2003 784
rect 2193 767 2213 787
rect 4110 1829 4130 1849
rect 4326 1832 4348 1853
rect 4534 1832 4555 1852
rect 4154 1770 4180 1796
rect 3005 1662 3024 1688
rect 3425 1665 3445 1684
rect 3097 1595 3117 1615
rect 3308 1596 3332 1616
rect 3521 1598 3542 1618
rect 4532 1683 4553 1703
rect 4089 1590 4109 1610
rect 3141 1536 3167 1562
rect 3519 1449 3540 1469
rect 3076 1356 3096 1376
rect 4109 1414 4129 1434
rect 4316 1415 4338 1436
rect 4533 1417 4554 1437
rect 4153 1355 4179 1381
rect 3047 1175 3067 1195
rect 3253 1179 3277 1196
rect 3471 1178 3492 1198
rect 4531 1268 4552 1288
rect 4088 1175 4108 1195
rect 3091 1116 3117 1142
rect 3469 1029 3490 1049
rect 3026 936 3046 956
rect 4115 848 4135 868
rect 4331 851 4353 872
rect 4539 851 4560 871
rect 4159 789 4185 815
rect 1081 581 1107 607
rect 706 525 727 545
rect 922 526 944 547
rect 1131 528 1151 548
rect 2164 586 2184 606
rect 1720 493 1741 513
rect 2093 400 2119 426
rect 1151 352 1171 372
rect 707 259 728 279
rect 1718 344 1739 364
rect 1928 346 1952 366
rect 2143 347 2163 367
rect 1815 278 1835 297
rect 2328 698 2348 716
rect 3430 684 3450 703
rect 3102 614 3122 634
rect 3312 616 3336 636
rect 3526 617 3547 637
rect 4537 702 4558 722
rect 4094 609 4114 629
rect 3146 555 3172 581
rect 3524 468 3545 488
rect 3081 375 3101 395
rect 4114 433 4134 453
rect 4321 434 4343 455
rect 4538 436 4559 456
rect 4158 374 4184 400
rect 2236 274 2255 300
rect 1080 166 1106 192
rect 705 110 726 130
rect 912 109 934 130
rect 1130 113 1150 133
rect 4536 287 4557 307
rect 4093 194 4113 214
rect 756 -15 779 7
rect 5089 -15 5112 7
rect 2554 -129 2574 -109
rect 2110 -222 2131 -202
rect 2651 -224 2679 -204
rect 2483 -315 2509 -289
rect 2108 -371 2129 -351
rect 2322 -373 2347 -351
rect 2533 -368 2553 -348
<< metal1 >>
rect 3914 7800 4323 7801
rect 3908 7771 4323 7800
rect 1111 7650 1143 7651
rect 1108 7645 1143 7650
rect 1108 7625 1115 7645
rect 1135 7625 1143 7645
rect 1108 7617 1143 7625
rect 3908 7620 3948 7771
rect 4282 7738 4323 7771
rect 4070 7733 4105 7734
rect 664 7552 696 7559
rect 664 7532 671 7552
rect 692 7532 696 7552
rect 664 7467 696 7532
rect 1034 7467 1074 7468
rect 664 7465 1076 7467
rect 664 7439 1044 7465
rect 1070 7439 1076 7465
rect 664 7431 1076 7439
rect 664 7403 696 7431
rect 1109 7411 1143 7617
rect 3385 7592 3948 7620
rect 4049 7726 4105 7733
rect 4049 7706 4078 7726
rect 4098 7706 4105 7726
rect 4049 7701 4105 7706
rect 4278 7730 4328 7738
rect 4278 7709 4294 7730
rect 4316 7709 4328 7730
rect 2964 7565 3311 7569
rect 2964 7539 2973 7565
rect 2992 7539 3311 7565
rect 3386 7564 3420 7592
rect 2964 7534 3311 7539
rect 3385 7561 3421 7564
rect 3385 7542 3393 7561
rect 3413 7542 3421 7561
rect 3385 7538 3421 7542
rect 3271 7504 3311 7534
rect 3057 7499 3092 7500
rect 664 7383 669 7403
rect 690 7383 696 7403
rect 664 7376 696 7383
rect 873 7405 913 7410
rect 873 7384 885 7405
rect 907 7384 913 7405
rect 873 7372 913 7384
rect 1087 7406 1143 7411
rect 1087 7386 1094 7406
rect 1114 7386 1143 7406
rect 1087 7379 1143 7386
rect 1200 7480 2157 7499
rect 3036 7492 3092 7499
rect 1087 7378 1122 7379
rect 879 7340 907 7372
rect 1200 7340 1231 7480
rect 2120 7464 2155 7480
rect 2120 7444 2127 7464
rect 2147 7444 2155 7464
rect 2120 7436 2155 7444
rect 879 7309 1231 7340
rect 1676 7371 1708 7378
rect 1676 7351 1683 7371
rect 1704 7351 1708 7371
rect 1676 7286 1708 7351
rect 2046 7286 2086 7287
rect 1676 7284 2088 7286
rect 1676 7258 2056 7284
rect 2082 7258 2088 7284
rect 1676 7250 2088 7258
rect 1110 7235 1142 7236
rect 1107 7230 1142 7235
rect 1107 7210 1114 7230
rect 1134 7210 1142 7230
rect 1107 7202 1142 7210
rect 663 7137 695 7144
rect 663 7117 670 7137
rect 691 7117 695 7137
rect 663 7052 695 7117
rect 1033 7052 1073 7053
rect 663 7050 1075 7052
rect 663 7024 1043 7050
rect 1069 7024 1075 7050
rect 663 7016 1075 7024
rect 663 6988 695 7016
rect 663 6968 668 6988
rect 689 6968 695 6988
rect 663 6961 695 6968
rect 863 6988 913 6997
rect 1108 6996 1142 7202
rect 1676 7222 1708 7250
rect 1676 7202 1681 7222
rect 1702 7202 1708 7222
rect 1676 7195 1708 7202
rect 1883 7223 1925 7231
rect 2121 7230 2155 7436
rect 1883 7203 1892 7223
rect 1916 7203 1925 7223
rect 1883 7191 1925 7203
rect 2099 7225 2155 7230
rect 2099 7205 2106 7225
rect 2126 7205 2155 7225
rect 3036 7472 3065 7492
rect 3085 7472 3092 7492
rect 3036 7467 3092 7472
rect 3268 7493 3311 7504
rect 3268 7473 3276 7493
rect 3300 7487 3311 7493
rect 3483 7495 3515 7502
rect 3300 7473 3310 7487
rect 3036 7261 3070 7467
rect 3268 7464 3310 7473
rect 3483 7475 3489 7495
rect 3510 7475 3515 7495
rect 3483 7447 3515 7475
rect 4049 7495 4083 7701
rect 4278 7700 4328 7709
rect 4496 7729 4528 7736
rect 4496 7709 4502 7729
rect 4523 7709 4528 7729
rect 4496 7681 4528 7709
rect 4116 7673 4528 7681
rect 4116 7647 4122 7673
rect 4148 7647 4528 7673
rect 4116 7645 4528 7647
rect 4118 7644 4158 7645
rect 4496 7580 4528 7645
rect 4496 7560 4500 7580
rect 4521 7560 4528 7580
rect 4496 7553 4528 7560
rect 4049 7487 4084 7495
rect 4049 7467 4057 7487
rect 4077 7467 4084 7487
rect 4049 7462 4084 7467
rect 4049 7461 4081 7462
rect 3103 7439 3515 7447
rect 3103 7413 3109 7439
rect 3135 7413 3515 7439
rect 3103 7411 3515 7413
rect 3105 7410 3145 7411
rect 3483 7346 3515 7411
rect 3483 7326 3487 7346
rect 3508 7326 3515 7346
rect 3483 7319 3515 7326
rect 3960 7357 4312 7388
rect 3036 7253 3071 7261
rect 3036 7233 3044 7253
rect 3064 7233 3071 7253
rect 3036 7217 3071 7233
rect 3960 7217 3991 7357
rect 4284 7325 4312 7357
rect 4069 7318 4104 7319
rect 2099 7198 2155 7205
rect 3034 7198 3991 7217
rect 4048 7311 4104 7318
rect 4048 7291 4077 7311
rect 4097 7291 4104 7311
rect 4048 7286 4104 7291
rect 4278 7313 4318 7325
rect 4278 7292 4284 7313
rect 4306 7292 4318 7313
rect 4278 7287 4318 7292
rect 4495 7314 4527 7321
rect 4495 7294 4501 7314
rect 4522 7294 4527 7314
rect 2099 7197 2134 7198
rect 1885 7162 1920 7191
rect 1885 7161 2195 7162
rect 1770 7155 1806 7159
rect 1770 7136 1778 7155
rect 1798 7136 1806 7155
rect 1770 7133 1806 7136
rect 1771 7105 1805 7133
rect 1885 7127 2212 7161
rect 863 6967 875 6988
rect 897 6967 913 6988
rect 863 6959 913 6967
rect 1086 6991 1142 6996
rect 1086 6971 1093 6991
rect 1113 6971 1142 6991
rect 1086 6964 1142 6971
rect 1243 7077 1806 7105
rect 1086 6963 1121 6964
rect 868 6926 909 6959
rect 1243 6926 1283 7077
rect 868 6897 1283 6926
rect 2172 6903 2212 7127
rect 2873 7146 2902 7148
rect 2873 7141 3246 7146
rect 2873 7123 2880 7141
rect 2900 7123 3246 7141
rect 2873 7118 3246 7123
rect 2878 7116 3246 7118
rect 3007 7079 3042 7080
rect 3222 7079 3246 7116
rect 868 6896 1277 6897
rect 2172 6883 2182 6903
rect 2202 6883 2212 6903
rect 2172 6873 2212 6883
rect 2986 7072 3042 7079
rect 2986 7052 3015 7072
rect 3035 7052 3042 7072
rect 2986 7047 3042 7052
rect 3217 7074 3254 7079
rect 3217 7055 3225 7074
rect 3248 7055 3254 7074
rect 3217 7049 3254 7055
rect 3433 7075 3465 7082
rect 3433 7055 3439 7075
rect 3460 7055 3465 7075
rect 1731 6810 1763 6817
rect 1731 6790 1738 6810
rect 1759 6790 1763 6810
rect 1731 6725 1763 6790
rect 2101 6725 2141 6726
rect 1731 6723 2143 6725
rect 1731 6697 2111 6723
rect 2137 6697 2143 6723
rect 1731 6689 2143 6697
rect 1116 6669 1148 6670
rect 1113 6664 1148 6669
rect 1113 6644 1120 6664
rect 1140 6644 1148 6664
rect 1113 6636 1148 6644
rect 669 6571 701 6578
rect 669 6551 676 6571
rect 697 6551 701 6571
rect 669 6486 701 6551
rect 1039 6486 1079 6487
rect 669 6484 1081 6486
rect 669 6458 1049 6484
rect 1075 6458 1081 6484
rect 669 6450 1081 6458
rect 669 6422 701 6450
rect 1114 6430 1148 6636
rect 1731 6661 1763 6689
rect 1731 6641 1736 6661
rect 1757 6641 1763 6661
rect 1731 6634 1763 6641
rect 1942 6660 1980 6672
rect 2176 6669 2210 6873
rect 2986 6843 3020 7047
rect 3433 7027 3465 7055
rect 4048 7080 4082 7286
rect 4495 7266 4527 7294
rect 4115 7258 4527 7266
rect 4115 7232 4121 7258
rect 4147 7232 4527 7258
rect 4115 7230 4527 7232
rect 4117 7229 4157 7230
rect 4495 7165 4527 7230
rect 4495 7145 4499 7165
rect 4520 7145 4527 7165
rect 4495 7138 4527 7145
rect 4048 7072 4083 7080
rect 4048 7052 4056 7072
rect 4076 7052 4083 7072
rect 4048 7047 4083 7052
rect 4048 7046 4080 7047
rect 3053 7019 3465 7027
rect 3053 6993 3059 7019
rect 3085 6993 3465 7019
rect 3053 6991 3465 6993
rect 3055 6990 3095 6991
rect 3433 6926 3465 6991
rect 3433 6906 3437 6926
rect 3458 6906 3465 6926
rect 3433 6899 3465 6906
rect 1942 6643 1951 6660
rect 1975 6643 1980 6660
rect 1942 6600 1980 6643
rect 2154 6664 2210 6669
rect 2154 6644 2161 6664
rect 2181 6644 2210 6664
rect 2154 6637 2210 6644
rect 2984 6833 3024 6843
rect 2984 6813 2994 6833
rect 3014 6813 3024 6833
rect 3919 6819 4328 6820
rect 2154 6636 2189 6637
rect 2288 6600 2372 6605
rect 1942 6571 2372 6600
rect 669 6402 674 6422
rect 695 6402 701 6422
rect 669 6395 701 6402
rect 878 6424 918 6429
rect 878 6403 890 6424
rect 912 6403 918 6424
rect 878 6391 918 6403
rect 1092 6425 1148 6430
rect 1092 6405 1099 6425
rect 1119 6405 1148 6425
rect 1092 6398 1148 6405
rect 1205 6499 2162 6518
rect 1092 6397 1127 6398
rect 884 6359 912 6391
rect 1205 6359 1236 6499
rect 2125 6483 2160 6499
rect 2125 6463 2132 6483
rect 2152 6463 2160 6483
rect 2125 6455 2160 6463
rect 884 6328 1236 6359
rect 1681 6390 1713 6397
rect 1681 6370 1688 6390
rect 1709 6370 1713 6390
rect 1681 6305 1713 6370
rect 2051 6305 2091 6306
rect 1681 6303 2093 6305
rect 1681 6277 2061 6303
rect 2087 6277 2093 6303
rect 1681 6269 2093 6277
rect 1115 6254 1147 6255
rect 1112 6249 1147 6254
rect 1112 6229 1119 6249
rect 1139 6229 1147 6249
rect 1112 6221 1147 6229
rect 668 6156 700 6163
rect 668 6136 675 6156
rect 696 6136 700 6156
rect 668 6071 700 6136
rect 1038 6071 1078 6072
rect 668 6069 1080 6071
rect 668 6043 1048 6069
rect 1074 6043 1080 6069
rect 668 6035 1080 6043
rect 668 6007 700 6035
rect 668 5987 673 6007
rect 694 5987 700 6007
rect 668 5980 700 5987
rect 868 6007 918 6016
rect 1113 6015 1147 6221
rect 1681 6241 1713 6269
rect 1681 6221 1686 6241
rect 1707 6221 1713 6241
rect 1886 6243 1928 6252
rect 2126 6249 2160 6455
rect 1886 6229 1896 6243
rect 1681 6214 1713 6221
rect 1885 6223 1896 6229
rect 1920 6223 1928 6243
rect 1885 6212 1928 6223
rect 2104 6244 2160 6249
rect 2104 6224 2111 6244
rect 2131 6224 2160 6244
rect 2104 6217 2160 6224
rect 2104 6216 2139 6217
rect 1885 6182 1925 6212
rect 1775 6174 1811 6178
rect 1775 6155 1783 6174
rect 1803 6155 1811 6174
rect 1775 6152 1811 6155
rect 1885 6177 2232 6182
rect 1776 6124 1810 6152
rect 1885 6151 2204 6177
rect 2223 6151 2232 6177
rect 1885 6147 2232 6151
rect 868 5986 880 6007
rect 902 5986 918 6007
rect 868 5978 918 5986
rect 1091 6010 1147 6015
rect 1091 5990 1098 6010
rect 1118 5990 1147 6010
rect 1091 5983 1147 5990
rect 1248 6096 1811 6124
rect 1091 5982 1126 5983
rect 873 5945 914 5978
rect 1248 5945 1288 6096
rect 2337 5977 2372 6571
rect 2984 6589 3024 6813
rect 3913 6790 4328 6819
rect 3913 6639 3953 6790
rect 4287 6757 4328 6790
rect 4075 6752 4110 6753
rect 3390 6611 3953 6639
rect 4054 6745 4110 6752
rect 4054 6725 4083 6745
rect 4103 6725 4110 6745
rect 4054 6720 4110 6725
rect 4283 6749 4333 6757
rect 4283 6728 4299 6749
rect 4321 6728 4333 6749
rect 2984 6555 3311 6589
rect 3391 6583 3425 6611
rect 3390 6580 3426 6583
rect 3390 6561 3398 6580
rect 3418 6561 3426 6580
rect 3390 6557 3426 6561
rect 3001 6554 3311 6555
rect 3276 6525 3311 6554
rect 3062 6518 3097 6519
rect 3041 6511 3097 6518
rect 3041 6491 3070 6511
rect 3090 6491 3097 6511
rect 3041 6486 3097 6491
rect 3271 6513 3313 6525
rect 3271 6493 3280 6513
rect 3304 6493 3313 6513
rect 3041 6280 3075 6486
rect 3271 6485 3313 6493
rect 3488 6514 3520 6521
rect 3488 6494 3494 6514
rect 3515 6494 3520 6514
rect 3488 6466 3520 6494
rect 4054 6514 4088 6720
rect 4283 6719 4333 6728
rect 4501 6748 4533 6755
rect 4501 6728 4507 6748
rect 4528 6728 4533 6748
rect 4501 6700 4533 6728
rect 4121 6692 4533 6700
rect 4121 6666 4127 6692
rect 4153 6666 4533 6692
rect 4121 6664 4533 6666
rect 4123 6663 4163 6664
rect 4501 6599 4533 6664
rect 4501 6579 4505 6599
rect 4526 6579 4533 6599
rect 4501 6572 4533 6579
rect 4054 6506 4089 6514
rect 4054 6486 4062 6506
rect 4082 6486 4089 6506
rect 4054 6481 4089 6486
rect 4054 6480 4086 6481
rect 3108 6458 3520 6466
rect 3108 6432 3114 6458
rect 3140 6432 3520 6458
rect 3108 6430 3520 6432
rect 3110 6429 3150 6430
rect 3488 6365 3520 6430
rect 3488 6345 3492 6365
rect 3513 6345 3520 6365
rect 3488 6338 3520 6345
rect 3965 6376 4317 6407
rect 3041 6272 3076 6280
rect 3041 6252 3049 6272
rect 3069 6252 3076 6272
rect 3041 6236 3076 6252
rect 3965 6236 3996 6376
rect 4289 6344 4317 6376
rect 4074 6337 4109 6338
rect 3039 6217 3996 6236
rect 4053 6330 4109 6337
rect 4053 6310 4082 6330
rect 4102 6310 4109 6330
rect 4053 6305 4109 6310
rect 4283 6332 4323 6344
rect 4283 6311 4289 6332
rect 4311 6311 4323 6332
rect 4283 6306 4323 6311
rect 4500 6333 4532 6340
rect 4500 6313 4506 6333
rect 4527 6313 4532 6333
rect 2749 6119 2786 6124
rect 2749 6113 3096 6119
rect 2749 6094 2757 6113
rect 2780 6094 3096 6113
rect 2749 6089 3096 6094
rect 2749 6083 2786 6089
rect 3066 6058 3096 6089
rect 4053 6099 4087 6305
rect 4500 6285 4532 6313
rect 4120 6277 4532 6285
rect 4120 6251 4126 6277
rect 4152 6251 4532 6277
rect 4120 6249 4532 6251
rect 4122 6248 4162 6249
rect 4500 6184 4532 6249
rect 4500 6164 4504 6184
rect 4525 6164 4532 6184
rect 4500 6157 4532 6164
rect 4053 6091 4088 6099
rect 4053 6071 4061 6091
rect 4081 6071 4088 6091
rect 4053 6066 4088 6071
rect 4053 6065 4085 6066
rect 2854 6051 2889 6052
rect 2833 6044 2889 6051
rect 2833 6024 2862 6044
rect 2882 6024 2889 6044
rect 2833 6019 2889 6024
rect 3064 6045 3103 6058
rect 3064 6026 3069 6045
rect 3092 6026 3103 6045
rect 3064 6020 3103 6026
rect 3280 6047 3312 6054
rect 3280 6027 3286 6047
rect 3307 6027 3312 6047
rect 2337 5971 2375 5977
rect 2337 5951 2347 5971
rect 2367 5951 2375 5971
rect 2337 5949 2375 5951
rect 873 5916 1288 5945
rect 2340 5943 2375 5949
rect 873 5915 1282 5916
rect 1896 5878 1928 5885
rect 1896 5858 1903 5878
rect 1924 5858 1928 5878
rect 1896 5793 1928 5858
rect 2266 5793 2306 5794
rect 1896 5791 2308 5793
rect 1896 5765 2276 5791
rect 2302 5765 2308 5791
rect 1896 5757 2308 5765
rect 1896 5729 1928 5757
rect 1896 5709 1901 5729
rect 1922 5709 1928 5729
rect 1896 5702 1928 5709
rect 2100 5734 2147 5740
rect 2341 5737 2375 5943
rect 2833 5813 2867 6019
rect 3280 5999 3312 6027
rect 2900 5991 3312 5999
rect 2900 5965 2906 5991
rect 2932 5965 3312 5991
rect 2900 5963 3312 5965
rect 2902 5962 2942 5963
rect 3280 5898 3312 5963
rect 3280 5878 3284 5898
rect 3305 5878 3312 5898
rect 3280 5871 3312 5878
rect 3926 5840 4335 5841
rect 2833 5807 2868 5813
rect 3920 5811 4335 5840
rect 2833 5805 2871 5807
rect 2833 5785 2841 5805
rect 2861 5785 2871 5805
rect 2833 5779 2871 5785
rect 2100 5708 2110 5734
rect 2135 5708 2147 5734
rect 2100 5706 2147 5708
rect 2319 5732 2375 5737
rect 2319 5712 2326 5732
rect 2346 5712 2375 5732
rect 1123 5690 1155 5691
rect 1120 5685 1155 5690
rect 1120 5665 1127 5685
rect 1147 5665 1155 5685
rect 1120 5657 1155 5665
rect 676 5592 708 5599
rect 676 5572 683 5592
rect 704 5572 708 5592
rect 676 5507 708 5572
rect 1046 5507 1086 5508
rect 676 5505 1088 5507
rect 676 5479 1056 5505
rect 1082 5479 1088 5505
rect 676 5471 1088 5479
rect 676 5443 708 5471
rect 1121 5451 1155 5657
rect 2105 5671 2142 5706
rect 2319 5705 2375 5712
rect 2319 5704 2354 5705
rect 2439 5671 2471 5673
rect 2105 5638 2475 5671
rect 676 5423 681 5443
rect 702 5423 708 5443
rect 676 5416 708 5423
rect 885 5445 925 5450
rect 885 5424 897 5445
rect 919 5424 925 5445
rect 885 5412 925 5424
rect 1099 5446 1155 5451
rect 1099 5426 1106 5446
rect 1126 5426 1155 5446
rect 1099 5419 1155 5426
rect 1212 5520 2169 5539
rect 1099 5418 1134 5419
rect 891 5380 919 5412
rect 1212 5380 1243 5520
rect 2132 5504 2167 5520
rect 2132 5484 2139 5504
rect 2159 5484 2167 5504
rect 2132 5476 2167 5484
rect 891 5349 1243 5380
rect 1688 5411 1720 5418
rect 1688 5391 1695 5411
rect 1716 5391 1720 5411
rect 1688 5326 1720 5391
rect 2058 5326 2098 5327
rect 1688 5324 2100 5326
rect 1688 5298 2068 5324
rect 2094 5298 2100 5324
rect 1688 5290 2100 5298
rect 1122 5275 1154 5276
rect 1119 5270 1154 5275
rect 1119 5250 1126 5270
rect 1146 5250 1154 5270
rect 1119 5242 1154 5250
rect 675 5177 707 5184
rect 675 5157 682 5177
rect 703 5157 707 5177
rect 675 5092 707 5157
rect 1045 5092 1085 5093
rect 675 5090 1087 5092
rect 675 5064 1055 5090
rect 1081 5064 1087 5090
rect 675 5056 1087 5064
rect 675 5028 707 5056
rect 675 5008 680 5028
rect 701 5008 707 5028
rect 675 5001 707 5008
rect 875 5028 925 5037
rect 1120 5036 1154 5242
rect 1688 5262 1720 5290
rect 1688 5242 1693 5262
rect 1714 5242 1720 5262
rect 1688 5235 1720 5242
rect 1895 5263 1937 5271
rect 2133 5270 2167 5476
rect 1895 5243 1904 5263
rect 1928 5243 1937 5263
rect 1895 5231 1937 5243
rect 2111 5265 2167 5270
rect 2111 5245 2118 5265
rect 2138 5245 2167 5265
rect 2111 5238 2167 5245
rect 2111 5237 2146 5238
rect 1897 5202 1932 5231
rect 1897 5201 2207 5202
rect 1782 5195 1818 5199
rect 1782 5176 1790 5195
rect 1810 5176 1818 5195
rect 1782 5173 1818 5176
rect 1783 5145 1817 5173
rect 1897 5167 2224 5201
rect 875 5007 887 5028
rect 909 5007 925 5028
rect 875 4999 925 5007
rect 1098 5031 1154 5036
rect 1098 5011 1105 5031
rect 1125 5011 1154 5031
rect 1098 5004 1154 5011
rect 1255 5117 1818 5145
rect 1098 5003 1133 5004
rect 880 4966 921 4999
rect 1255 4966 1295 5117
rect 880 4937 1295 4966
rect 2184 4943 2224 5167
rect 880 4936 1289 4937
rect 2184 4923 2194 4943
rect 2214 4923 2224 4943
rect 2184 4913 2224 4923
rect 1743 4850 1775 4857
rect 1743 4830 1750 4850
rect 1771 4830 1775 4850
rect 1743 4765 1775 4830
rect 2113 4765 2153 4766
rect 1743 4763 2155 4765
rect 1743 4737 2123 4763
rect 2149 4737 2155 4763
rect 1743 4729 2155 4737
rect 1128 4709 1160 4710
rect 1125 4704 1160 4709
rect 1125 4684 1132 4704
rect 1152 4684 1160 4704
rect 1125 4676 1160 4684
rect 681 4611 713 4618
rect 681 4591 688 4611
rect 709 4591 713 4611
rect 681 4526 713 4591
rect 1051 4526 1091 4527
rect 681 4524 1093 4526
rect 681 4498 1061 4524
rect 1087 4498 1093 4524
rect 681 4490 1093 4498
rect 681 4462 713 4490
rect 1126 4470 1160 4676
rect 1743 4701 1775 4729
rect 2188 4709 2222 4913
rect 1743 4681 1748 4701
rect 1769 4681 1775 4701
rect 1743 4674 1775 4681
rect 1954 4701 1991 4707
rect 1954 4682 1960 4701
rect 1983 4682 1991 4701
rect 1954 4677 1991 4682
rect 2166 4704 2222 4709
rect 2166 4684 2173 4704
rect 2193 4684 2222 4704
rect 2166 4677 2222 4684
rect 1962 4640 1986 4677
rect 2166 4676 2201 4677
rect 1962 4638 2330 4640
rect 1962 4633 2335 4638
rect 1962 4615 2308 4633
rect 2328 4615 2335 4633
rect 1962 4610 2335 4615
rect 2306 4608 2335 4610
rect 681 4442 686 4462
rect 707 4442 713 4462
rect 681 4435 713 4442
rect 890 4464 930 4469
rect 890 4443 902 4464
rect 924 4443 930 4464
rect 890 4431 930 4443
rect 1104 4465 1160 4470
rect 1104 4445 1111 4465
rect 1131 4445 1160 4465
rect 1104 4438 1160 4445
rect 1217 4539 2174 4558
rect 1104 4437 1139 4438
rect 896 4399 924 4431
rect 1217 4399 1248 4539
rect 2137 4523 2172 4539
rect 2137 4503 2144 4523
rect 2164 4503 2172 4523
rect 2137 4495 2172 4503
rect 896 4368 1248 4399
rect 1693 4430 1725 4437
rect 1693 4410 1700 4430
rect 1721 4410 1725 4430
rect 1693 4345 1725 4410
rect 2063 4345 2103 4346
rect 1693 4343 2105 4345
rect 1693 4317 2073 4343
rect 2099 4317 2105 4343
rect 1693 4309 2105 4317
rect 1127 4294 1159 4295
rect 1124 4289 1159 4294
rect 1124 4269 1131 4289
rect 1151 4269 1159 4289
rect 1124 4261 1159 4269
rect 680 4196 712 4203
rect 680 4176 687 4196
rect 708 4176 712 4196
rect 680 4111 712 4176
rect 1050 4111 1090 4112
rect 680 4109 1092 4111
rect 680 4083 1060 4109
rect 1086 4083 1092 4109
rect 680 4075 1092 4083
rect 680 4047 712 4075
rect 680 4027 685 4047
rect 706 4027 712 4047
rect 680 4020 712 4027
rect 880 4047 930 4056
rect 1125 4055 1159 4261
rect 1693 4281 1725 4309
rect 1693 4261 1698 4281
rect 1719 4261 1725 4281
rect 1898 4283 1940 4292
rect 2138 4289 2172 4495
rect 1898 4269 1908 4283
rect 1693 4254 1725 4261
rect 1897 4263 1908 4269
rect 1932 4263 1940 4283
rect 1897 4252 1940 4263
rect 2116 4284 2172 4289
rect 2116 4264 2123 4284
rect 2143 4264 2172 4284
rect 2116 4257 2172 4264
rect 2116 4256 2151 4257
rect 1897 4222 1937 4252
rect 1787 4214 1823 4218
rect 1787 4195 1795 4214
rect 1815 4195 1823 4214
rect 1787 4192 1823 4195
rect 1897 4217 2244 4222
rect 1788 4164 1822 4192
rect 1897 4191 2216 4217
rect 2235 4191 2244 4217
rect 1897 4187 2244 4191
rect 880 4026 892 4047
rect 914 4026 930 4047
rect 880 4018 930 4026
rect 1103 4050 1159 4055
rect 1103 4030 1110 4050
rect 1130 4030 1159 4050
rect 1103 4023 1159 4030
rect 1260 4136 1823 4164
rect 1103 4022 1138 4023
rect 885 3985 926 4018
rect 1260 3985 1300 4136
rect 2439 3985 2471 5638
rect 2836 5185 2871 5779
rect 3920 5660 3960 5811
rect 4294 5778 4335 5811
rect 4082 5773 4117 5774
rect 3397 5632 3960 5660
rect 4061 5766 4117 5773
rect 4061 5746 4090 5766
rect 4110 5746 4117 5766
rect 4061 5741 4117 5746
rect 4290 5770 4340 5778
rect 4290 5749 4306 5770
rect 4328 5749 4340 5770
rect 2976 5605 3323 5609
rect 2976 5579 2985 5605
rect 3004 5579 3323 5605
rect 3398 5604 3432 5632
rect 2976 5574 3323 5579
rect 3397 5601 3433 5604
rect 3397 5582 3405 5601
rect 3425 5582 3433 5601
rect 3397 5578 3433 5582
rect 3283 5544 3323 5574
rect 3069 5539 3104 5540
rect 3048 5532 3104 5539
rect 3048 5512 3077 5532
rect 3097 5512 3104 5532
rect 3048 5507 3104 5512
rect 3280 5533 3323 5544
rect 3280 5513 3288 5533
rect 3312 5527 3323 5533
rect 3495 5535 3527 5542
rect 3312 5513 3322 5527
rect 3048 5301 3082 5507
rect 3280 5504 3322 5513
rect 3495 5515 3501 5535
rect 3522 5515 3527 5535
rect 3495 5487 3527 5515
rect 4061 5535 4095 5741
rect 4290 5740 4340 5749
rect 4508 5769 4540 5776
rect 4508 5749 4514 5769
rect 4535 5749 4540 5769
rect 4508 5721 4540 5749
rect 4128 5713 4540 5721
rect 4128 5687 4134 5713
rect 4160 5687 4540 5713
rect 4128 5685 4540 5687
rect 4130 5684 4170 5685
rect 4508 5620 4540 5685
rect 4508 5600 4512 5620
rect 4533 5600 4540 5620
rect 4508 5593 4540 5600
rect 4061 5527 4096 5535
rect 4061 5507 4069 5527
rect 4089 5507 4096 5527
rect 4061 5502 4096 5507
rect 4061 5501 4093 5502
rect 3115 5479 3527 5487
rect 3115 5453 3121 5479
rect 3147 5453 3527 5479
rect 3115 5451 3527 5453
rect 3117 5450 3157 5451
rect 3495 5386 3527 5451
rect 3495 5366 3499 5386
rect 3520 5366 3527 5386
rect 3495 5359 3527 5366
rect 3972 5397 4324 5428
rect 3048 5293 3083 5301
rect 3048 5273 3056 5293
rect 3076 5273 3083 5293
rect 3048 5257 3083 5273
rect 3972 5257 4003 5397
rect 4296 5365 4324 5397
rect 4081 5358 4116 5359
rect 3046 5238 4003 5257
rect 4060 5351 4116 5358
rect 4060 5331 4089 5351
rect 4109 5331 4116 5351
rect 4060 5326 4116 5331
rect 4290 5353 4330 5365
rect 4290 5332 4296 5353
rect 4318 5332 4330 5353
rect 4290 5327 4330 5332
rect 4507 5354 4539 5361
rect 4507 5334 4513 5354
rect 4534 5334 4539 5354
rect 2836 5156 3266 5185
rect 2836 5151 2920 5156
rect 3019 5119 3054 5120
rect 2998 5112 3054 5119
rect 2998 5092 3027 5112
rect 3047 5092 3054 5112
rect 2998 5087 3054 5092
rect 3228 5113 3266 5156
rect 3228 5096 3233 5113
rect 3257 5096 3266 5113
rect 2998 4883 3032 5087
rect 3228 5084 3266 5096
rect 3445 5115 3477 5122
rect 3445 5095 3451 5115
rect 3472 5095 3477 5115
rect 3445 5067 3477 5095
rect 4060 5120 4094 5326
rect 4507 5306 4539 5334
rect 4127 5298 4539 5306
rect 4127 5272 4133 5298
rect 4159 5272 4539 5298
rect 4127 5270 4539 5272
rect 4129 5269 4169 5270
rect 4507 5205 4539 5270
rect 4507 5185 4511 5205
rect 4532 5185 4539 5205
rect 4507 5178 4539 5185
rect 4060 5112 4095 5120
rect 4060 5092 4068 5112
rect 4088 5092 4095 5112
rect 4060 5087 4095 5092
rect 4060 5086 4092 5087
rect 3065 5059 3477 5067
rect 3065 5033 3071 5059
rect 3097 5033 3477 5059
rect 3065 5031 3477 5033
rect 3067 5030 3107 5031
rect 3445 4966 3477 5031
rect 3445 4946 3449 4966
rect 3470 4946 3477 4966
rect 3445 4939 3477 4946
rect 2996 4873 3036 4883
rect 2996 4853 3006 4873
rect 3026 4853 3036 4873
rect 3931 4859 4340 4860
rect 2996 4629 3036 4853
rect 3925 4830 4340 4859
rect 3925 4679 3965 4830
rect 4299 4797 4340 4830
rect 4087 4792 4122 4793
rect 3402 4651 3965 4679
rect 4066 4785 4122 4792
rect 4066 4765 4095 4785
rect 4115 4765 4122 4785
rect 4066 4760 4122 4765
rect 4295 4789 4345 4797
rect 4295 4768 4311 4789
rect 4333 4768 4345 4789
rect 2996 4595 3323 4629
rect 3403 4623 3437 4651
rect 3402 4620 3438 4623
rect 3402 4601 3410 4620
rect 3430 4601 3438 4620
rect 3402 4597 3438 4601
rect 3013 4594 3323 4595
rect 3288 4565 3323 4594
rect 3074 4558 3109 4559
rect 3053 4551 3109 4558
rect 3053 4531 3082 4551
rect 3102 4531 3109 4551
rect 3053 4526 3109 4531
rect 3283 4553 3325 4565
rect 3283 4533 3292 4553
rect 3316 4533 3325 4553
rect 3053 4320 3087 4526
rect 3283 4525 3325 4533
rect 3500 4554 3532 4561
rect 3500 4534 3506 4554
rect 3527 4534 3532 4554
rect 3500 4506 3532 4534
rect 4066 4554 4100 4760
rect 4295 4759 4345 4768
rect 4513 4788 4545 4795
rect 4513 4768 4519 4788
rect 4540 4768 4545 4788
rect 4513 4740 4545 4768
rect 4133 4732 4545 4740
rect 4133 4706 4139 4732
rect 4165 4706 4545 4732
rect 4133 4704 4545 4706
rect 4135 4703 4175 4704
rect 4513 4639 4545 4704
rect 4513 4619 4517 4639
rect 4538 4619 4545 4639
rect 4513 4612 4545 4619
rect 4066 4546 4101 4554
rect 4066 4526 4074 4546
rect 4094 4526 4101 4546
rect 4066 4521 4101 4526
rect 4066 4520 4098 4521
rect 3120 4498 3532 4506
rect 3120 4472 3126 4498
rect 3152 4472 3532 4498
rect 3120 4470 3532 4472
rect 3122 4469 3162 4470
rect 3500 4405 3532 4470
rect 3500 4385 3504 4405
rect 3525 4385 3532 4405
rect 3500 4378 3532 4385
rect 3977 4416 4329 4447
rect 3053 4312 3088 4320
rect 3053 4292 3061 4312
rect 3081 4292 3088 4312
rect 3053 4276 3088 4292
rect 3977 4276 4008 4416
rect 4301 4384 4329 4416
rect 4086 4377 4121 4378
rect 3051 4257 4008 4276
rect 4065 4370 4121 4377
rect 4065 4350 4094 4370
rect 4114 4350 4121 4370
rect 4065 4345 4121 4350
rect 4295 4372 4335 4384
rect 4295 4351 4301 4372
rect 4323 4351 4335 4372
rect 4295 4346 4335 4351
rect 4512 4373 4544 4380
rect 4512 4353 4518 4373
rect 4539 4353 4544 4373
rect 2649 4200 2734 4203
rect 2642 4196 2734 4200
rect 2642 4195 3023 4196
rect 2642 4165 2649 4195
rect 2686 4166 3023 4195
rect 2686 4165 2734 4166
rect 2642 4163 2734 4165
rect 2642 4160 2727 4163
rect 2988 4128 3023 4166
rect 4065 4139 4099 4345
rect 4512 4325 4544 4353
rect 4132 4317 4544 4325
rect 4132 4291 4138 4317
rect 4164 4291 4544 4317
rect 4132 4289 4544 4291
rect 4134 4288 4174 4289
rect 4512 4224 4544 4289
rect 4512 4204 4516 4224
rect 4537 4204 4544 4224
rect 4512 4197 4544 4204
rect 4065 4131 4100 4139
rect 2779 4126 2814 4127
rect 885 3956 1300 3985
rect 2438 3984 2471 3985
rect 2435 3979 2471 3984
rect 2435 3959 2442 3979
rect 2462 3959 2471 3979
rect 885 3955 1294 3956
rect 2435 3954 2471 3959
rect 2758 4119 2814 4126
rect 2758 4099 2787 4119
rect 2807 4099 2814 4119
rect 2758 4094 2814 4099
rect 2983 4119 3032 4128
rect 2983 4100 2991 4119
rect 3017 4100 3032 4119
rect 2435 3951 2470 3954
rect 1991 3886 2023 3893
rect 1991 3866 1998 3886
rect 2019 3866 2023 3886
rect 1991 3801 2023 3866
rect 2361 3801 2401 3802
rect 1991 3799 2403 3801
rect 1991 3773 2371 3799
rect 2397 3773 2403 3799
rect 1991 3765 2403 3773
rect 1991 3737 2023 3765
rect 1131 3733 1163 3734
rect 1128 3728 1163 3733
rect 1128 3708 1135 3728
rect 1155 3708 1163 3728
rect 1991 3717 1996 3737
rect 2017 3717 2023 3737
rect 1991 3710 2023 3717
rect 2196 3739 2245 3749
rect 2436 3745 2470 3951
rect 2758 3888 2792 4094
rect 2983 4090 3032 4100
rect 3205 4122 3237 4129
rect 3205 4102 3211 4122
rect 3232 4102 3237 4122
rect 4065 4111 4073 4131
rect 4093 4111 4100 4131
rect 4065 4106 4100 4111
rect 4065 4105 4097 4106
rect 3205 4074 3237 4102
rect 2825 4066 3237 4074
rect 2825 4040 2831 4066
rect 2857 4040 3237 4066
rect 2825 4038 3237 4040
rect 2827 4037 2867 4038
rect 3205 3973 3237 4038
rect 3205 3953 3209 3973
rect 3230 3953 3237 3973
rect 3205 3946 3237 3953
rect 2758 3885 2793 3888
rect 2196 3720 2211 3739
rect 2237 3720 2245 3739
rect 2196 3711 2245 3720
rect 2414 3740 2470 3745
rect 2414 3720 2421 3740
rect 2441 3720 2470 3740
rect 2414 3713 2470 3720
rect 2757 3880 2793 3885
rect 3934 3883 4343 3884
rect 2757 3860 2766 3880
rect 2786 3860 2793 3880
rect 2757 3855 2793 3860
rect 2757 3854 2790 3855
rect 3928 3854 4343 3883
rect 2414 3712 2449 3713
rect 1128 3700 1163 3708
rect 684 3635 716 3642
rect 684 3615 691 3635
rect 712 3615 716 3635
rect 684 3550 716 3615
rect 1054 3550 1094 3551
rect 684 3548 1096 3550
rect 684 3522 1064 3548
rect 1090 3522 1096 3548
rect 684 3514 1096 3522
rect 684 3486 716 3514
rect 1129 3494 1163 3700
rect 2205 3673 2240 3711
rect 2463 3673 2586 3678
rect 2205 3672 2586 3673
rect 2205 3644 2548 3672
rect 2582 3671 2586 3672
rect 2582 3644 2587 3671
rect 2205 3643 2587 3644
rect 2463 3638 2587 3643
rect 684 3466 689 3486
rect 710 3466 716 3486
rect 684 3459 716 3466
rect 893 3488 933 3493
rect 893 3467 905 3488
rect 927 3467 933 3488
rect 893 3455 933 3467
rect 1107 3489 1163 3494
rect 1107 3469 1114 3489
rect 1134 3469 1163 3489
rect 1107 3462 1163 3469
rect 1220 3563 2177 3582
rect 1107 3461 1142 3462
rect 899 3423 927 3455
rect 1220 3423 1251 3563
rect 2140 3547 2175 3563
rect 2140 3527 2147 3547
rect 2167 3527 2175 3547
rect 2140 3519 2175 3527
rect 899 3392 1251 3423
rect 1696 3454 1728 3461
rect 1696 3434 1703 3454
rect 1724 3434 1728 3454
rect 1696 3369 1728 3434
rect 2066 3369 2106 3370
rect 1696 3367 2108 3369
rect 1696 3341 2076 3367
rect 2102 3341 2108 3367
rect 1696 3333 2108 3341
rect 1130 3318 1162 3319
rect 1127 3313 1162 3318
rect 1127 3293 1134 3313
rect 1154 3293 1162 3313
rect 1127 3285 1162 3293
rect 683 3220 715 3227
rect 683 3200 690 3220
rect 711 3200 715 3220
rect 683 3135 715 3200
rect 1053 3135 1093 3136
rect 683 3133 1095 3135
rect 683 3107 1063 3133
rect 1089 3107 1095 3133
rect 683 3099 1095 3107
rect 683 3071 715 3099
rect 683 3051 688 3071
rect 709 3051 715 3071
rect 683 3044 715 3051
rect 883 3071 933 3080
rect 1128 3079 1162 3285
rect 1696 3305 1728 3333
rect 1696 3285 1701 3305
rect 1722 3285 1728 3305
rect 1696 3278 1728 3285
rect 1903 3306 1945 3314
rect 2141 3313 2175 3519
rect 1903 3286 1912 3306
rect 1936 3286 1945 3306
rect 1903 3274 1945 3286
rect 2119 3308 2175 3313
rect 2119 3288 2126 3308
rect 2146 3288 2175 3308
rect 2119 3281 2175 3288
rect 2119 3280 2154 3281
rect 1905 3245 1940 3274
rect 1905 3244 2215 3245
rect 1790 3238 1826 3242
rect 1790 3219 1798 3238
rect 1818 3219 1826 3238
rect 1790 3216 1826 3219
rect 1791 3188 1825 3216
rect 1905 3210 2232 3244
rect 883 3050 895 3071
rect 917 3050 933 3071
rect 883 3042 933 3050
rect 1106 3074 1162 3079
rect 1106 3054 1113 3074
rect 1133 3054 1162 3074
rect 1106 3047 1162 3054
rect 1263 3160 1826 3188
rect 1106 3046 1141 3047
rect 888 3009 929 3042
rect 1263 3009 1303 3160
rect 888 2980 1303 3009
rect 2192 2986 2232 3210
rect 888 2979 1297 2980
rect 2192 2966 2202 2986
rect 2222 2966 2232 2986
rect 2192 2956 2232 2966
rect 1751 2893 1783 2900
rect 1751 2873 1758 2893
rect 1779 2873 1783 2893
rect 1751 2808 1783 2873
rect 2121 2808 2161 2809
rect 1751 2806 2163 2808
rect 1751 2780 2131 2806
rect 2157 2780 2163 2806
rect 1751 2772 2163 2780
rect 1136 2752 1168 2753
rect 1133 2747 1168 2752
rect 1133 2727 1140 2747
rect 1160 2727 1168 2747
rect 1133 2719 1168 2727
rect 689 2654 721 2661
rect 689 2634 696 2654
rect 717 2634 721 2654
rect 689 2569 721 2634
rect 1059 2569 1099 2570
rect 689 2567 1101 2569
rect 689 2541 1069 2567
rect 1095 2541 1101 2567
rect 689 2533 1101 2541
rect 689 2505 721 2533
rect 1134 2513 1168 2719
rect 1751 2744 1783 2772
rect 1751 2724 1756 2744
rect 1777 2724 1783 2744
rect 1751 2717 1783 2724
rect 1962 2743 2000 2755
rect 2196 2752 2230 2956
rect 1962 2726 1971 2743
rect 1995 2726 2000 2743
rect 1962 2683 2000 2726
rect 2174 2747 2230 2752
rect 2174 2727 2181 2747
rect 2201 2727 2230 2747
rect 2174 2720 2230 2727
rect 2174 2719 2209 2720
rect 2308 2683 2392 2688
rect 1962 2654 2392 2683
rect 689 2485 694 2505
rect 715 2485 721 2505
rect 689 2478 721 2485
rect 898 2507 938 2512
rect 898 2486 910 2507
rect 932 2486 938 2507
rect 898 2474 938 2486
rect 1112 2508 1168 2513
rect 1112 2488 1119 2508
rect 1139 2488 1168 2508
rect 1112 2481 1168 2488
rect 1225 2582 2182 2601
rect 1112 2480 1147 2481
rect 904 2442 932 2474
rect 1225 2442 1256 2582
rect 2145 2566 2180 2582
rect 2145 2546 2152 2566
rect 2172 2546 2180 2566
rect 2145 2538 2180 2546
rect 904 2411 1256 2442
rect 1701 2473 1733 2480
rect 1701 2453 1708 2473
rect 1729 2453 1733 2473
rect 1701 2388 1733 2453
rect 2071 2388 2111 2389
rect 1701 2386 2113 2388
rect 1701 2360 2081 2386
rect 2107 2360 2113 2386
rect 1701 2352 2113 2360
rect 1135 2337 1167 2338
rect 1132 2332 1167 2337
rect 1132 2312 1139 2332
rect 1159 2312 1167 2332
rect 1132 2304 1167 2312
rect 688 2239 720 2246
rect 688 2219 695 2239
rect 716 2219 720 2239
rect 688 2154 720 2219
rect 1058 2154 1098 2155
rect 688 2152 1100 2154
rect 688 2126 1068 2152
rect 1094 2126 1100 2152
rect 688 2118 1100 2126
rect 688 2090 720 2118
rect 688 2070 693 2090
rect 714 2070 720 2090
rect 688 2063 720 2070
rect 888 2090 938 2099
rect 1133 2098 1167 2304
rect 1701 2324 1733 2352
rect 1701 2304 1706 2324
rect 1727 2304 1733 2324
rect 1906 2326 1948 2335
rect 2146 2332 2180 2538
rect 1906 2312 1916 2326
rect 1701 2297 1733 2304
rect 1905 2306 1916 2312
rect 1940 2306 1948 2326
rect 1905 2295 1948 2306
rect 2124 2327 2180 2332
rect 2124 2307 2131 2327
rect 2151 2307 2180 2327
rect 2124 2300 2180 2307
rect 2124 2299 2159 2300
rect 1905 2265 1945 2295
rect 1795 2257 1831 2261
rect 1795 2238 1803 2257
rect 1823 2238 1831 2257
rect 1795 2235 1831 2238
rect 1905 2260 2252 2265
rect 1796 2207 1830 2235
rect 1905 2234 2224 2260
rect 2243 2234 2252 2260
rect 1905 2230 2252 2234
rect 888 2069 900 2090
rect 922 2069 938 2090
rect 888 2061 938 2069
rect 1111 2093 1167 2098
rect 1111 2073 1118 2093
rect 1138 2073 1167 2093
rect 1111 2066 1167 2073
rect 1268 2179 1831 2207
rect 1111 2065 1146 2066
rect 893 2028 934 2061
rect 1268 2028 1308 2179
rect 2357 2060 2392 2654
rect 2757 2201 2789 3854
rect 3928 3703 3968 3854
rect 4302 3821 4343 3854
rect 4090 3816 4125 3817
rect 3405 3675 3968 3703
rect 4069 3809 4125 3816
rect 4069 3789 4098 3809
rect 4118 3789 4125 3809
rect 4069 3784 4125 3789
rect 4298 3813 4348 3821
rect 4298 3792 4314 3813
rect 4336 3792 4348 3813
rect 2984 3648 3331 3652
rect 2984 3622 2993 3648
rect 3012 3622 3331 3648
rect 3406 3647 3440 3675
rect 2984 3617 3331 3622
rect 3405 3644 3441 3647
rect 3405 3625 3413 3644
rect 3433 3625 3441 3644
rect 3405 3621 3441 3625
rect 3291 3587 3331 3617
rect 3077 3582 3112 3583
rect 3056 3575 3112 3582
rect 3056 3555 3085 3575
rect 3105 3555 3112 3575
rect 3056 3550 3112 3555
rect 3288 3576 3331 3587
rect 3288 3556 3296 3576
rect 3320 3570 3331 3576
rect 3503 3578 3535 3585
rect 3320 3556 3330 3570
rect 3056 3344 3090 3550
rect 3288 3547 3330 3556
rect 3503 3558 3509 3578
rect 3530 3558 3535 3578
rect 3503 3530 3535 3558
rect 4069 3578 4103 3784
rect 4298 3783 4348 3792
rect 4516 3812 4548 3819
rect 4516 3792 4522 3812
rect 4543 3792 4548 3812
rect 4516 3764 4548 3792
rect 4136 3756 4548 3764
rect 4136 3730 4142 3756
rect 4168 3730 4548 3756
rect 4136 3728 4548 3730
rect 4138 3727 4178 3728
rect 4516 3663 4548 3728
rect 4516 3643 4520 3663
rect 4541 3643 4548 3663
rect 4516 3636 4548 3643
rect 4069 3570 4104 3578
rect 4069 3550 4077 3570
rect 4097 3550 4104 3570
rect 4069 3545 4104 3550
rect 4069 3544 4101 3545
rect 3123 3522 3535 3530
rect 3123 3496 3129 3522
rect 3155 3496 3535 3522
rect 3123 3494 3535 3496
rect 3125 3493 3165 3494
rect 3503 3429 3535 3494
rect 3503 3409 3507 3429
rect 3528 3409 3535 3429
rect 3503 3402 3535 3409
rect 3980 3440 4332 3471
rect 3056 3336 3091 3344
rect 3056 3316 3064 3336
rect 3084 3316 3091 3336
rect 3056 3300 3091 3316
rect 3980 3300 4011 3440
rect 4304 3408 4332 3440
rect 4089 3401 4124 3402
rect 3054 3281 4011 3300
rect 4068 3394 4124 3401
rect 4068 3374 4097 3394
rect 4117 3374 4124 3394
rect 4068 3369 4124 3374
rect 4298 3396 4338 3408
rect 4298 3375 4304 3396
rect 4326 3375 4338 3396
rect 4298 3370 4338 3375
rect 4515 3397 4547 3404
rect 4515 3377 4521 3397
rect 4542 3377 4547 3397
rect 2893 3229 2922 3231
rect 2893 3224 3266 3229
rect 2893 3206 2900 3224
rect 2920 3206 3266 3224
rect 2893 3201 3266 3206
rect 2898 3199 3266 3201
rect 3027 3162 3062 3163
rect 3242 3162 3266 3199
rect 3006 3155 3062 3162
rect 3006 3135 3035 3155
rect 3055 3135 3062 3155
rect 3006 3130 3062 3135
rect 3237 3157 3274 3162
rect 3237 3138 3245 3157
rect 3268 3138 3274 3157
rect 3237 3132 3274 3138
rect 3453 3158 3485 3165
rect 3453 3138 3459 3158
rect 3480 3138 3485 3158
rect 3006 2926 3040 3130
rect 3453 3110 3485 3138
rect 4068 3163 4102 3369
rect 4515 3349 4547 3377
rect 4135 3341 4547 3349
rect 4135 3315 4141 3341
rect 4167 3315 4547 3341
rect 4135 3313 4547 3315
rect 4137 3312 4177 3313
rect 4515 3248 4547 3313
rect 4515 3228 4519 3248
rect 4540 3228 4547 3248
rect 4515 3221 4547 3228
rect 4068 3155 4103 3163
rect 4068 3135 4076 3155
rect 4096 3135 4103 3155
rect 4068 3130 4103 3135
rect 4068 3129 4100 3130
rect 3073 3102 3485 3110
rect 3073 3076 3079 3102
rect 3105 3076 3485 3102
rect 3073 3074 3485 3076
rect 3075 3073 3115 3074
rect 3453 3009 3485 3074
rect 3453 2989 3457 3009
rect 3478 2989 3485 3009
rect 3453 2982 3485 2989
rect 3004 2916 3044 2926
rect 3004 2896 3014 2916
rect 3034 2896 3044 2916
rect 3939 2902 4348 2903
rect 3004 2672 3044 2896
rect 3933 2873 4348 2902
rect 3933 2722 3973 2873
rect 4307 2840 4348 2873
rect 4095 2835 4130 2836
rect 3410 2694 3973 2722
rect 4074 2828 4130 2835
rect 4074 2808 4103 2828
rect 4123 2808 4130 2828
rect 4074 2803 4130 2808
rect 4303 2832 4353 2840
rect 4303 2811 4319 2832
rect 4341 2811 4353 2832
rect 3004 2638 3331 2672
rect 3411 2666 3445 2694
rect 3410 2663 3446 2666
rect 3410 2644 3418 2663
rect 3438 2644 3446 2663
rect 3410 2640 3446 2644
rect 3021 2637 3331 2638
rect 3296 2608 3331 2637
rect 3082 2601 3117 2602
rect 3061 2594 3117 2601
rect 3061 2574 3090 2594
rect 3110 2574 3117 2594
rect 3061 2569 3117 2574
rect 3291 2596 3333 2608
rect 3291 2576 3300 2596
rect 3324 2576 3333 2596
rect 3061 2363 3095 2569
rect 3291 2568 3333 2576
rect 3508 2597 3540 2604
rect 3508 2577 3514 2597
rect 3535 2577 3540 2597
rect 3508 2549 3540 2577
rect 4074 2597 4108 2803
rect 4303 2802 4353 2811
rect 4521 2831 4553 2838
rect 4521 2811 4527 2831
rect 4548 2811 4553 2831
rect 4521 2783 4553 2811
rect 4141 2775 4553 2783
rect 4141 2749 4147 2775
rect 4173 2749 4553 2775
rect 4141 2747 4553 2749
rect 4143 2746 4183 2747
rect 4521 2682 4553 2747
rect 4521 2662 4525 2682
rect 4546 2662 4553 2682
rect 4521 2655 4553 2662
rect 4074 2589 4109 2597
rect 4074 2569 4082 2589
rect 4102 2569 4109 2589
rect 4074 2564 4109 2569
rect 4074 2563 4106 2564
rect 3128 2541 3540 2549
rect 3128 2515 3134 2541
rect 3160 2515 3540 2541
rect 3128 2513 3540 2515
rect 3130 2512 3170 2513
rect 3508 2448 3540 2513
rect 3508 2428 3512 2448
rect 3533 2428 3540 2448
rect 3508 2421 3540 2428
rect 3985 2459 4337 2490
rect 3061 2355 3096 2363
rect 3061 2335 3069 2355
rect 3089 2335 3096 2355
rect 3061 2319 3096 2335
rect 3985 2319 4016 2459
rect 4309 2427 4337 2459
rect 4094 2420 4129 2421
rect 3059 2300 4016 2319
rect 4073 2413 4129 2420
rect 4073 2393 4102 2413
rect 4122 2393 4129 2413
rect 4073 2388 4129 2393
rect 4303 2415 4343 2427
rect 4303 2394 4309 2415
rect 4331 2394 4343 2415
rect 4303 2389 4343 2394
rect 4520 2416 4552 2423
rect 4520 2396 4526 2416
rect 4547 2396 4552 2416
rect 2753 2168 3123 2201
rect 2757 2166 2789 2168
rect 2874 2134 2909 2135
rect 2853 2127 2909 2134
rect 3086 2133 3123 2168
rect 4073 2182 4107 2388
rect 4520 2368 4552 2396
rect 4140 2360 4552 2368
rect 4140 2334 4146 2360
rect 4172 2334 4552 2360
rect 4140 2332 4552 2334
rect 4142 2331 4182 2332
rect 4520 2267 4552 2332
rect 4520 2247 4524 2267
rect 4545 2247 4552 2267
rect 4520 2240 4552 2247
rect 4073 2174 4108 2182
rect 4073 2154 4081 2174
rect 4101 2154 4108 2174
rect 4073 2149 4108 2154
rect 4073 2148 4105 2149
rect 2853 2107 2882 2127
rect 2902 2107 2909 2127
rect 2853 2102 2909 2107
rect 3081 2131 3128 2133
rect 3081 2105 3093 2131
rect 3118 2105 3128 2131
rect 2357 2054 2395 2060
rect 2357 2034 2367 2054
rect 2387 2034 2395 2054
rect 2357 2032 2395 2034
rect 893 1999 1308 2028
rect 2360 2026 2395 2032
rect 893 1998 1302 1999
rect 1916 1961 1948 1968
rect 1916 1941 1923 1961
rect 1944 1941 1948 1961
rect 1916 1876 1948 1941
rect 2286 1876 2326 1877
rect 1916 1874 2328 1876
rect 1916 1848 2296 1874
rect 2322 1848 2328 1874
rect 1916 1840 2328 1848
rect 1916 1812 1948 1840
rect 2361 1820 2395 2026
rect 2853 1896 2887 2102
rect 3081 2099 3128 2105
rect 3300 2130 3332 2137
rect 3300 2110 3306 2130
rect 3327 2110 3332 2130
rect 3300 2082 3332 2110
rect 2920 2074 3332 2082
rect 2920 2048 2926 2074
rect 2952 2048 3332 2074
rect 2920 2046 3332 2048
rect 2922 2045 2962 2046
rect 3300 1981 3332 2046
rect 3300 1961 3304 1981
rect 3325 1961 3332 1981
rect 3300 1954 3332 1961
rect 3946 1923 4355 1924
rect 2853 1890 2888 1896
rect 3940 1894 4355 1923
rect 2853 1888 2891 1890
rect 2853 1868 2861 1888
rect 2881 1868 2891 1888
rect 2853 1862 2891 1868
rect 1916 1792 1921 1812
rect 1942 1792 1948 1812
rect 1916 1785 1948 1792
rect 2125 1813 2164 1819
rect 2125 1794 2136 1813
rect 2159 1794 2164 1813
rect 2125 1781 2164 1794
rect 2339 1815 2395 1820
rect 2339 1795 2346 1815
rect 2366 1795 2395 1815
rect 2339 1788 2395 1795
rect 2339 1787 2374 1788
rect 1143 1773 1175 1774
rect 1140 1768 1175 1773
rect 1140 1748 1147 1768
rect 1167 1748 1175 1768
rect 1140 1740 1175 1748
rect 696 1675 728 1682
rect 696 1655 703 1675
rect 724 1655 728 1675
rect 696 1590 728 1655
rect 1066 1590 1106 1591
rect 696 1588 1108 1590
rect 696 1562 1076 1588
rect 1102 1562 1108 1588
rect 696 1554 1108 1562
rect 696 1526 728 1554
rect 1141 1534 1175 1740
rect 2132 1750 2162 1781
rect 2442 1750 2479 1756
rect 2132 1745 2479 1750
rect 2132 1726 2448 1745
rect 2471 1726 2479 1745
rect 2132 1720 2479 1726
rect 2442 1715 2479 1720
rect 696 1506 701 1526
rect 722 1506 728 1526
rect 696 1499 728 1506
rect 905 1528 945 1533
rect 905 1507 917 1528
rect 939 1507 945 1528
rect 905 1495 945 1507
rect 1119 1529 1175 1534
rect 1119 1509 1126 1529
rect 1146 1509 1175 1529
rect 1119 1502 1175 1509
rect 1232 1603 2189 1622
rect 1119 1501 1154 1502
rect 911 1463 939 1495
rect 1232 1463 1263 1603
rect 2152 1587 2187 1603
rect 2152 1567 2159 1587
rect 2179 1567 2187 1587
rect 2152 1559 2187 1567
rect 911 1432 1263 1463
rect 1708 1494 1740 1501
rect 1708 1474 1715 1494
rect 1736 1474 1740 1494
rect 1708 1409 1740 1474
rect 2078 1409 2118 1410
rect 1708 1407 2120 1409
rect 1708 1381 2088 1407
rect 2114 1381 2120 1407
rect 1708 1373 2120 1381
rect 1142 1358 1174 1359
rect 1139 1353 1174 1358
rect 1139 1333 1146 1353
rect 1166 1333 1174 1353
rect 1139 1325 1174 1333
rect 695 1260 727 1267
rect 695 1240 702 1260
rect 723 1240 727 1260
rect 695 1175 727 1240
rect 1065 1175 1105 1176
rect 695 1173 1107 1175
rect 695 1147 1075 1173
rect 1101 1147 1107 1173
rect 695 1139 1107 1147
rect 695 1111 727 1139
rect 695 1091 700 1111
rect 721 1091 727 1111
rect 695 1084 727 1091
rect 895 1111 945 1120
rect 1140 1119 1174 1325
rect 1708 1345 1740 1373
rect 1708 1325 1713 1345
rect 1734 1325 1740 1345
rect 1708 1318 1740 1325
rect 1915 1346 1957 1354
rect 2153 1353 2187 1559
rect 1915 1326 1924 1346
rect 1948 1326 1957 1346
rect 1915 1314 1957 1326
rect 2131 1348 2187 1353
rect 2131 1328 2138 1348
rect 2158 1328 2187 1348
rect 2131 1321 2187 1328
rect 2131 1320 2166 1321
rect 1917 1285 1952 1314
rect 1917 1284 2227 1285
rect 1802 1278 1838 1282
rect 1802 1259 1810 1278
rect 1830 1259 1838 1278
rect 1802 1256 1838 1259
rect 1803 1228 1837 1256
rect 1917 1250 2244 1284
rect 895 1090 907 1111
rect 929 1090 945 1111
rect 895 1082 945 1090
rect 1118 1114 1174 1119
rect 1118 1094 1125 1114
rect 1145 1094 1174 1114
rect 1118 1087 1174 1094
rect 1275 1200 1838 1228
rect 1118 1086 1153 1087
rect 900 1049 941 1082
rect 1275 1049 1315 1200
rect 900 1020 1315 1049
rect 2204 1026 2244 1250
rect 2856 1268 2891 1862
rect 3940 1743 3980 1894
rect 4314 1861 4355 1894
rect 4102 1856 4137 1857
rect 3417 1715 3980 1743
rect 4081 1849 4137 1856
rect 4081 1829 4110 1849
rect 4130 1829 4137 1849
rect 4081 1824 4137 1829
rect 4310 1853 4360 1861
rect 4310 1832 4326 1853
rect 4348 1832 4360 1853
rect 2996 1688 3343 1692
rect 2996 1662 3005 1688
rect 3024 1662 3343 1688
rect 3418 1687 3452 1715
rect 2996 1657 3343 1662
rect 3417 1684 3453 1687
rect 3417 1665 3425 1684
rect 3445 1665 3453 1684
rect 3417 1661 3453 1665
rect 3303 1627 3343 1657
rect 3089 1622 3124 1623
rect 3068 1615 3124 1622
rect 3068 1595 3097 1615
rect 3117 1595 3124 1615
rect 3068 1590 3124 1595
rect 3300 1616 3343 1627
rect 3300 1596 3308 1616
rect 3332 1610 3343 1616
rect 3515 1618 3547 1625
rect 3332 1596 3342 1610
rect 3068 1384 3102 1590
rect 3300 1587 3342 1596
rect 3515 1598 3521 1618
rect 3542 1598 3547 1618
rect 3515 1570 3547 1598
rect 4081 1618 4115 1824
rect 4310 1823 4360 1832
rect 4528 1852 4560 1859
rect 4528 1832 4534 1852
rect 4555 1832 4560 1852
rect 4528 1804 4560 1832
rect 4148 1796 4560 1804
rect 4148 1770 4154 1796
rect 4180 1770 4560 1796
rect 4148 1768 4560 1770
rect 4150 1767 4190 1768
rect 4528 1703 4560 1768
rect 4528 1683 4532 1703
rect 4553 1683 4560 1703
rect 4528 1676 4560 1683
rect 4081 1610 4116 1618
rect 4081 1590 4089 1610
rect 4109 1590 4116 1610
rect 4081 1585 4116 1590
rect 4081 1584 4113 1585
rect 3135 1562 3547 1570
rect 3135 1536 3141 1562
rect 3167 1536 3547 1562
rect 3135 1534 3547 1536
rect 3137 1533 3177 1534
rect 3515 1469 3547 1534
rect 3515 1449 3519 1469
rect 3540 1449 3547 1469
rect 3515 1442 3547 1449
rect 3992 1480 4344 1511
rect 3068 1376 3103 1384
rect 3068 1356 3076 1376
rect 3096 1356 3103 1376
rect 3068 1340 3103 1356
rect 3992 1340 4023 1480
rect 4316 1448 4344 1480
rect 4101 1441 4136 1442
rect 3066 1321 4023 1340
rect 4080 1434 4136 1441
rect 4080 1414 4109 1434
rect 4129 1414 4136 1434
rect 4080 1409 4136 1414
rect 4310 1436 4350 1448
rect 4310 1415 4316 1436
rect 4338 1415 4350 1436
rect 4310 1410 4350 1415
rect 4527 1437 4559 1444
rect 4527 1417 4533 1437
rect 4554 1417 4559 1437
rect 2856 1239 3286 1268
rect 2856 1234 2940 1239
rect 3039 1202 3074 1203
rect 900 1019 1309 1020
rect 2204 1006 2214 1026
rect 2234 1006 2244 1026
rect 2204 996 2244 1006
rect 3018 1195 3074 1202
rect 3018 1175 3047 1195
rect 3067 1175 3074 1195
rect 3018 1170 3074 1175
rect 3248 1196 3286 1239
rect 3248 1179 3253 1196
rect 3277 1179 3286 1196
rect 1763 933 1795 940
rect 1763 913 1770 933
rect 1791 913 1795 933
rect 1763 848 1795 913
rect 2133 848 2173 849
rect 1763 846 2175 848
rect 1763 820 2143 846
rect 2169 820 2175 846
rect 1763 812 2175 820
rect 1148 792 1180 793
rect 1145 787 1180 792
rect 1145 767 1152 787
rect 1172 767 1180 787
rect 1145 759 1180 767
rect 701 694 733 701
rect 701 674 708 694
rect 729 674 733 694
rect 701 609 733 674
rect 1071 609 1111 610
rect 701 607 1113 609
rect 701 581 1081 607
rect 1107 581 1113 607
rect 701 573 1113 581
rect 701 545 733 573
rect 1146 553 1180 759
rect 1763 784 1795 812
rect 2208 792 2242 996
rect 3018 966 3052 1170
rect 3248 1167 3286 1179
rect 3465 1198 3497 1205
rect 3465 1178 3471 1198
rect 3492 1178 3497 1198
rect 3465 1150 3497 1178
rect 4080 1203 4114 1409
rect 4527 1389 4559 1417
rect 4147 1381 4559 1389
rect 4147 1355 4153 1381
rect 4179 1355 4559 1381
rect 4147 1353 4559 1355
rect 4149 1352 4189 1353
rect 4527 1288 4559 1353
rect 4527 1268 4531 1288
rect 4552 1268 4559 1288
rect 4527 1261 4559 1268
rect 4080 1195 4115 1203
rect 4080 1175 4088 1195
rect 4108 1175 4115 1195
rect 4080 1170 4115 1175
rect 4080 1169 4112 1170
rect 3085 1142 3497 1150
rect 3085 1116 3091 1142
rect 3117 1116 3497 1142
rect 3085 1114 3497 1116
rect 3087 1113 3127 1114
rect 3465 1049 3497 1114
rect 3465 1029 3469 1049
rect 3490 1029 3497 1049
rect 3465 1022 3497 1029
rect 1763 764 1768 784
rect 1789 764 1795 784
rect 1763 757 1795 764
rect 1974 784 2011 790
rect 1974 765 1980 784
rect 2003 765 2011 784
rect 1974 760 2011 765
rect 2186 787 2242 792
rect 2186 767 2193 787
rect 2213 767 2242 787
rect 2186 760 2242 767
rect 3016 956 3056 966
rect 3016 936 3026 956
rect 3046 936 3056 956
rect 3951 942 4360 943
rect 1982 723 2006 760
rect 2186 759 2221 760
rect 1982 721 2350 723
rect 1982 716 2355 721
rect 1982 698 2328 716
rect 2348 698 2355 716
rect 1982 693 2355 698
rect 2326 691 2355 693
rect 3016 712 3056 936
rect 3945 913 4360 942
rect 3945 762 3985 913
rect 4319 880 4360 913
rect 4107 875 4142 876
rect 3422 734 3985 762
rect 4086 868 4142 875
rect 4086 848 4115 868
rect 4135 848 4142 868
rect 4086 843 4142 848
rect 4315 872 4365 880
rect 4315 851 4331 872
rect 4353 851 4365 872
rect 3016 678 3343 712
rect 3423 706 3457 734
rect 3422 703 3458 706
rect 3422 684 3430 703
rect 3450 684 3458 703
rect 3422 680 3458 684
rect 3033 677 3343 678
rect 3308 648 3343 677
rect 3094 641 3129 642
rect 701 525 706 545
rect 727 525 733 545
rect 701 518 733 525
rect 910 547 950 552
rect 910 526 922 547
rect 944 526 950 547
rect 910 514 950 526
rect 1124 548 1180 553
rect 1124 528 1131 548
rect 1151 528 1180 548
rect 1124 521 1180 528
rect 1237 622 2194 641
rect 3073 634 3129 641
rect 1124 520 1159 521
rect 916 482 944 514
rect 1237 482 1268 622
rect 2157 606 2192 622
rect 2157 586 2164 606
rect 2184 586 2192 606
rect 2157 578 2192 586
rect 916 451 1268 482
rect 1713 513 1745 520
rect 1713 493 1720 513
rect 1741 493 1745 513
rect 1713 428 1745 493
rect 2083 428 2123 429
rect 1713 426 2125 428
rect 1713 400 2093 426
rect 2119 400 2125 426
rect 1713 392 2125 400
rect 1147 377 1179 378
rect 1144 372 1179 377
rect 1144 352 1151 372
rect 1171 352 1179 372
rect 1144 344 1179 352
rect 700 279 732 286
rect 700 259 707 279
rect 728 259 732 279
rect 700 194 732 259
rect 1070 194 1110 195
rect 700 192 1112 194
rect 700 166 1080 192
rect 1106 166 1112 192
rect 700 158 1112 166
rect 700 130 732 158
rect 700 110 705 130
rect 726 110 732 130
rect 700 103 732 110
rect 900 130 950 139
rect 1145 138 1179 344
rect 1713 364 1745 392
rect 1713 344 1718 364
rect 1739 344 1745 364
rect 1918 366 1960 375
rect 2158 372 2192 578
rect 1918 352 1928 366
rect 1713 337 1745 344
rect 1917 346 1928 352
rect 1952 346 1960 366
rect 1917 335 1960 346
rect 2136 367 2192 372
rect 2136 347 2143 367
rect 2163 347 2192 367
rect 3073 614 3102 634
rect 3122 614 3129 634
rect 3073 609 3129 614
rect 3303 636 3345 648
rect 3303 616 3312 636
rect 3336 616 3345 636
rect 3073 403 3107 609
rect 3303 608 3345 616
rect 3520 637 3552 644
rect 3520 617 3526 637
rect 3547 617 3552 637
rect 3520 589 3552 617
rect 4086 637 4120 843
rect 4315 842 4365 851
rect 4533 871 4565 878
rect 4533 851 4539 871
rect 4560 851 4565 871
rect 4533 823 4565 851
rect 4153 815 4565 823
rect 4153 789 4159 815
rect 4185 789 4565 815
rect 4153 787 4565 789
rect 4155 786 4195 787
rect 4533 722 4565 787
rect 4533 702 4537 722
rect 4558 702 4565 722
rect 4533 695 4565 702
rect 4086 629 4121 637
rect 4086 609 4094 629
rect 4114 609 4121 629
rect 4086 604 4121 609
rect 4086 603 4118 604
rect 3140 581 3552 589
rect 3140 555 3146 581
rect 3172 555 3552 581
rect 3140 553 3552 555
rect 3142 552 3182 553
rect 3520 488 3552 553
rect 3520 468 3524 488
rect 3545 468 3552 488
rect 3520 461 3552 468
rect 3997 499 4349 530
rect 3073 395 3108 403
rect 3073 375 3081 395
rect 3101 375 3108 395
rect 3073 359 3108 375
rect 3997 359 4028 499
rect 4321 467 4349 499
rect 4106 460 4141 461
rect 2136 340 2192 347
rect 3071 340 4028 359
rect 4085 453 4141 460
rect 4085 433 4114 453
rect 4134 433 4141 453
rect 4085 428 4141 433
rect 4315 455 4355 467
rect 4315 434 4321 455
rect 4343 434 4355 455
rect 4315 429 4355 434
rect 4532 456 4564 463
rect 4532 436 4538 456
rect 4559 436 4564 456
rect 2136 339 2171 340
rect 1917 305 1957 335
rect 1807 297 1843 301
rect 1807 278 1815 297
rect 1835 278 1843 297
rect 1807 275 1843 278
rect 1917 300 2264 305
rect 1808 247 1842 275
rect 1917 274 2236 300
rect 2255 274 2264 300
rect 1917 270 2264 274
rect 900 109 912 130
rect 934 109 950 130
rect 900 101 950 109
rect 1123 133 1179 138
rect 1123 113 1130 133
rect 1150 113 1179 133
rect 1123 106 1179 113
rect 1280 219 1843 247
rect 4085 222 4119 428
rect 4532 408 4564 436
rect 4152 400 4564 408
rect 4152 374 4158 400
rect 4184 374 4564 400
rect 4152 372 4564 374
rect 4154 371 4194 372
rect 4532 307 4564 372
rect 4532 287 4536 307
rect 4557 287 4564 307
rect 4532 280 4564 287
rect 1123 105 1158 106
rect 905 68 946 101
rect 1280 68 1320 219
rect 4085 214 4120 222
rect 4085 194 4093 214
rect 4113 194 4120 214
rect 4085 189 4120 194
rect 4085 188 4117 189
rect 905 39 1320 68
rect 905 38 1314 39
rect 747 10 787 15
rect 694 7 5119 10
rect 694 -15 756 7
rect 779 -15 5089 7
rect 5112 -15 5119 7
rect 694 -20 5119 -15
rect 747 -30 787 -20
rect 2543 -62 2592 -58
rect 2543 -63 2553 -62
rect 2543 -92 2552 -63
rect 2584 -92 2592 -62
rect 2543 -93 2592 -92
rect 2542 -101 2592 -93
rect 2542 -109 2591 -101
rect 2542 -129 2554 -109
rect 2574 -129 2591 -109
rect 2542 -136 2591 -129
rect 2646 -110 2694 -107
rect 2547 -137 2582 -136
rect 2103 -202 2135 -195
rect 2103 -222 2110 -202
rect 2131 -222 2135 -202
rect 2103 -287 2135 -222
rect 2473 -287 2513 -286
rect 2103 -289 2515 -287
rect 2103 -315 2483 -289
rect 2509 -315 2515 -289
rect 2103 -323 2515 -315
rect 2103 -351 2135 -323
rect 2548 -343 2582 -137
rect 2646 -137 2649 -110
rect 2684 -137 2694 -110
rect 2646 -204 2694 -137
rect 2646 -224 2651 -204
rect 2679 -224 2694 -204
rect 2646 -234 2694 -224
rect 2103 -371 2108 -351
rect 2129 -371 2135 -351
rect 2103 -378 2135 -371
rect 2311 -351 2355 -344
rect 2311 -373 2322 -351
rect 2347 -373 2355 -351
rect 2311 -381 2355 -373
rect 2526 -348 2582 -343
rect 2526 -368 2533 -348
rect 2553 -368 2582 -348
rect 2526 -375 2582 -368
rect 2526 -376 2561 -375
rect 2317 -411 2342 -381
rect 2317 -444 2748 -411
<< via1 >>
rect 2649 4165 2686 4195
rect 2548 3644 2582 3672
rect 2553 -63 2584 -62
rect 2552 -92 2584 -63
rect 2649 -137 2684 -110
<< metal2 >>
rect 2644 4195 2693 4201
rect 2644 4165 2649 4195
rect 2686 4165 2693 4195
rect 2542 3672 2587 3678
rect 2542 3644 2548 3672
rect 2582 3644 2587 3672
rect 2542 34 2587 3644
rect 2644 65 2693 4165
rect 2548 -58 2586 34
rect 2543 -62 2592 -58
rect 2543 -63 2553 -62
rect 2543 -92 2552 -63
rect 2584 -92 2592 -62
rect 2543 -101 2592 -92
rect 2646 -110 2692 65
rect 2646 -137 2649 -110
rect 2684 -137 2692 -110
rect 2646 -152 2692 -137
<< labels >>
rlabel locali 304 7629 333 7635 1 vdd
rlabel locali 517 7626 546 7632 1 vdd
rlabel locali 250 7441 272 7456 1 d0
rlabel nwell 671 7596 694 7599 1 vdd
rlabel locali 301 7330 330 7336 1 gnd
rlabel locali 514 7330 543 7336 1 gnd
rlabel space 611 7325 640 7334 1 gnd
rlabel locali 303 7214 332 7220 1 vdd
rlabel locali 516 7211 545 7217 1 vdd
rlabel locali 249 7026 271 7041 1 d0
rlabel nwell 670 7181 693 7184 1 vdd
rlabel locali 300 6915 329 6921 1 gnd
rlabel locali 513 6915 542 6921 1 gnd
rlabel space 610 6910 639 6919 1 gnd
rlabel locali 1316 7448 1345 7454 1 vdd
rlabel locali 1529 7445 1558 7451 1 vdd
rlabel nwell 1683 7415 1706 7418 1 vdd
rlabel locali 1313 7149 1342 7155 1 gnd
rlabel locali 1526 7149 1555 7155 1 gnd
rlabel space 1623 7144 1652 7153 1 gnd
rlabel locali 1254 7259 1301 7280 1 d1
rlabel locali 116 7821 141 7830 1 vref
rlabel locali 309 6648 338 6654 1 vdd
rlabel locali 522 6645 551 6651 1 vdd
rlabel locali 255 6460 277 6475 1 d0
rlabel nwell 676 6615 699 6618 1 vdd
rlabel locali 306 6349 335 6355 1 gnd
rlabel locali 519 6349 548 6355 1 gnd
rlabel space 616 6344 645 6353 1 gnd
rlabel locali 308 6233 337 6239 1 vdd
rlabel locali 521 6230 550 6236 1 vdd
rlabel locali 254 6045 276 6060 1 d0
rlabel nwell 675 6200 698 6203 1 vdd
rlabel locali 305 5934 334 5940 1 gnd
rlabel locali 518 5934 547 5940 1 gnd
rlabel locali 1321 6467 1350 6473 1 vdd
rlabel locali 1534 6464 1563 6470 1 vdd
rlabel nwell 1688 6434 1711 6437 1 vdd
rlabel locali 1318 6168 1347 6174 1 gnd
rlabel locali 1531 6168 1560 6174 1 gnd
rlabel space 1628 6163 1657 6172 1 gnd
rlabel locali 1259 6278 1306 6299 1 d1
rlabel locali 1371 6887 1400 6893 1 vdd
rlabel locali 1584 6884 1613 6890 1 vdd
rlabel nwell 1738 6854 1761 6857 1 vdd
rlabel locali 1368 6588 1397 6594 1 gnd
rlabel locali 1581 6588 1610 6594 1 gnd
rlabel space 1678 6583 1707 6592 1 gnd
rlabel locali 1314 6699 1337 6714 1 d2
rlabel space 615 5929 644 5938 1 gnd
rlabel locali 1326 4739 1349 4754 1 d2
rlabel space 1690 4623 1719 4632 1 gnd
rlabel locali 1593 4628 1622 4634 1 gnd
rlabel locali 1380 4628 1409 4634 1 gnd
rlabel nwell 1750 4894 1773 4897 1 vdd
rlabel locali 1596 4924 1625 4930 1 vdd
rlabel locali 1383 4927 1412 4933 1 vdd
rlabel locali 1271 4318 1318 4339 1 d1
rlabel space 1640 4203 1669 4212 1 gnd
rlabel locali 1543 4208 1572 4214 1 gnd
rlabel locali 1330 4208 1359 4214 1 gnd
rlabel nwell 1700 4474 1723 4477 1 vdd
rlabel locali 1546 4504 1575 4510 1 vdd
rlabel locali 1333 4507 1362 4513 1 vdd
rlabel space 627 3969 656 3978 1 gnd
rlabel locali 530 3974 559 3980 1 gnd
rlabel locali 317 3974 346 3980 1 gnd
rlabel nwell 687 4240 710 4243 1 vdd
rlabel locali 266 4085 288 4100 1 d0
rlabel locali 533 4270 562 4276 1 vdd
rlabel locali 320 4273 349 4279 1 vdd
rlabel space 628 4384 657 4393 1 gnd
rlabel locali 531 4389 560 4395 1 gnd
rlabel locali 318 4389 347 4395 1 gnd
rlabel nwell 688 4655 711 4658 1 vdd
rlabel locali 267 4500 289 4515 1 d0
rlabel locali 534 4685 563 4691 1 vdd
rlabel locali 321 4688 350 4694 1 vdd
rlabel locali 1266 5299 1313 5320 1 d1
rlabel space 1635 5184 1664 5193 1 gnd
rlabel locali 1538 5189 1567 5195 1 gnd
rlabel locali 1325 5189 1354 5195 1 gnd
rlabel nwell 1695 5455 1718 5458 1 vdd
rlabel locali 1541 5485 1570 5491 1 vdd
rlabel locali 1328 5488 1357 5494 1 vdd
rlabel space 622 4950 651 4959 1 gnd
rlabel locali 525 4955 554 4961 1 gnd
rlabel locali 312 4955 341 4961 1 gnd
rlabel nwell 682 5221 705 5224 1 vdd
rlabel locali 261 5066 283 5081 1 d0
rlabel locali 528 5251 557 5257 1 vdd
rlabel locali 315 5254 344 5260 1 vdd
rlabel space 623 5365 652 5374 1 gnd
rlabel locali 526 5370 555 5376 1 gnd
rlabel locali 313 5370 342 5376 1 gnd
rlabel nwell 683 5636 706 5639 1 vdd
rlabel locali 262 5481 284 5496 1 d0
rlabel locali 529 5666 558 5672 1 vdd
rlabel locali 316 5669 345 5675 1 vdd
rlabel locali 1536 5955 1565 5961 1 vdd
rlabel locali 1749 5952 1778 5958 1 vdd
rlabel nwell 1903 5922 1926 5925 1 vdd
rlabel locali 1533 5656 1562 5662 1 gnd
rlabel locali 1746 5656 1775 5662 1 gnd
rlabel space 1843 5651 1872 5660 1 gnd
rlabel locali 1474 5765 1506 5784 1 d3
rlabel locali 1494 1848 1526 1867 1 d3
rlabel space 1863 1734 1892 1743 1 gnd
rlabel locali 1766 1739 1795 1745 1 gnd
rlabel locali 1553 1739 1582 1745 1 gnd
rlabel nwell 1923 2005 1946 2008 1 vdd
rlabel locali 1769 2035 1798 2041 1 vdd
rlabel locali 1556 2038 1585 2044 1 vdd
rlabel locali 336 1752 365 1758 1 vdd
rlabel locali 549 1749 578 1755 1 vdd
rlabel locali 282 1564 304 1579 1 d0
rlabel nwell 703 1719 726 1722 1 vdd
rlabel locali 333 1453 362 1459 1 gnd
rlabel locali 546 1453 575 1459 1 gnd
rlabel space 643 1448 672 1457 1 gnd
rlabel locali 335 1337 364 1343 1 vdd
rlabel locali 548 1334 577 1340 1 vdd
rlabel locali 281 1149 303 1164 1 d0
rlabel nwell 702 1304 725 1307 1 vdd
rlabel locali 332 1038 361 1044 1 gnd
rlabel locali 545 1038 574 1044 1 gnd
rlabel space 642 1033 671 1042 1 gnd
rlabel locali 1348 1571 1377 1577 1 vdd
rlabel locali 1561 1568 1590 1574 1 vdd
rlabel nwell 1715 1538 1738 1541 1 vdd
rlabel locali 1345 1272 1374 1278 1 gnd
rlabel locali 1558 1272 1587 1278 1 gnd
rlabel space 1655 1267 1684 1276 1 gnd
rlabel locali 1286 1382 1333 1403 1 d1
rlabel locali 341 771 370 777 1 vdd
rlabel locali 554 768 583 774 1 vdd
rlabel locali 287 583 309 598 1 d0
rlabel nwell 708 738 731 741 1 vdd
rlabel locali 338 472 367 478 1 gnd
rlabel locali 551 472 580 478 1 gnd
rlabel space 648 467 677 476 1 gnd
rlabel locali 340 356 369 362 1 vdd
rlabel locali 553 353 582 359 1 vdd
rlabel locali 286 168 308 183 1 d0
rlabel nwell 707 323 730 326 1 vdd
rlabel locali 337 57 366 63 1 gnd
rlabel locali 550 57 579 63 1 gnd
rlabel space 647 52 676 61 1 gnd
rlabel locali 1353 590 1382 596 1 vdd
rlabel locali 1566 587 1595 593 1 vdd
rlabel nwell 1720 557 1743 560 1 vdd
rlabel locali 1350 291 1379 297 1 gnd
rlabel locali 1563 291 1592 297 1 gnd
rlabel space 1660 286 1689 295 1 gnd
rlabel locali 1291 401 1338 422 1 d1
rlabel locali 1403 1010 1432 1016 1 vdd
rlabel locali 1616 1007 1645 1013 1 vdd
rlabel nwell 1770 977 1793 980 1 vdd
rlabel locali 1400 711 1429 717 1 gnd
rlabel locali 1613 711 1642 717 1 gnd
rlabel space 1710 706 1739 715 1 gnd
rlabel locali 1346 822 1369 837 1 d2
rlabel space 635 2012 664 2021 1 gnd
rlabel locali 1334 2782 1357 2797 1 d2
rlabel space 1698 2666 1727 2675 1 gnd
rlabel locali 1601 2671 1630 2677 1 gnd
rlabel locali 1388 2671 1417 2677 1 gnd
rlabel nwell 1758 2937 1781 2940 1 vdd
rlabel locali 1604 2967 1633 2973 1 vdd
rlabel locali 1391 2970 1420 2976 1 vdd
rlabel locali 1279 2361 1326 2382 1 d1
rlabel space 1648 2246 1677 2255 1 gnd
rlabel locali 1551 2251 1580 2257 1 gnd
rlabel locali 1338 2251 1367 2257 1 gnd
rlabel nwell 1708 2517 1731 2520 1 vdd
rlabel locali 1554 2547 1583 2553 1 vdd
rlabel locali 1341 2550 1370 2556 1 vdd
rlabel locali 538 2017 567 2023 1 gnd
rlabel locali 325 2017 354 2023 1 gnd
rlabel nwell 695 2283 718 2286 1 vdd
rlabel locali 274 2128 296 2143 1 d0
rlabel locali 541 2313 570 2319 1 vdd
rlabel locali 328 2316 357 2322 1 vdd
rlabel space 636 2427 665 2436 1 gnd
rlabel locali 539 2432 568 2438 1 gnd
rlabel locali 326 2432 355 2438 1 gnd
rlabel nwell 696 2698 719 2701 1 vdd
rlabel locali 275 2543 297 2558 1 d0
rlabel locali 542 2728 571 2734 1 vdd
rlabel locali 329 2731 358 2737 1 vdd
rlabel locali 1274 3342 1321 3363 1 d1
rlabel space 1643 3227 1672 3236 1 gnd
rlabel locali 1546 3232 1575 3238 1 gnd
rlabel locali 1333 3232 1362 3238 1 gnd
rlabel nwell 1703 3498 1726 3501 1 vdd
rlabel locali 1549 3528 1578 3534 1 vdd
rlabel locali 1336 3531 1365 3537 1 vdd
rlabel space 630 2993 659 3002 1 gnd
rlabel locali 533 2998 562 3004 1 gnd
rlabel locali 320 2998 349 3004 1 gnd
rlabel nwell 690 3264 713 3267 1 vdd
rlabel locali 269 3109 291 3124 1 d0
rlabel locali 536 3294 565 3300 1 vdd
rlabel locali 323 3297 352 3303 1 vdd
rlabel space 631 3408 660 3417 1 gnd
rlabel locali 534 3413 563 3419 1 gnd
rlabel locali 321 3413 350 3419 1 gnd
rlabel nwell 691 3679 714 3682 1 vdd
rlabel locali 270 3524 292 3539 1 d0
rlabel locali 537 3709 566 3715 1 vdd
rlabel locali 324 3712 353 3718 1 vdd
rlabel locali 1631 3963 1660 3969 1 vdd
rlabel locali 1844 3960 1873 3966 1 vdd
rlabel nwell 1998 3930 2021 3933 1 vdd
rlabel locali 1628 3664 1657 3670 1 gnd
rlabel locali 1841 3664 1870 3670 1 gnd
rlabel space 1938 3659 1967 3668 1 gnd
rlabel locali 1573 3769 1595 3793 1 d4
rlabel locali 4895 204 4924 210 5 vdd
rlabel locali 4682 207 4711 213 5 vdd
rlabel locali 4956 383 4978 398 5 d0
rlabel nwell 4534 240 4557 243 5 vdd
rlabel locali 4898 503 4927 509 5 gnd
rlabel locali 4685 503 4714 509 5 gnd
rlabel space 4588 505 4617 514 5 gnd
rlabel locali 4896 619 4925 625 5 vdd
rlabel locali 4683 622 4712 628 5 vdd
rlabel locali 4957 798 4979 813 5 d0
rlabel nwell 4535 655 4558 658 5 vdd
rlabel locali 4899 918 4928 924 5 gnd
rlabel locali 4686 918 4715 924 5 gnd
rlabel space 4589 920 4618 929 5 gnd
rlabel locali 3883 385 3912 391 5 vdd
rlabel locali 3670 388 3699 394 5 vdd
rlabel nwell 3522 421 3545 424 5 vdd
rlabel locali 3886 684 3915 690 5 gnd
rlabel locali 3673 684 3702 690 5 gnd
rlabel space 3576 686 3605 695 5 gnd
rlabel locali 3927 559 3974 580 5 d1
rlabel locali 4890 1185 4919 1191 5 vdd
rlabel locali 4677 1188 4706 1194 5 vdd
rlabel locali 4951 1364 4973 1379 5 d0
rlabel nwell 4529 1221 4552 1224 5 vdd
rlabel locali 4893 1484 4922 1490 5 gnd
rlabel locali 4680 1484 4709 1490 5 gnd
rlabel space 4583 1486 4612 1495 5 gnd
rlabel locali 4891 1600 4920 1606 5 vdd
rlabel locali 4678 1603 4707 1609 5 vdd
rlabel locali 4952 1779 4974 1794 5 d0
rlabel nwell 4530 1636 4553 1639 5 vdd
rlabel locali 4894 1899 4923 1905 5 gnd
rlabel locali 4681 1899 4710 1905 5 gnd
rlabel locali 3878 1366 3907 1372 5 vdd
rlabel locali 3665 1369 3694 1375 5 vdd
rlabel nwell 3517 1402 3540 1405 5 vdd
rlabel locali 3881 1665 3910 1671 5 gnd
rlabel locali 3668 1665 3697 1671 5 gnd
rlabel space 3571 1667 3600 1676 5 gnd
rlabel locali 3922 1540 3969 1561 5 d1
rlabel locali 3828 946 3857 952 5 vdd
rlabel locali 3615 949 3644 955 5 vdd
rlabel nwell 3467 982 3490 985 5 vdd
rlabel locali 3831 1245 3860 1251 5 gnd
rlabel locali 3618 1245 3647 1251 5 gnd
rlabel space 3521 1247 3550 1256 5 gnd
rlabel locali 3891 1125 3914 1140 5 d2
rlabel space 4584 1901 4613 1910 5 gnd
rlabel locali 3879 3085 3902 3100 5 d2
rlabel space 3509 3207 3538 3216 5 gnd
rlabel locali 3606 3205 3635 3211 5 gnd
rlabel locali 3819 3205 3848 3211 5 gnd
rlabel nwell 3455 2942 3478 2945 5 vdd
rlabel locali 3603 2909 3632 2915 5 vdd
rlabel locali 3816 2906 3845 2912 5 vdd
rlabel locali 3910 3500 3957 3521 5 d1
rlabel space 3559 3627 3588 3636 5 gnd
rlabel locali 3656 3625 3685 3631 5 gnd
rlabel locali 3869 3625 3898 3631 5 gnd
rlabel nwell 3505 3362 3528 3365 5 vdd
rlabel locali 3653 3329 3682 3335 5 vdd
rlabel locali 3866 3326 3895 3332 5 vdd
rlabel space 4572 3861 4601 3870 5 gnd
rlabel locali 4669 3859 4698 3865 5 gnd
rlabel locali 4882 3859 4911 3865 5 gnd
rlabel nwell 4518 3596 4541 3599 5 vdd
rlabel locali 4940 3739 4962 3754 5 d0
rlabel locali 4666 3563 4695 3569 5 vdd
rlabel locali 4879 3560 4908 3566 5 vdd
rlabel space 4571 3446 4600 3455 5 gnd
rlabel locali 4668 3444 4697 3450 5 gnd
rlabel locali 4881 3444 4910 3450 5 gnd
rlabel nwell 4517 3181 4540 3184 5 vdd
rlabel locali 4939 3324 4961 3339 5 d0
rlabel locali 4665 3148 4694 3154 5 vdd
rlabel locali 4878 3145 4907 3151 5 vdd
rlabel locali 3915 2519 3962 2540 5 d1
rlabel space 3564 2646 3593 2655 5 gnd
rlabel locali 3661 2644 3690 2650 5 gnd
rlabel locali 3874 2644 3903 2650 5 gnd
rlabel nwell 3510 2381 3533 2384 5 vdd
rlabel locali 3658 2348 3687 2354 5 vdd
rlabel locali 3871 2345 3900 2351 5 vdd
rlabel space 4577 2880 4606 2889 5 gnd
rlabel locali 4674 2878 4703 2884 5 gnd
rlabel locali 4887 2878 4916 2884 5 gnd
rlabel nwell 4523 2615 4546 2618 5 vdd
rlabel locali 4945 2758 4967 2773 5 d0
rlabel locali 4671 2582 4700 2588 5 vdd
rlabel locali 4884 2579 4913 2585 5 vdd
rlabel space 4576 2465 4605 2474 5 gnd
rlabel locali 4673 2463 4702 2469 5 gnd
rlabel locali 4886 2463 4915 2469 5 gnd
rlabel nwell 4522 2200 4545 2203 5 vdd
rlabel locali 4944 2343 4966 2358 5 d0
rlabel locali 4670 2167 4699 2173 5 vdd
rlabel locali 4883 2164 4912 2170 5 vdd
rlabel locali 3663 1878 3692 1884 5 vdd
rlabel locali 3450 1881 3479 1887 5 vdd
rlabel nwell 3302 1914 3325 1917 5 vdd
rlabel locali 3666 2177 3695 2183 5 gnd
rlabel locali 3453 2177 3482 2183 5 gnd
rlabel space 3356 2179 3385 2188 5 gnd
rlabel locali 3722 2055 3754 2074 5 d3
rlabel locali 3702 5972 3734 5991 5 d3
rlabel space 3336 6096 3365 6105 5 gnd
rlabel locali 3433 6094 3462 6100 5 gnd
rlabel locali 3646 6094 3675 6100 5 gnd
rlabel nwell 3282 5831 3305 5834 5 vdd
rlabel locali 3430 5798 3459 5804 5 vdd
rlabel locali 3643 5795 3672 5801 5 vdd
rlabel locali 4863 6081 4892 6087 5 vdd
rlabel locali 4650 6084 4679 6090 5 vdd
rlabel locali 4924 6260 4946 6275 5 d0
rlabel nwell 4502 6117 4525 6120 5 vdd
rlabel locali 4866 6380 4895 6386 5 gnd
rlabel locali 4653 6380 4682 6386 5 gnd
rlabel space 4556 6382 4585 6391 5 gnd
rlabel locali 4864 6496 4893 6502 5 vdd
rlabel locali 4651 6499 4680 6505 5 vdd
rlabel locali 4925 6675 4947 6690 5 d0
rlabel nwell 4503 6532 4526 6535 5 vdd
rlabel locali 4867 6795 4896 6801 5 gnd
rlabel locali 4654 6795 4683 6801 5 gnd
rlabel space 4557 6797 4586 6806 5 gnd
rlabel locali 3851 6262 3880 6268 5 vdd
rlabel locali 3638 6265 3667 6271 5 vdd
rlabel nwell 3490 6298 3513 6301 5 vdd
rlabel locali 3854 6561 3883 6567 5 gnd
rlabel locali 3641 6561 3670 6567 5 gnd
rlabel space 3544 6563 3573 6572 5 gnd
rlabel locali 3895 6436 3942 6457 5 d1
rlabel locali 4858 7062 4887 7068 5 vdd
rlabel locali 4645 7065 4674 7071 5 vdd
rlabel locali 4919 7241 4941 7256 5 d0
rlabel nwell 4497 7098 4520 7101 5 vdd
rlabel locali 4861 7361 4890 7367 5 gnd
rlabel locali 4648 7361 4677 7367 5 gnd
rlabel space 4551 7363 4580 7372 5 gnd
rlabel locali 4859 7477 4888 7483 5 vdd
rlabel locali 4646 7480 4675 7486 5 vdd
rlabel locali 4920 7656 4942 7671 5 d0
rlabel nwell 4498 7513 4521 7516 5 vdd
rlabel locali 4862 7776 4891 7782 5 gnd
rlabel locali 4649 7776 4678 7782 5 gnd
rlabel space 4552 7778 4581 7787 5 gnd
rlabel locali 3846 7243 3875 7249 5 vdd
rlabel locali 3633 7246 3662 7252 5 vdd
rlabel nwell 3485 7279 3508 7282 5 vdd
rlabel locali 3849 7542 3878 7548 5 gnd
rlabel locali 3636 7542 3665 7548 5 gnd
rlabel space 3539 7544 3568 7553 5 gnd
rlabel locali 3890 7417 3937 7438 5 d1
rlabel locali 5043 7818 5070 7831 5 gnd
rlabel locali 3796 6823 3825 6829 5 vdd
rlabel locali 3583 6826 3612 6832 5 vdd
rlabel nwell 3435 6859 3458 6862 5 vdd
rlabel locali 3799 7122 3828 7128 5 gnd
rlabel locali 3586 7122 3615 7128 5 gnd
rlabel space 3489 7124 3518 7133 5 gnd
rlabel locali 3859 7002 3882 7017 5 d2
rlabel space 4564 5818 4593 5827 5 gnd
rlabel locali 3871 5042 3894 5057 5 d2
rlabel space 3501 5164 3530 5173 5 gnd
rlabel locali 3598 5162 3627 5168 5 gnd
rlabel locali 3811 5162 3840 5168 5 gnd
rlabel nwell 3447 4899 3470 4902 5 vdd
rlabel locali 3595 4866 3624 4872 5 vdd
rlabel locali 3808 4863 3837 4869 5 vdd
rlabel locali 3902 5457 3949 5478 5 d1
rlabel space 3551 5584 3580 5593 5 gnd
rlabel locali 3648 5582 3677 5588 5 gnd
rlabel locali 3861 5582 3890 5588 5 gnd
rlabel nwell 3497 5319 3520 5322 5 vdd
rlabel locali 3645 5286 3674 5292 5 vdd
rlabel locali 3858 5283 3887 5289 5 vdd
rlabel locali 4661 5816 4690 5822 5 gnd
rlabel locali 4874 5816 4903 5822 5 gnd
rlabel nwell 4510 5553 4533 5556 5 vdd
rlabel locali 4932 5696 4954 5711 5 d0
rlabel locali 4658 5520 4687 5526 5 vdd
rlabel locali 4871 5517 4900 5523 5 vdd
rlabel space 4563 5403 4592 5412 5 gnd
rlabel locali 4660 5401 4689 5407 5 gnd
rlabel locali 4873 5401 4902 5407 5 gnd
rlabel nwell 4509 5138 4532 5141 5 vdd
rlabel locali 4931 5281 4953 5296 5 d0
rlabel locali 4657 5105 4686 5111 5 vdd
rlabel locali 4870 5102 4899 5108 5 vdd
rlabel locali 3907 4476 3954 4497 5 d1
rlabel space 3556 4603 3585 4612 5 gnd
rlabel locali 3653 4601 3682 4607 5 gnd
rlabel locali 3866 4601 3895 4607 5 gnd
rlabel nwell 3502 4338 3525 4341 5 vdd
rlabel locali 3650 4305 3679 4311 5 vdd
rlabel locali 3863 4302 3892 4308 5 vdd
rlabel space 4569 4837 4598 4846 5 gnd
rlabel locali 4666 4835 4695 4841 5 gnd
rlabel locali 4879 4835 4908 4841 5 gnd
rlabel nwell 4515 4572 4538 4575 5 vdd
rlabel locali 4937 4715 4959 4730 5 d0
rlabel locali 4663 4539 4692 4545 5 vdd
rlabel locali 4876 4536 4905 4542 5 vdd
rlabel space 4568 4422 4597 4431 5 gnd
rlabel locali 4665 4420 4694 4426 5 gnd
rlabel locali 4878 4420 4907 4426 5 gnd
rlabel nwell 4514 4157 4537 4160 5 vdd
rlabel locali 4936 4300 4958 4315 5 d0
rlabel locali 4662 4124 4691 4130 5 vdd
rlabel locali 4875 4121 4904 4127 5 vdd
rlabel locali 3568 3870 3597 3876 5 vdd
rlabel locali 3355 3873 3384 3879 5 vdd
rlabel nwell 3207 3906 3230 3909 5 vdd
rlabel locali 3571 4169 3600 4175 5 gnd
rlabel locali 3358 4169 3387 4175 5 gnd
rlabel space 3261 4171 3290 4180 5 gnd
rlabel locali 3633 4046 3655 4070 5 d4
rlabel locali 1743 -125 1772 -119 1 vdd
rlabel locali 1956 -128 1985 -122 1 vdd
rlabel nwell 2110 -158 2133 -155 1 vdd
rlabel locali 1740 -424 1769 -418 1 gnd
rlabel locali 1953 -424 1982 -418 1 gnd
rlabel space 2050 -429 2079 -420 1 gnd
rlabel locali 2319 -278 2341 -263 1 vout
rlabel locali 1685 -316 1709 -299 1 d5
<< end >>
