magic
tech sky130A
timestamp 1616448691
<< metal1 >>
rect -984 12417 -496 12449
rect -984 11818 12410 12417
rect -984 -1163 12375 11818
rect -984 -1226 -464 -1163
rect 11855 -1226 12375 -1163
<< metal3 >>
rect -984 12417 -496 12449
rect -984 11818 12410 12417
rect -984 -1163 12375 11818
rect -984 -1226 -464 -1163
rect 11855 -1226 12375 -1163
<< mimcap >>
rect -260 -442 11803 11706
<< end >>
