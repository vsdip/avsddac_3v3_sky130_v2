* SPICE3 file created from 4bit_DAC.ext - technology: sky130A

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_852_1280# a_1583_1590# a_1791_1590# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1 a_433_731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_118_n1178# a_118_n1365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3 a_117_n262# a_646_n372# a_854_n372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_432_177# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5 a_1584_487# a_1371_487# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_116_1485# a_644_1280# a_852_1280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7 a_118_n1365# a_118_n1594# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8 a_852_1280# a_431_1280# a_116_1485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9 a_118_n1594# a_647_n1475# a_855_n1475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X10 a_1725_n1208# a_1512_n1208# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X11 a_853_1834# a_432_1834# a_116_1944# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X12 a_1803_n92# a_1512_n1208# a_1792_n616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X13 a_117_382# a_117_n75# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X14 a_1511_998# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_1808_27# a_1511_998# a_1792_487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_645_n926# a_432_n926# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 a_116_1944# a_645_1834# a_853_1834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_646_n372# a_433_n372# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X19 a_1372_n1719# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X20 a_432_n926# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X21 a_117_n75# a_117_n262# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X22 a_855_n1475# a_434_n1475# a_118_n1365# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X23 a_118_n1824# a_646_n2029# a_854_n2029# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_1481_n92# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X25 a_433_731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X26 a_433_n372# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X27 a_1724_998# a_1511_998# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X28 vout a_1481_n92# a_1808_27# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X29 a_1584_n616# a_1371_n616# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X30 a_1511_998# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X31 a_1583_1590# a_1370_1590# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X32 a_1371_n616# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X33 a_117_612# a_117_382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X34 a_1585_n1719# a_1372_n1719# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X35 a_118_n1365# a_647_n1475# a_855_n1475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X36 a_1370_1590# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X37 a_647_n1475# a_434_n1475# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X38 a_1791_1590# a_1370_1590# a_852_1280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 gnd a_646_n2029# a_854_n2029# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X40 a_854_n2029# a_433_n2029# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X41 a_853_n926# a_432_n926# a_117_n721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X42 vout a_1481_n92# a_1803_n92# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X43 a_1481_n92# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X44 a_1793_n1719# a_1372_n1719# a_855_n1475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X45 a_853_177# a_432_177# a_117_n75# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X46 a_117_1028# a_644_1280# a_852_1280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X47 a_1792_n616# a_1371_n616# a_853_n926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_117_382# a_645_177# a_853_177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_116_1715# a_645_1834# a_853_1834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X50 a_855_n1475# a_1585_n1719# a_1793_n1719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_645_177# a_432_177# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_1791_1590# a_1724_998# a_1808_27# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X53 a_646_n372# a_433_n372# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_117_n491# a_117_n721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X55 a_855_n1475# a_434_n1475# a_118_n1594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X56 a_644_1280# a_431_1280# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X57 a_433_n372# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X58 a_646_n2029# a_433_n2029# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X59 a_854_n2029# a_433_n2029# a_118_n1824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X60 a_853_1834# a_1583_1590# a_1791_1590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X61 a_431_1280# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X62 a_853_n926# a_1584_n616# a_1792_n616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X63 a_1803_n92# a_1694_n92# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X64 a_1792_n616# a_1725_n1208# a_1803_n92# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 a_853_177# a_1584_487# a_1792_487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X66 a_1694_n92# a_1481_n92# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X67 a_117_1028# a_117_841# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X68 a_1512_n1208# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X69 a_854_731# a_433_731# a_117_612# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X70 a_1792_487# a_1371_487# a_853_177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X71 a_1371_487# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_647_n1475# a_434_n1475# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 a_853_177# a_432_177# a_117_382# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X74 a_1584_487# a_1371_487# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X75 a_853_n926# a_432_n926# a_118_n1178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X76 a_117_841# a_646_731# a_854_731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 a_645_1834# a_432_1834# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 a_646_n2029# a_433_n2029# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X79 a_117_n721# a_118_n1178# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X80 a_854_n372# a_433_n372# a_117_n262# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X81 a_1808_27# a_1694_n92# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X82 a_117_n75# a_645_177# a_853_177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X83 a_646_731# a_433_731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X84 a_432_1834# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X85 a_1725_n1208# a_1512_n1208# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X86 a_645_177# a_432_177# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X87 a_116_1944# a_116_1715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X88 a_118_n1178# a_645_n926# a_853_n926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X89 a_1803_n92# a_1512_n1208# a_1793_n1719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_1724_998# a_1511_998# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X91 a_1372_n1719# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_854_731# a_433_731# a_117_841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X93 a_1583_1590# a_1370_1590# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 a_644_1280# a_431_1280# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X95 a_117_n262# a_117_n491# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X96 a_434_n1475# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X97 a_117_612# a_646_731# a_854_731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X98 a_645_1834# a_432_1834# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X99 a_431_1280# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X100 a_1370_1590# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_116_1485# a_117_1028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X102 a_646_731# a_433_731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X103 a_1584_n616# a_1371_n616# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X104 a_432_1834# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X105 a_118_n1594# a_118_n1824# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X106 a_854_n372# a_433_n372# a_117_n491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X107 a_1792_487# a_1724_998# a_1808_27# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X108 a_1371_n616# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X109 a_1585_n1719# a_1372_n1719# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X110 a_852_1280# a_431_1280# a_117_1028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_117_n721# a_645_n926# a_853_n926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X112 a_1808_27# a_1511_998# a_1791_1590# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X113 a_117_n491# a_646_n372# a_854_n372# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X114 a_433_n2029# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X115 a_1793_n1719# a_1372_n1719# a_854_n2029# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X116 a_1792_n616# a_1371_n616# a_854_n372# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X117 a_1694_n92# a_1481_n92# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 a_432_177# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X119 a_854_n2029# a_1585_n1719# a_1793_n1719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X120 a_116_1715# a_116_1485# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X121 a_1791_1590# a_1370_1590# a_853_1834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X122 a_118_n1824# gnd gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X123 a_853_1834# a_432_1834# a_116_1715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X124 a_434_n1475# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X125 a_433_n2029# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X126 a_645_n926# a_432_n926# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X127 vref a_116_1944# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X128 a_1793_n1719# a_1725_n1208# a_1803_n92# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X129 a_854_n372# a_1584_n616# a_1792_n616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_117_841# a_117_612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X131 a_1512_n1208# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X132 a_432_n926# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X133 a_854_731# a_1584_487# a_1792_487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X134 a_1792_487# a_1371_487# a_854_731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X135 a_1371_487# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
C0 d0 gnd 2.90fF
C1 a_118_n1824# gnd 2.75fF
C2 a_854_n2029# gnd 2.79fF
C3 a_118_n1594# gnd 2.38fF
C4 a_855_n1475# gnd 2.18fF
C5 a_118_n1365# gnd 2.28fF
C6 a_118_n1178# gnd 2.49fF
C7 a_117_n721# gnd 2.23fF
C8 a_853_n926# gnd 2.52fF
C9 a_117_n491# gnd 2.38fF
C10 a_854_n372# gnd 2.45fF
C11 a_117_n262# gnd 2.28fF
C12 a_1803_n92# gnd 2.28fF
C13 a_117_n75# gnd 2.49fF
C14 a_117_382# gnd 2.23fF
C15 a_853_177# gnd 2.52fF
C16 a_117_612# gnd 2.38fF
C17 a_854_731# gnd 2.18fF
C18 a_117_841# gnd 2.28fF
C19 a_117_1028# gnd 2.49fF
C20 a_116_1485# gnd 2.23fF
C21 a_852_1280# gnd 2.52fF
C22 a_116_1715# gnd 2.38fF
C23 a_853_1834# gnd 2.38fF
C24 a_116_1944# gnd 2.22fF
C25 vdd gnd 21.37fF

Vdd vdd 0 dc 3.3
Vin1 vref 0 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5us 10us)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10us 20us)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20us 40us)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40us 80us)

.tran 0.1us 80us
.control
run
plot V(vout) V(d0) V(d1) V(d2) V(d3)
.endc
.end
