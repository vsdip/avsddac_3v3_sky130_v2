magic
tech sky130A
timestamp 1616081794
<< ndiffc >>
rect -46 16 -28 34
rect -48 -83 -30 -65
<< ndiffres >>
rect -64 34 -7 53
rect -64 16 -46 34
rect -28 31 -7 34
rect -28 16 87 31
rect -64 -7 87 16
rect 45 -43 87 -7
rect -12 -44 88 -43
rect -68 -65 88 -44
rect -68 -83 -48 -65
rect -30 -83 88 -65
rect -68 -87 88 -83
rect -68 -103 -7 -87
<< locali >>
rect -55 34 -18 43
rect -55 16 -46 34
rect -28 16 -18 34
rect -55 6 -18 16
rect -58 -65 -21 -56
rect -58 -83 -48 -65
rect -30 -83 -21 -65
rect -58 -93 -21 -83
<< labels >>
rlabel ndiffc -37 27 -37 27 1 b
rlabel ndiffc -39 -75 -39 -75 3 a
<< end >>
