* SPICE3 file created from 10bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_33949_5530# a_33567_5972# a_32976_6153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1 a_19071_4304# a_20132_3933# a_20087_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2 a_23203_n8061# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3 a_21645_1643# a_21643_1429# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4 vdd d1 a_24856_8015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5 a_16359_3223# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_35381_n3789# a_35638_n3805# a_35335_n3181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7 gnd d2 a_35588_n3385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_30922_3343# a_31175_3330# a_29909_3109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9 gnd d0 a_20442_n4047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X10 a_34195_359# a_33982_359# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X11 a_23139_2047# a_22926_2047# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 a_136_4399# a_136_4117# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X13 a_16760_7140# a_17564_6959# a_17723_7379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X14 vdd a_24962_n6733# a_24754_n6733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X15 gnd a_24578_4642# a_24370_4642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_11270_6746# a_11057_6746# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X17 a_13786_6105# a_14039_6092# a_13736_5685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_481_n9764# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X19 a_13802_2365# a_14863_1994# a_14814_2184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 a_20080_6318# a_20076_6495# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X21 a_13656_n8247# a_13870_n7331# a_13821_n7315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X22 gnd a_25958_n9908# a_25750_n9908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X23 a_16080_4005# a_16566_3789# a_16774_3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 vdd a_20337_4909# a_20129_4909# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X25 vdd a_41937_n3037# a_41729_n3037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X26 a_17614_7379# a_17401_7379# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X27 a_5987_n7783# a_5774_n7783# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X28 a_33069_n6387# a_32648_n6387# a_32378_n6021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_27393_5143# a_27180_5143# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X30 a_16169_n5434# a_16174_n5048# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X31 gnd d3 a_24653_6567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X32 a_11064_5767# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X33 vdd a_9781_n4039# a_9573_n4039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X34 a_10811_2661# a_11290_2829# a_11498_2829# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X35 a_5999_n4430# a_5786_n4430# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X36 a_2906_6786# a_3120_5664# a_3075_5677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X37 a_230_n4847# a_719_n4866# a_927_n4866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_4131_7310# a_4384_7297# a_3118_7076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 vdd d0 a_9780_n3624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X40 a_6710_3034# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X41 a_13895_n3630# a_14953_n4068# a_14904_n4052# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X42 a_1654_1095# a_1441_1095# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X43 a_3063_7637# a_3316_7624# a_2910_6609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X44 a_26924_1126# a_27413_1226# a_27621_1226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X45 gnd d0 a_25963_n8927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X46 vdd d0 a_15160_n3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X47 a_38261_4736# a_37840_4736# a_37570_4571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_23050_n7033# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_16660_n4438# a_16447_n4438# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X50 vdd d1 a_30258_n3776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X51 a_37824_8092# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_22323_4188# a_21902_4188# a_21626_4088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X53 vdd a_40907_n5744# a_40699_n5744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X54 a_32768_6153# a_32555_6153# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X55 a_37394_271# a_37285_271# a_31994_256# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X56 a_901_n9349# a_480_n9349# a_212_n8978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X57 vdd d1 a_8756_n5765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X58 a_10900_n3495# a_10905_n3109# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X59 a_32548_7132# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X60 a_5424_3611# a_5422_3397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X61 a_26921_2008# a_26926_1622# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X62 gnd d1 a_30149_6034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X63 a_29766_n8189# a_29980_n7273# a_29931_n7257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X64 gnd a_9786_n3058# a_9578_n3058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 gnd a_4403_2965# a_4195_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X66 a_14893_n6800# a_15146_n7004# a_13880_n6566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X67 a_6105_5738# a_5684_5738# a_5416_5568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X68 a_33780_5972# a_33567_5972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X69 a_30986_n8475# a_30998_n7723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X70 gnd d1 a_14044_5111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X71 a_26909_4563# a_26907_4349# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X72 a_38158_n3845# a_37945_n3845# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 vdd d4 a_13838_n6338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X74 a_5781_n5411# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X75 vdd a_24806_7595# a_24598_7595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X76 a_28666_n5055# a_28284_n5616# a_27692_n5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 a_16097_1659# a_16095_1445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X78 a_33622_5411# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_38950_n4643# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X80 a_24674_n3173# a_24769_n3797# a_24724_n3593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X81 a_41674_n3587# a_41684_n2833# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X82 a_23742_351# a_23321_351# a_23643_351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X83 a_37642_n8440# a_37644_n8341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X84 a_32375_n6997# a_32373_n6783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X85 a_2808_n10402# a_2969_n6330# a_2920_n6314# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X86 a_35272_6253# a_35529_6063# a_35226_5656# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X87 a_7510_n6077# a_7089_n6077# a_7415_n8069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X88 a_28924_330# a_28815_330# a_26733_263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X89 a_11490_4786# a_11069_4786# a_10796_5002# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X90 a_6985_1494# a_6772_1494# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X91 a_23321_351# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_39566_n8048# a_39145_n8048# a_39413_n7020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 a_38942_n6600# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X94 a_1731_n4685# a_1518_n4685# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X95 a_33085_n3866# a_32664_n3866# a_32388_n3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X96 vdd a_20422_n7964# a_20214_n7964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X97 a_24396_6757# a_24653_6567# a_24325_4655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X98 a_22411_n5403# a_23216_n5637# a_23385_n5076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X99 a_17834_5419# a_17413_5419# a_17740_5538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X100 a_13469_n10410# a_13630_n6338# a_13581_n6322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 gnd d2 a_14086_n5374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 a_39473_4426# a_39076_2501# a_39344_1473# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X103 gnd a_35554_1165# a_35346_1165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X104 a_8504_n4768# a_9565_n4603# a_9516_n4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X105 a_35331_n3369# a_35588_n3385# a_35166_n4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X106 a_10782_7343# a_10782_7061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X107 a_8407_5272# a_9468_4901# a_9419_5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X108 a_3075_5677# a_3170_6084# a_3121_6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X109 a_11278_6182# a_11065_6182# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 a_36284_6072# a_36541_5882# a_35272_6253# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X111 a_14875_n9326# a_14871_n9514# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X112 a_37570_3976# a_37575_3590# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X113 a_5491_n8743# a_5491_n8461# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X114 a_22416_n4422# a_21995_n4422# a_21729_n4236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X115 a_23531_4439# a_23134_2514# a_23390_3446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X116 a_5518_n3847# a_6007_n3866# a_6215_n3866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 a_412_4217# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 vdd d1 a_40887_n9661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X119 a_10866_n9753# a_11355_n9772# a_11563_n9772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X120 a_4223_n7961# a_4226_n7358# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X121 a_21638_2410# a_22127_2228# a_22335_2228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X122 a_23620_n5892# a_23511_n6069# a_23719_n6069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X123 a_713_n5432# a_500_n5432# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X124 a_4215_n8525# a_4227_n7773# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X125 a_41590_2372# a_41843_2359# a_40577_2138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X126 vdd a_19414_n6749# a_19206_n6749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X127 a_32390_n3466# a_32395_n3080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X128 a_18750_n10389# a_18911_n6317# a_18866_n6113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X129 a_20093_3380# a_20089_3557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X130 a_22339_832# a_21918_832# a_21645_1048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X131 a_29989_n5720# a_30246_n5736# a_29943_n5112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X132 gnd d0 a_15128_n9530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X133 a_28577_3544# a_28463_3425# a_28671_3425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X134 a_30918_3520# a_31175_3330# a_29909_3109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X135 a_902_n9764# a_1706_n9583# a_1875_n9022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_36387_n5002# a_36644_n5018# a_35378_n4580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X137 a_25636_3126# a_25893_2936# a_24624_3307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X138 a_12132_5440# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_29579_n10352# a_29740_n6280# a_29691_n6264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X140 vdd a_24578_4642# a_24370_4642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X141 a_22189_n8754# a_21976_n8754# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X142 a_617_6174# a_404_6174# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X143 a_5974_n9328# a_5761_n9328# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 a_29000_n6048# a_28579_n6048# a_28901_n5871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X145 a_832_3802# a_1637_4036# a_1806_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X146 vdd d0 a_4391_6318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X147 gnd a_24856_8015# a_24648_8015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X148 a_11594_n3480# a_11173_n3480# a_10905_n3109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X149 a_2041_4468# a_1932_4468# a_2140_4468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X150 vdd d0 a_31251_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X151 a_27284_n3837# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X152 a_19017_5664# a_19112_6071# a_19063_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 a_1801_3475# a_1429_3055# a_837_2821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 a_36371_n8731# a_36624_n8935# a_35358_n8497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X155 gnd d1 a_19333_3133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 gnd a_14064_1194# a_13856_1194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X157 a_24397_n10373# a_24347_n10389# a_24298_n10373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X158 a_40662_n3768# a_40919_n3784# a_40616_n3160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X159 a_6118_2800# a_5697_2800# a_5424_3016# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X160 a_7054_n7041# a_6841_n7041# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X161 vdd d0 a_31263_n4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X162 gnd d1 a_3492_n2845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X163 vdd a_36635_n6560# a_36427_n6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X164 a_27589_7103# a_27168_7103# a_26892_7285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X165 a_38911_3433# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_30916_3909# a_31169_3896# a_29900_4267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X167 vdd a_30243_n6712# a_30035_n6712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X168 a_22931_1066# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X169 a_38359_n4824# a_37938_n4824# a_37662_n4805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X170 a_7270_n5084# a_6849_n5084# a_7176_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X171 vdd a_4485_n6996# a_4277_n6996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X172 a_40580_n9225# a_40684_n8680# a_40635_n8664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 a_3059_7814# a_3316_7624# a_2910_6609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X174 a_16656_n5834# a_16443_n5834# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X175 a_17943_n3132# a_17888_n4160# a_18072_n5908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X176 gnd a_19340_2154# a_19132_2154# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X177 gnd a_31239_n9887# a_31031_n9887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X178 vdd d5 a_19007_n10405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X179 a_39477_6418# a_39056_6418# a_39312_7350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X180 a_37580_2397# a_37580_2115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X181 a_21709_n8153# a_22188_n8339# a_22396_n8339# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X182 a_37639_n9917# a_41643_n9879# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X183 vdd d0 a_41827_4880# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X184 a_29892_6224# a_30953_5853# a_30908_5866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X185 a_11367_n7812# a_11154_n7812# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X186 a_20100_2401# a_20353_2388# a_19087_2167# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X187 a_16863_n5419# a_17668_n5653# a_17837_n5092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X188 a_32299_2136# a_32788_2236# a_32996_2236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X189 a_26899_6306# a_26899_6024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X190 a_11583_n5855# a_11162_n5855# a_10886_n5836# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X191 vdd d1 a_30149_6034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X192 a_30909_5062# a_30917_4324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X193 a_22302_7690# a_23107_7924# a_23276_7482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X194 a_33001_1255# a_32580_1255# a_32304_1155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X195 a_32279_6335# a_32279_6053# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X196 a_27704_n3422# a_27283_n3422# a_27015_n3051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X197 a_12642_n7070# a_12221_n7070# a_12543_n6893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X198 gnd a_9685_3359# a_9477_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_21700_n8735# a_21700_n8453# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 vdd a_3455_n9703# a_3247_n9703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X201 gnd d0 a_41822_5861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X202 a_13787_5301# a_14848_4930# a_14803_4943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X203 a_27603_3752# a_27182_3752# a_26909_3968# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X204 a_22120_3207# a_21907_3207# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X205 a_19164_n5569# a_19417_n5773# a_19114_n5149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 a_24713_n4760# a_25774_n4595# a_25729_n4391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X207 a_5503_n6501# a_5992_n6802# a_6200_n6802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X208 vdd d1 a_14044_5111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X209 a_23380_n4899# a_23271_n5076# a_23479_n5076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X210 a_1801_3475# a_1692_3475# a_1900_3475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X211 a_1857_2543# a_1644_2543# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X212 a_33937_7490# a_33555_7932# a_32963_7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X213 a_18072_n5908# a_17963_n6085# a_18171_n6085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X214 a_21734_n3072# a_22215_n3443# a_22423_n3443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X215 a_13782_6282# a_14843_5911# a_14794_6101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X216 a_33877_n5645# a_33664_n5645# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X217 a_16786_1829# a_17591_2063# a_17760_1621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X218 a_17728_7498# a_17614_7379# a_17822_7379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X219 a_9527_n3420# a_9523_n3608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X220 a_14788_7495# a_14791_6903# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X221 gnd a_8664_5082# a_8456_5082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 a_33072_n5411# a_32651_n5411# a_32383_n5040# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X223 a_16060_7922# a_16546_7706# a_16754_7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X224 vdd d2 a_40837_n9241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X225 a_35269_7055# a_35522_7042# a_35210_7793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X226 a_20174_n6779# a_20427_n6983# a_19161_n6545# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X227 a_28815_330# a_28602_330# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X228 a_41590_2372# a_41586_2549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X229 a_27477_n7754# a_27264_n7754# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X230 a_8520_n2620# a_9578_n3058# a_9533_n2854# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X231 a_17421_3462# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X232 a_12365_1523# a_12152_1523# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X233 a_21608_7906# a_22094_7690# a_22302_7690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X234 a_20848_n805# a_21446_n10615# a_21397_n10599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X235 a_16184_n2592# a_16186_n2493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X236 gnd d0 a_31174_2915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X237 a_27693_n5797# a_27272_n5797# a_26996_n5778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X238 vdd a_35554_1165# a_35346_1165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X239 a_16149_n9946# a_16147_n9732# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X240 a_3075_5677# a_3170_6084# a_3125_6097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X241 gnd a_3437_n3406# a_3229_n3406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X242 a_36385_n5380# a_36638_n5584# a_35369_n5749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X243 a_24697_n8489# a_25755_n8927# a_25706_n8911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X244 a_13891_n3818# a_14952_n3653# a_14907_n3449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X245 a_39314_n6843# a_38942_n6600# a_38350_n6366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 gnd a_31181_1936# a_30973_1936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 a_22303_8105# a_21882_8105# a_21606_8005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 a_32862_n6802# a_32649_n6802# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X249 a_3113_8057# a_3366_8044# a_3063_7637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X250 a_38891_7350# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X251 gnd a_25962_n8512# a_25754_n8512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X252 a_1887_n7062# a_1505_n7623# a_913_n7389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X253 a_40545_8015# a_41603_8236# a_41554_8426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X254 vdd a_36529_7842# a_36321_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X255 a_219_n7404# a_705_n7389# a_913_n7389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X256 a_8453_n5141# a_8548_n5765# a_8503_n5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X257 a_11511_1284# a_11090_1284# a_10814_1184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X258 a_41582_2936# a_41578_3113# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X259 a_24573_3691# a_24826_3678# a_24420_2663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 a_35150_n8030# a_35348_n9262# a_35303_n9058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X261 a_5991_n6387# a_5778_n6387# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X262 a_33069_n6387# a_33874_n6621# a_34033_n6864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X263 a_40612_n3348# a_40869_n3364# a_40447_n4280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X264 gnd d0 a_25906_1391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X265 a_29850_3847# a_29954_3096# a_29909_3109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X266 a_26995_n6968# a_27476_n7339# a_27684_n7339# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X267 vdd a_9785_n2643# a_9577_n2643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X268 a_32996_2236# a_33800_2055# a_33969_1613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X269 a_33932_7371# a_33560_6951# a_32969_7132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X270 a_10880_n8190# a_10878_n7793# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X271 a_21645_1048# a_21652_847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X272 a_1548_n9022# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X273 vdd d0 a_41919_n5563# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X274 a_16787_2244# a_16366_2244# a_16090_2144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 a_41655_n7919# a_41912_n7935# a_40646_n7497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X276 a_12447_7519# a_12065_7961# a_11473_7727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X277 a_16161_n8169# a_16640_n8355# a_16848_n8355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X278 a_14883_n7554# a_14893_n6800# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X279 a_35370_n6537# a_35623_n6741# a_35311_n7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 a_6183_n9743# a_5762_n9743# a_5486_n9442# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X281 gnd a_4479_n7562# a_4271_n7562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X282 a_26926_1622# a_27407_1792# a_27615_1792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X283 a_16849_n8770# a_16428_n8770# a_16152_n8751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X284 a_3134_3336# a_4195_2965# a_4146_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 gnd a_19007_n10405# a_18799_n10405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X286 a_23132_3026# a_22919_3026# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X287 a_25627_5887# a_25623_6064# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X288 a_13744_3728# a_13997_3715# a_13591_2700# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X289 a_27271_n5382# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 a_37565_5051# a_38054_5151# a_38262_5151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X291 gnd d3 a_8464_2658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X292 a_13779_7084# a_14032_7071# a_13720_7822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X293 a_32363_n8957# a_32844_n9328# a_33052_n9328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X294 vdd a_24856_8015# a_24648_8015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X295 gnd d2 a_35479_5643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_1786_7511# a_1404_7953# a_813_8134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X297 a_6965_5411# a_6752_5411# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X298 a_205_n9463# a_694_n9764# a_902_n9764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X299 a_19017_5664# a_19112_6071# a_19067_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X300 a_27010_n4215# a_27489_n4401# a_27697_n4401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X301 vdd d1 a_19333_3133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X302 a_23003_n5637# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X303 a_23221_n4656# a_23008_n4656# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X304 a_5488_n9938# a_9749_n9916# a_8483_n9478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X305 a_2140_4468# a_2044_380# a_2252_380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X306 a_41668_n4981# a_41925_n4997# a_40659_n4559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X307 a_19055_8044# a_19308_8031# a_19005_7624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X308 a_17849_n3132# a_17467_n3693# a_16876_n3874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X309 a_5399_7914# a_5404_7528# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X310 a_7421_4447# a_7000_4447# a_7326_6439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X311 a_14823_1026# a_14819_1203# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X312 a_19114_n5149# a_19367_n5353# a_18961_n4121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X313 a_12372_n8610# a_12159_n8610# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X314 a_38338_n8326# a_37917_n8326# a_37651_n8140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X315 a_5409_6053# a_5898_6153# a_6106_6153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X316 a_35369_n5749# a_36430_n5584# a_36385_n5380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X317 vdd a_19340_2154# a_19132_2154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X318 vdd a_15039_7871# a_14831_7871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X319 a_17401_7379# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X320 a_19055_8044# a_20113_8265# a_20064_8455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X321 a_27180_5143# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X322 a_3222_n5582# a_4280_n6020# a_4235_n5816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X323 a_24396_6757# a_24610_5635# a_24561_5825# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X324 a_5794_n3866# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 a_41594_976# a_41847_963# a_40578_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X326 a_32761_7132# a_32548_7132# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X327 a_1738_n3706# a_1525_n3706# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X328 a_41651_n8295# a_41647_n8483# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X329 gnd d2 a_40760_5622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X330 gnd a_20341_4348# a_20133_4348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X331 a_32876_n3451# a_32663_n3451# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X332 a_32555_6153# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X333 a_1493_n9583# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X334 a_7094_1494# a_6722_1074# a_6131_1255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X335 a_128_6356# a_617_6174# a_825_6174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_17812_n8832# a_17440_n8589# a_16848_n8355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 a_6012_n2885# a_5799_n2885# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X338 a_162_876# a_641_861# a_849_861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X339 a_29943_n5112# a_30196_n5316# a_29790_n4084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 a_34041_n4907# a_33932_n5084# a_34140_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X341 gnd d2 a_13989_5672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X342 vdd a_3252_n8255# a_3044_n8255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X343 vdd a_8664_5082# a_8456_5082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X344 a_18961_n4121# a_19214_n4325# a_18862_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X345 a_22429_n2877# a_22008_n2877# a_21732_n2576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X346 a_1902_n2968# a_1530_n2725# a_939_n2906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X347 a_31885_256# a_31672_256# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X348 a_7181_3454# a_6760_3454# a_7087_3573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X349 a_5424_3016# a_5431_2632# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X350 a_27464_n9299# a_27251_n9299# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X351 a_8300_n4113# a_8498_n5345# a_8453_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X352 a_6219_n2470# a_7024_n2704# a_7183_n2947# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X353 a_1459_7392# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X354 a_36302_3372# a_36298_3549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X355 a_39069_3994# a_38856_3994# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X356 a_35265_7232# a_35522_7042# a_35210_7793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X357 gnd a_14044_5111# a_13836_5111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X358 a_726_n3887# a_513_n3887# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X359 vdd d0 a_36567_1399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X360 a_824_5759# a_1629_5993# a_1798_5551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X361 gnd a_25889_4332# a_25681_4332# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X362 a_38138_n7762# a_37925_n7762# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X363 a_21907_3207# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X364 a_8520_n2620# a_8773_n2824# a_8461_n3369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_22911_4983# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X366 a_30896_7826# a_31149_7813# a_29880_8184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X367 a_33843_3454# a_33630_3454# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X368 a_17675_n4160# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X369 a_481_n9764# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X370 a_19172_n3797# a_20233_n3632# a_20188_n3428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X371 a_6772_1494# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 a_32775_3781# a_32562_3781# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X373 vdd a_25975_n6967# a_25767_n6967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X374 a_20104_1005# a_20357_992# a_19088_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 a_11271_7161# a_11058_7161# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X376 a_21975_n8339# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X377 a_3109_8234# a_3366_8044# a_3063_7637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X378 a_39193_n8980# a_38980_n8980# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X379 a_40545_8015# a_41603_8236# a_41558_8249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X380 a_39054_6930# a_38841_6930# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X381 a_17660_n7610# a_17447_n7610# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X382 a_17455_n5653# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X383 a_30001_n3760# a_31062_n3595# a_31013_n3579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X384 a_24640_1170# a_25698_1391# a_25653_1404# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X385 a_11153_n7397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X386 a_16443_n5834# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X387 a_11065_6182# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 a_38056_3760# a_37843_3760# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 a_12607_n4181# a_12394_n4181# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X390 a_10802_3426# a_11291_3244# a_11499_3244# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X391 a_3148_n9267# a_3252_n8722# a_3207_n8518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X392 a_38351_n6781# a_37930_n6781# a_37654_n6762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X393 a_3152_n9079# a_3405_n9283# a_2999_n8051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X394 vdd a_20414_n8528# a_20206_n8528# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X395 a_36403_n2854# a_36656_n3058# a_35390_n2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X396 a_41666_n5359# a_41919_n5563# a_40650_n5728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 vdd a_24945_n9674# a_24737_n9674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X398 a_5779_n6802# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X399 a_21625_5560# a_21623_5346# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X400 a_1781_7392# a_1672_7392# a_1880_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X401 a_2910_6609# a_3163_6596# a_2835_4684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X402 gnd a_31243_n8491# a_31035_n8491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X403 a_22002_n3443# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X404 a_22220_n2462# a_22007_n2462# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X405 a_27375_7669# a_27162_7669# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X406 a_13740_3905# a_13997_3715# a_13591_2700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X407 a_13775_7261# a_14032_7071# a_13720_7822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X408 a_610_7153# a_397_7153# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X409 a_40431_n8009# a_40629_n9241# a_40584_n9037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X410 a_11371_n6416# a_11158_n6416# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X411 vdd d0 a_15077_1428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X412 a_20177_n5803# a_20430_n6007# a_19164_n5569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X413 a_22099_6709# a_21886_6709# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X414 vdd d2 a_35479_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X415 gnd d2 a_8617_3686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X416 a_34172_n6077# a_33959_n6077# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X417 a_7094_1494# a_6985_1494# a_7193_1494# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X418 a_36298_3549# a_36301_2957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X419 a_27010_n4215# a_27008_n3818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X420 a_32568_3215# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X421 vdd a_14098_n3414# a_13890_n3414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X422 a_19051_8221# a_19308_8031# a_19005_7624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X423 a_40651_n6516# a_40904_n6720# a_40592_n7265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 a_404_6174# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X425 a_9423_4914# a_9419_5091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X426 a_27001_n4515# a_27003_n4416# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X427 a_16546_7706# a_16333_7706# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_141_3136# a_630_3236# a_838_3236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X429 a_14892_n6012# a_15149_n6028# a_13883_n5590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X430 vdd d0 a_4383_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X431 a_25736_n3412# a_25732_n3600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X432 a_40546_7211# a_41607_6840# a_41558_7030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_205_n9745# a_205_n9463# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X434 a_19055_8044# a_20113_8265# a_20068_8278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X435 a_17868_n8077# a_17655_n8077# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X436 a_12454_n3153# a_12241_n3153# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X437 gnd a_19333_3133# a_19125_3133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X438 a_38950_n4643# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X439 a_24396_6757# a_24610_5635# a_24565_5648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X440 a_23377_n7033# a_22995_n7594# a_22403_n7360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 a_25621_7281# a_25874_7268# a_24608_7047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X442 a_11491_5201# a_11070_5201# a_10794_5101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X443 a_33085_n3866# a_32664_n3866# a_32388_n3565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X444 a_10868_n9967# a_15129_n9945# a_13863_n9507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X445 vdd a_35631_n4784# a_35423_n4784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X446 vdd d2 a_40760_5622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X447 a_33661_n6621# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X448 a_18852_6596# a_19105_6583# a_18777_4671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X449 a_22412_n5818# a_23216_n5637# a_23385_n5076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X450 vdd a_25989_n3616# a_25781_n3616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X451 a_4146_4374# a_4399_4361# a_3133_4140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X452 a_27481_n6358# a_27268_n6358# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X453 a_24623_4111# a_24876_4098# a_24573_3691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X454 a_16636_n9751# a_16423_n9751# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X455 vdd d0 a_9768_n5584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X456 a_37587_1035# a_38073_819# a_38281_819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X457 a_39344_1473# a_38923_1473# a_39245_1473# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X458 vdd a_15140_n7570# a_14932_n7570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X459 a_40650_n5728# a_41711_n5563# a_41666_n5359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X460 a_25653_1404# a_25649_1581# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X461 a_15660_n10477# a_15917_n10493# a_10399_n10484# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X462 a_38276_1800# a_37855_1800# a_37587_1630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X463 vdd a_41827_4880# a_41619_4880# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X464 a_34120_n9001# a_34077_n8069# a_34285_n8069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X465 a_4145_3959# a_4141_4136# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X466 a_3215_n6746# a_4276_n6581# a_4227_n6565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X467 a_11174_n3895# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_6118_2800# a_6923_3034# a_7082_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X469 gnd a_25969_n7533# a_25761_n7533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X470 a_8445_n7098# a_8540_n7722# a_8495_n7518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X471 vdd d2 a_13989_5672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X472 a_16179_n3573# a_16181_n3474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X473 a_39143_n8560# a_38930_n8560# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X474 a_10903_n2613# a_11392_n2914# a_11600_n2914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X475 gnd a_41822_5861# a_41614_5861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 a_16779_2808# a_17584_3042# a_17743_3462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X477 a_41648_n8898# a_41651_n8295# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X478 a_713_n5432# a_500_n5432# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 a_27595_5709# a_27174_5709# a_26906_5539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 a_28564_n3095# a_28351_n3095# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X481 a_25616_8262# a_26887_8266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X482 a_5402_7314# a_5402_7032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X483 a_11078_3244# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X484 vdd a_14044_5111# a_13836_5111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X485 a_13587_2877# a_13844_2687# a_13492_4869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X486 gnd d1 a_35529_6063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X487 a_830_5193# a_409_5193# a_133_5375# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X488 a_6905_6439# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X489 vdd a_25889_4332# a_25681_4332# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X490 a_27620_811# a_27199_811# a_26926_1027# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X491 a_32361_n8743# a_32361_n8461# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X492 gnd d1 a_35643_n2824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X493 gnd a_19030_4658# a_18822_4658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_22189_n8754# a_21976_n8754# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X495 a_829_4778# a_408_4778# a_135_4994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X496 a_8445_n7098# a_8698_n7302# a_8276_n8218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X497 a_29909_3109# a_30967_3330# a_30918_3520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X498 a_24700_n7698# a_24957_n7714# a_24654_n7090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X499 gnd d2 a_24907_n7294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X500 a_12152_1523# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 gnd a_31174_2915# a_30966_2915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X502 a_32636_n8347# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X503 a_30892_8003# a_30902_7260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X504 a_20076_6495# a_20333_6305# a_19067_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X505 a_27284_n3837# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X506 a_37550_7893# a_37555_7507# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X507 a_24565_5648# a_24660_6055# a_24611_6245# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X508 a_18866_n6113# a_18986_n8242# a_18941_n8038# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X509 a_39378_n4131# a_39165_n4131# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X510 a_10811_2661# a_10809_2447# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X511 a_27013_n2555# a_27502_n2856# a_27710_n2856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X512 a_21638_2128# a_21640_2029# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X513 a_6119_3215# a_5698_3215# a_5422_3115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X514 gnd d0 a_15060_4369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X515 a_38359_n4824# a_37938_n4824# a_37662_n4523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X516 a_7074_5411# a_6702_4991# a_6111_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X517 vdd a_31256_n6946# a_31048_n6946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X518 a_23119_5964# a_22906_5964# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 a_16780_3223# a_16359_3223# a_16083_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X520 a_22216_n3858# a_22003_n3858# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_25649_1581# a_25652_989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X522 vdd a_8667_4106# a_8459_4106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X523 a_33719_n5084# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X524 a_21918_832# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X525 a_37150_n10448# a_37407_n10464# a_31889_n10455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X526 a_11367_n7812# a_11154_n7812# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 gnd a_25906_1391# a_25698_1391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_5678_7132# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X529 a_16864_n5834# a_17668_n5653# a_17837_n5092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X530 a_32381_n4544# a_32870_n4845# a_33078_n4845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X531 a_38256_5717# a_37835_5717# a_37562_5933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X532 gnd d1 a_14039_6092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X533 a_901_n9349# a_480_n9349# a_207_n9364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X534 a_11583_n5855# a_11162_n5855# a_10886_n5554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X535 a_6811_n2704# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X536 a_23271_n5076# a_23058_n5076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X537 vdd d2 a_8617_3686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X538 gnd a_31182_2351# a_30974_2351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X539 a_41684_n2833# a_41937_n3037# a_40671_n2599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X540 vdd a_30226_n9653# a_30018_n9653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X541 gnd d0 a_25989_n3616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 vdd a_4468_n9937# a_4260_n9937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X543 a_7270_n5084# a_7227_n4152# a_7411_n5900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X544 vdd a_36624_n8935# a_36416_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X545 a_5503_n6783# a_5992_n6802# a_6200_n6802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X546 gnd a_8464_2658# a_8256_2658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X547 a_36298_3549# a_36555_3359# a_35289_3138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X548 a_4243_n4044# a_4500_n4060# a_3234_n3622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X549 a_23531_4439# a_23422_4439# a_23630_4439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X550 a_13875_n7547# a_14128_n7751# a_13825_n7127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_3234_n3622# a_4292_n4060# a_4243_n4044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 a_21729_n3458# a_22215_n3443# a_22423_n3443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X553 a_6752_5411# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X554 a_8276_n8218# a_8490_n7302# a_8445_n7098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X555 gnd a_14136_n5794# a_13928_n5794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X556 vdd a_19333_3133# a_19125_3133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X557 a_17576_4999# a_17363_4999# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X558 a_26489_n10440# a_29628_n10368# a_29000_n6048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X559 a_5897_5738# a_5684_5738# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X560 a_10880_n7412# a_11366_n7397# a_11574_n7397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_34192_4447# a_33795_2522# a_34051_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X562 a_27477_n7754# a_27264_n7754# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_39104_7350# a_38891_7350# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X564 a_17963_n6085# a_17750_n6085# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X565 a_24549_7785# a_24806_7595# a_24400_6580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X566 a_138_4018# a_143_3632# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X567 a_9501_n8731# a_9497_n8919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X568 a_18848_6773# a_19105_6583# a_18777_4671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X569 a_4142_4551# a_4399_4361# a_3133_4140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X570 vdd d0 a_25886_5308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X571 a_8205_n6105# a_8458_n6309# a_8089_n10381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X572 a_36272_8032# a_36282_7289# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X573 a_32294_3016# a_32780_2800# a_32988_2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X574 a_37924_n7347# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X575 a_38142_n6366# a_37929_n6366# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X576 a_36398_n2627# a_36655_n2643# a_35386_n2808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X577 vdd a_40497_n10376# a_40289_n10376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X578 gnd a_30208_n3356# a_30000_n3356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_30006_n2779# a_30263_n2795# a_29951_n3340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X580 a_19152_n7714# a_19409_n7730# a_19106_n7106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X581 a_8414_4119# a_9472_4340# a_9423_4530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X582 vdd d1 a_24888_2138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X583 a_22404_n7775# a_21983_n7775# a_21707_n7756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X584 a_23162_7363# a_22949_7363# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X585 a_25725_n4579# a_25737_n3827# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X586 a_31006_n5766# a_31259_n5970# a_29993_n5532# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_24658_n5321# a_24915_n5337# a_24509_n4105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X588 a_21613_6925# a_22099_6709# a_22307_6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X589 a_7188_n3124# a_7074_n3124# a_7282_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X590 a_16563_4765# a_16350_4765# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X591 a_141_3136# a_143_3037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X592 a_16760_7140# a_16339_7140# a_16063_7322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X593 a_33070_n6802# a_33874_n6621# a_34033_n6864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X594 a_28408_3986# a_28195_3986# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X595 a_23291_3446# a_23182_3446# a_23390_3446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X596 a_7004_n6621# a_6791_n6621# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X597 a_3164_n7119# a_3259_n7743# a_3214_n7539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X598 vdd d1 a_35529_6063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X599 vdd a_20421_n7549# a_20213_n7549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X600 vdd d0 a_25900_1957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X601 a_10799_4026# a_11285_3810# a_11493_3810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X602 gnd d1 a_8667_4106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X603 a_37669_n3544# a_38158_n3845# a_38366_n3845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X604 a_21623_5064# a_21625_4965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X605 a_16154_n8370# a_16640_n8355# a_16848_n8355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 a_9511_n5568# a_9521_n4814# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X607 vdd d1 a_19422_n4792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X608 gnd a_40919_n3784# a_40711_n3784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X609 vdd a_10656_n10500# a_10448_n10500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X610 a_37285_271# a_37072_271# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X611 vdd d6 a_26746_n10456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X612 gnd d1 a_8768_n3805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X613 vdd a_36567_1399# a_36359_1399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X614 a_29909_3109# a_30967_3330# a_30922_3343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X615 a_5974_n9328# a_5761_n9328# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X616 gnd d1 a_14116_n9711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X617 a_3125_6097# a_4183_6318# a_4138_6331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X618 a_25706_n8911# a_25963_n8927# a_24697_n8489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X619 a_205_n9745# a_694_n9764# a_902_n9764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X620 a_8508_n4580# a_9566_n5018# a_9517_n5002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X621 a_27003_n4416# a_27489_n4401# a_27697_n4401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X622 a_24565_5648# a_24660_6055# a_24615_6068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X623 a_9509_n6959# a_9766_n6975# a_8500_n6537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X624 a_33630_3454# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X625 a_23003_n5637# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 a_23221_n4656# a_23008_n4656# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_32562_3781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X628 vdd a_41830_3904# a_41622_3904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X629 a_26978_n9314# a_26983_n8928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X630 a_8089_n10381# a_8250_n6309# a_8205_n6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X631 a_148_2439# a_148_2157# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X632 vdd d0 a_9672_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X633 a_35272_6253# a_36333_5882# a_36284_6072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_16181_n3474# a_16667_n3459# a_16875_n3459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X635 a_24603_8028# a_24856_8015# a_24553_7608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X636 gnd d0 a_36554_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X637 a_143_3632# a_624_3802# a_832_3802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X638 a_37550_7893# a_38036_7677# a_38244_7677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X639 a_33864_n8069# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X640 vdd a_5256_n10485# a_5048_n10485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X641 a_17799_2530# a_17586_2530# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X642 a_14896_n4616# a_15153_n4632# a_13884_n4797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X643 a_13825_n7127# a_14078_n7331# a_13656_n8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X644 gnd d2 a_30188_n7273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X645 a_29993_n5532# a_31051_n5970# a_31006_n5766# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X646 a_39175_n2683# a_38962_n2683# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X647 a_32281_6549# a_32760_6717# a_32968_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X648 a_135_4994# a_138_4613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X649 vdd d0 a_20346_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X650 a_21881_7690# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X651 a_21899_5164# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X652 gnd a_14086_n5374# a_13878_n5374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 gnd a_36561_1965# a_36353_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X654 a_23382_5403# a_22961_5403# a_23288_5522# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X655 a_10866_n9753# a_10866_n9471# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X656 a_1738_n3706# a_1525_n3706# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X657 a_27678_n8733# a_27257_n8733# a_26981_n8714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X658 a_33000_840# a_32579_840# a_32306_1056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X659 vdd a_31182_2351# a_30974_2351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X660 vdd a_41899_n9480# a_41691_n9480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X661 a_34053_n2947# a_33681_n2704# a_33090_n2885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X662 a_24624_3307# a_25685_2936# a_25636_3126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X663 a_27162_7669# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_16640_n8355# a_16427_n8355# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X665 a_24410_n6285# a_24667_n6301# a_24298_n10373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X666 a_32996_2236# a_32575_2236# a_32299_2418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X667 a_1837_6460# a_1624_6460# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X668 vdd a_40887_n9661# a_40679_n9661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X669 a_25717_n7744# a_25970_n7948# a_24704_n7510# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X670 gnd d0 a_4473_n8956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 a_37150_n10448# a_40289_n10376# a_39661_n6056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X672 a_15795_300# a_15582_300# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X673 a_37567_5547# a_37565_5333# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X674 a_21625_4965# a_21628_4584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X675 a_19102_n7294# a_19359_n7310# a_18937_n8226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X676 vdd a_15077_1428# a_14869_1428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X677 a_35331_n3369# a_35435_n2824# a_35386_n2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X678 gnd d0 a_36562_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 a_4246_n3441# a_4499_n3645# a_3230_n3810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X680 a_10784_7557# a_11265_7727# a_11473_7727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X681 a_37553_7293# a_37553_7011# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X682 gnd d0 a_31169_3896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X683 a_26887_7984# a_26889_7885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X684 a_1902_n2968# a_1530_n2725# a_938_n2491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X685 a_28911_4418# a_28490_4418# a_28816_6410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X686 a_6220_n2885# a_7024_n2704# a_7183_n2947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X687 a_8479_n9666# a_9540_n9501# a_9491_n9485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X688 vdd a_32146_n10471# a_31938_n10471# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X689 a_16333_7706# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 a_14907_n3449# a_15160_n3653# a_13891_n3818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X691 a_26899_6024# a_27388_6124# a_27596_6124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X692 a_33932_n5084# a_33719_n5084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X693 a_17723_n5092# a_17510_n5092# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X694 gnd d0 a_15064_2973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X695 a_31005_n5351# a_31001_n5539# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X696 a_38138_n7762# a_37925_n7762# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X697 a_35234_3699# a_35487_3686# a_35081_2671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X698 gnd a_13933_n4346# a_13725_n4346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X699 a_22391_n9320# a_21970_n9320# a_21702_n8949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X700 a_37671_n4223# a_37669_n3826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X701 a_24635_2151# a_25693_2372# a_25644_2562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X702 gnd d0 a_9753_n8520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 a_8414_4119# a_9472_4340# a_9427_4353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X704 a_37662_n4523# a_37664_n4424# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X705 a_518_n2906# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X706 gnd a_4504_n2664# a_4296_n2664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X707 gnd a_15071_1994# a_14863_1994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 gnd a_40869_n3364# a_40661_n3364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X709 a_850_1276# a_1654_1095# a_1813_1515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X710 a_16095_1445# a_16095_1163# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X711 a_36397_n3420# a_36393_n3608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X712 a_17455_n5653# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X713 a_32657_n4845# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X714 a_17779_6447# a_17566_6447# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X715 gnd d2 a_14066_n9291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X716 a_28584_1465# a_28212_1045# a_27621_1226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X717 a_25704_n9289# a_25957_n9493# a_24688_n9658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X718 a_41563_7268# a_41559_7445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X719 gnd d2 a_24818_5635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X720 a_16443_n5834# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X721 a_37659_n5405# a_38145_n5390# a_38353_n5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X722 a_12166_n7631# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X723 a_13845_n3210# a_13940_n3834# a_13895_n3630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X724 gnd d0 a_31275_n2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 vdd d2 a_8597_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X726 a_11506_2265# a_11085_2265# a_10809_2447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X727 a_16759_6725# a_16338_6725# a_16072_6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 a_29919_n9217# a_30023_n8672# a_29978_n8468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X729 a_21397_n10599# a_31938_n10471# a_31889_n10455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 vdd a_19214_n4325# a_19006_n4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X731 a_3207_n8518# a_4265_n8956# a_4220_n8752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X732 a_7014_n4152# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X733 a_5779_n6802# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X734 a_5511_n4826# a_5511_n4544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X735 a_28671_3425# a_28250_3425# a_28577_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X736 a_28760_n5055# a_28717_n4123# a_28901_n5871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X737 a_7250_n9001# a_6829_n9001# a_7151_n8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 a_4243_n4044# a_4246_n3441# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X739 a_22002_n3443# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 a_22220_n2462# a_22007_n2462# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X741 a_40491_7772# a_40595_7021# a_40546_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X742 a_3230_n3810# a_4291_n3645# a_4246_n3441# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X743 a_33969_1613# a_33587_2055# a_32995_1821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X744 a_6740_7371# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X745 gnd a_41925_n4997# a_41717_n4997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X746 vdd a_8773_n2824# a_8565_n2824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X747 a_1684_5432# a_1471_5432# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X748 a_938_n2491# a_517_n2491# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X749 a_23127_4007# a_22914_4007# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X750 a_9509_n6959# a_9512_n6356# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X751 a_11371_n6416# a_11158_n6416# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X752 a_11166_n4459# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X753 gnd a_9769_n5999# a_9561_n5999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X754 a_35057_6765# a_35271_5643# a_35222_5833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X755 a_18862_n6301# a_19119_n6317# a_18750_n10389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X756 a_29955_n3152# a_30050_n3776# a_30005_n3572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X757 a_37585_1134# a_37587_1035# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X758 gnd d3 a_24762_n4309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X759 a_11290_2829# a_11077_2829# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X760 a_32976_6153# a_33780_5972# a_33949_5530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X761 a_13720_7822# a_13824_7071# a_13775_7261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X762 vdd d0 a_36636_n6975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X763 a_24599_8205# a_24856_8015# a_24553_7608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X764 vdd a_4472_n8541# a_4264_n8541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X765 gnd a_9671_5882# a_9463_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X766 a_14804_5358# a_14800_5535# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X767 a_28276_n7573# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X768 gnd d3 a_13913_n8263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X769 a_22203_n5403# a_21990_n5403# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X770 a_41590_1153# a_41847_963# a_40578_1334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X771 a_36276_7855# a_36529_7842# a_35260_8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X772 a_27413_1226# a_27200_1226# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 a_8372_1916# a_8476_1165# a_8427_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X774 a_28905_n8040# a_28792_n6048# a_29000_n6048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 a_23112_6943# a_22899_6943# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_23365_n8993# a_23251_n8993# a_23459_n8993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X777 a_14897_n5031# a_14900_n4428# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X778 gnd d0 a_4484_n6581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X779 a_20996_141# a_31672_256# a_31994_256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X780 a_40642_n7685# a_40899_n7701# a_40596_n7077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X781 a_6861_n3124# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_30893_8418# a_31150_8228# a_29884_8007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X783 a_927_n4866# a_506_n4866# a_230_n4847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X784 a_25710_n8723# a_25706_n8911# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X785 a_22114_3773# a_21901_3773# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 gnd d1 a_3472_n6762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X787 a_33661_n6621# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X788 a_12795_n8098# a_12374_n8098# a_12630_n9030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X789 a_38339_n8741# a_37918_n8741# a_37642_n8722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X790 a_32756_8113# a_32543_8113# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X791 a_28388_7903# a_28175_7903# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X792 a_24400_6580# a_24653_6567# a_24325_4655# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X793 a_19157_n6733# a_20218_n6568# a_20173_n6364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X794 a_41559_7445# a_41562_6853# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X795 a_16636_n9751# a_16423_n9751# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X796 a_38163_n2864# a_37950_n2864# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X797 a_3019_n4134# a_3217_n5366# a_3168_n5350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X798 vdd d2 a_40780_1705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X799 gnd d1 a_8647_8023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X800 a_20177_n4595# a_20434_n4611# a_19165_n4776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X801 a_7188_n3124# a_6806_n3685# a_6215_n3866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X802 a_28661_n4878# a_28289_n4635# a_27698_n4816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X803 a_12479_1642# a_12097_2084# a_11505_1850# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X804 a_12536_n9030# a_12154_n9591# a_11563_n9772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X805 a_41667_n5774# a_41663_n5962# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X806 a_20853_n686# a_20739_n805# vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 a_29986_n6696# a_31047_n6531# a_30998_n6515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X808 a_20068_7059# a_20080_6318# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X809 a_34304_359# a_35031_4650# a_34982_4840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X810 a_230_n4565# a_232_n4466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X811 vdd d0 a_36562_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X812 a_31010_n4370# a_31263_n4574# a_29994_n4739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 a_21902_4188# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X814 a_8495_n7518# a_9553_n7956# a_9508_n7752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X815 a_6093_7698# a_5672_7698# a_5399_7914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X816 a_10903_n2895# a_11392_n2914# a_11600_n2914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_6935_1074# a_6722_1074# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X818 a_13813_n9087# a_13908_n9711# a_13859_n9695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X819 a_8344_7616# a_8597_7603# a_8191_6588# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X820 a_21717_n6013# a_21715_n5799# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X821 a_19144_n9486# a_19397_n9690# a_19094_n9066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X822 a_5890_6717# a_5677_6717# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X823 a_25720_n5560# a_25730_n4806# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X824 a_13676_n4330# a_13890_n3414# a_13845_n3210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X825 a_19126_n3189# a_19221_n3813# a_19172_n3797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X826 gnd d0 a_41931_n3603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X827 a_35230_3876# a_35487_3686# a_35081_2671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X828 a_16454_n3459# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X829 a_9438_1978# a_9434_2155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X830 a_38256_5717# a_39061_5951# a_39230_5509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X831 a_6973_3454# a_6760_3454# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X832 a_14786_7884# a_15039_7871# a_13770_8242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 a_3198_n9687# a_4259_n9522# a_4210_n9506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X834 a_17363_4999# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X835 a_25632_4522# a_25635_3930# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X836 a_5684_5738# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 gnd a_8741_n8701# a_8533_n8701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X838 a_24635_2151# a_25693_2372# a_25648_2385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X839 a_38074_1234# a_37861_1234# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X840 gnd d0 a_4415_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 a_14800_5535# a_14803_4943# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X842 a_7151_n8824# a_6779_n8581# a_6187_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X843 a_17824_n6872# a_17715_n7049# a_17923_n7049# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X844 a_25636_4345# a_25889_4332# a_24623_4111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 vdd d1 a_24881_3117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X846 a_28393_6922# a_28180_6922# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X847 a_812_7719# a_391_7719# a_123_7549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X848 a_32636_n8347# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X849 gnd d0 a_4391_6318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X850 a_38265_4175# a_39069_3994# a_39238_3552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 gnd a_19402_n8709# a_19194_n8709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X852 a_20188_n3428# a_20441_n3632# a_19172_n3797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 a_11266_8142# a_11053_8142# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X854 a_29901_5066# a_30154_5053# a_29842_5804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X855 vdd d2 a_24818_5635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X856 a_27013_n2837# a_27502_n2856# a_27710_n2856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 a_16672_n2478# a_16459_n2478# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_28187_5943# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X859 vdd d0 a_15134_n8964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X860 a_22334_1813# a_21913_1813# a_21645_1643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X861 vdd d0 a_31154_6832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X862 a_27608_2771# a_28413_3005# a_28572_3425# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X863 a_1880_7392# a_1459_7392# a_1781_7392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X864 a_14913_n2883# a_14909_n3071# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X865 a_21626_4088# a_22115_4188# a_22323_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X866 a_16350_4765# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_3207_n8518# a_3460_n8722# a_3148_n9267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X868 a_34281_n5900# a_33884_n4152# a_34152_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X869 gnd d1 a_40830_2125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X870 a_1644_2543# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 a_40491_7772# a_40595_7021# a_40550_7034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X872 a_28195_3986# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 gnd d0 a_4500_n4060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X874 gnd d0 a_31149_7813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X875 vdd a_31161_5853# a_30953_5853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X876 a_39364_4426# a_39151_4426# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X877 a_32381_n4826# a_32870_n4845# a_33078_n4845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X878 a_6199_n6387# a_5778_n6387# a_5505_n6402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X879 a_6811_n2704# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X880 a_38257_6132# a_37836_6132# a_37560_6032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X881 a_39165_n4131# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X882 a_2835_4684# a_2955_6596# a_2906_6786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X883 a_35057_6765# a_35271_5643# a_35226_5656# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X884 vdd a_25885_4893# a_25677_4893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X885 a_40527_1718# a_40780_1705# a_40358_2827# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X886 a_36293_4914# a_36289_5091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X887 vdd d0 a_15161_n4068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X888 a_16661_n4853# a_16448_n4853# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X889 a_14786_7884# a_14782_8061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X890 a_37676_n2464# a_37332_n2231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X891 a_637_2257# a_424_2257# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X892 a_13720_7822# a_13824_7071# a_13779_7084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X893 a_5518_n3847# a_5518_n3565# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X894 a_26914_2987# a_27400_2771# a_27608_2771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X895 a_18872_2679# a_19070_3694# a_19021_3884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X896 a_8484_n8685# a_8741_n8701# a_8429_n9246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X897 vdd a_14153_n2853# a_13945_n2853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X898 gnd a_15051_5911# a_14843_5911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 a_830_5193# a_1634_5012# a_1793_5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X900 a_8372_1916# a_8476_1165# a_8431_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X901 a_35077_2848# a_35334_2658# a_34982_4840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X902 a_3114_7253# a_4175_6882# a_4130_6895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X903 gnd a_25994_n2635# a_25786_n2635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X904 a_7089_n6077# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X905 a_34026_n9001# a_33912_n9001# a_34120_n9001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X906 a_39086_1053# a_38873_1053# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X907 a_13660_n8059# a_13858_n9291# a_13809_n9275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 gnd a_36554_2944# a_36346_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X909 gnd d3 a_30043_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 a_34152_n3124# a_33731_n3124# a_34053_n2947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X911 a_22131_832# a_21918_832# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X912 vdd d0 a_9664_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X913 a_38150_n4409# a_37937_n4409# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X914 vdd d0 a_41917_n6954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X915 a_17586_2530# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X916 a_3109_8234# a_4170_7863# a_4121_8053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X917 a_11486_6182# a_11065_6182# a_10789_6364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X918 gnd d0 a_20429_n5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X919 a_18957_n4309# a_19171_n3393# a_19122_n3377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X920 a_5513_n4445# a_5520_n4244# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X921 gnd d1 a_24868_6055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 a_37924_n7347# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 a_38142_n6366# a_37929_n6366# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X924 a_5697_2800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X925 a_39661_n6056# a_39240_n6056# a_39566_n8048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X926 vdd d1 a_8647_8023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X927 vdd a_20346_3367# a_20138_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X928 a_37639_n9322# a_37644_n8936# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X929 a_28504_n4123# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X930 a_22404_n7775# a_21983_n7775# a_21707_n7474# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X931 a_33882_n4664# a_33669_n4664# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X932 a_12890_n6106# a_12469_n6106# a_12791_n5929# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X933 gnd d0 a_9659_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X934 a_34304_359# a_35031_4650# a_34986_4663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X935 a_4126_8291# a_4122_8468# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X936 a_22323_4188# a_23127_4007# a_23296_3565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X937 gnd d0 a_9766_n6975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X938 a_22314_5730# a_21893_5730# a_21620_5946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X939 gnd a_41811_8236# a_41603_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X940 gnd a_8369_4650# a_8161_4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X941 a_7207_n8069# a_6994_n8069# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X942 vdd d0 a_15148_n5613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X943 a_17591_2063# a_17378_2063# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X944 a_41570_5070# a_41827_4880# a_40558_5251# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X945 a_1624_6460# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X946 a_21628_4584# a_21626_4370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X947 a_7004_n6621# a_6791_n6621# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X948 a_12315_1103# a_12102_1103# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X949 a_38270_3194# a_37849_3194# a_37573_3094# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X950 gnd d0 a_25977_n5576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X951 a_37937_n4409# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_38125_n9307# a_37912_n9307# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X953 vdd d0 a_36639_n5999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X954 a_24410_n6285# a_24554_n4309# a_24505_n4293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X955 a_10816_1680# a_10814_1466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X956 gnd a_36562_2380# a_36354_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X957 a_37669_n3826# a_38158_n3845# a_38366_n3845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X958 gnd a_24957_n7714# a_24749_n7714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X959 a_35370_n6537# a_36428_n6975# a_36383_n6771# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X960 a_12587_n8098# a_12374_n8098# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_41569_5874# a_41822_5861# a_40553_6232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X962 vdd d2 a_19278_3694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X963 a_13879_n5778# a_14940_n5613# a_14891_n5597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X964 a_13585_n6134# a_13705_n8263# a_13656_n8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_16849_n8770# a_17653_n8589# a_17812_n8832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X966 a_1882_n6885# a_1510_n6642# a_919_n6823# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X967 a_18941_n8038# a_19194_n8242# a_18866_n6113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_11568_n8791# a_11147_n8791# a_10871_n8490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X969 a_5436_1056# a_5443_855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X970 a_12353_3483# a_12140_3483# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X971 a_25718_n6951# a_25721_n6348# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X972 a_28579_n6048# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 a_938_n2491# a_1743_n2725# a_1902_n2968# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X974 a_19037_1747# a_19290_1734# a_18868_2856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_25632_4522# a_25889_4332# a_24623_4111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X976 vdd d1 a_14133_n6770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X977 a_6114_4196# a_5693_4196# a_5417_4096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X978 gnd a_15064_2973# a_14856_2973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X979 a_9512_n6356# a_9765_n6560# a_8496_n6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X980 gnd d2 a_30087_7574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X981 a_242_n2605# a_731_n2906# a_939_n2906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X982 a_4138_5112# a_4395_4922# a_3126_5293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X983 a_29897_5243# a_30154_5053# a_29842_5804# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X984 gnd a_9773_n4603# a_9565_n4603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X985 a_28351_n3095# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X986 gnd d1 a_24962_n6733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X987 a_12241_n3153# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X988 vdd a_29836_n10368# a_29628_n10368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X989 a_21714_n6394# a_22200_n6379# a_22408_n6379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X990 a_3145_2180# a_4203_2401# a_4158_2414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X991 a_27187_2771# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X992 vdd a_20410_n9924# a_20202_n9924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X993 vdd a_4493_n5039# a_4285_n5039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X994 a_39066_4970# a_38853_4970# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X995 gnd a_14121_n8730# a_13913_n8730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X996 a_41667_n4566# a_41679_n3814# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X997 a_4240_n4835# a_4493_n5039# a_3227_n4601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X998 a_40573_2315# a_41634_1944# a_41589_1957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X999 a_12459_5559# a_12077_6001# a_11485_5767# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1000 a_17566_6447# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1001 gnd a_25886_5308# a_25678_5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1002 vdd d1 a_40830_2125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1003 a_32983_3781# a_33788_4015# a_33957_3573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1004 a_28697_n8040# a_28484_n8040# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 a_1989_n5105# a_1568_n5105# a_1890_n4928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1006 vdd d0 a_36542_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1007 a_22216_n3858# a_22003_n3858# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1008 gnd a_24818_5635# a_24610_5635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1009 a_29695_n6076# a_29815_n8205# a_29766_n8189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 a_16097_1064# a_16104_863# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1011 a_16058_8021# a_16060_7922# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1012 a_32272_7314# a_32761_7132# a_32969_7132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1013 a_16775_4204# a_16354_4204# a_16078_4386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1014 a_21722_n4437# a_21729_n4236# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1015 a_21882_8105# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 a_33952_3454# a_33580_3034# a_32988_2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1017 a_4122_8468# a_4125_7876# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1018 a_40342_6567# a_40540_7582# a_40491_7772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1019 a_27678_n8733# a_27257_n8733# a_26981_n8432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1020 vdd d0 a_31264_n4989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1021 a_6915_4991# a_6702_4991# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1022 a_32772_4757# a_32559_4757# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1023 a_41578_3113# a_41590_2372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1024 a_41646_n9276# a_41899_n9480# a_40630_n9645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1025 a_12650_n5113# a_12229_n5113# a_12551_n4936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1026 vdd d0 a_20415_n8943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1027 a_10784_7557# a_10782_7343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1028 a_34053_n2947# a_33681_n2704# a_33089_n2470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1029 a_20079_5903# a_20332_5890# a_19063_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 a_40662_n3768# a_41723_n3603# a_41674_n3587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1031 a_17571_5980# a_17358_5980# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1032 a_16640_n8355# a_16427_n8355# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_25653_1404# a_25906_1391# a_24640_1170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1034 a_21700_n8453# a_22189_n8754# a_22397_n8754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1035 a_35210_7793# a_35467_7603# a_35061_6588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1036 gnd a_40768_3665# a_40560_3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1037 a_37585_1416# a_38074_1234# a_38282_1234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1038 a_1471_5432# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1039 a_40451_n4092# a_40704_n4296# a_40352_n6272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_24615_6068# a_25673_6289# a_25628_6302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1041 a_1806_3594# a_1424_4036# a_832_3802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1042 gnd a_9664_6861# a_9456_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 gnd d0 a_4395_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1044 vdd d1 a_35611_n8701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1045 vdd a_35606_n9682# a_35398_n9682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1046 a_17502_n7049# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1047 a_10777_8324# a_11266_8142# a_11474_8142# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1048 a_32289_3997# a_32775_3781# a_32983_3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1049 a_14892_n6385# a_14888_n6573# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1050 a_13469_n10410# a_13726_n10426# a_13568_n10410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1051 a_38245_8092# a_39049_7911# a_39218_7469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1052 a_7163_n6864# a_7054_n7041# a_7262_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1053 vdd d6 a_37407_n10464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1054 vdd a_14078_n7331# a_13870_n7331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1055 a_16856_n7791# a_16435_n7791# a_16159_n7490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1056 a_24717_n4572# a_25775_n5010# a_25730_n4806# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1057 vdd d0 a_20442_n4047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1058 a_26919_2389# a_26919_2107# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1059 a_5429_2418# a_5918_2236# a_6126_2236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1060 gnd a_24915_n5337# a_24707_n5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 a_25631_4107# a_25641_3364# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1062 a_19083_2344# a_20144_1973# a_20099_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1063 a_13868_n8526# a_14926_n8964# a_14881_n8760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1064 a_27200_1226# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1065 vdd d1 a_24868_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1066 a_28760_n5055# a_28339_n5055# a_28661_n4878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1067 a_17986_367# a_17773_367# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1068 a_30934_1383# a_31187_1370# a_29921_1149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1069 a_7000_4447# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1070 a_38930_n8560# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1071 a_34008_2522# a_33795_2522# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1072 a_21618_6327# a_21618_6045# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1073 a_10878_n7511# a_11367_n7812# a_11575_n7812# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1074 a_518_n2906# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1075 a_9427_3134# a_9684_2944# a_8415_3315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1076 a_16772_5180# a_17576_4999# a_17735_5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1077 a_12462_3483# a_12090_3063# a_11498_2829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1078 a_32988_2800# a_32567_2800# a_32301_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 vdd a_41811_8236# a_41603_8236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1080 vdd a_8369_4650# a_8161_4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1081 a_28175_7903# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1082 a_32657_n4845# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 a_1880_7392# a_1837_6460# a_2045_6460# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1084 gnd a_19409_n7730# a_19201_n7730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1085 a_9528_n3835# a_9781_n4039# a_8515_n3601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1086 vdd d0 a_4499_n3645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1087 a_25717_n6536# a_25974_n6552# a_24705_n6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1088 gnd d0 a_25990_n4031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1089 a_1409_6972# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1090 a_35386_n2808# a_35643_n2824# a_35331_n3369# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1091 a_116_8034# a_605_8134# a_813_8134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1092 a_26988_n7453# a_26990_n7354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1093 a_40630_n9645# a_41691_n9480# a_41646_n9276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1094 a_12166_n7631# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1095 a_17748_3581# a_17366_4023# a_16774_3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1096 a_16558_5746# a_16345_5746# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1097 a_40507_5635# a_40760_5622# a_40338_6744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_36386_n5795# a_36639_n5999# a_35373_n5561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1099 a_13895_n3630# a_14953_n4068# a_14908_n3864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1100 vdd a_36562_2380# a_36354_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1101 a_30929_2364# a_30925_2541# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1102 a_6722_1074# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1103 a_18852_6596# a_19050_7611# a_19001_7801# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 a_3075_5677# a_3328_5664# a_2906_6786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_37656_n6976# a_37654_n6762# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1106 vdd a_9697_1399# a_9489_1399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1107 a_1890_n4928# a_1518_n4685# a_926_n4451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1108 a_19033_1924# a_19290_1734# a_18868_2856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1109 a_26901_6520# a_26899_6306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1110 a_41590_1153# a_37594_834# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1111 vdd a_9786_n3058# a_9578_n3058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1112 a_26988_n7453# a_27477_n7754# a_27685_n7754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1113 a_33699_n9001# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 vdd d2 a_30087_7574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1115 a_32281_6549# a_32279_6335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1116 gnd d0 a_31258_n5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1117 gnd d0 a_15077_1428# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1118 a_6760_3454# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1119 vdd d0 a_41920_n5978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1120 a_32542_7698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1121 gnd a_36630_n7541# a_36422_n7541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1122 gnd d0 a_36635_n6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1123 a_16075_5362# a_16075_5080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1124 gnd a_30238_n7693# a_30030_n7693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_12551_n4936# a_12179_n4693# a_11587_n4459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1126 a_40651_n6516# a_41709_n6954# a_41664_n6750# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1127 a_32381_n4826# a_32381_n4544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1128 a_30997_n7308# a_30993_n7496# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1129 gnd a_4480_n7977# a_4272_n7977# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1130 a_22340_1247# a_23144_1066# a_23303_1486# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1131 gnd a_4415_1005# a_4207_1005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1132 a_6093_7698# a_6898_7932# a_7067_7490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1133 a_34959_n10381# a_35216_n10397# a_35058_n10381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1134 a_30921_2928# a_30917_3105# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1135 a_12518_2551# a_12305_2551# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1136 a_10789_6082# a_10791_5983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1137 a_28276_n7573# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1138 vdd a_40912_n4763# a_40704_n4763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1139 a_28180_6922# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1140 a_14880_n8345# a_14876_n8533# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1141 a_16186_n3088# a_16667_n3459# a_16875_n3459# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1142 a_22203_n5403# a_21990_n5403# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 a_32356_n9442# a_32845_n9743# a_33053_n9743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1144 gnd d0 a_9769_n5999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1145 a_17943_n3132# a_17522_n3132# a_17844_n2955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1146 a_11053_8142# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1147 vdd a_8756_n5765# a_8548_n5765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1148 a_37654_n6480# a_37656_n6381# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1149 vdd d1 a_8761_n4784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1150 a_20853_n686# a_20674_141# a_10603_285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1151 vdd a_24818_5635# a_24610_5635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1152 a_10797_4125# a_10799_4026# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1153 vdd a_35556_n9262# a_35348_n9262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1154 a_25628_5083# a_25636_4345# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1155 gnd a_15153_n4632# a_14945_n4632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1156 a_927_n4866# a_506_n4866# a_230_n4565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1157 a_40342_6567# a_40540_7582# a_40495_7595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1158 a_11511_1284# a_12315_1103# a_12474_1523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1159 vdd a_31154_6832# a_30946_6832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1160 a_38339_n8741# a_37918_n8741# a_37642_n8440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1161 gnd a_37407_n10464# a_37199_n10464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1162 a_207_n9364# a_693_n9349# a_901_n9349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1163 a_12442_7400# a_12070_6980# a_11479_7161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1164 a_24708_n5741# a_25769_n5576# a_25720_n5560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1165 a_33912_n9001# a_33699_n9001# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1166 a_35373_n5561# a_36431_n5999# a_36386_n5795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1167 a_38250_7111# a_37829_7111# a_37553_7011# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1168 a_32968_6717# a_32547_6717# a_32274_6933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1169 a_28494_n6592# a_28281_n6592# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1170 vdd d1 a_3475_n5786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1171 a_38163_n2864# a_37950_n2864# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1172 a_30897_8241# a_30893_8418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1173 a_33057_n8347# a_33862_n8581# a_34021_n8824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1174 a_11599_n2499# a_11178_n2499# a_10905_n2514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1175 a_28661_n4878# a_28289_n4635# a_27697_n4401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1176 a_10905_n3109# a_10903_n2895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1177 a_39151_4426# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1178 vdd a_40768_3665# a_40560_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1179 a_5503_n6783# a_5503_n6501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1180 gnd a_20320_7850# a_20112_7850# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1181 a_630_3236# a_417_3236# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1182 a_24670_n3361# a_24774_n2816# a_24729_n2612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1183 a_24674_n3173# a_24927_n3377# a_24505_n4293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1184 a_2044_380# a_1831_380# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1185 a_17728_7498# a_17346_7940# a_16755_8121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1186 a_23372_n6856# a_23000_n6613# a_22409_n6794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1187 a_7062_n5084# a_6849_n5084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1188 a_837_2821# a_416_2821# a_143_3037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1189 a_33090_n2885# a_32669_n2885# a_32393_n2866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1190 a_13821_n7315# a_13925_n6770# a_13880_n6566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1191 a_7421_4447# a_7325_359# a_5243_292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1192 a_6094_8113# a_5673_8113# a_5397_8013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1193 a_28455_5382# a_28242_5382# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1194 a_424_2257# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1195 a_36373_n7525# a_36630_n7541# a_35361_n7706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1196 a_29000_n6048# a_29836_n10368# a_26489_n10440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1197 a_24650_n7278# a_24754_n6733# a_24705_n6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1198 gnd d1 a_30137_7994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1199 a_8364_3699# a_8617_3686# a_8211_2671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1200 a_4223_n7961# a_4480_n7977# a_3214_n7539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1201 a_29862_1887# a_29966_1136# a_29917_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1202 a_21987_n6379# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1203 a_24717_n4572# a_24970_n4776# a_24658_n5321# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1204 a_41684_n2833# a_41680_n3021# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1205 a_39205_n7020# a_38992_n7020# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1206 a_30930_1560# a_31187_1370# a_29921_1149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1207 a_22391_n9320# a_21970_n9320# a_21697_n9335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1208 gnd d1 a_24861_7034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1209 a_2995_n8239# a_3209_n7323# a_3164_n7119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1210 a_39421_n5063# a_39000_n5063# a_39322_n4886# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1211 a_29862_1887# a_30119_1697# a_29697_2819# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1212 a_10791_5983# a_10796_5597# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1213 vdd d1 a_40892_n8680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1214 a_29978_n8468# a_31036_n8906# a_30987_n8890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 a_6849_n5084# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1216 gnd a_41936_n2622# a_41728_n2622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1217 a_39332_3433# a_38911_3433# a_39238_3552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1218 a_30985_n9268# a_30981_n9456# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1219 a_844_1842# a_1649_2076# a_1818_1634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1220 a_33649_n8581# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1221 a_30998_n6515# a_31255_n6531# a_29986_n6696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1222 gnd a_9780_n3624# a_9572_n3624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1223 gnd a_24868_6055# a_24660_6055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1224 a_11478_6746# a_11057_6746# a_10784_6962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1225 a_36273_8447# a_36530_8257# a_35264_8036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1226 gnd d0 a_15133_n8549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1227 gnd d0 a_36651_n4039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1228 a_1813_1515# a_1441_1095# a_849_861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1229 a_40495_7595# a_40590_8002# a_40541_8192# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1230 a_17510_n5092# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1231 gnd d1 a_19345_1173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1232 a_40503_5812# a_40760_5622# a_40338_6744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1233 a_41574_4509# a_41577_3917# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1234 gnd a_30188_n7273# a_29980_n7273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1235 a_5443_855# a_5922_840# a_6130_840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1236 a_4251_n2460# a_4247_n2648# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1237 a_21976_n8754# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1238 a_5506_n5525# a_5995_n5826# a_6203_n5826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1239 a_11490_4786# a_12295_5020# a_12454_5440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1240 a_36377_n7337# a_36373_n7525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1241 a_1981_n7062# a_1560_n7062# a_1882_n6885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1242 a_38923_1473# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1243 a_32294_3611# a_32292_3397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1244 a_18852_6596# a_19050_7611# a_19005_7624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1245 a_37855_1800# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1246 a_12387_n5674# a_12174_n5674# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1247 a_30005_n3572# a_31063_n4010# a_31014_n3994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_3071_5854# a_3328_5664# a_2906_6786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1249 a_26978_n9314# a_27464_n9299# a_27672_n9299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1250 a_222_n6522# a_224_n6423# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1251 a_35299_n9246# a_35403_n8701# a_35358_n8497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1252 a_38345_n7347# a_39150_n7581# a_39319_n7020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1253 a_12102_1103# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1254 a_19156_n7526# a_20214_n7964# a_20165_n7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1255 a_4210_n9506# a_4467_n9522# a_3198_n9687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1256 a_40667_n2787# a_40924_n2803# a_40612_n3348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1257 vdd a_40615_2637# a_40407_2637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1258 a_8187_6765# a_8401_5643# a_8352_5833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1259 vdd a_3065_n10418# a_2857_n10418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1260 a_40511_3855# a_40615_3104# a_40570_3117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1261 a_11166_n4459# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1262 a_37567_4952# a_38053_4736# a_38261_4736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 vdd a_19278_3694# a_19070_3694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1264 a_31889_n10455# a_37199_n10464# a_37150_n10448# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1265 a_5488_n9938# a_5486_n9724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1266 a_38281_819# a_37860_819# a_37594_834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1267 a_22314_5730# a_23119_5964# a_23288_5522# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1268 a_6207_n4430# a_7012_n4664# a_7171_n4907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1269 a_30987_n8890# a_30990_n8287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1270 a_16661_n4853# a_16448_n4853# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1271 a_19063_6261# a_20124_5890# a_20079_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1272 a_39150_n7581# a_38937_n7581# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1273 a_4214_n9318# a_4210_n9506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1274 gnd a_19119_n6317# a_18911_n6317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 gnd d2 a_19379_n3393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1276 a_22132_1247# a_21919_1247# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1277 a_11285_3810# a_11072_3810# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1278 gnd a_8629_1726# a_8421_1726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1279 a_36302_3372# a_36555_3359# a_35289_3138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_11372_n6831# a_11159_n6831# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1281 a_14815_2599# a_14818_2007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1282 a_33949_5530# a_33567_5972# a_32975_5738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1283 a_40263_4819# a_40520_4629# a_39585_338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1284 gnd d0 a_31276_n3029# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1285 a_19102_n7294# a_19206_n6749# a_19157_n6733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1286 a_12662_n3153# a_12607_n4181# a_12791_n5929# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1287 a_27408_2207# a_27195_2207# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1288 gnd d0 a_41916_n6539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1289 a_27179_4728# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1290 a_26998_n5397# a_27003_n5011# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1291 a_16072_5962# a_16558_5746# a_16766_5746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1292 a_19169_n4588# a_19422_n4792# a_19110_n5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1293 a_35281_5095# a_35534_5082# a_35222_5833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1294 a_16161_n8169# a_16159_n7772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1295 a_16860_n6395# a_16439_n6395# a_16169_n6029# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1296 a_35315_n7098# a_35410_n7722# a_35361_n7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1297 a_10799_4621# a_11282_4786# a_11490_4786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1298 vdd a_36542_6297# a_36334_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1299 a_14877_n8948# a_14880_n8345# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1300 a_17703_n9009# a_17490_n9009# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1301 a_29884_8007# a_30942_8228# a_30897_8241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1302 vdd d0 a_9684_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1303 a_38937_n7581# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1304 a_5698_3215# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1305 vdd d0 a_36534_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1306 a_33882_n4664# a_33669_n4664# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1307 a_6702_4991# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1308 gnd d1 a_24888_2138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1309 a_10886_n5836# a_10886_n5554# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1310 a_23422_4439# a_23209_4439# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1311 gnd a_29948_n6280# a_29740_n6280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1312 vdd a_31186_955# a_30978_955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1313 a_3125_6097# a_3378_6084# a_3075_5677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1314 a_22315_6145# a_21894_6145# a_21618_6045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1315 gnd d0 a_9679_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 a_27482_n6773# a_27269_n6773# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1317 vdd d3 a_3272_n4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1318 vdd a_36541_5882# a_36333_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1319 gnd d0 a_36529_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1320 a_40557_6055# a_41615_6276# a_41566_6466# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1321 a_24729_n2612# a_25787_n3050# a_25738_n3034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 a_40654_n5540# a_41712_n5978# a_41667_n5774# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1323 a_35366_n6725# a_36427_n6560# a_36378_n6544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1324 gnd d0 a_15149_n6028# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1325 a_36308_1978# a_36304_2155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1326 a_11359_n8376# a_11146_n8376# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1327 a_29931_n7257# a_30035_n6712# a_29986_n6696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 a_12561_3483# a_12518_2551# a_12702_4476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1329 vdd d0 a_4378_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1330 a_38125_n9307# a_37912_n9307# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1331 a_8431_1178# a_9489_1399# a_9444_1412# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1332 a_2134_n8090# a_1713_n8090# a_1969_n9022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1333 a_8360_3876# a_8617_3686# a_8211_2671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1334 a_36390_n4399# a_36643_n4603# a_35374_n4768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1335 a_5885_7698# a_5672_7698# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1336 a_493_n7804# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1337 a_29862_1887# a_29966_1136# a_29921_1149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1338 gnd a_4395_4922# a_4187_4922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1339 a_24604_7224# a_25665_6853# a_25620_6866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1340 a_14812_3401# a_15065_3388# a_13799_3167# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1341 gnd a_25970_n7948# a_25762_n7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1342 a_12563_n2976# a_12454_n3153# a_12662_n3153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1343 a_16454_n3459# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1344 a_19056_7240# a_20117_6869# a_20068_7059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1345 a_37565_5333# a_37565_5051# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1346 a_1882_n6885# a_1510_n6642# a_918_n6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1347 vdd d1 a_24861_7034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1348 a_26899_6024# a_26901_5925# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1349 a_21697_n9930# a_21695_n9716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1350 a_8449_n5329# a_8553_n4784# a_8508_n4580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1351 a_35246_1739# a_35341_2146# a_35292_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1352 a_8453_n5141# a_8706_n5345# a_8300_n4113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1353 a_939_n2906# a_1743_n2725# a_1902_n2968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1354 a_23144_1066# a_22931_1066# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1355 a_32279_6053# a_32281_5954# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1356 a_24599_8205# a_25660_7834# a_25611_8024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1357 gnd d0 a_31250_n7512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_5436_1651# a_5434_1437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1359 a_242_n2887# a_731_n2906# a_939_n2906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1360 a_3125_6097# a_4183_6318# a_4134_6508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1361 vdd a_24868_6055# a_24660_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1362 a_3152_n9079# a_3247_n9703# a_3198_n9687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1363 gnd a_20409_n9509# a_20201_n9509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1364 a_5422_3397# a_5422_3115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1365 a_28740_n8972# a_28319_n8972# a_28646_n8972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1366 a_33795_2522# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1367 vdd d1 a_19345_1173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1368 a_23182_3446# a_22969_3446# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1369 gnd a_4484_n6581# a_4276_n6581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 a_16551_6725# a_16338_6725# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1371 vdd d1 a_24965_n5757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1372 a_913_n7389# a_492_n7389# a_224_n7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1373 a_32637_n8762# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1374 a_17435_n9570# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1375 a_34083_4447# a_33870_4447# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1376 a_28673_n2918# a_28564_n3095# a_28772_n3095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1377 gnd d0 a_15039_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1378 a_19067_6084# a_20125_6305# a_20076_6495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1379 gnd d0 a_20346_3367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1380 a_33800_2055# a_33587_2055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1381 gnd d0 a_20414_n8528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1382 a_16092_2640# a_16571_2808# a_16779_2808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1383 gnd d0 a_41932_n4018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1384 a_8187_6765# a_8401_5643# a_8356_5656# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1385 a_32773_5172# a_32560_5172# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1386 a_13891_n3818# a_14148_n3834# a_13845_n3210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1387 a_12801_4476# a_12705_388# a_12913_388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 a_23624_n8061# a_23203_n8061# a_23471_n7033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1389 a_9412_7289# a_9665_7276# a_8399_7055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 a_609_6738# a_396_6738# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1391 a_37649_n7461# a_37651_n7362# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1392 vdd d0 a_31186_955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1393 a_21700_n8735# a_22189_n8754# a_22397_n8754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1394 a_25643_2147# a_25900_1957# a_24631_2328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1395 a_27604_4167# a_27183_4167# a_26907_4067# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1396 a_8414_4119# a_8667_4106# a_8364_3699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1397 vdd a_8629_1726# a_8421_1726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1398 a_30910_5477# a_31167_5287# a_29901_5066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1399 a_12553_5440# a_12498_6468# a_12706_6468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1400 a_902_n9764# a_481_n9764# a_205_n9745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1401 a_9529_n3042# a_9532_n2439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1402 a_25628_5083# a_25885_4893# a_24616_5264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1403 gnd a_15077_1428# a_14869_1428# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1404 a_9415_6487# a_9418_5895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1405 a_6110_4757# a_5689_4757# a_5419_4592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1406 a_1743_n2725# a_1530_n2725# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1407 a_37829_7111# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1408 a_22328_3207# a_21907_3207# a_21631_3389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1409 a_26901_5925# a_26906_5539# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1410 a_5404_7528# a_5402_7314# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1411 a_29912_2307# a_30169_2117# a_29866_1710# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1412 a_39421_n5063# a_39378_n4131# a_39562_n5879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1413 a_37654_n6762# a_38143_n6781# a_38351_n6781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1414 a_8516_n2808# a_9577_n2643# a_9528_n2627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1415 a_32881_n2470# a_32668_n2470# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1416 a_12305_2551# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1417 a_13864_n8714# a_14925_n8549# a_14876_n8533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1418 a_5498_n7764# a_5498_n7482# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1419 a_35385_n3601# a_36443_n4039# a_36394_n4023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1420 a_35277_5272# a_35534_5082# a_35222_5833# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1421 a_23643_351# a_23534_351# a_23742_351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1422 a_38150_n4409# a_37937_n4409# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1423 a_21727_n3839# a_22216_n3858# a_22424_n3858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1424 a_4222_n7546# a_4232_n6792# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1425 a_5782_n5826# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1426 a_21919_1247# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1427 a_7411_n5900# a_7014_n4152# a_7270_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1428 a_10878_n7793# a_11367_n7812# a_11575_n7812# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1429 a_6841_n7041# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1430 a_7415_n8069# a_7302_n6077# a_7510_n6077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1431 a_23471_n7033# a_23050_n7033# a_23372_n6856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1432 a_38048_5717# a_37835_5717# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1433 a_32787_1821# a_32574_1821# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1434 a_9492_n9900# a_9495_n9297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1435 a_21714_n6394# a_21717_n6013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1436 a_32864_n5411# a_32651_n5411# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1437 a_3121_6274# a_3378_6084# a_3075_5677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1438 a_5493_n8362# a_5500_n8161# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1439 a_40557_6055# a_41615_6276# a_41570_6289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1440 a_39066_4970# a_38853_4970# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1441 a_22961_5403# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1442 a_37925_n7762# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1443 a_2999_n8051# a_3197_n9283# a_3148_n9267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1444 a_38143_n6781# a_37930_n6781# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1445 vdd a_31270_n3595# a_31062_n3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1446 a_36399_n3042# a_36656_n3058# a_35390_n2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1447 gnd a_9692_2380# a_9484_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1448 gnd d2 a_40748_7582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1449 gnd d0 a_15146_n7004# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1450 a_6799_n4664# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1451 a_8356_5656# a_8451_6063# a_8402_6253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1452 a_7322_4447# a_6925_2522# a_7193_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1453 a_16559_6161# a_16346_6161# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1454 a_37937_n4409# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1455 a_10814_1466# a_11303_1284# a_11511_1284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1456 a_38265_4175# a_37844_4175# a_37568_4357# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1457 a_12333_7400# a_12120_7400# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1458 gnd a_9677_5316# a_9469_5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1459 a_20080_5099# a_20088_4361# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1460 a_22417_n4837# a_21996_n4837# a_21720_n4818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1461 a_29697_2819# a_29911_1697# a_29862_1887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1462 a_38980_n8980# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1463 a_17460_n4672# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1464 a_35246_1739# a_35341_2146# a_35296_2159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1465 a_13571_6617# a_13769_7632# a_13720_7822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1466 a_26919_2389# a_27408_2207# a_27616_2207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 a_1969_n9022# a_1548_n9022# a_1875_n9022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1468 gnd a_8679_2146# a_8471_2146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 gnd a_30137_7994# a_29929_7994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1470 a_22303_8105# a_23107_7924# a_23276_7482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1471 a_26988_n7735# a_27477_n7754# a_27685_n7754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1472 a_35369_n5749# a_35626_n5765# a_35323_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1473 a_17571_5980# a_17358_5980# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1474 a_40647_n6704# a_41708_n6539# a_41659_n6523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1475 a_16152_n8751# a_16641_n8770# a_16849_n8770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1476 a_7282_n3124# a_6861_n3124# a_7188_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1477 a_41671_n4378# a_41924_n4582# a_40655_n4747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_13841_n3398# a_14098_n3414# a_13676_n4330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1479 a_32543_8113# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1480 a_40592_n7265# a_40696_n6720# a_40647_n6704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1481 gnd a_31251_n7927# a_31043_n7927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1482 a_5906_4196# a_5693_4196# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1483 a_14814_2184# a_14824_1441# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1484 a_6910_5972# a_6697_5972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1485 a_34063_1494# a_33642_1494# a_33969_1613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1486 a_32356_n9724# a_32845_n9743# a_33053_n9743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1487 a_22899_6943# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1488 a_5975_n9743# a_5762_n9743# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1489 a_21707_n7756# a_21707_n7474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1490 a_2924_n6126# a_3044_n8255# a_2995_n8239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1491 a_7322_4447# a_7213_4447# a_7421_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1492 a_40558_5251# a_41619_4880# a_41570_5070# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1493 gnd a_19345_1173# a_19137_1173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1494 vdd a_3467_n7743# a_3259_n7743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1495 a_30897_8241# a_31150_8228# a_29884_8007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1496 a_25733_n4015# a_25990_n4031# a_24724_n3593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1497 a_13883_n5590# a_14941_n6028# a_14892_n6012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1498 a_25633_5321# a_25886_5308# a_24620_5087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1499 a_33957_3573# a_33575_4015# a_32984_4196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1500 gnd a_36619_n9916# a_36411_n9916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1501 a_23392_n2939# a_23283_n3116# a_23491_n3116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1502 a_9408_7466# a_9665_7276# a_8399_7055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1503 gnd d0 a_4390_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1504 a_24565_5648# a_24818_5635# a_24396_6757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1505 vdd d1 a_30246_n5736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1506 a_15904_300# a_17773_367# a_18095_367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1507 a_32969_7132# a_32548_7132# a_32272_7032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1508 a_33889_n3685# a_33676_n3685# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1509 a_1704_1515# a_1491_1515# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1510 a_21702_n8354# a_21709_n8153# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1511 a_8427_1355# a_9488_984# a_9443_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1512 a_32294_3016# a_32301_2632# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1513 a_8205_n6105# a_8325_n8234# a_8280_n8030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1514 a_37580_2115# a_38069_2215# a_38277_2215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1515 a_7326_6439# a_6905_6439# a_7161_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1516 a_23372_n6856# a_23000_n6613# a_22408_n6379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1517 gnd a_9774_n5018# a_9566_n5018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1518 a_13794_4148# a_14047_4135# a_13744_3728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1519 a_14881_n8760# a_15134_n8964# a_13868_n8526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1520 a_3126_5293# a_4187_4922# a_4138_5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1521 a_27583_7669# a_28388_7903# a_28557_7461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1522 a_27705_n3837# a_27284_n3837# a_27008_n3818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1523 a_5404_6933# a_5890_6717# a_6098_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1524 a_33932_7371# a_33560_6951# a_32968_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1525 vdd d0 a_9773_n4603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1526 vdd a_15145_n6589# a_14937_n6589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1527 a_27401_3186# a_27188_3186# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1528 a_11072_3810# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1529 a_26832_263# a_26411_263# a_26733_263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1530 a_32373_n6783# a_32373_n6501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1531 a_30005_n3572# a_30258_n3776# a_29955_n3152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1532 a_20674_141# d8 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1533 vdd d1 a_19325_5090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1534 a_32983_3781# a_32562_3781# a_32294_3611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1535 a_7082_3454# a_6973_3454# a_7181_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1536 a_29846_5627# a_30099_5614# a_29677_6736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1537 a_26411_263# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1538 a_24662_n5133# a_24757_n5757# a_24712_n5553# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1539 gnd a_25974_n6552# a_25766_n6552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_38371_n2864# a_39175_n2683# a_39334_n2926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1541 a_27195_2207# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1542 a_38930_n8560# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1543 a_33073_n5826# a_32652_n5826# a_32376_n5807# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1544 a_1786_7511# a_1404_7953# a_812_7719# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1545 a_34132_n7041# a_33711_n7041# a_34033_n6864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1546 gnd d1 a_24881_3117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1547 a_35319_n5329# a_35576_n5345# a_35170_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1548 a_12467_3602# a_12085_4044# a_11494_4225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1549 a_40666_n3580# a_41724_n4018# a_41675_n4002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1550 a_29921_1149# a_30979_1370# a_30930_1560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1551 gnd a_31186_955# a_30978_955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1552 a_3118_7076# a_3371_7063# a_3059_7814# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1553 a_11479_7161# a_11058_7161# a_10782_7061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 vdd a_36534_6861# a_36326_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1555 a_6195_n7783# a_5774_n7783# a_5498_n7482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1556 a_37659_n5405# a_37664_n5019# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1557 vdd a_9692_2380# a_9484_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1558 vdd d2 a_40748_7582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1559 a_8356_5656# a_8451_6063# a_8406_6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1560 gnd d1 a_19417_n5773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1561 gnd a_35643_n2824# a_35435_n2824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1562 a_21976_n8754# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1563 a_5506_n5807# a_5995_n5826# a_6203_n5826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1564 a_40515_3678# a_40610_4085# a_40561_4275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1565 vdd a_9677_5316# a_9469_5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1566 a_12795_n8098# a_12682_n6106# a_12890_n6106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1567 gnd d0 a_15072_2409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1568 a_33001_1255# a_33805_1074# a_33964_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1569 a_8394_8036# a_8647_8023# a_8344_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1570 a_24705_n6717# a_24962_n6733# a_24650_n7278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1571 a_12387_n5674# a_12174_n5674# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1572 a_13571_6617# a_13769_7632# a_13724_7645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1573 a_217_n7503# a_706_n7804# a_914_n7804# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1574 a_16792_1263# a_16371_1263# a_16095_1163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1575 a_21697_n9930# a_25958_n9908# a_24692_n9470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1576 a_12442_7400# a_12070_6980# a_11478_6746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1577 vdd a_8679_2146# a_8471_2146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1578 a_30981_n9456# a_31238_n9472# a_29969_n9637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1579 vdd a_4378_7863# a_4170_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1580 a_8201_n6293# a_8345_n4317# a_8296_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1581 a_41680_n3021# a_41937_n3037# a_40671_n2599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1582 a_21640_2624# a_21638_2410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1583 a_5672_7698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1584 a_35280_4296# a_35537_4106# a_35234_3699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1585 a_38277_2215# a_39081_2034# a_39250_1592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 gnd d0 a_20427_n6983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 a_1946_n4173# a_1733_n4173# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1588 a_7173_5411# a_6752_5411# a_7079_5530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1589 a_6208_n4845# a_7012_n4664# a_7171_n4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_17728_7498# a_17346_7940# a_16754_7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1591 a_1781_7392# a_1409_6972# a_818_7153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1592 a_22003_n3858# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1593 a_818_7153# a_397_7153# a_121_7335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1594 a_14895_n5409# a_15148_n5613# a_13879_n5778# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_3234_n3622# a_4292_n4060# a_4247_n3856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1596 a_8415_3315# a_9476_2944# a_9427_3134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1597 a_25738_n3034# a_25741_n2431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1598 a_28413_3005# a_28200_3005# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1599 a_30902_7260# a_30898_7437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1600 a_918_n6408# a_1723_n6642# a_1882_n6885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1601 a_22334_1813# a_23139_2047# a_23308_1605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1602 a_11372_n6831# a_11159_n6831# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1603 vdd d0 a_31239_n9887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1604 a_11286_4225# a_11073_4225# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1605 a_19060_7063# a_19313_7050# a_19001_7801# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_33835_5411# a_33622_5411# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1607 a_12290_6001# a_12077_6001# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1608 a_40650_n5728# a_40907_n5744# a_40604_n5120# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1609 a_28331_n7012# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1610 a_35081_2671# a_35334_2658# a_34982_4840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1611 a_32358_n9938# a_32356_n9724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1612 vdd a_19345_1173# a_19137_1173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1613 a_28207_2026# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1614 vdd a_4473_n8956# a_4265_n8956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1615 gnd a_3480_n4805# a_3272_n4805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1616 a_30006_n2779# a_31067_n2614# a_31022_n2410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1617 a_23208_n7594# a_22995_n7594# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1618 a_39116_5390# a_38903_5390# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1619 a_13880_n6566# a_14938_n7004# a_14889_n6988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1620 a_11505_1850# a_12310_2084# a_12479_1642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1621 a_24561_5825# a_24818_5635# a_24396_6757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1622 a_212_n8978# a_693_n9349# a_901_n9349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1623 a_13880_n6566# a_14133_n6770# a_13821_n7315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1624 a_28289_n4635# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1625 a_20188_n3428# a_20184_n3616# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1626 a_10794_5383# a_11283_5201# a_11491_5201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1627 a_21913_1813# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1628 a_14788_7495# a_15045_7305# a_13779_7084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1629 gnd a_20346_3367# a_20138_3367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1630 vdd d5 a_35216_n10397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1631 a_1793_n3145# a_1580_n3145# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1632 a_26924_1126# a_26926_1027# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1633 a_8426_2159# a_9484_2380# a_9435_2570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1634 a_20076_6495# a_20079_5903# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1635 a_32560_5172# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1636 a_40577_2138# a_40830_2125# a_40527_1718# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1637 a_13790_4325# a_14047_4135# a_13744_3728# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1638 a_24692_n9470# a_25750_n9908# a_21697_n9930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1639 a_625_4217# a_412_4217# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1640 a_12630_n9030# a_12209_n9030# a_12531_n8853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1641 a_27692_n5382# a_27271_n5382# a_27003_n5011# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1642 a_396_6738# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1643 a_27482_n6773# a_27269_n6773# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1644 a_6829_n9001# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1645 a_21625_4965# a_22111_4749# a_22319_4749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1646 a_3218_n5770# a_4279_n5605# a_4234_n5401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1647 a_39339_n3103# a_38957_n3664# a_38366_n3845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1648 gnd d0 a_41905_n8914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_32877_n3866# a_32664_n3866# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1650 a_19025_3707# a_19120_4114# a_19071_4304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1651 a_20178_n5010# a_20435_n5026# a_19169_n4588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1652 a_11359_n8376# a_11146_n8376# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1653 a_16772_5180# a_16351_5180# a_16075_5362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1654 a_9523_n3608# a_9533_n2854# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1655 a_40431_n8009# a_40684_n8213# a_40356_n6084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1656 a_493_n7804# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 a_227_n5447# a_232_n5061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1658 gnd d2 a_19367_n5353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1659 a_3180_n3390# a_3437_n3406# a_3015_n4322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1660 a_10811_2066# a_11297_1850# a_11505_1850# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1661 a_29842_5804# a_30099_5614# a_29677_6736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1662 a_39074_3013# a_38861_3013# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1663 a_5886_8113# a_5673_8113# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1664 a_31011_n4785# a_31264_n4989# a_29998_n4551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1665 vdd d0 a_4398_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1666 a_133_5093# a_622_5193# a_830_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1667 a_30898_7437# a_30901_6845# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1668 a_16078_4386# a_16078_4104# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1669 a_20162_n8739# a_20415_n8943# a_19149_n8505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1670 a_27465_n9714# a_27252_n9714# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1671 a_30901_6845# a_31154_6832# a_29885_7203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1672 a_16147_n9732# a_16147_n9450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1673 a_36282_7289# a_36278_7466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1674 a_20190_n3050# a_20193_n2447# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1675 a_18171_n6085# a_19007_n10405# a_15660_n10477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1676 a_29900_4267# a_30961_3896# a_30916_3909# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1677 a_3164_n7119# a_3417_n7323# a_2995_n8239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1678 a_3160_n7307# a_3264_n6762# a_3219_n6558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1679 vdd d0 a_41835_2923# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1680 vdd a_20426_n6568# a_20218_n6568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1681 a_29921_1149# a_30979_1370# a_30934_1383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1682 a_23327_6431# a_23114_6431# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1683 a_29923_n9029# a_30018_n9653# a_29969_n9637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1684 a_3223_n4789# a_3480_n4805# a_3168_n5350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1685 a_3114_7253# a_3371_7063# a_3059_7814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1686 a_28740_n8972# a_28319_n8972# a_28641_n8795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1687 gnd a_3425_n5366# a_3217_n5366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1688 a_10777_8324# a_10777_8042# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1689 gnd a_31255_n6531# a_31047_n6531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1690 gnd a_40924_n2803# a_40716_n2803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1691 a_37835_5717# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1692 a_1875_n9022# a_1493_n9583# a_901_n9349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1693 a_32574_1821# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1694 a_1818_1634# a_1436_2076# a_845_2257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1695 a_24615_6068# a_24868_6055# a_24565_5648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1696 a_16552_7140# a_16339_7140# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_40515_3678# a_40610_4085# a_40565_4098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1698 gnd d0 a_36566_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1699 a_32637_n8762# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1700 gnd a_8768_n3805# a_8560_n3805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1701 a_8390_8213# a_8647_8023# a_8344_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1702 a_5342_292# a_10395_285# a_10603_285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1703 a_10878_n7793# a_10878_n7511# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1704 a_5525_n2485# a_6011_n2470# a_6219_n2470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1705 gnd a_35568_n7302# a_35360_n7302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1706 a_27008_n3536# a_27010_n3437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1707 a_32289_4592# a_32772_4757# a_32980_4757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1708 vdd d0 a_20340_3933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1709 a_21893_5730# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1710 gnd d3 a_19214_n4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 gnd a_8672_3125# a_8464_3125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1712 vdd d2 a_30119_1697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1713 a_27380_6688# a_27167_6688# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1714 a_20088_4361# a_20084_4538# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1715 a_16083_3405# a_16572_3223# a_16780_3223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1716 a_41643_n9879# a_41900_n9895# a_40634_n9457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1717 a_9427_3134# a_9439_2393# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1718 a_12120_7400# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1719 gnd a_4467_n9522# a_4259_n9522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1720 a_34031_7371# a_33610_7371# a_33932_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1721 vdd d1 a_24876_4098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1722 a_24636_1347# a_25697_976# a_25648_1166# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1723 a_8191_6588# a_8444_6575# a_8116_4663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1724 a_38962_n2683# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1725 a_20072_6882# a_20068_7059# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1726 vdd a_25881_6289# a_25673_6289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1727 a_10873_n8391# a_10880_n8190# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1728 a_902_n9764# a_481_n9764# a_205_n9463# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1729 gnd a_35216_n10397# a_35008_n10397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1730 a_2252_380# a_5134_292# a_5342_292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1731 a_19056_7240# a_19313_7050# a_19001_7801# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1732 a_1743_n2725# a_1530_n2725# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 a_7325_359# a_7112_359# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1734 a_34097_n4152# a_33884_n4152# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1735 gnd d0 a_25881_6289# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1736 a_10796_5597# a_11277_5767# a_11485_5767# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1737 a_26995_n6968# a_26993_n6754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1738 a_207_n9364# a_212_n8978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1739 a_27288_n2441# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1740 vdd a_41904_n8499# a_41696_n8499# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1741 a_17837_n5092# a_17455_n5653# a_16864_n5834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1742 a_31017_n3391# a_31013_n3579# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1743 a_5693_4196# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 a_36278_7466# a_36281_6874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1745 a_17634_3462# a_17421_3462# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1746 gnd d0 a_25868_7834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1747 vdd a_9748_n9501# a_9540_n9501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1748 a_11574_n7397# a_11153_n7397# a_10880_n7412# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1749 a_14913_n2883# a_15166_n3087# a_13900_n2649# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1750 a_16345_5746# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1751 a_20176_n5388# a_20429_n5592# a_19160_n5757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1752 gnd d3 a_24673_2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1753 gnd d2 a_3405_n9283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1754 a_2926_2869# a_3140_1747# a_3095_1760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1755 vdd a_3383_5103# a_3175_5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1756 a_5782_n5826# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1757 a_12469_n6106# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1758 gnd d0 a_15052_6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1759 a_37639_n9917# a_37637_n9703# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1760 a_8426_2159# a_9484_2380# a_9439_2393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1761 a_40573_2315# a_40830_2125# a_40527_1718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1762 a_32368_n7764# a_32368_n7482# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1763 a_32864_n5411# a_32651_n5411# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1764 gnd d0 a_20430_n6007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_37925_n7762# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_1491_1515# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_19025_3707# a_19120_4114# a_19075_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1768 a_6799_n4664# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_23436_n4144# a_23223_n4144# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1770 gnd a_35328_n6309# a_35120_n6309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1771 a_27600_4728# a_27179_4728# a_26909_4563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1772 a_39358_n8048# a_39145_n8048# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1773 vdd d0 a_25994_n2635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1774 a_16063_7040# a_16552_7140# a_16760_7140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1775 a_22417_n4837# a_21996_n4837# a_21720_n4536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1776 a_6125_1821# a_5704_1821# a_5436_1651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1777 a_37582_2611# a_38061_2779# a_38269_2779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1778 a_5417_4096# a_5906_4196# a_6114_4196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1779 a_17460_n4672# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1780 a_28683_1465# a_28262_1465# a_28589_1584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1781 a_32363_n8362# a_32370_n8161# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1782 a_714_n5847# a_501_n5847# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1783 a_12682_n6106# a_12469_n6106# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1784 a_25709_n8308# a_25962_n8512# a_24693_n8677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1785 a_10816_1085# a_11302_869# a_11510_869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1786 a_13799_3167# a_14857_3388# a_14808_3578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1787 a_16359_3223# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1788 gnd d0 a_25978_n5991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1789 a_4153_2176# a_4410_1986# a_3141_2357# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1790 a_38126_n9722# a_37913_n9722# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1791 vdd a_14141_n4813# a_13933_n4813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1792 vdd a_19325_5090# a_19117_5090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1793 a_23139_2047# a_22926_2047# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1794 a_10603_285# a_10182_285# a_5342_292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1795 a_19160_n5757# a_20221_n5592# a_20176_n5388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1796 gnd a_24970_n4776# a_24762_n4776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1797 a_10182_285# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1798 a_24611_6245# a_24868_6055# a_24565_5648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1799 a_7262_n7041# a_7207_n8069# a_7415_n8069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1800 a_29989_n5720# a_31050_n5555# a_31001_n5539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1801 a_16876_n3874# a_17680_n3693# a_17849_n3132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1802 a_5975_n9743# a_5762_n9743# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1803 a_1429_3055# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1804 a_136_4399# a_625_4217# a_833_4217# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1805 a_11595_n3895# a_11174_n3895# a_10898_n3594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1806 a_17435_n9570# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1807 a_23283_n3116# a_23070_n3116# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1808 a_32272_7032# a_32274_6933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1809 a_16578_1829# a_16365_1829# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1810 a_29846_5627# a_29941_6034# a_29892_6224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1811 a_23124_4983# a_22911_4983# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1812 a_6182_n9328# a_6987_n9562# a_7156_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1813 a_36391_n4814# a_36644_n5018# a_35378_n4580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1814 a_37644_n8936# a_38125_n9307# a_38333_n9307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1815 vdd a_8672_3125# a_8464_3125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1816 gnd a_24762_n4309# a_24554_n4309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 a_28792_n6048# a_28579_n6048# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1818 a_41586_2549# a_41589_1957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1819 a_30905_6458# a_31162_6268# a_29896_6047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1820 vdd a_36636_n6975# a_36428_n6975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1821 a_12630_n9030# a_12587_n8098# a_12795_n8098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1822 gnd a_15072_2409# a_14864_2409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1823 a_25623_6064# a_25880_5874# a_24611_6245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1824 a_28281_n6592# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1825 a_38270_3194# a_39074_3013# a_39233_3433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1826 a_38261_4736# a_37840_4736# a_37567_4952# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1827 a_239_n4265# a_237_n3868# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1828 a_32768_6153# a_32555_6153# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1829 a_21990_n5403# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1830 a_8483_n9478# a_8736_n9682# a_8433_n9058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_1887_n7062# a_1773_n7062# a_1981_n7062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1832 a_8187_6765# a_8444_6575# a_8116_4663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1833 gnd a_14148_n3834# a_13940_n3834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1834 a_242_n2605# a_244_n2506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1835 a_9508_n7752# a_9504_n7940# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1836 a_10399_n10484# a_15709_n10493# a_13568_n10410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1837 a_27008_n3818# a_27008_n3536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1838 a_11146_n8376# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1839 gnd d1 a_19320_6071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1840 a_5508_n6021# a_5506_n5807# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1841 a_6114_4196# a_6918_4015# a_7087_3573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1842 a_6105_5738# a_5684_5738# a_5411_5954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1843 a_27705_n3837# a_27284_n3837# a_27008_n3536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1844 a_27251_n9299# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1845 a_25732_n3600# a_25742_n2846# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1846 a_29901_5066# a_30959_5287# a_30914_5300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1847 a_16641_n8770# a_16428_n8770# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1848 a_31007_n4973# a_31010_n4370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1849 a_37950_n2864# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1850 a_28200_3005# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1851 a_32881_n2470# a_32668_n2470# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1852 a_5902_4757# a_5689_4757# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1853 gnd d2 a_19359_n7310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 a_4234_n5401# a_4230_n5589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1855 a_35061_6588# a_35259_7603# a_35210_7793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1856 vdd d3 a_24673_2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1857 a_11073_4225# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1858 a_33622_5411# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1859 vdd a_19429_n3813# a_19221_n3813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1860 a_9500_n8316# a_9496_n8504# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1861 a_23742_351# a_23321_351# a_23630_4439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1862 a_21727_n3557# a_22216_n3858# a_22424_n3858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1863 a_12434_n7070# a_12221_n7070# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1864 vdd d0 a_15052_6326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1865 a_23321_351# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1866 a_33073_n5826# a_32652_n5826# a_32376_n5525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1867 a_36399_n3042# a_36402_n2439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1868 a_3079_3897# a_3336_3707# a_2930_2692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1869 a_5798_n2470# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1870 vdd a_25977_n5576# a_25769_n5576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1871 a_39473_4426# a_39076_2501# a_39332_3433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1872 vdd d1 a_24893_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1873 a_28405_4962# a_28192_4962# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1874 gnd a_9672_6297# a_9464_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1875 a_32274_6933# a_32281_6549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1876 a_824_5759# a_403_5759# a_135_5589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1877 a_16166_n6410# a_16652_n6395# a_16860_n6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1878 a_36277_8270# a_36530_8257# a_35264_8036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1879 a_3203_n8706# a_4264_n8541# a_4215_n8525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1880 vdd d1 a_30169_2117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1881 a_22428_n2462# a_23233_n2696# a_23392_n2939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1882 a_28816_6410# a_28395_6410# a_28651_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1883 gnd d1 a_24977_n3797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1884 a_412_4217# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1885 vdd d0 a_31166_4872# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1886 vdd d0 a_4500_n4060# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1887 a_21638_2128# a_22127_2228# a_22335_2228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1888 gnd d1 a_14128_n7751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1889 a_28552_n5055# a_28339_n5055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1890 vdd a_36650_n3624# a_36442_n3624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1891 gnd d0 a_25885_4893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1892 a_217_n7785# a_706_n7804# a_914_n7804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1893 a_25718_n6951# a_25975_n6967# a_24709_n6529# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1894 a_38249_6696# a_39054_6930# a_39213_7350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1895 a_23233_n2696# a_23020_n2696# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1896 a_41562_6853# a_41558_7030# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1897 gnd a_40615_2637# a_40407_2637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1898 gnd d0 a_31161_5853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1899 a_28572_3425# a_28463_3425# a_28671_3425# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1900 a_28658_n7012# a_28544_n7012# a_28752_n7012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 vdd a_3492_n2845# a_3284_n2845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1902 vdd d2 a_8718_n3385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1903 a_5673_8113# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1904 a_12179_n4693# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1905 a_8484_n8685# a_9545_n8520# a_9500_n8316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1906 gnd a_40609_n6288# a_40401_n6288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1907 vdd a_4398_3946# a_4190_3946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1908 a_16434_n7376# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1909 a_16152_n8469# a_16641_n8770# a_16849_n8770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1910 a_14908_n2656# a_15165_n2672# a_13896_n2837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1911 gnd d4 a_8458_n6309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1912 gnd d0 a_15056_4930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1913 a_8433_n9058# a_8686_n9262# a_8280_n8030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1914 a_3019_n4134# a_3272_n4338# a_2920_n6314# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1915 gnd d2 a_24895_n9254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1916 a_24688_n9658# a_24945_n9674# a_24642_n9050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1917 a_919_n6823# a_1723_n6642# a_1882_n6885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1918 a_35226_5656# a_35479_5643# a_35057_6765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1919 a_485_n8368# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 vdd d1 a_30263_n2795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1921 a_27272_n5797# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1922 a_8296_n4301# a_8510_n3385# a_8461_n3369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1923 vdd a_41835_2923# a_41627_2923# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1924 a_1801_3475# a_1429_3055# a_838_3236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1925 a_3095_1760# a_3190_2167# a_3145_2180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1926 a_23114_6431# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1927 a_11498_2829# a_11077_2829# a_10811_2661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1928 a_24608_7047# a_24861_7034# a_24549_7785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1929 a_8406_6076# a_9464_6297# a_9419_6310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1930 a_27001_n4515# a_27490_n4816# a_27698_n4816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1931 a_29846_5627# a_29941_6034# a_29896_6047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1932 a_40267_4642# a_40520_4629# a_39585_338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1933 a_5434_1437# a_5434_1155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1934 a_14787_8299# a_15040_8286# a_13774_8065# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1935 a_23459_n8993# a_23038_n8993# a_23365_n8993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1936 a_38911_3433# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1937 a_1733_n4173# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1938 a_33855_1494# a_33642_1494# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1939 gnd a_30251_n4755# a_30043_n4755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1940 a_5525_n2485# a_5181_n2252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1941 vdd d0 a_4487_n5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1942 a_36309_1174# a_32313_855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1943 a_22204_n5818# a_21991_n5818# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1944 a_16179_n3573# a_16668_n3874# a_16876_n3874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1945 gnd a_36566_984# a_36358_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1946 a_8296_n4301# a_8553_n4317# a_8201_n6293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1947 vdd a_31150_8228# a_30942_8228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1948 a_3121_6274# a_4182_5903# a_4133_6093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1949 a_28289_n4635# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1950 a_21620_6541# a_21618_6327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1951 a_14807_3163# a_14819_2422# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1952 vdd a_19379_n3393# a_19171_n3393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1953 gnd d0 a_41816_7255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1954 a_29884_8007# a_30942_8228# a_30893_8418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1955 a_5399_7914# a_5885_7698# a_6093_7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1956 gnd d1 a_35606_n9682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1957 a_37562_6528# a_38041_6696# a_38249_6696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1958 a_8491_n7706# a_9552_n7541# a_9503_n7525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1959 gnd d0 a_9671_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1960 a_28663_5382# a_28242_5382# a_28569_5501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1961 a_33001_1255# a_32580_1255# a_32304_1437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1962 gnd d1 a_40818_4085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1963 a_20162_n8739# a_20158_n8927# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1964 vdd d1 a_19320_6071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1965 a_17735_n3132# a_17522_n3132# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1966 a_39339_n3103# a_38957_n3664# a_38365_n3430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 a_8280_n8030# a_8533_n8234# a_8205_n6105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1968 a_37669_n3544# a_37671_n3445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1969 vdd a_24876_4098# a_24668_4098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1970 a_32877_n3866# a_32664_n3866# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1971 a_34986_4663# a_35239_4650# a_34304_359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_6130_840# a_5709_840# a_5436_1056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1973 a_25732_n3600# a_25989_n3616# a_24720_n3781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1974 a_3146_1376# a_4207_1005# a_4162_1018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1975 a_13744_3728# a_13839_4135# a_13790_4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1976 a_3222_n5582# a_4280_n6020# a_4231_n6004# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1977 a_33084_n3451# a_33889_n3685# a_34058_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1978 a_29951_n3340# a_30208_n3356# a_29786_n4272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1979 gnd d0 a_20321_8265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1980 a_17723_7379# a_17614_7379# a_17822_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1981 a_30917_4324# a_30913_4501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1982 a_27167_6688# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1983 a_16065_7536# a_16546_7706# a_16754_7706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1984 a_6994_n8069# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1985 a_17467_n3693# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1986 a_1580_n3145# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1987 a_20173_n6364# a_20169_n6552# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1988 vdd d0 a_15153_n4632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1989 gnd d2 a_14078_n7331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1990 a_28752_n7012# a_28697_n8040# a_28905_n8040# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1991 a_17421_3462# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1992 a_27465_n9714# a_27252_n9714# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1993 a_17626_5419# a_17413_5419# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 a_25716_n7329# a_25969_n7533# a_24700_n7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1995 a_36374_n7940# a_36631_n7956# a_35365_n7518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1996 a_12365_1523# a_12152_1523# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1997 gnd a_25868_7834# a_25660_7834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1998 a_35385_n3601# a_35638_n3805# a_35335_n3181# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1999 a_6774_n9562# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2000 a_10399_n10484# a_10656_n10500# a_10498_n10484# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2001 a_33089_n2470# a_32668_n2470# a_31952_n2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2002 a_38130_n8326# a_37917_n8326# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2003 a_37912_n9307# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2004 a_27690_n6773# a_28494_n6592# a_28653_n6835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2005 a_29994_n4739# a_30251_n4755# a_29939_n5300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2006 a_22392_n9735# a_21971_n9735# a_21695_n9716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2007 a_4236_n5023# a_4493_n5039# a_3227_n4601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2008 gnd a_15052_6326# a_14844_6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2009 a_22106_5730# a_21893_5730# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2010 a_22303_8105# a_21882_8105# a_21606_8287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2011 a_9508_n6544# a_9516_n5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2012 a_24638_n9238# a_24895_n9254# a_24489_n8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2013 a_6131_1255# a_6935_1074# a_7094_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2014 a_11178_n2499# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2015 vdd d1 a_40919_n3784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2016 a_4999_n10469# a_5256_n10485# a_5098_n10469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2017 a_39213_n5063# a_39000_n5063# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2018 a_32995_1821# a_33800_2055# a_33969_1613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2019 a_41585_2134# a_41595_1391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2020 a_12442_n5113# a_12229_n5113# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2021 a_37657_n5504# a_38146_n5805# a_38354_n5805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2022 a_16787_2244# a_16366_2244# a_16090_2426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2023 a_21894_6145# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2024 a_32284_5354# a_32773_5172# a_32981_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2025 a_23360_n8816# a_22988_n8573# a_22397_n8754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2026 a_33964_1494# a_33592_1074# a_33000_840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2027 a_25640_2949# a_25636_3126# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2028 gnd d0 a_15160_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2029 a_39319_n7020# a_39205_n7020# a_39413_n7020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2030 gnd a_40907_n5744# a_40699_n5744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2031 a_23132_3026# a_22919_3026# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2032 vdd a_3417_n7323# a_3209_n7323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2033 a_219_n7404# a_224_n7018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2034 a_36361_n9485# a_36618_n9501# a_35349_n9666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2035 a_40352_n6272# a_40496_n4296# a_40447_n4280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2036 a_19122_n3377# a_19226_n2832# a_19181_n2628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2037 gnd a_31244_n8906# a_31036_n8906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2038 gnd d1 a_8756_n5765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2039 a_22003_n3858# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2040 a_22221_n2877# a_22008_n2877# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2041 vdd d0 a_41936_n2622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2042 a_6965_5411# a_6752_5411# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2043 a_35222_5833# a_35479_5643# a_35057_6765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2044 gnd a_40780_1705# a_40572_1705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2045 a_4127_7487# a_4384_7297# a_3118_7076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2046 a_30913_4501# a_30916_3909# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2047 a_32981_5172# a_33785_4991# a_33944_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2048 a_939_n2906# a_518_n2906# a_242_n2887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2049 a_28408_3986# a_28195_3986# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2050 a_1773_n7062# a_1560_n7062# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2051 vdd d2 a_30196_n5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2052 a_11167_n4874# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2053 a_24604_7224# a_24861_7034# a_24549_7785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2054 gnd a_9676_4901# a_9468_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2055 a_12801_4476# a_12380_4476# a_12702_4476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2056 a_38358_n4409# a_39163_n4643# a_39322_n4886# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2057 a_35335_n3181# a_35430_n3805# a_35385_n3601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2058 a_17837_n5092# a_17455_n5653# a_16863_n5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2059 a_27288_n2441# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2060 a_3129_4317# a_3386_4127# a_3083_3720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2061 a_29916_2130# a_30169_2117# a_29866_1710# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2062 a_10789_6364# a_11278_6182# a_11486_6182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2063 a_19025_3707# a_19278_3694# a_18872_2679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2064 a_16648_n7791# a_16435_n7791# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2065 a_32378_n6021# a_32861_n6387# a_33069_n6387# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2066 a_14783_8476# a_15040_8286# a_13774_8065# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2067 a_36281_6874# a_36534_6861# a_35265_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2068 a_16169_n5434# a_16655_n5419# a_16863_n5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2069 a_40565_4098# a_41623_4319# a_41578_4332# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2070 a_16571_2808# a_16358_2808# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2071 a_38257_6132# a_39061_5951# a_39230_5509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2072 a_20189_n2635# a_20446_n2651# a_19177_n2816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2073 gnd d4 a_13838_n6338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2074 a_12548_n7070# a_12166_n7631# a_11575_n7812# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2075 a_39269_6418# a_39056_6418# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2076 gnd d4 a_29859_4621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2077 a_31889_n10455# a_32146_n10471# a_21397_n10599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2078 a_11582_n5440# a_12387_n5674# a_12556_n5113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2079 a_24674_n3173# a_24769_n3797# a_24720_n3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2080 gnd d0 a_25888_3917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2081 a_9407_7051# a_9419_6310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2082 vdd d0 a_41816_7255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2083 vdd d8 a_21654_n10615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2084 a_16365_1829# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2085 a_32761_7132# a_32548_7132# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2086 a_28393_6922# a_28180_6922# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2087 gnd a_20422_n7964# a_20214_n7964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2088 a_4125_7876# a_4378_7863# a_3109_8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2089 a_9524_n4023# a_9781_n4039# a_8515_n3601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2090 gnd d1 a_8652_7042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2091 vdd d1 a_40818_4085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2092 a_41666_n5359# a_41662_n5547# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2093 a_27395_3752# a_27182_3752# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2094 a_16861_n6810# a_16440_n6810# a_16164_n6509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2095 a_35335_n3181# a_35588_n3385# a_35166_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2096 a_39661_n6056# a_40497_n10376# a_37150_n10448# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2097 a_11587_n4459# a_11166_n4459# a_10900_n4273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2098 vdd a_25990_n4031# a_25782_n4031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2099 a_13779_7084# a_14837_7305# a_14792_7318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2100 a_32555_6153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2101 a_28187_5943# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2102 a_35285_3315# a_36346_2944# a_36301_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2103 a_29681_6559# a_29934_6546# a_29606_4634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2104 a_14896_n5824# a_15149_n6028# a_13883_n5590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2105 a_22119_2792# a_21906_2792# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2106 a_128_6074# a_617_6174# a_825_6174# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2107 a_34982_4840# a_35239_4650# a_34304_359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2108 vdd a_15141_n7985# a_14933_n7985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2109 a_19090_n9254# a_19347_n9270# a_18941_n8038# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2110 a_13744_3728# a_13839_4135# a_13794_4148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2111 a_9438_1978# a_9691_1965# a_8422_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2112 a_17760_1621# a_17378_2063# a_16786_1829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2113 a_12561_3483# a_12140_3483# a_12462_3483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2114 a_3219_n6558# a_4277_n6996# a_4228_n6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2115 gnd d1 a_40887_n9661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2116 vdd d0 a_20321_8265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2117 a_35280_4296# a_36341_3925# a_36292_4115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2118 a_28658_n7012# a_28276_n7573# a_27685_n7754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2119 a_4125_7876# a_4121_8053# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2120 a_32648_n6387# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2121 a_31001_n5539# a_31011_n4785# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2122 a_37573_3376# a_38062_3194# a_38270_3194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2123 gnd a_19414_n6749# a_19206_n6749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2124 a_18848_6773# a_19062_5651# a_19013_5841# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2125 vdd d2 a_40869_n3364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2126 a_714_n5847# a_501_n5847# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2127 a_14791_6903# a_15044_6890# a_13775_7261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2128 a_34285_n8069# a_33864_n8069# a_34120_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2129 a_19075_4127# a_20133_4348# a_20088_4361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2130 a_13790_4325# a_14851_3954# a_14806_3967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2131 a_21907_3207# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2132 a_38126_n9722# a_37913_n9722# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2133 a_12171_n6650# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2134 a_24416_2840# a_24630_1718# a_24585_1731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2135 a_28319_n8972# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2136 a_40523_1895# a_40627_1144# a_40578_1334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2137 a_13492_4869# a_13636_2687# a_13587_2877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2138 a_25641_3364# a_25894_3351# a_24628_3130# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2139 a_34026_n9001# a_33644_n9562# a_33053_n9743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2140 a_23223_n4144# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2141 a_16455_n3874# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2142 a_11386_n3480# a_11173_n3480# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2143 gnd a_19290_1734# a_19082_1734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2144 a_9511_n5568# a_9768_n5584# a_8499_n5749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2145 gnd a_4492_n4624# a_4284_n4624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2146 a_36393_n3608# a_36403_n2854# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2147 vdd a_15052_6326# a_14844_6326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2148 a_29885_7203# a_30946_6832# a_30897_7022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2149 gnd a_40857_n5324# a_40649_n5324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2150 a_11271_7161# a_11058_7161# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2151 a_6105_5738# a_6910_5972# a_7079_5530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2152 vdd d0 a_20434_n4611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2153 a_27188_3186# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2154 a_29919_n9217# a_30176_n9233# a_29770_n8001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2155 a_20170_n6967# a_20173_n6364# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2156 a_32393_n2866# a_32882_n2885# a_33090_n2885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2157 vdd a_24893_1157# a_24685_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2158 vdd d0 a_25869_8249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2159 a_28192_4962# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2160 a_2021_n6098# a_1808_n6098# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2161 a_40666_n3580# a_40919_n3784# a_40616_n3160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2162 a_16154_n8965# a_16152_n8751# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2163 gnd d0 a_31263_n4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2164 a_136_4117# a_138_4018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2165 a_5181_n2252# a_6011_n2470# a_6219_n2470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2166 a_36297_3134# a_36309_2393# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2167 a_10802_3144# a_11291_3244# a_11499_3244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2168 gnd a_36635_n6560# a_36427_n6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2169 a_6183_n9743# a_6987_n9562# a_7156_n9001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2170 a_35166_n4301# a_35380_n3385# a_35335_n3181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2171 a_10880_n8190# a_11359_n8376# a_11567_n8376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2172 gnd a_30243_n6712# a_30035_n6712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2173 a_37639_n9322# a_38125_n9307# a_38333_n9307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2174 vdd a_31166_4872# a_30958_4872# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2175 gnd d5 a_19007_n10405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2176 a_21618_6045# a_21620_5946# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2177 a_8496_n6725# a_8753_n6741# a_8441_n7286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2178 a_27375_7669# a_27162_7669# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2179 a_21990_n5403# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2180 a_38262_5151# a_37841_5151# a_37565_5051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2181 a_40495_7595# a_40748_7582# a_40342_6567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2182 a_33676_n3685# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2183 a_16875_n3459# a_16454_n3459# a_16186_n3088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2184 a_6925_2522# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2185 a_39572_4426# a_39476_338# a_37394_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2186 a_36371_n8731# a_36367_n8919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2187 a_13884_n4797# a_14945_n4632# a_14900_n4428# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2188 a_12479_1642# a_12365_1523# a_12573_1523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2189 a_10885_n7026# a_10883_n6812# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2190 a_4138_6331# a_4134_6508# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2191 a_642_1276# a_429_1276# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2192 a_28484_n8040# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2193 a_11146_n8376# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2194 a_23070_n3116# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2195 a_17740_5538# a_17358_5980# a_16767_6161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2196 a_29981_n7677# a_31042_n7512# a_30997_n7308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2197 gnd a_3455_n9703# a_3247_n9703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2198 a_5342_292# a_4921_292# a_5243_292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 a_7213_4447# a_7000_4447# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2200 a_212_n8383# a_698_n8368# a_906_n8368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2201 a_24713_n4760# a_25774_n4595# a_25725_n4579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2202 gnd d0 a_20441_n3632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2203 a_16546_7706# a_16333_7706# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2204 gnd a_15056_4930# a_14848_4930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2205 a_29766_n8189# a_30023_n8205# a_29695_n6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2206 a_6106_6153# a_5685_6153# a_5409_6053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2207 a_28264_n9533# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2208 a_37950_n2864# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2209 a_20096_2578# a_20353_2388# a_19087_2167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2210 a_6930_2055# a_6717_2055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2211 a_33894_n2704# a_33681_n2704# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2212 a_22919_3026# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2213 vdd d4 a_29859_4621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2214 a_23416_n8061# a_23203_n8061# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2215 a_16080_4005# a_16085_3619# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2216 a_40630_n9645# a_40887_n9661# a_40584_n9037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2217 gnd d2 a_40837_n9241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2218 a_8395_7232# a_9456_6861# a_9411_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2219 a_30924_2126# a_31181_1936# a_29912_2307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2220 a_11491_5201# a_11070_5201# a_10794_5383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2221 gnd d1 a_3460_n8722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2222 a_32378_n6021# a_32376_n5807# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2223 a_40616_n3160# a_40711_n3784# a_40666_n3580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2224 gnd d1 a_24873_5074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2225 vdd d1 a_8652_7042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2226 a_2926_2869# a_3183_2679# a_2831_4861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2227 a_16075_5080# a_16077_4981# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2228 a_37843_3760# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2229 a_36381_n5568# a_36391_n4814# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2230 vdd d0 a_36651_n4039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2231 a_37594_834# a_38073_819# a_38281_819# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2232 a_39155_n6600# a_38942_n6600# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2233 a_237_n3868# a_237_n3586# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2234 a_39344_1473# a_38923_1473# a_39250_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2235 a_38151_n4824# a_37938_n4824# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2236 a_7176_n5084# a_6794_n5645# a_6203_n5826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2237 a_32579_840# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2238 a_8390_8213# a_9451_7842# a_9402_8032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2239 a_29677_6736# a_29934_6546# a_29606_4634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2240 a_39562_n5879# a_39165_n4131# a_39421_n5063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2241 gnd a_41816_7255# a_41608_7255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2242 a_11499_3244# a_12303_3063# a_12462_3483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2243 a_38992_n7020# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2244 a_13891_n3818# a_14952_n3653# a_14903_n3637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2245 a_39566_n8048# a_39453_n6056# a_39661_n6056# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_16083_3123# a_16085_3024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2247 a_13680_n4142# a_13933_n4346# a_13581_n6322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2248 gnd a_40818_4085# a_40610_4085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2249 vdd d3 a_40704_n4296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2250 a_8453_n5141# a_8548_n5765# a_8499_n5749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2251 a_40667_n2787# a_41728_n2622# a_41683_n2418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2252 vdd a_24907_n7294# a_24699_n7294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2253 a_10395_285# a_10182_285# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2254 a_37548_8274# a_37548_7992# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2255 a_27595_5709# a_27174_5709# a_26901_5925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2256 gnd a_9679_3925# a_9471_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2257 a_35150_n8030# a_35348_n9262# a_35299_n9246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2258 a_16339_7140# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2259 gnd a_40760_5622# a_40552_5622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2260 a_40616_n3160# a_40869_n3364# a_40447_n4280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2261 a_18848_6773# a_19062_5651# a_19017_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2262 gnd a_9785_n2643# a_9577_n2643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2263 vdd a_31271_n4010# a_31063_n4010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2264 a_23263_n7033# a_23050_n7033# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2265 a_6905_6439# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2266 a_5500_n8161# a_5498_n7764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2267 gnd d0 a_41919_n5563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2268 a_18076_n8077# a_17655_n8077# a_17923_n7049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 a_17596_1082# a_17383_1082# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2270 a_19005_7624# a_19258_7611# a_18852_6596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2271 a_6200_n6802# a_5779_n6802# a_5503_n6783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2272 a_37938_n4824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2273 a_5917_1821# a_5704_1821# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2274 a_30999_n6930# a_31002_n6327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2275 a_12454_5440# a_12345_5440# a_12553_5440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2276 a_10796_5597# a_10794_5383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2277 a_40523_1895# a_40627_1144# a_40582_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2278 a_25637_3541# a_25894_3351# a_24628_3130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2279 a_16434_n7376# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2280 a_41591_1568# a_41594_976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2281 gnd d0 a_31181_1936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2282 a_18171_n6085# a_17750_n6085# a_18076_n8077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2283 vdd a_19290_1734# a_19082_1734# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2284 a_30912_4086# a_30922_3343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2285 a_5500_n7383# a_5986_n7368# a_6194_n7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2286 a_12392_n4693# a_12179_n4693# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2287 a_17413_5419# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2288 vdd d0 a_36638_n5584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2289 a_12152_1523# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2290 a_16167_n5815# a_16167_n5533# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2291 a_28901_n5871# a_28504_n4123# a_28772_n3095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2292 a_16090_2426# a_16090_2144# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2293 a_35071_n6293# a_35215_n4317# a_35170_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2294 a_11297_1850# a_11084_1850# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2295 a_36314_1412# a_36567_1399# a_35301_1178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2296 a_28443_7342# a_28230_7342# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2297 a_27001_n4797# a_27490_n4816# a_27698_n4816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2298 a_26889_7885# a_26894_7499# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2299 a_41672_n4793# a_41925_n4997# a_40659_n4559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2300 vdd d1 a_40798_8002# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2301 a_9419_5091# a_9676_4901# a_8407_5272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2302 a_41558_8249# a_41554_8426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2303 a_12454_5440# a_12082_5020# a_11490_4786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2304 a_6119_3215# a_5698_3215# a_5422_3397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2305 a_16077_4981# a_16080_4600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2306 a_16447_n4438# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2307 a_35369_n5749# a_36430_n5584# a_36381_n5568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2308 a_16179_n3855# a_16668_n3874# a_16876_n3874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2309 a_4151_3393# a_4147_3570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2310 a_16780_3223# a_16359_3223# a_16083_3405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2311 a_5134_292# a_4921_292# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2312 a_21918_832# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2313 a_40491_7772# a_40748_7582# a_40342_6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2314 vdd d1 a_35623_n6741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2315 a_38264_3760# a_39069_3994# a_39238_3552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2316 vdd d0 a_41810_7821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2317 a_29896_6047# a_30954_6268# a_30909_6281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2318 a_6187_n8347# a_5766_n8347# a_5493_n8362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2319 a_11478_6746# a_12283_6980# a_12442_7400# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2320 a_37553_7293# a_38042_7111# a_38250_7111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2321 a_3141_2357# a_4202_1986# a_4153_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2322 a_1409_6972# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2323 gnd d3 a_40595_6554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2324 a_40447_n4280# a_40661_n3364# a_40616_n3160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2325 a_24729_n2612# a_25787_n3050# a_25742_n2846# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2326 a_121_7335# a_121_7053# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2327 a_39145_n8048# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2328 a_17653_n8589# a_17440_n8589# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2329 vdd a_41900_n9895# a_41692_n9895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2330 a_838_3236# a_417_3236# a_141_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2331 a_25737_n3827# a_25733_n4015# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2332 a_37580_2115# a_37582_2016# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2333 gnd d0 a_9691_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2334 a_28772_n3095# a_28351_n3095# a_28673_n2918# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2335 gnd d0 a_36541_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2336 a_16641_n8770# a_16428_n8770# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2337 a_38942_n6600# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2338 a_1969_n9022# a_1926_n8090# a_2134_n8090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2339 a_24585_1731# a_24680_2138# a_24635_2151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2340 a_14799_6339# a_14795_6516# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2341 a_6752_5411# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2342 a_38250_7111# a_39054_6930# a_39213_7350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2343 a_28195_3986# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2344 gnd a_3252_n8255# a_3044_n8255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2345 a_7019_n3685# a_6806_n3685# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2346 a_5897_5738# a_5684_5738# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2347 a_8300_n4113# a_8498_n5345# a_8449_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2348 a_27168_7103# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2349 a_6214_n3451# a_5793_n3451# a_5520_n3466# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2350 a_32669_n2885# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2351 a_16058_8303# a_16547_8121# a_16755_8121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2352 a_37570_3976# a_38056_3760# a_38264_3760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2353 a_27015_n3051# a_27013_n2837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2354 a_13756_1768# a_14009_1755# a_13587_2877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2355 a_19068_5280# a_20129_4909# a_20080_5099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2356 vdd d1 a_24873_5074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2357 vdd d0 a_9774_n5018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2358 a_10814_1184# a_10816_1085# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2359 a_8483_n9478# a_9541_n9916# a_9492_n9900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2360 a_5798_n2470# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2361 a_17680_n3693# a_17467_n3693# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2362 a_39056_6418# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2363 vdd a_31169_3896# a_30961_3896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2364 a_6774_n9562# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2365 a_21633_3008# a_21640_2624# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2366 a_24611_6245# a_25672_5874# a_25623_6064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2367 a_38130_n8326# a_37917_n8326# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2368 a_37912_n9307# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2369 a_6094_8113# a_6898_7932# a_7067_7490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2370 a_26889_7885# a_27375_7669# a_27583_7669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2371 vdd a_41816_7255# a_41608_7255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2372 a_14791_6903# a_14787_7080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2373 a_28180_6922# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2374 a_22392_n9735# a_21971_n9735# a_21695_n9434# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2375 gnd a_25975_n6967# a_25767_n6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2376 vdd a_8533_n8234# a_8325_n8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2377 gnd d0 a_9754_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2378 a_36379_n6959# a_36382_n6356# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2379 a_4147_3570# a_4150_2978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2380 a_23194_1486# a_22981_1486# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2381 a_21620_6541# a_22099_6709# a_22307_6709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2382 vdd a_40818_4085# a_40610_4085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2383 a_27182_3752# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2384 a_17743_3462# a_17371_3042# a_16779_2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2385 vdd a_36530_8257# a_36322_8257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2386 a_16563_4765# a_16350_4765# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2387 a_14814_2184# a_15071_1994# a_13802_2365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2388 a_32844_n9328# a_32631_n9328# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2389 vdd a_14116_n9711# a_13908_n9711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2390 a_32388_n3847# a_32388_n3565# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2391 a_40545_8015# a_40798_8002# a_40495_7595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2392 vdd a_40760_5622# a_40552_5622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2393 a_6992_n8581# a_6779_n8581# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2394 vdd d0 a_36566_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2395 a_17923_n7049# a_17502_n7049# a_17829_n7049# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2396 gnd d0 a_25889_4332# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 gnd a_24945_n9674# a_24737_n9674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2398 a_37657_n5786# a_38146_n5805# a_38354_n5805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2399 gnd d0 a_20358_1407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2400 a_23360_n8816# a_22988_n8573# a_22396_n8339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2401 a_36309_1174# a_36566_984# a_35297_1355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2402 a_19001_7801# a_19258_7611# a_18852_6596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2403 vdd d1 a_24970_n4776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2404 a_34140_n5084# a_33719_n5084# a_34046_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2405 a_22221_n2877# a_22008_n2877# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2406 a_8356_5656# a_8609_5643# a_8187_6765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2407 a_40431_n8009# a_40629_n9241# a_40580_n9225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2408 a_9500_n8316# a_9753_n8520# a_8484_n8685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2409 a_32383_n4445# a_32390_n4244# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2410 a_35269_7055# a_36327_7276# a_36278_7466# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2411 a_30982_n9871# a_31239_n9887# a_29973_n9449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2412 a_939_n2906# a_518_n2906# a_242_n2605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2413 a_485_n8368# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2414 a_11167_n4874# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2415 a_38359_n4824# a_39163_n4643# a_39322_n4886# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2416 a_35234_3699# a_35329_4106# a_35280_4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2417 gnd a_14098_n3414# a_13890_n3414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2418 a_35385_n3601# a_36443_n4039# a_36398_n3835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2419 a_37555_7507# a_38036_7677# a_38244_7677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2420 gnd a_9696_984# a_9488_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2421 a_41578_3113# a_41835_2923# a_40566_3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2422 a_13568_n10410# a_13518_n10426# a_12890_n6106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2423 a_12548_n7070# a_12166_n7631# a_11574_n7397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2424 vdd a_40520_4629# a_40312_4629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2425 a_19114_n5149# a_19209_n5773# a_19164_n5569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2426 a_20739_n805# a_20526_n805# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2427 a_41565_6051# a_41575_5308# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2428 a_22204_n5818# a_21991_n5818# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2429 a_11583_n5855# a_12387_n5674# a_12556_n5113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2430 a_16652_n6395# a_16439_n6395# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2431 a_2926_2869# a_3140_1747# a_3091_1937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2432 a_13774_8065# a_14832_8286# a_14783_8476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2433 vdd a_40899_n7701# a_40691_n7701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2434 gnd d0 a_4485_n6996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2435 a_512_n3472# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2436 gnd a_35631_n4784# a_35423_n4784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2437 vdd d1 a_8748_n7722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2438 gnd a_8553_n4317# a_8345_n4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2439 vdd d3 a_40595_6554# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2440 a_12209_n9030# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2441 a_5505_n6402# a_5508_n6021# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2442 a_30010_n2591# a_31068_n3029# a_31023_n2825# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2443 gnd d0 a_9768_n5584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2444 a_27162_7669# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2445 gnd a_15140_n7570# a_14932_n7570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2446 a_40650_n5728# a_41711_n5563# a_41662_n5547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2447 a_17723_7379# a_17351_6959# a_16760_7140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2448 a_13568_n10410# a_15917_n10493# a_10399_n10484# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2449 a_19161_n6545# a_20219_n6983# a_20174_n6779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2450 a_29905_3286# a_30162_3096# a_29850_3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2451 a_13496_4692# a_13616_6604# a_13571_6617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2452 a_10504_285# a_15582_300# a_15904_300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2453 a_39433_n3103# a_39012_n3103# a_39334_n2926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2454 a_29990_n6508# a_31048_n6946# a_30999_n6930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2455 a_5773_n7368# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2456 a_23491_n3116# a_23436_n4144# a_23620_n5892# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2457 a_17490_n9009# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2458 a_15582_300# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 a_28658_n7012# a_28276_n7573# a_27684_n7339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2460 a_32306_1651# a_32304_1437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2461 a_26912_3368# a_26912_3086# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2462 a_24619_4288# a_24876_4098# a_24573_3691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2463 a_12345_5440# a_12132_5440# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2464 a_32292_3397# a_32292_3115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2465 vdd a_14066_n9291# a_13858_n9291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2466 a_13752_1945# a_14009_1755# a_13587_2877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2467 a_16333_7706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2468 a_36294_5329# a_36547_5316# a_35281_5095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2469 a_37930_n6781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2470 vdd a_31275_n2614# a_31067_n2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2471 a_20088_3142# a_20345_2952# a_19076_3323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2472 a_21611_7306# a_21611_7024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2473 a_22315_6145# a_23119_5964# a_23288_5522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2474 a_22403_n7360# a_23208_n7594# a_23377_n7033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2475 vdd d5 a_40497_n10376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2476 a_28319_n8972# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2477 a_33089_n2470# a_32668_n2470# a_32395_n2485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2478 a_1441_1095# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2479 a_32780_2800# a_32567_2800# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2480 a_35296_2159# a_35549_2146# a_35246_1739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2481 a_34026_n9001# a_33644_n9562# a_33052_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2482 a_16455_n3874# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2483 gnd d5 a_13726_n10426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2484 a_9520_n4399# a_9516_n4587# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2485 a_25615_7847# a_25868_7834# a_24599_8205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2486 a_9418_5895# a_9414_6072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2487 a_12399_n3714# a_12186_n3714# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2488 gnd a_24873_5074# a_24665_5074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2489 a_20087_3946# a_20340_3933# a_19071_4304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2490 a_24704_n7510# a_24957_n7714# a_24654_n7090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2491 a_24420_2663# a_24673_2650# a_24321_4832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2492 gnd d4 a_35239_4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2493 a_35311_n7286# a_35415_n6741# a_35370_n6537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2494 a_35058_n10381# a_35008_n10397# a_34380_n6077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2495 a_4222_n7546# a_4479_n7562# a_3210_n7727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2496 a_38061_2779# a_37848_2779# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2497 a_18866_n6113# a_18986_n8242# a_18937_n8226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2498 a_5486_n9442# a_5488_n9343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2499 a_35374_n4768# a_35631_n4784# a_35319_n5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2500 vdd a_4487_n5605# a_4279_n5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2501 a_12154_n9591# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2502 a_41658_n7316# a_41654_n7504# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2503 a_16759_6725# a_16338_6725# a_16065_6941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2504 vdd d0 a_25889_4332# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2505 a_10873_n8391# a_11359_n8376# a_11567_n8376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2506 a_14883_n7554# a_15140_n7570# a_13871_n7735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2507 a_6113_3781# a_5692_3781# a_5419_3997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2508 a_16673_n2893# a_16460_n2893# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2509 a_30909_6281# a_31162_6268# a_29896_6047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2510 vdd a_13913_n8263# a_13705_n8263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2511 a_5910_2800# a_5697_2800# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2512 a_37676_n2464# a_38162_n2449# a_38370_n2449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2513 a_25621_7281# a_25617_7458# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2514 a_16771_4765# a_17576_4999# a_17735_5419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2515 a_1713_n8090# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2516 a_18961_n4121# a_19159_n5353# a_19114_n5149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2517 a_33969_1613# a_33587_2055# a_32996_2236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2518 a_23643_351# a_24370_4642# a_24321_4832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2519 a_35058_n10381# a_37407_n10464# a_31889_n10455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2520 a_16880_n2478# a_17685_n2712# a_17844_n2955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2521 a_5980_n8762# a_5767_n8762# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2522 a_27376_8084# a_27163_8084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2523 a_8352_5833# a_8609_5643# a_8187_6765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2524 a_11600_n2914# a_11179_n2914# a_10903_n2895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2525 vdd a_40849_n7281# a_40641_n7281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2526 a_26976_n9413# a_27465_n9714# a_27673_n9714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2527 a_35269_7055# a_36327_7276# a_36282_7289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2528 a_39218_7469# a_39104_7350# a_39312_7350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2529 a_14804_5358# a_15057_5345# a_13791_5124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2530 a_28509_n3656# a_28296_n3656# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2531 a_17383_1082# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2532 a_5704_1821# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2533 vdd a_3472_n6762# a_3264_n6762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2534 gnd d0 a_36623_n8520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2535 a_19181_n2628# a_19434_n2832# a_19122_n3377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2536 gnd a_30226_n9653# a_30018_n9653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2537 gnd a_4468_n9937# a_4260_n9937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2538 a_13806_2188# a_14059_2175# a_13756_1768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2539 a_11290_2829# a_11077_2829# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2540 vdd d6 a_5256_n10485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2541 a_27595_5709# a_28400_5943# a_28569_5501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2542 a_832_3802# a_411_3802# a_143_3632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2543 vdd d0 a_31255_n6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2544 a_28264_n9533# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2545 a_16174_n5048# a_16655_n5419# a_16863_n5419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2546 a_16547_8121# a_16334_8121# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2547 a_5416_4973# a_5902_4757# a_6110_4757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 a_33944_5411# a_33572_4991# a_32980_4757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2549 a_33894_n2704# a_33681_n2704# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2550 a_17931_n5092# a_17510_n5092# a_17832_n4915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2551 a_27413_1226# a_27200_1226# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2552 vdd d2 a_24838_1718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2553 a_16566_3789# a_16353_3789# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2554 a_27677_n8318# a_28482_n8552# a_28641_n8795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2555 a_8276_n8218# a_8490_n7302# a_8441_n7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2556 a_11084_1850# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2557 a_26489_n10440# a_29628_n10368# a_29579_n10352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2558 a_699_n8783# a_486_n8783# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2559 a_20996_141# a_31672_256# a_26832_263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2560 a_28230_7342# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2561 a_13774_8065# a_14832_8286# a_14787_8299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2562 a_23174_5403# a_22961_5403# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2563 vdd a_40798_8002# a_40590_8002# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2564 a_16080_4600# a_16078_4386# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2565 a_27604_4167# a_28408_3986# a_28577_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2566 a_22114_3773# a_21901_3773# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2567 gnd d0 a_9781_n4039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2568 a_11510_869# a_11089_869# a_10823_884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2569 a_27710_n2856# a_27289_n2856# a_27013_n2837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2570 vdd a_9749_n9916# a_9541_n9916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2571 a_1798_5551# a_1416_5993# a_824_5759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2572 vdd d0 a_4467_n9522# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2573 a_37844_4175# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2574 a_38151_n4824# a_37938_n4824# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2575 a_36402_n2439# a_36655_n2643# a_35386_n2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2576 a_32788_2236# a_32575_2236# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2577 a_9407_8270# a_10777_8324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2578 a_16861_n6810# a_16440_n6810# a_16164_n6791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2579 a_7176_n5084# a_6794_n5645# a_6202_n5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2580 gnd d1 a_24893_1157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2581 gnd d0 a_20338_5324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2582 a_11587_n4459# a_11166_n4459# a_10893_n4474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2583 a_30010_n2591# a_30263_n2795# a_29951_n3340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2584 vdd d3 a_24742_n8226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2585 a_3184_n3202# a_3279_n3826# a_3234_n3622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2586 a_22320_5164# a_21899_5164# a_21623_5064# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2587 a_24662_n5133# a_24915_n5337# a_24509_n4105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2588 a_24658_n5321# a_24762_n4776# a_24717_n4572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2589 a_11473_7727# a_11052_7727# a_10784_7557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2590 a_3130_5116# a_3383_5103# a_3071_5854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2591 a_10871_n8772# a_10871_n8490# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2592 gnd d1 a_30169_2117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2593 a_40562_5074# a_41620_5295# a_41571_5485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2594 a_25617_7458# a_25620_6866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2595 a_921_n5432# a_1726_n5666# a_1895_n5105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2596 a_28703_4418# a_28490_4418# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2597 vdd d7 a_32146_n10471# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2598 a_34152_n3124# a_34097_n4152# a_34281_n5900# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2599 a_33064_n7368# a_32643_n7368# a_32375_n6997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2600 a_5890_6717# a_5677_6717# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2601 a_8406_6076# a_8659_6063# a_8356_5656# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2602 a_27596_6124# a_27175_6124# a_26899_6024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2603 a_3164_n7119# a_3259_n7743# a_3210_n7727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2604 gnd a_20421_n7549# a_20213_n7549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2605 a_36290_5506# a_36547_5316# a_35281_5095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2606 a_16060_7922# a_16065_7536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2607 a_35214_7616# a_35309_8023# a_35260_8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2608 a_3222_n5582# a_3475_n5786# a_3172_n5162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2609 a_6200_n6802# a_5779_n6802# a_5503_n6501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2610 a_37938_n4824# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2611 a_39193_n8980# a_38980_n8980# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2612 a_12171_n6650# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2613 gnd d1 a_19422_n4792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2614 a_5684_5738# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2615 a_35292_2336# a_35549_2146# a_35246_1739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2616 a_34403_359# a_33982_359# a_34304_359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2617 a_33969_1613# a_33855_1494# a_34063_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2618 gnd a_10656_n10500# a_10448_n10500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2619 a_13775_7261# a_14836_6890# a_14787_7080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2620 a_2808_n10402# a_3065_n10418# a_2907_n10402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2621 a_17447_n7610# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2622 a_32649_n6802# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2623 a_2130_n5921# a_2021_n6098# a_2229_n6098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2624 a_17740_5538# a_17358_5980# a_16766_5746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2625 vdd a_24873_5074# a_24665_5074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2626 a_24416_2840# a_24673_2650# a_24321_4832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2627 a_812_7719# a_391_7719# a_118_7935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2628 vdd d4 a_35239_4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2629 a_40604_n5120# a_40699_n5744# a_40654_n5540# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2630 a_28425_1045# a_28212_1045# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2631 a_30986_n8475# a_31243_n8491# a_29974_n8656# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2632 a_8427_1355# a_9488_984# a_9439_1174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2633 a_32370_n8161# a_32368_n7764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2634 a_9513_n6771# a_9766_n6975# a_8500_n6537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2635 a_14896_n5824# a_14892_n6012# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2636 a_3095_1760# a_3190_2167# a_3141_2357# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2637 a_11298_2265# a_11085_2265# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2638 a_19072_5103# a_19325_5090# a_19013_5841# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2639 a_36304_2155# a_36561_1965# a_35292_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2640 a_20089_3557# a_20092_2965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2641 gnd a_30176_n9233# a_29968_n9233# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2642 a_8089_n10381# a_8250_n6309# a_8201_n6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2643 a_19164_n5569# a_20222_n6007# a_20177_n5803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2644 a_22334_1813# a_21913_1813# a_21640_2029# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2645 a_39413_n7020# a_39358_n8048# a_39566_n8048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2646 gnd a_5256_n10485# a_5048_n10485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2647 a_19106_n7106# a_19201_n7730# a_19156_n7526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2648 a_21712_n6775# a_22201_n6794# a_22409_n6794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2649 a_34053_n2947# a_33944_n3124# a_34152_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2650 a_28463_3425# a_28250_3425# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2651 a_33768_7932# a_33555_7932# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2652 vdd d0 a_41911_n7520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2653 a_9528_n2627# a_10462_n2231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2654 a_16350_4765# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2655 a_29993_n5532# a_31051_n5970# a_31002_n5954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2656 a_1644_2543# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2657 a_914_n7804# a_493_n7804# a_217_n7785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2658 a_23643_351# a_24370_4642# a_24325_4655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2659 gnd a_31150_8228# a_30942_8228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2660 a_39364_4426# a_39151_4426# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2661 a_38333_n9307# a_39138_n9541# a_39307_n8980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2662 a_20156_n9305# a_20152_n9493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2663 a_19144_n9486# a_20202_n9924# a_20153_n9908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2664 a_40655_n4747# a_40912_n4763# a_40600_n5308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2665 a_16875_n3459# a_16454_n3459# a_16181_n3474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2666 a_6187_n8347# a_5766_n8347# a_5500_n8161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2667 a_27263_n7339# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2668 a_14800_5535# a_15057_5345# a_13791_5124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2669 gnd a_20358_1407# a_20150_1407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2670 a_38257_6132# a_37836_6132# a_37560_6314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2671 a_37637_n9421# a_38126_n9722# a_38334_n9722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2672 gnd a_41899_n9480# a_41691_n9480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2673 a_20164_n7533# a_20421_n7549# a_19152_n7714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2674 vdd a_30043_n4288# a_29835_n4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2675 a_13802_2365# a_14059_2175# a_13756_1768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2676 a_22995_n7594# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2677 a_24414_n6097# a_24667_n6301# a_24298_n10373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2678 gnd a_40887_n9661# a_40679_n9661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2679 a_9444_1412# a_9440_1589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2680 a_637_2257# a_424_2257# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2681 a_408_4778# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2682 a_219_n8182# a_698_n8368# a_906_n8368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2683 vdd d0 a_4411_2401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2684 a_26921_2603# a_27400_2771# a_27608_2771# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2685 a_239_n3487# a_244_n3101# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2686 a_19106_n7106# a_19359_n7310# a_18937_n8226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2687 a_23624_n8061# a_23511_n6069# a_23719_n6069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 a_19037_1747# a_19132_2154# a_19083_2344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2689 vdd d4 a_13749_4679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2690 a_9491_n9485# a_9501_n8731# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2691 a_829_4778# a_1634_5012# a_1793_5432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2692 a_11147_n8791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2693 a_30925_2541# a_30928_1949# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2694 a_6214_n3451# a_5793_n3451# a_5525_n3080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_39086_1053# a_38873_1053# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2696 a_5898_6153# a_5685_6153# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2697 a_35146_n8218# a_35403_n8234# a_35075_n6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2698 a_27609_3186# a_27188_3186# a_26912_3368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2699 gnd a_32146_n10471# a_31938_n10471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2700 a_3223_n4789# a_4284_n4624# a_4239_n4420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2701 a_39334_n2926# a_38962_n2683# a_38371_n2864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2702 a_32882_n2885# a_32669_n2885# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2703 a_12278_7961# a_12065_7961# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2704 a_30913_4885# a_31166_4872# a_29897_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2705 a_20526_n805# d9 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2706 a_16583_848# a_16370_848# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2707 a_244_n3101# a_725_n3472# a_933_n3472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2708 vdd d0 a_20338_5324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2709 a_20194_n2862# a_20447_n3066# a_19181_n2628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2710 a_29912_2307# a_30973_1936# a_30928_1949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2711 vdd d1 a_14148_n3834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2712 a_6910_5972# a_6697_5972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2713 a_2831_4861# a_2975_2679# a_2930_2692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2714 a_22899_6943# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2715 a_22322_3773# a_23127_4007# a_23296_3565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2716 a_17472_n2712# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2717 vdd d0 a_25970_n7948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2718 a_38353_n5390# a_37932_n5390# a_37659_n5405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2719 a_17591_2063# a_17378_2063# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2720 gnd a_3371_7063# a_3163_7063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2721 a_21611_7306# a_22100_7124# a_22308_7124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2722 a_27470_n8733# a_27257_n8733# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2723 gnd d0 a_41842_1944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2724 a_41563_7268# a_41816_7255# a_40550_7034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2725 a_16564_5180# a_16351_5180# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2726 a_8402_6253# a_8659_6063# a_8356_5656# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2727 a_17931_n5092# a_17888_n4160# a_18072_n5908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2728 a_35354_n8685# a_36415_n8520# a_36366_n8504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2729 vdd d1 a_14064_1194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2730 a_16164_n6791# a_16653_n6810# a_16861_n6810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2731 a_29919_n9217# a_30023_n8672# a_29974_n8656# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2732 a_41683_n2418# a_41936_n2622# a_40667_n2787# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2733 a_34031_7371# a_33988_6439# a_34196_6439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2734 a_40634_n9457# a_41692_n9895# a_37639_n9917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2735 a_35214_7616# a_35309_8023# a_35264_8036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2736 a_40565_4098# a_40818_4085# a_40515_3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2737 vdd d0 a_20352_1973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2738 a_21645_1048# a_22131_832# a_22339_832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2739 vdd d0 a_20409_n9509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2740 gnd a_8684_1165# a_8476_1165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2741 a_18937_n8226# a_19151_n7310# a_19106_n7106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2742 a_9440_1589# a_9443_997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2743 a_32368_n7764# a_32857_n7783# a_33065_n7783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2744 a_11479_7161# a_12283_6980# a_12442_7400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2745 a_12132_5440# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2746 a_3230_n3810# a_4291_n3645# a_4242_n3629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2747 a_35289_3138# a_35542_3125# a_35230_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2748 a_9414_6072# a_9671_5882# a_8402_6253# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2749 a_21722_n5032# a_21720_n4818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2750 a_39476_338# a_39263_338# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2751 a_21628_3989# a_22114_3773# a_22322_3773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2752 a_4252_n2875# a_4505_n3079# a_3239_n2641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2753 a_5505_n6997# a_5986_n7368# a_6194_n7368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2754 a_35260_8213# a_36321_7842# a_36276_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2755 a_27584_8084# a_28388_7903# a_28557_7461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2756 a_34986_4663# a_35106_6575# a_35057_6765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2757 a_817_6738# a_1622_6972# a_1781_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2758 a_16435_n7791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2759 gnd a_36631_n7956# a_36423_n7956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 gnd d0 a_36636_n6975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2761 gnd a_4472_n8541# a_4264_n8541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2762 a_35170_n4113# a_35423_n4317# a_35071_n6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2763 a_14909_n3071# a_15166_n3087# a_13900_n2649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2764 vdd a_41831_4319# a_41623_4319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2765 a_3133_4140# a_3386_4127# a_3083_3720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2766 vdd d0 a_25957_n9493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2767 a_40565_4098# a_41623_4319# a_41574_4509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2768 vdd a_36549_3925# a_36341_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2769 a_24414_n6097# a_24534_n8226# a_24489_n8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2770 a_14806_3967# a_14802_4144# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2771 a_28752_n7012# a_28331_n7012# a_28658_n7012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2772 a_16447_n4438# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2773 a_37548_8274# a_38037_8092# a_38245_8092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 a_12459_5559# a_12077_6001# a_11486_6182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2775 a_8511_n3789# a_9572_n3624# a_9527_n3420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2776 a_13859_n9695# a_14920_n9530# a_14875_n9326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2777 a_17849_n3132# a_17735_n3132# a_17943_n3132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2778 a_30901_6845# a_30897_7022# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2779 a_40646_n7497# a_40899_n7701# a_40596_n7077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2780 a_20073_7297# a_20326_7284# a_19060_7063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2781 a_32272_7032# a_32761_7132# a_32969_7132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2782 a_1513_n5666# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2783 a_21882_8105# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2784 a_2229_n6098# a_1808_n6098# a_2130_n5921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2785 a_33952_3454# a_33580_3034# a_32989_3215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2786 a_33884_n4152# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2787 a_512_n3472# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2788 a_17832_n4915# a_17460_n4672# a_16869_n4853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2789 a_40507_5635# a_40602_6042# a_40553_6232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2790 a_13879_n5778# a_14136_n5794# a_13833_n5170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2791 a_28628_2493# a_28415_2493# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2792 a_19157_n6733# a_20218_n6568# a_20169_n6552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2793 vdd d0 a_4488_n6020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2794 vdd a_9753_n8520# a_9545_n8520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2795 a_20181_n4407# a_20434_n4611# a_19165_n4776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2796 a_27484_n5382# a_27271_n5382# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2797 a_27163_8084# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2798 a_37585_1134# a_38074_1234# a_38282_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2799 vdd d2 a_30107_3657# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2800 a_13799_3167# a_14052_3154# a_13740_3905# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2801 gnd d2 a_35499_1726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2802 a_33949_5530# a_33835_5411# a_34043_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2803 a_1806_3594# a_1424_4036# a_833_4217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2804 a_1808_n6098# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2805 a_19037_1747# a_19132_2154# a_19087_2167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2806 a_20153_n9908# a_20156_n9305# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2807 a_730_n2491# a_517_n2491# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2808 a_10777_8042# a_11266_8142# a_11474_8142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2809 a_19075_4127# a_19328_4114# a_19025_3707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2810 a_32375_n6402# a_32378_n6021# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2811 a_14907_n3449# a_14903_n3637# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2812 a_1719_4468# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2813 a_28815_330# a_28602_330# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2814 a_5429_2136# a_5918_2236# a_6126_2236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2815 a_16334_8121# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2816 a_13676_n4330# a_13890_n3414# a_13841_n3398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2817 a_5523_n2866# a_5523_n2584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2818 vdd a_15059_3954# a_14851_3954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2819 a_19075_4127# a_20133_4348# a_20084_4538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2820 a_21715_n5799# a_22204_n5818# a_22412_n5818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2821 a_27200_1226# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2822 vdd a_24838_1718# a_24630_1718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2823 a_16353_3789# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2824 a_1781_7392# a_1409_6972# a_817_6738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2825 a_24416_2840# a_24630_1718# a_24581_1908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2826 a_21988_n6794# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2827 a_40642_n7685# a_41703_n7520# a_41658_n7316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2828 a_32781_3215# a_32568_3215# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2829 a_1926_n8090# a_1713_n8090# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2830 a_39477_6418# a_39364_4426# a_39572_4426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2831 a_12399_n3714# a_12186_n3714# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2832 a_12462_3483# a_12090_3063# a_11499_3244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2833 a_40596_n7077# a_40691_n7701# a_40646_n7497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2834 a_4142_4935# a_4138_5112# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2835 vdd a_3371_7063# a_3163_7063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2836 a_32575_2236# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2837 a_41559_7445# a_41816_7255# a_40550_7034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2838 a_36281_6874# a_36277_7051# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2839 a_1706_n9583# a_1493_n9583# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2840 gnd a_24893_1157# a_24685_1157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2841 gnd d0 a_25869_8249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2842 gnd a_20338_5324# a_20130_5324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2843 a_38131_n8741# a_37918_n8741# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2844 a_37913_n9722# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2845 vdd a_31258_n5555# a_31050_n5555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2846 a_32844_n9328# a_32631_n9328# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2847 a_17748_3581# a_17366_4023# a_16775_4204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2848 gnd d0 a_15134_n8964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2849 a_8399_7055# a_8652_7042# a_8340_7793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2850 a_40561_4275# a_40818_4085# a_40515_3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2851 a_13782_6282# a_14039_6092# a_13736_5685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2852 a_11568_n8791# a_12372_n8610# a_12531_n8853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2853 gnd d2 a_14009_1755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2854 a_13802_2365# a_14863_1994# a_14818_2007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2855 vdd a_8684_1165# a_8476_1165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2856 a_28490_4418# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 vdd a_4383_6882# a_4175_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2858 a_1479_3475# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2859 a_5980_n8762# a_5767_n8762# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2860 gnd d1 a_30258_n3776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2861 a_16881_n2893# a_17685_n2712# a_17844_n2955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2862 a_35285_3315# a_35542_3125# a_35230_3876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2863 a_38282_1234# a_39086_1053# a_39245_1473# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2864 a_37560_6314# a_37560_6032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2865 a_32356_n9442# a_32358_n9343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2866 a_27588_6688# a_27167_6688# a_26901_6520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2867 a_11600_n2914# a_11179_n2914# a_10903_n2613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2868 a_27199_811# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2869 a_17440_n8589# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2870 a_26976_n9695# a_27465_n9714# a_27673_n9714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2871 a_28509_n3656# a_28296_n3656# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2872 a_14794_6101# a_15051_5911# a_13782_6282# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2873 vdd a_9659_7842# a_9451_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2874 a_34986_4663# a_35106_6575# a_35061_6588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2875 vdd d5 a_29836_n10368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2876 a_26976_n9695# a_26976_n9413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2877 a_13829_n5358# a_14086_n5374# a_13680_n4142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2878 a_19176_n3609# a_20234_n4047# a_20185_n4031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2879 a_31019_n3013# a_31022_n2410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2880 a_22339_832# a_23144_1066# a_23303_1486# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2881 a_5417_4378# a_5417_4096# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2882 a_2153_380# a_2044_380# a_2252_380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2883 a_11291_3244# a_11078_3244# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2884 vdd d2 a_35576_n5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2885 a_17987_6447# a_17874_4455# a_18082_4455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2886 a_36362_n9900# a_36619_n9916# a_35353_n9478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2887 a_23397_n3116# a_23015_n3677# a_22424_n3858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2888 a_6126_2236# a_6930_2055# a_7099_1613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2889 a_8488_n8497# a_8741_n8701# a_8429_n9246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2890 a_10794_5383# a_10794_5101# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2891 gnd a_14153_n2853# a_13945_n2853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2892 a_28212_1045# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2893 a_30924_2126# a_30934_1383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2894 a_27678_n8733# a_28482_n8552# a_28641_n8795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2895 vdd d1 a_3487_n3826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2896 a_16567_4204# a_16354_4204# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2897 a_11085_2265# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2898 a_20069_7474# a_20326_7284# a_19060_7063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2899 a_24704_n7510# a_25762_n7948# a_25717_n7744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2900 a_22949_7363# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2901 a_11510_869# a_12315_1103# a_12474_1523# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2902 a_40507_5635# a_40602_6042# a_40557_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2903 a_28250_3425# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2904 gnd d0 a_41917_n6954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2905 a_17675_n4160# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2906 a_27710_n2856# a_27289_n2856# a_27013_n2555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2907 a_33555_7932# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2908 a_20190_n3050# a_20447_n3066# a_19181_n2628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2909 a_3091_1937# a_3348_1747# a_2926_2869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2910 a_38250_7111# a_37829_7111# a_37553_7293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2911 a_2930_2692# a_3183_2679# a_2831_4861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2912 vdd d0 a_31238_n9472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2913 a_29834_7587# a_29929_7994# a_29880_8184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2914 vdd d0 a_20332_5890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2915 a_39151_4426# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2916 a_13795_3344# a_14052_3154# a_13740_3905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2917 a_630_3236# a_417_3236# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2918 vdd a_19434_n2832# a_19226_n2832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2919 vdd d2 a_35499_1726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2920 a_36289_6310# a_36542_6297# a_35276_6076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2921 gnd d0 a_15148_n5613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2922 a_20189_n2635# a_21123_n2239# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2923 vdd d0 a_9749_n9916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2924 a_922_n5847# a_1726_n5666# a_1895_n5105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2925 a_7434_359# a_7325_359# a_5243_292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2926 a_5773_n7368# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2927 a_1831_380# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_3150_1199# a_3403_1186# a_3091_1937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 a_6094_8113# a_5673_8113# a_5397_8295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2930 a_4247_n2648# a_4504_n2664# a_3235_n2829# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2931 a_19071_4304# a_19328_4114# a_19025_3707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2932 a_424_2257# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2933 a_4126_8291# a_5397_8295# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2934 a_17748_3581# a_17634_3462# a_17842_3462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2935 a_26906_4944# a_27392_4728# a_27600_4728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2936 a_5891_7132# a_5678_7132# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2937 vdd a_15133_n8549# a_14925_n8549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2938 gnd d0 a_36639_n5999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2939 a_38261_4736# a_39066_4970# a_39225_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2940 a_3235_n2829# a_3492_n2845# a_3180_n3390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2941 vdd d0 a_4403_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2942 a_35370_n6537# a_36428_n6975# a_36379_n6959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2943 a_40566_3294# a_41627_2923# a_41578_3113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2944 a_29993_n5532# a_30246_n5736# a_29943_n5112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2945 a_31672_256# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2946 a_24688_n9658# a_25749_n9493# a_25704_n9289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2947 a_15660_n10477# a_18799_n10405# a_18171_n6085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2948 a_5685_6153# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2949 a_32649_n6802# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2950 vdd a_4410_1986# a_4202_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2951 gnd d1 a_14133_n6770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2952 a_18872_2679# a_19125_2666# a_18773_4848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2953 a_34120_n9001# a_33699_n9001# a_34021_n8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2954 a_813_8134# a_392_8134# a_116_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2955 a_12065_7961# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2956 a_22408_n6379# a_21987_n6379# a_21714_n6394# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2957 a_23020_n2696# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2958 vdd a_20338_5324# a_20130_5324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2959 vdd d0 a_25905_976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2960 a_37840_4736# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2961 vdd a_8718_n3385# a_8510_n3385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2962 a_28608_6410# a_28395_6410# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2963 a_24620_5087# a_24873_5074# a_24561_5825# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2964 a_9427_4353# a_9423_4530# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2965 gnd a_29836_n10368# a_29628_n10368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2966 a_38056_3760# a_37843_3760# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2967 a_11387_n3895# a_11174_n3895# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2968 a_8395_7232# a_8652_7042# a_8340_7793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2969 a_9512_n5983# a_9769_n5999# a_8503_n5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2970 vdd d2 a_14009_1755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2971 vdd a_41847_963# a_41639_963# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2972 vdd d0 a_31155_7247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2973 a_38923_1473# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2974 gnd a_4485_n6996# a_4277_n6996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2975 vdd d0 a_20435_n5026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2976 a_24693_n8677# a_24950_n8693# a_24638_n9238# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2977 gnd a_41842_1944# a_41634_1944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2978 a_36390_n4399# a_36386_n4587# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2979 a_16351_5180# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2980 a_914_n7804# a_493_n7804# a_217_n7503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2981 gnd d0 a_20325_6869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2982 vdd d1 a_30157_4077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2983 vdd d2 a_3437_n3406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2984 a_37332_n2231# a_38162_n2449# a_38370_n2449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2985 a_26993_n6472# a_26995_n6373# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2986 vdd a_14064_1194# a_13856_1194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2987 a_38334_n9722# a_39138_n9541# a_39307_n8980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2988 a_23298_n6069# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2989 gnd d1 a_35549_2146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2990 a_5905_3781# a_5692_3781# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2991 gnd d0 a_31264_n4989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2992 a_5523_n2584# a_6012_n2885# a_6220_n2885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2993 a_29896_6047# a_30954_6268# a_30905_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2994 gnd d0 a_41828_5295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2995 a_10871_n8490# a_11360_n8791# a_11568_n8791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2996 vdd a_41916_n6539# a_41708_n6539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2997 a_37637_n9703# a_38126_n9722# a_38334_n9722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2998 vdd a_20352_1973# a_20144_1973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2999 a_37570_4571# a_38053_4736# a_38261_4736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3000 a_19076_3323# a_20137_2952# a_20088_3142# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 gnd d0 a_20415_n8943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3002 a_33731_n3124# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3003 a_32792_840# a_32579_840# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3004 a_26995_n6373# a_27481_n6358# a_27689_n6358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3005 a_38281_819# a_37860_819# a_37587_1035# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3006 vdd a_9760_n7541# a_9552_n7541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3007 vdd a_25886_5308# a_25678_5308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3008 vdd d0 a_4492_n4624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3009 a_21991_n5818# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3010 gnd d2 a_3417_n7323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3011 vdd d2 a_40857_n5324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3012 a_10905_n3109# a_11386_n3480# a_11594_n3480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3013 a_13791_5124# a_14849_5345# a_14800_5535# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3014 a_906_n8368# a_1711_n8602# a_1870_n8845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3015 vdd a_24888_2138# a_24680_2138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3016 a_11360_n8791# a_11147_n8791# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3017 a_36362_n9900# a_36365_n9297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3018 gnd d1 a_35611_n8701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3019 gnd a_35606_n9682# a_35398_n9682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3020 a_24585_1731# a_24680_2138# a_24631_2328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3021 a_29985_n7489# a_31043_n7927# a_30998_n7723# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3022 gnd d0 a_25873_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3023 gnd d0 a_20333_6305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3024 a_27179_4728# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3025 gnd d6 a_37407_n10464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3026 a_16077_5576# a_16558_5746# a_16766_5746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3027 a_24717_n4572# a_25775_n5010# a_25726_n4994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3028 a_29994_n4739# a_31055_n4574# a_31010_n4370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3029 a_23196_n9554# a_22983_n9554# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3030 a_13868_n8526# a_14926_n8964# a_14877_n8948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3031 a_20153_n9908# a_20410_n9924# a_19144_n9486# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3032 gnd a_25880_5874# a_25672_5874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3033 a_13868_n8526# a_14121_n8730# a_13809_n9275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3034 a_239_n3487# a_725_n3472# a_933_n3472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3035 a_19094_n9066# a_19189_n9690# a_19144_n9486# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3036 a_9423_4530# a_9426_3938# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3037 a_5698_3215# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3038 a_38276_1800# a_37855_1800# a_37582_2016# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3039 gnd d1 a_14059_2175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3040 a_1781_n5105# a_1568_n5105# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3041 a_23422_4439# a_23209_4439# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3042 a_17472_n2712# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3043 a_629_2821# a_416_2821# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3044 a_28415_2493# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3045 gnd d0 a_4499_n3645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3046 a_22315_6145# a_21894_6145# a_21618_6327# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3047 a_27470_n8733# a_27257_n8733# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3048 a_25721_n6348# a_25974_n6552# a_24705_n6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3049 a_3146_1376# a_3403_1186# a_3091_1937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3050 a_39327_n5063# a_38945_n5624# a_38354_n5805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3051 gnd a_36530_8257# a_36322_8257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3052 a_40630_n9645# a_41691_n9480# a_41642_n9464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3053 a_41553_8011# a_41810_7821# a_40541_8192# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3054 a_32865_n5826# a_32652_n5826# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3055 vdd a_30107_3657# a_29899_3657# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3056 a_33064_n7368# a_32643_n7368# a_32370_n7383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3057 a_12573_1523# a_12518_2551# a_12702_4476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3058 a_33924_n7041# a_33711_n7041# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3059 a_19145_n8693# a_19402_n8709# a_19090_n9254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3060 a_27709_n2441# a_27288_n2441# a_27015_n2456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3061 a_23058_n5076# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3062 a_3168_n5350# a_3425_n5366# a_3019_n4134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3063 a_23471_n7033# a_23416_n8061# a_23624_n8061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3064 a_32281_5954# a_32767_5738# a_32975_5738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3065 gnd d0 a_15166_n3087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3066 a_5987_n7783# a_5774_n7783# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3067 a_23144_1066# a_22931_1066# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3068 a_39124_3433# a_38911_3433# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3069 a_17447_n7610# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3070 a_18868_2856# a_19125_2666# a_18773_4848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3071 a_32304_1437# a_32304_1155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3072 a_39000_n5063# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3073 vdd d0 a_25906_1391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3074 a_18777_4671# a_18897_6583# a_18848_6773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3075 a_6194_n7368# a_6999_n7602# a_7168_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3076 gnd d0 a_41920_n5978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3077 a_38350_n6366# a_39155_n6600# a_39314_n6843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3078 a_11374_n5440# a_11161_n5440# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3079 a_4252_n2875# a_4248_n3063# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3080 a_40651_n6516# a_41709_n6954# a_41660_n6938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3081 a_4139_5527# a_4396_5337# a_3130_5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3082 a_34380_n6077# a_35216_n10397# a_35058_n10381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3083 a_24616_5264# a_24873_5074# a_24561_5825# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3084 a_23182_3446# a_22969_3446# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3085 gnd a_40912_n4763# a_40704_n4763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3086 a_8495_n7518# a_8748_n7722# a_8445_n7098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3087 a_3141_2357# a_3398_2167# a_3095_1760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3088 a_36293_4914# a_36546_4901# a_35277_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3089 a_36366_n8504# a_36623_n8520# a_35354_n8685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3090 a_40577_2138# a_41635_2359# a_41590_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3091 gnd a_8756_n5765# a_8548_n5765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3092 gnd d1 a_8761_n4784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3093 gnd a_40520_4629# a_40312_4629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3094 a_5513_n4445# a_5999_n4430# a_6207_n4430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3095 gnd a_15040_8286# a_14832_8286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3096 a_28569_5501# a_28455_5382# a_28663_5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3097 gnd a_35556_n9262# a_35348_n9262# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3098 a_5506_n5525# a_5508_n5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3099 a_20063_8040# a_20320_7850# a_19051_8221# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3100 a_17665_n6629# a_17452_n6629# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3101 a_1513_n5666# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3102 vdd d1 a_35549_2146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3103 vdd d5 a_3065_n10418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3104 a_41678_n3399# a_41674_n3587# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3105 a_17832_n4915# a_17460_n4672# a_16868_n4438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3106 a_32773_5172# a_32560_5172# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3107 a_28405_4962# a_28192_4962# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3108 a_27263_n7339# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3109 a_28717_n4123# a_28504_n4123# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3110 a_35373_n5561# a_36431_n5999# a_36382_n5983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3111 a_36314_1412# a_36310_1589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3112 a_609_6738# a_396_6738# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3113 gnd d1 a_8664_5082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3114 a_4227_n7773# a_4223_n7961# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3115 a_27407_1792# a_27194_1792# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3116 a_27604_4167# a_27183_4167# a_26907_4349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3117 a_13791_5124# a_14849_5345# a_14804_5358# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3118 a_36398_n2627# a_37332_n2231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3119 a_6188_n8762# a_5767_n8762# a_5491_n8743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3120 a_6110_4757# a_5689_4757# a_5416_4973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3121 a_1731_n4685# a_1518_n4685# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3122 vdd a_35423_n4317# a_35215_n4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3123 a_13821_n7315# a_13925_n6770# a_13876_n6754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3124 a_31013_n3579# a_31023_n2825# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3125 a_36277_8270# a_37548_8274# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3126 a_5397_8013# a_5399_7914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3127 a_27276_n4401# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3128 a_25737_n3827# a_25990_n4031# a_24724_n3593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3129 a_35292_2336# a_36353_1965# a_36304_2155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3130 a_36377_n7337# a_36630_n7541# a_35361_n7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3131 a_2920_n6314# a_3177_n6330# a_2808_n10402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3132 a_11562_n9357# a_11141_n9357# a_10868_n9372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3133 a_4227_n7773# a_4480_n7977# a_3214_n7539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3134 a_4219_n8337# a_4215_n8525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3135 a_14901_n4843# a_15154_n5047# a_13888_n4609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3136 a_39104_7350# a_38891_7350# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3137 gnd a_35403_n8234# a_35195_n8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3138 vdd a_15146_n7004# a_14938_n7004# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3139 a_37637_n9703# a_37637_n9421# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3140 a_32301_2632# a_32780_2800# a_32988_2800# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3141 a_16354_4204# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3142 a_4239_n4420# a_4492_n4624# a_3223_n4789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3143 a_21919_1247# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3144 a_849_861# a_428_861# a_162_876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3145 a_30917_4324# a_31170_4311# a_29904_4090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3146 gnd d1 a_40892_n8680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3147 a_17837_n5092# a_17723_n5092# a_17931_n5092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3148 a_23402_1486# a_22981_1486# a_23308_1605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3149 a_28653_n6835# a_28281_n6592# a_27690_n6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3150 vdd d1 a_14059_2175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3151 a_428_861# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3152 a_38048_5717# a_37835_5717# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3153 a_9428_3549# a_9685_3359# a_8419_3138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3154 a_16092_2640# a_16090_2426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3155 a_29897_5243# a_30958_4872# a_30909_5062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3156 a_26919_2107# a_26921_2008# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3157 vdd d2 a_24927_n3377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3158 a_5799_n2885# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3159 a_38131_n8741# a_37918_n8741# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3160 a_37913_n9722# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3161 vdd a_20332_5890# a_20124_5890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3162 a_8496_n6725# a_9557_n6560# a_9512_n6356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3163 a_7322_4447# a_6925_2522# a_7181_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3164 a_16559_6161# a_16346_6161# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3165 a_34021_n8824# a_33649_n8581# a_33058_n8762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3166 a_16164_n6509# a_16653_n6810# a_16861_n6810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3167 a_16460_n2893# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3168 a_10804_3640# a_11285_3810# a_11493_3810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3169 a_40451_n4092# a_40649_n5324# a_40604_n5120# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3170 a_11391_n2499# a_11178_n2499# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3171 a_36310_1589# a_36313_997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3172 a_10891_n4855# a_10891_n4573# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3173 a_9516_n4587# a_9773_n4603# a_8504_n4768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3174 a_20100_1182# a_20357_992# a_19088_1363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3175 a_27672_n9299# a_27251_n9299# a_26978_n9314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3176 vdd d0 a_25982_n4595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3177 a_1498_n8602# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3178 a_5424_3016# a_5910_2800# a_6118_2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3179 a_497_n6408# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3180 a_35299_n9246# a_35403_n8701# a_35354_n8685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3181 a_26919_2107# a_27408_2207# a_27616_2207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3182 a_40671_n2599# a_40924_n2803# a_40612_n3348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3183 vdd a_4403_2965# a_4195_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3184 a_31994_256# a_37072_271# a_37394_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3185 a_138_4613# a_136_4399# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3186 a_18777_4671# a_18897_6583# a_18852_6596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3187 a_37072_271# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3188 a_123_7549# a_121_7335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3189 a_2130_n5921# a_1733_n4173# a_2001_n3145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3190 a_32543_8113# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3191 a_2906_6786# a_3163_6596# a_2835_4684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3192 a_21702_n8949# a_21700_n8735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3193 a_23397_n3116# a_23015_n3677# a_22423_n3443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3194 a_39324_5390# a_38903_5390# a_39230_5509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3195 a_24420_2663# a_24618_3678# a_24573_3691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3196 a_20169_n7760# a_20165_n7948# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3197 a_12706_6468# a_12593_4476# a_12801_4476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3198 a_17799_2530# a_17586_2530# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3199 gnd d1 a_35618_n7722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3200 a_486_n8783# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3201 gnd d2 a_24838_1718# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3202 gnd d0 a_4384_7297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3203 a_4157_1999# a_4153_2176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3204 vdd a_15040_8286# a_14832_8286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3205 a_28395_6410# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3206 a_16779_2808# a_16358_2808# a_16092_2640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3207 a_9527_n3420# a_9780_n3624# a_8511_n3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3208 a_41668_n4981# a_41671_n4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3209 vdd a_31155_7247# a_30947_7247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3210 a_5414_5354# a_5414_5072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3211 a_34033_n6864# a_33924_n7041# a_34132_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3212 gnd a_25989_n3616# a_25781_n3616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3213 a_22327_2792# a_21906_2792# a_21640_2624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3214 a_9422_4115# a_9432_3372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3215 a_22969_3446# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3216 vdd d1 a_8664_5082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3217 a_32969_7132# a_32548_7132# a_32272_7314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3218 a_15904_300# a_17773_367# a_18082_4455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3219 gnd a_20325_6869# a_20117_6869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3220 a_41647_n8483# a_41904_n8499# a_40635_n8664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3221 vdd a_30157_4077# a_29949_4077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3222 a_1875_n9022# a_1761_n9022# a_1969_n9022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3223 a_1704_1515# a_1491_1515# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3224 gnd d1 a_40823_3104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3225 a_5692_3781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3226 a_12706_6468# a_12285_6468# a_12553_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3227 a_8402_6253# a_9463_5882# a_9414_6072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3228 a_40635_n8664# a_40892_n8680# a_40580_n9225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3229 a_13900_n2649# a_14958_n3087# a_14909_n3071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3230 a_14787_7080# a_14799_6339# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3231 gnd a_41828_5295# a_41620_5295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3232 vdd d0 a_15165_n2672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3233 a_35077_2848# a_35291_1726# a_35242_1916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3234 gnd d3 a_3272_n4338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3235 a_23124_4983# a_22911_4983# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3236 a_28816_6410# a_28703_4418# a_28911_4418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3237 a_906_n8368# a_485_n8368# a_219_n8182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3238 a_13740_3905# a_13844_3154# a_13795_3344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3239 a_5411_6549# a_5890_6717# a_6098_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3240 a_6786_n7602# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3241 a_40654_n5540# a_41712_n5978# a_41663_n5962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3242 a_27693_n5797# a_27272_n5797# a_26996_n5496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3243 a_4230_n5589# a_4240_n4835# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3244 a_27616_2207# a_28420_2026# a_28589_1584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3245 gnd a_9691_1965# a_9483_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3246 a_30904_6043# a_30914_5300# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3247 a_12467_3602# a_12353_3483# a_12561_3483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3248 a_7171_n4907# a_6799_n4664# a_6208_n4845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3249 a_26832_263# a_26411_263# a_23742_351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3250 a_36296_3938# a_36549_3925# a_35280_4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3251 a_37587_1035# a_37594_834# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3252 a_20674_141# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3253 vdd a_19417_n5773# a_19209_n5773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3254 a_26411_263# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3255 a_20084_4538# a_20087_3946# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3256 a_21715_n5517# a_22204_n5818# a_22412_n5818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3257 a_12422_n9030# a_12209_n9030# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3258 gnd a_25873_6853# a_25665_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3259 a_2835_4684# a_3088_4671# a_2153_380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3260 a_30913_4501# a_31170_4311# a_29904_4090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3261 vdd a_26746_n10456# a_26538_n10456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3262 vdd a_40704_n4296# a_40496_n4296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3263 gnd a_20333_6305# a_20125_6305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3264 a_8449_n5329# a_8553_n4784# a_8504_n4768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3265 a_14887_n7366# a_14883_n7554# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3266 a_5991_n6387# a_5778_n6387# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3267 a_5786_n4430# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3268 vdd d3 a_8553_n4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3269 a_32776_4196# a_32563_4196# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3270 a_24581_1908# a_24838_1718# a_24416_2840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3271 a_39225_n3103# a_39012_n3103# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3272 a_41658_n7316# a_41911_n7520# a_40642_n7685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3273 vdd a_31276_n3029# a_31068_n3029# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3274 a_14808_3578# a_15065_3388# a_13799_3167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3275 a_123_6954# a_609_6738# a_817_6738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3276 a_11479_7161# a_11058_7161# a_10782_7343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3277 a_38249_6696# a_37828_6696# a_37562_6528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3278 vdd a_20427_n6983# a_20219_n6983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3279 a_4227_n6565# a_4235_n5816# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3280 a_705_n7389# a_492_n7389# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3281 a_22416_n4422# a_23221_n4656# a_23380_n4899# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3282 gnd d3 a_8533_n8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3283 a_38057_4175# a_37844_4175# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3284 gnd d1 a_24965_n5757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3285 a_4163_1433# a_4416_1420# a_3150_1199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3286 a_416_2821# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3287 a_21631_3389# a_21631_3107# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3288 a_39061_5951# a_38848_5951# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3289 a_29981_n7677# a_30238_n7693# a_29935_n7069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3290 a_11567_n8376# a_12372_n8610# a_12531_n8853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3291 gnd a_31256_n6946# a_31048_n6946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3292 a_27584_8084# a_27163_8084# a_26887_8266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3293 a_35277_5272# a_36338_4901# a_36293_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3294 a_33000_840# a_33805_1074# a_33964_1494# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3295 vdd a_36638_n5584# a_36430_n5584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3296 vdd d0 a_36643_n4603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3297 a_16792_1263# a_16371_1263# a_16095_1445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3298 vdd a_4488_n6020# a_4280_n6020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3299 vdd d2 a_30208_n3356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3300 a_11179_n2914# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3301 a_9419_5091# a_9427_4353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3302 a_12553_5440# a_12132_5440# a_12454_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3303 a_41577_3917# a_41573_4094# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3304 a_17849_n3132# a_17467_n3693# a_16875_n3459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3305 a_2001_n3145# a_1580_n3145# a_1907_n3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3306 vdd d2 a_8706_n5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3307 a_38276_1800# a_39081_2034# a_39250_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3308 vdd d0 a_41822_5861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3309 a_14806_3967# a_15059_3954# a_13790_4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3310 a_718_n4451# a_505_n4451# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3311 a_14889_n6988# a_14892_n6385# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3312 a_30998_n7723# a_30994_n7911# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3313 a_16422_n9336# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3314 a_150_2058# a_155_1672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3315 a_28413_3005# a_28200_3005# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3316 a_11594_n3480# a_12399_n3714# a_12568_n3153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3317 a_36284_6072# a_36294_5329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3318 a_907_n8783# a_1711_n8602# a_1870_n8845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3319 a_13782_6282# a_14843_5911# a_14798_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3320 vdd d1 a_30251_n4755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3321 vdd d1 a_19397_n9690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3322 vdd a_25906_1391# a_25698_1391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3323 a_11286_4225# a_11073_4225# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3324 vdd a_35623_n6741# a_35415_n6741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3325 a_29921_1149# a_30174_1136# a_29862_1887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3326 a_11057_6746# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3327 vdd d1 a_14039_6092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3328 a_26914_3582# a_26912_3368# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3329 gnd d4 a_13749_4679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3330 vdd d0 a_9760_n7541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3331 a_38262_5151# a_39066_4970# a_39225_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3332 a_28207_2026# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3333 a_24505_n4293# a_24719_n3377# a_24674_n3173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3334 vdd d0 a_31174_2915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3335 a_1900_3475# a_1479_3475# a_1801_3475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3336 a_30990_n8287# a_30986_n8475# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3337 a_11599_n2499# a_11178_n2499# a_10462_n2231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3338 a_27289_n2856# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3339 a_33788_4015# a_33575_4015# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3340 vdd a_41905_n8914# a_41697_n8914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3341 a_16070_6343# a_16559_6161# a_16767_6161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3342 gnd d0 a_36650_n3624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3343 a_153_1176# a_155_1077# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3344 gnd d0 a_25893_2936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3345 a_21613_7520# a_21611_7306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3346 a_23196_n9554# a_22983_n9554# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3347 a_16167_n5533# a_16656_n5834# a_16864_n5834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3348 a_17829_n7049# a_17715_n7049# a_17923_n7049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3349 a_21712_n6775# a_21712_n6493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3350 a_14818_2007# a_14814_2184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3351 a_4130_6895# a_4383_6882# a_3114_7253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3352 a_10794_5101# a_11283_5201# a_11491_5201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3353 vdd a_31181_1936# a_30973_1936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3354 vdd a_19367_n5353# a_19159_n5353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3355 a_21913_1813# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3356 a_6106_6153# a_6910_5972# a_7079_5530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3357 vdd d0 a_9685_3359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3358 gnd a_40497_n10376# a_40289_n10376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3359 a_27400_2771# a_27187_2771# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3360 a_14871_n9514# a_15128_n9530# a_13859_n9695# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3361 a_10498_n10484# a_10448_n10500# a_5098_n10469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3362 gnd a_25900_1957# a_25692_1957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3363 a_12140_3483# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3364 a_38277_2215# a_37856_2215# a_37580_2115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3365 a_7118_6439# a_6905_6439# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3366 vdd a_20441_n3632# a_20233_n3632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3367 a_32560_5172# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3368 a_28192_4962# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3369 a_2831_4861# a_2975_2679# a_2926_2869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3370 a_37860_819# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3371 a_27704_n3422# a_28509_n3656# a_28678_n3095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3372 a_35077_2848# a_35291_1726# a_35246_1739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3373 a_40561_4275# a_41622_3904# a_41573_4094# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3374 a_726_n3887# a_513_n3887# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3375 a_9406_7855# a_9659_7842# a_8390_8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3376 a_396_6738# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3377 a_39302_n8803# a_39193_n8980# a_39401_n8980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3378 gnd a_30087_7574# a_29879_7574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3379 a_21628_4584# a_22111_4749# a_22319_4749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3380 a_39327_n5063# a_38945_n5624# a_38353_n5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3381 a_16868_n4438# a_17673_n4672# a_17832_n4915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3382 a_13740_3905# a_13844_3154# a_13799_3167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3383 gnd a_31270_n3595# a_31062_n3595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3384 a_17755_1502# a_17383_1082# a_16791_848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3385 a_27194_1792# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3386 a_32865_n5826# a_32652_n5826# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3387 vdd a_41932_n4018# a_41724_n4018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3388 a_11588_n4874# a_11167_n4874# a_10891_n4855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3389 a_25720_n5560# a_25977_n5576# a_24708_n5741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3390 a_34038_n7041# a_33656_n7602# a_33065_n7783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3391 a_27709_n2441# a_27288_n2441# a_26671_n2223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3392 vdd a_3460_n8722# a_3252_n8722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3393 a_5098_n10469# a_5048_n10485# a_2907_n10402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3394 gnd d0 a_25901_2372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3395 a_5886_8113# a_5673_8113# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3396 a_3134_3336# a_4195_2965# a_4150_2978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3397 a_20169_n6552# a_20177_n5803# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3398 a_33072_n5411# a_33877_n5645# a_34046_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3399 a_24608_7047# a_25666_7268# a_25621_7281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3400 vdd d0 a_20446_n2651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3401 a_2831_4861# a_3088_4671# a_2153_380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3402 a_29931_n7257# a_30188_n7273# a_29766_n8189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3403 gnd a_41912_n7935# a_41704_n7935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3404 a_32395_n2485# a_31952_n2202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3405 gnd d6 a_26746_n10456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3406 a_11153_n7397# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3407 a_21123_n2239# a_22220_n2462# a_22428_n2462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3408 a_35373_n5561# a_35626_n5765# a_35323_n5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3409 a_12607_n4181# a_12394_n4181# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3410 a_121_7053# a_123_6954# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3411 a_3129_4317# a_4190_3946# a_4141_4136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3412 a_7434_359# a_8161_4650# a_8112_4840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3413 a_12298_4044# a_12085_4044# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3414 a_38351_n6781# a_37930_n6781# a_37654_n6480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3415 a_38041_6696# a_37828_6696# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3416 a_6195_n7783# a_6999_n7602# a_7168_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3417 a_33077_n4430# a_32656_n4430# a_32390_n4244# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3418 a_10888_n6050# a_11371_n6416# a_11579_n6416# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3419 a_23327_6431# a_23114_6431# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3420 vdd d1 a_8667_4106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3421 a_13845_n3210# a_14098_n3414# a_13676_n4330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3422 a_29697_2819# a_29911_1697# a_29866_1710# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3423 a_33711_n7041# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3424 a_34281_n5900# a_34172_n6077# a_34380_n6077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3425 vdd a_3487_n3826# a_3279_n3826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3426 a_18773_4848# a_18917_2666# a_18868_2856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3427 a_36378_n7752# a_36374_n7940# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3428 vout a_20526_n805# a_20848_n805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3429 a_37835_5717# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3430 gnd a_41831_4319# a_41623_4319# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3431 a_4159_1610# a_4416_1420# a_3150_1199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3432 gnd d1 a_40803_7021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3433 a_7510_n6077# a_7089_n6077# a_7411_n5900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3434 vdd d2 a_19347_n9270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3435 vdd d3 a_13933_n4346# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3436 a_30987_n8890# a_31244_n8906# a_29978_n8468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3437 a_13896_n2837# a_14957_n2672# a_14912_n2468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3438 a_16092_2045# a_16097_1659# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3439 a_39218_7469# a_38836_7911# a_38245_8092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3440 a_5422_3115# a_5424_3016# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3441 gnd a_3467_n7743# a_3259_n7743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3442 a_224_n6423# a_710_n6408# a_918_n6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3443 gnd a_40810_6042# a_40602_6042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3444 a_16083_3123# a_16572_3223# a_16780_3223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3445 a_24725_n2800# a_25786_n2635# a_25737_n2619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3446 a_31013_n3579# a_31270_n3595# a_30001_n3760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3447 a_41589_1957# a_41842_1944# a_40573_2315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3448 a_34031_7371# a_33610_7371# a_33937_7490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3449 a_36370_n8316# a_36366_n8504# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3450 a_26998_n5992# a_27481_n6358# a_27689_n6358# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3451 a_12543_n6893# a_12171_n6650# a_11579_n6416# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3452 a_41652_n8710# a_41648_n8898# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3453 a_7207_n8069# a_6994_n8069# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3454 vdd a_3405_n9283# a_3197_n9283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3455 a_19110_n5337# a_19214_n4792# a_19169_n4588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3456 a_21991_n5818# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3457 vdd d0 a_41924_n4582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3458 a_32376_n5525# a_32378_n5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3459 gnd d2 a_30107_3657# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3460 a_37150_n10448# a_40289_n10376# a_40240_n10360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3461 gnd d1 a_8684_1165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3462 a_23620_n5892# a_23223_n4144# a_23479_n5076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3463 a_16876_n3874# a_16455_n3874# a_16179_n3855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3464 a_6188_n8762# a_5767_n8762# a_5491_n8461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3465 vdd a_40904_n6720# a_40696_n6720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3466 a_22195_n7360# a_21982_n7360# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3467 a_29917_1326# a_30174_1136# a_29862_1887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3468 a_32755_7698# a_32542_7698# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3469 a_1761_n9022# a_1548_n9022# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3470 a_7325_359# a_7112_359# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3471 a_25629_5498# a_25886_5308# a_24620_5087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3472 a_6111_5172# a_5690_5172# a_5414_5072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3473 vdd a_8748_n7722# a_8540_n7722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3474 a_27276_n4401# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3475 vdd d2 a_30176_n9233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3476 a_32370_n8161# a_32849_n8347# a_33057_n8347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3477 gnd d0 a_9773_n4603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3478 a_24631_2328# a_24888_2138# a_24585_1731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3479 a_11562_n9357# a_11141_n9357# a_10873_n8986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3480 gnd a_15145_n6589# a_14937_n6589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3481 a_210_n8482# a_699_n8783# a_907_n8783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3482 a_20099_1986# a_20095_2163# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3483 a_5429_2418# a_5429_2136# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3484 vdd d3 a_19194_n8242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3485 a_16345_5746# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3486 a_30998_n7723# a_31251_n7927# a_29985_n7489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3487 a_41663_n6335# a_41659_n6523# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3488 a_30892_8003# a_31149_7813# a_29880_8184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3489 a_41575_5308# a_41571_5485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3490 a_36293_4530# a_36296_3938# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3491 a_23008_n4656# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3492 a_17586_2530# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3493 a_24662_n5133# a_24757_n5757# a_24708_n5741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3494 gnd a_24838_1718# a_24630_1718# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3495 a_38365_n3430# a_37944_n3430# a_37676_n3059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3496 a_32292_3397# a_32781_3215# a_32989_3215# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3497 a_40362_2650# a_40560_3665# a_40511_3855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3498 a_5416_4973# a_5419_4592# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3499 a_32980_4757# a_33785_4991# a_33944_5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3500 a_35374_n4768# a_36435_n4603# a_36390_n4399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3501 a_5498_n7482# a_5500_n7383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3502 a_38049_6132# a_37836_6132# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3503 a_20099_1986# a_20352_1973# a_19083_2344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3504 a_35323_n5141# a_35576_n5345# a_35170_n4113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3505 a_32395_n3080# a_32876_n3451# a_33084_n3451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3506 a_7054_n7041# a_6841_n7041# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3507 vdd a_25978_n5991# a_25770_n5991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3508 vdd a_30087_7574# a_29879_7574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3509 a_30998_n6515# a_31006_n5766# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3510 a_8207_2848# a_8464_2658# a_8112_4840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3511 a_2930_2692# a_3128_3707# a_3079_3897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3512 a_28905_n8040# a_28484_n8040# a_28740_n8972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3513 a_1491_1515# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3514 a_23491_n3116# a_23070_n3116# a_23397_n3116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3515 gnd a_40823_3104# a_40615_3104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3516 vdd a_15129_n9945# a_14921_n9945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3517 gnd a_9684_2944# a_9476_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3518 a_27600_4728# a_27179_4728# a_26906_4944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3519 a_25706_n8911# a_25709_n8308# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3520 a_3207_n8518# a_4265_n8956# a_4216_n8940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3521 vdd a_15071_1994# a_14863_1994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3522 gnd d2 a_35467_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3523 a_10797_4407# a_11286_4225# a_11494_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3524 vdd d3 a_30023_n8205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3525 a_20152_n9493# a_20409_n9509# a_19140_n9674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3526 vdd d0 a_25901_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3527 a_12404_n2733# a_12191_n2733# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3528 a_1498_n8602# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3529 a_28646_n8972# a_28264_n9533# a_27673_n9714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3530 a_6125_1821# a_5704_1821# a_5431_2037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3531 a_1793_5432# a_1421_5012# a_829_4778# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3532 a_4227_n6565# a_4484_n6581# a_3215_n6746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3533 a_30985_n9268# a_31238_n9472# a_29969_n9637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3534 a_10823_884# a_11302_869# a_11510_869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3535 a_7434_359# a_8161_4650# a_8116_4663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3536 a_32975_5738# a_32554_5738# a_32286_5568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3537 a_27469_n8318# a_27256_n8318# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3538 a_25730_n4806# a_25726_n4994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3539 a_39230_5509# a_39116_5390# a_39324_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3540 a_35381_n3789# a_36442_n3624# a_36393_n3608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3541 vdd d0 a_15072_2409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3542 a_22094_7690# a_21881_7690# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3543 a_23385_n5076# a_23271_n5076# a_23479_n5076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3544 a_11374_n5440# a_11161_n5440# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3545 a_29955_n3152# a_30050_n3776# a_30001_n3760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3546 a_24400_6580# a_24598_7595# a_24549_7785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3547 a_8488_n8497# a_9546_n8935# a_9501_n8731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3548 a_18773_4848# a_18917_2666# a_18872_2679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3549 a_17502_n7049# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3550 a_40546_7211# a_41607_6840# a_41562_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3551 a_41571_5485# a_41574_4893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3552 a_37656_n6976# a_38137_n7347# a_38345_n7347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3553 a_32563_4196# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3554 a_26912_3086# a_26914_2987# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3555 a_844_1842# a_423_1842# a_155_1672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3556 a_1900_3475# a_1857_2543# a_2041_4468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3557 a_16152_n8751# a_16152_n8469# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3558 gnd d0 a_31239_n9887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3559 vdd d1 a_40803_7021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3560 a_5498_n7482# a_5987_n7783# a_6195_n7783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3561 a_1429_3055# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3562 a_136_4117# a_625_4217# a_833_4217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3563 a_40654_n5540# a_40907_n5744# a_40604_n5120# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3564 a_36297_4353# a_36550_4340# a_35284_4119# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3565 a_28514_n2675# a_28301_n2675# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3566 vdd d0 a_9781_n4039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3567 a_40541_8192# a_41602_7821# a_41553_8011# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3568 a_5520_n4244# a_5999_n4430# a_6207_n4430# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3569 a_16578_1829# a_16365_1829# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3570 a_4138_5112# a_4146_4374# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3571 gnd a_36623_n8520# a_36415_n8520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3572 a_28812_4418# a_28415_2493# a_28671_3425# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3573 a_21611_7024# a_21613_6925# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3574 a_28242_5382# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3575 a_17665_n6629# a_17452_n6629# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3576 a_30006_n2779# a_31067_n2614# a_31018_n2598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3577 vdd a_40810_6042# a_40602_6042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3578 vdd d0 a_25958_n9908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3579 a_38269_2779# a_39074_3013# a_39233_3433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3580 a_16448_n4853# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3581 a_3095_1760# a_3348_1747# a_2926_2869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3582 a_16863_n5419# a_16442_n5419# a_16174_n5048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3583 a_10883_n6812# a_10883_n6530# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3584 a_33664_n5645# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3585 gnd d5 a_35216_n10397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3586 vdd a_24950_n8693# a_24742_n8693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3587 a_27013_n2555# a_27015_n2456# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3588 vdd d1 a_8684_1165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3589 a_25644_2562# a_25647_1970# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3590 vdd a_8346_n10397# a_8138_n10397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3591 vdd a_41822_5861# a_41614_5861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3592 a_24692_n9470# a_25750_n9908# a_25701_n9892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3593 a_11485_5767# a_11064_5767# a_10796_5597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3594 a_29969_n9637# a_31030_n9472# a_30985_n9268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3595 a_22007_n2462# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3596 a_23370_7363# a_23327_6431# a_23535_6431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3597 a_8495_n7518# a_9553_n7956# a_9504_n7940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3598 a_3218_n5770# a_4279_n5605# a_4230_n5589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3599 a_6113_3781# a_6918_4015# a_7087_3573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3600 a_12913_388# a_12492_388# a_12801_4476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3601 a_6786_n7602# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3602 a_28200_3005# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3603 a_5402_7314# a_5891_7132# a_6099_7132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3604 a_12492_388# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3605 a_7171_n4907# a_6799_n4664# a_6207_n4430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3606 a_19056_7240# a_20117_6869# a_20072_6882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3607 a_5902_4757# a_5689_4757# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3608 a_33959_n6077# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3609 a_36378_n6544# a_36386_n5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3610 a_11073_4225# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3611 vdd a_24742_n8226# a_24534_n8226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3612 a_29790_n4084# a_29988_n5316# a_29943_n5112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3613 gnd a_3177_n6330# a_2969_n6330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3614 vdd a_24977_n3797# a_24769_n3797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3615 a_29866_1710# a_29961_2117# a_29916_2130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3616 a_27412_811# a_27199_811# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3617 a_40362_2650# a_40560_3665# a_40515_3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3618 a_13581_n6322# a_13725_n4346# a_13680_n4142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3619 vdd a_31174_2915# a_30966_2915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3620 a_19051_8221# a_20112_7850# a_20063_8040# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3621 vdd a_14128_n7751# a_13920_n7751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3622 a_9402_8032# a_9412_7289# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3623 a_8340_7793# a_8597_7603# a_8191_6588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3624 a_33575_4015# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3625 gnd a_25893_2936# a_25685_2936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3626 a_3160_n7307# a_3264_n6762# a_3215_n6746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3627 a_17773_367# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3628 a_32988_2800# a_32567_2800# a_32294_3016# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3629 gnd a_20426_n6568# a_20218_n6568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3630 a_1892_5432# a_1837_6460# a_2045_6460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3631 a_29770_n8001# a_29968_n9233# a_29919_n9217# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3632 a_824_5759# a_403_5759# a_130_5975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3633 a_29904_4090# a_30962_4311# a_30913_4501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3634 a_5419_3997# a_5905_3781# a_6113_3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3635 a_41660_n6938# a_41663_n6335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3636 a_3227_n4601# a_3480_n4805# a_3168_n5350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3637 gnd a_20340_3933# a_20132_3933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3638 a_38980_n8980# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3639 a_27003_n5011# a_27484_n5382# a_27692_n5382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3640 a_22417_n4837# a_23221_n4656# a_23380_n4899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3641 a_37644_n8936# a_37642_n8722# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3642 vdd d0 a_4415_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3643 vdd a_8458_n6309# a_8250_n6309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3644 a_38269_2779# a_37848_2779# a_37582_2611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3645 a_40655_n4747# a_41716_n4582# a_41671_n4378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3646 gnd d0 a_31155_7247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3647 vdd a_24895_n9254# a_24687_n9254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3648 a_33857_n9562# a_33644_n9562# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3649 a_26901_6520# a_27380_6688# a_27588_6688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3650 a_28475_1465# a_28262_1465# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3651 a_39307_n8980# a_38925_n9541# a_38334_n9722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3652 a_497_n6408# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3653 a_40604_n5120# a_40857_n5324# a_40451_n4092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3654 a_11179_n2914# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3655 a_16065_7536# a_16063_7322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3656 vdd a_31259_n5970# a_31051_n5970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3657 gnd d1 a_30157_4077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3658 a_32845_n9743# a_32632_n9743# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3659 a_39170_n3664# a_38957_n3664# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3660 a_29691_n6264# a_29835_n4288# a_29790_n4084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3661 vdd a_4379_8278# a_4171_8278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3662 a_37639_n9917# a_41900_n9895# a_40634_n9457# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3663 a_718_n4451# a_505_n4451# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3664 a_5673_8113# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3665 a_17723_7379# a_17351_6959# a_16759_6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3666 a_24325_4655# a_24578_4642# a_23643_351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3667 a_16422_n9336# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3668 a_17646_1502# a_17433_1502# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3669 a_16774_3789# a_16353_3789# a_16085_3619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3670 a_5488_n9343# a_5974_n9328# a_6182_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3671 a_11595_n3895# a_12399_n3714# a_12568_n3153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3672 a_25620_6866# a_25616_7043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3673 a_20080_5099# a_20337_4909# a_19068_5280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3674 a_12085_4044# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3675 a_16880_n2478# a_16459_n2478# a_16186_n2493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3676 gnd a_24888_2138# a_24680_2138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3677 a_23114_6431# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3678 a_11498_2829# a_11077_2829# a_10804_3045# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3679 a_2045_6460# a_1624_6460# a_1892_5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3680 a_36293_4530# a_36550_4340# a_35284_4119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3681 a_153_1458# a_642_1276# a_850_1276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3682 a_35075_n6105# a_35195_n8234# a_35150_n8030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3683 a_2835_4684# a_2955_6596# a_2910_6609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3684 a_39413_n7020# a_38992_n7020# a_39319_n7020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3685 gnd a_41904_n8499# a_41696_n8499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3686 a_40523_1895# a_40780_1705# a_40358_2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3687 a_32663_n3451# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3688 a_3118_7076# a_4176_7297# a_4127_7487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3689 a_10603_285# a_20887_141# a_20853_n686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3690 a_36292_4115# a_36302_3372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3691 a_2910_6609# a_3108_7624# a_3059_7814# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3692 a_27289_n2856# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3693 gnd a_9748_n9501# a_9540_n9501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3694 a_16167_n5815# a_16656_n5834# a_16864_n5834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3695 a_38053_4736# a_37840_4736# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3696 gnd a_40803_7021# a_40595_7021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3697 a_22115_4188# a_21902_4188# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3698 a_18872_2679# a_19070_3694# a_19025_3707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3699 gnd d0 a_9665_7276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3700 vdd d0 a_25881_6289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3701 a_8207_2848# a_8421_1726# a_8372_1916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3702 a_4150_2978# a_4403_2965# a_3134_3336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3703 a_38145_n5390# a_37932_n5390# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3704 a_27705_n3837# a_28509_n3656# a_28678_n3095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3705 a_397_7153# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3706 a_16869_n4853# a_17673_n4672# a_17832_n4915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3707 gnd a_20442_n4047# a_20234_n4047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3708 a_4235_n5816# a_4231_n6004# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3709 a_244_n3101# a_242_n2887# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3710 a_21623_5346# a_22112_5164# a_22320_5164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3711 vdd a_25982_n4595# a_25774_n4595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3712 a_906_n8368# a_485_n8368# a_212_n8383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3713 a_11588_n4874# a_11167_n4874# a_10891_n4573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3714 a_41575_5308# a_41828_5295# a_40562_5074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3715 gnd a_30107_3657# a_29899_3657# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3716 a_34038_n7041# a_33656_n7602# a_33064_n7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3717 a_9513_n6771# a_9509_n6959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3718 a_24624_3307# a_24881_3117# a_24569_3868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3719 vdd a_30231_n8672# a_30023_n8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3720 a_33073_n5826# a_33877_n5645# a_34046_n5084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3721 a_20079_5903# a_20075_6080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3722 a_11282_4786# a_11069_4786# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3723 a_7007_n5645# a_6794_n5645# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3724 a_14803_4559# a_15060_4369# a_13794_4148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3725 a_6202_n5411# a_5781_n5411# a_5508_n5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3726 a_37562_6528# a_37560_6314# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3727 a_21620_5946# a_21625_5560# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3728 a_5774_n7783# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3729 a_5513_n5040# a_5511_n4826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3730 a_4248_n3063# a_4505_n3079# a_3239_n2641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3731 a_22320_5164# a_23124_4983# a_23283_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3732 a_3239_n2641# a_4297_n3079# a_4248_n3063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3733 a_16092_2045# a_16578_1829# a_16786_1829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3734 a_24325_4655# a_24445_6567# a_24400_6580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3735 a_21734_n2477# a_22220_n2462# a_22428_n2462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3736 a_25737_n2619# a_26671_n2223# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3737 a_17626_5419# a_17413_5419# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3738 a_34172_n6077# a_33959_n6077# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3739 a_39289_2501# a_39076_2501# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3740 a_38245_8092# a_37824_8092# a_37548_8274# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3741 a_35301_1178# a_35554_1165# a_35242_1916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3742 gnd a_14141_n4813# a_13933_n4813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3743 a_5786_n4430# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3744 gnd a_25990_n4031# a_25782_n4031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3745 a_25701_n9892# a_25704_n9289# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3746 a_24650_n7278# a_24907_n7294# a_24485_n8210# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3747 a_4239_n4420# a_4235_n4608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3748 a_4158_2414# a_4411_2401# a_3145_2180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3749 a_29677_6736# a_29891_5614# a_29842_5804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3750 a_10885_n6431# a_11371_n6416# a_11579_n6416# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3751 a_25620_6866# a_25873_6853# a_24604_7224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3752 a_16070_6061# a_16072_5962# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3753 a_933_n3472# a_512_n3472# a_239_n3487# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3754 a_38042_7111# a_37829_7111# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3755 a_29904_4090# a_30962_4311# a_30917_4324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3756 vdd d0 a_41836_3338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3757 a_35272_6253# a_36333_5882# a_36288_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3758 a_4134_6508# a_4137_5916# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3759 a_37657_n5786# a_37657_n5504# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3760 a_27596_6124# a_28400_5943# a_28569_5501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3761 a_5419_4592# a_5417_4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3762 a_19160_n5757# a_20221_n5592# a_20172_n5576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3763 vdd d0 a_36554_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3764 gnd a_25963_n8927# a_25755_n8927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3765 a_4143_5350# a_4396_5337# a_3130_5116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3766 vdd a_30258_n3776# a_30050_n3776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3767 a_17868_n8077# a_17655_n8077# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3768 vdd a_15917_n10493# a_15709_n10493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3769 a_12454_n3153# a_12241_n3153# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3770 a_28544_n7012# a_28331_n7012# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3771 a_16078_4104# a_16080_4005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3772 a_5992_n6802# a_5779_n6802# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3773 a_6130_840# a_6935_1074# a_7094_1494# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3774 a_37929_n6366# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3775 a_37836_6132# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3776 a_13799_3167# a_14857_3388# a_14812_3401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3777 a_22335_2228# a_21914_2228# a_21638_2128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3778 a_3145_2180# a_3398_2167# a_3095_1760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3779 vdd a_36561_1965# a_36353_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3780 a_36289_5091# a_36297_4353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3781 gnd d0 a_36549_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3782 a_21722_n5032# a_22203_n5403# a_22411_n5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3783 a_40577_2138# a_41635_2359# a_41586_2549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3784 a_17963_n6085# a_17750_n6085# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3785 a_22409_n6794# a_21988_n6794# a_21712_n6775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3786 a_37855_1800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3787 a_17911_n9009# a_17490_n9009# a_17817_n9009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3788 gnd d2 a_19270_5651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3789 a_32274_7528# a_32755_7698# a_32963_7698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3790 a_32284_5072# a_32773_5172# a_32981_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3791 vdd d0 a_20341_4348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3792 a_21894_6145# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3793 a_35361_n7706# a_35618_n7722# a_35315_n7098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3794 gnd a_36636_n6975# a_36428_n6975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3795 a_24624_3307# a_25685_2936# a_25640_2949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3796 a_33964_1494# a_33592_1074# a_33001_1255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3797 gnd a_35467_7603# a_35259_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3798 vdd d0 a_25962_n8512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3799 a_24321_4832# a_24578_4642# a_23643_351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3800 vdd a_13838_n6338# a_13630_n6338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3801 a_9403_8447# a_9660_8257# a_8394_8036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3802 a_26990_n7354# a_26995_n6968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3803 a_25643_2147# a_25653_1404# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3804 a_37674_n2563# a_38163_n2864# a_38371_n2864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3805 a_24619_4288# a_25680_3917# a_25631_4107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3806 a_28924_330# a_29651_4621# a_29602_4811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3807 a_16876_n3874# a_16455_n3874# a_16179_n3573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3808 a_10399_n10484# a_15709_n10493# a_15660_n10477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3809 a_13811_1207# a_14064_1194# a_13752_1945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3810 a_26912_3368# a_27401_3186# a_27609_3186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3811 a_27600_4728# a_28405_4962# a_28564_5382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3812 a_12801_4476# a_12380_4476# a_12706_6468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3813 vdd a_15072_2409# a_14864_2409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3814 a_13884_n4797# a_14141_n4813# a_13829_n5358# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3815 vdd a_9761_n7956# a_9553_n7956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3816 a_32363_n8362# a_32849_n8347# a_33057_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3817 vdd d0 a_15064_2973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3818 a_5979_n8347# a_5766_n8347# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3819 a_10898_n3594# a_11387_n3895# a_11595_n3895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3820 a_16571_2808# a_16358_2808# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3821 a_7188_n3124# a_6806_n3685# a_6214_n3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3822 a_25649_1581# a_25906_1391# a_24640_1170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3823 a_2910_6609# a_3108_7624# a_3063_7637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3824 a_12536_n9030# a_12154_n9591# a_11562_n9357# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3825 a_16072_5962# a_16077_5576# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3826 vdd a_40803_7021# a_40595_7021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3827 a_39269_6418# a_39056_6418# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3828 a_23008_n4656# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3829 a_16346_6161# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3830 vdd d0 a_9665_7276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3831 gnd a_19429_n3813# a_19221_n3813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3832 vdd d0 a_15140_n7570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3833 gnd d0 a_15059_3954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3834 a_19087_2167# a_20145_2388# a_20096_2578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3835 a_25737_n2619# a_25994_n2635# a_24725_n2800# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3836 a_16365_1829# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3837 a_40356_n6084# a_40476_n8213# a_40431_n8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3838 a_500_n5432# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3839 a_23276_7482# a_22894_7924# a_22303_8105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3840 a_8207_2848# a_8421_1726# a_8376_1739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3841 gnd d0 a_25969_n7533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3842 vdd d1 a_8736_n9682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3843 a_32793_1255# a_32580_1255# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3844 a_29998_n4551# a_31056_n4989# a_31011_n4785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3845 a_27395_3752# a_27182_3752# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3846 a_9432_3372# a_9685_3359# a_8419_3138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3847 a_32390_n3466# a_32876_n3451# a_33084_n3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3848 gnd a_15128_n9530# a_14920_n9530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3849 a_6006_n3451# a_5793_n3451# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3850 a_3234_n3622# a_3487_n3826# a_3184_n3202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3851 a_19149_n8505# a_20207_n8943# a_20162_n8739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3852 a_116_8316# a_116_8034# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3853 gnd d1 a_19434_n2832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3854 a_20181_n4407# a_20177_n4595# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3855 a_33768_7932# a_33555_7932# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3856 a_17760_1621# a_17378_2063# a_16787_2244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3857 a_41554_8426# a_41557_7834# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3858 a_17822_7379# a_17401_7379# a_17723_7379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3859 a_8411_5095# a_8664_5082# a_8352_5833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3860 a_27601_5143# a_27180_5143# a_26904_5043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3861 a_5761_n9328# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3862 a_12404_n2733# a_12191_n2733# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3863 a_37849_3194# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3864 a_16754_7706# a_16333_7706# a_16065_7536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3865 a_28646_n8972# a_28264_n9533# a_27672_n9299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3866 a_30933_968# a_30929_1145# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3867 a_32368_n7482# a_32370_n7383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3868 a_25722_n6763# a_25975_n6967# a_24709_n6529# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3869 a_35210_7793# a_35314_7042# a_35265_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3870 vdd a_9672_6297# a_9464_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3871 a_20063_8040# a_20073_7297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3872 gnd d2 a_35487_3686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3873 a_37674_n2563# a_37676_n2464# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3874 a_22302_7690# a_21881_7690# a_21613_7520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3875 a_33065_n7783# a_32644_n7783# a_32368_n7764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3876 vdd a_31263_n4574# a_31055_n4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3877 a_35297_1355# a_35554_1165# a_35242_1916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3878 a_8511_n3789# a_8768_n3805# a_8465_n3181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3879 gnd d2 a_8718_n3385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3880 gnd a_3492_n2845# a_3284_n2845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3881 a_22391_n9320# a_23196_n9554# a_23365_n8993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3882 a_29677_6736# a_29891_5614# a_29846_5627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3883 a_19176_n3609# a_20234_n4047# a_20189_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3884 a_10809_2165# a_10811_2066# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3885 a_33077_n4430# a_32656_n4430# a_32383_n4445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3886 a_35311_n7286# a_35568_n7302# a_35146_n8218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3887 vdd a_9671_5882# a_9463_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3888 a_14912_n2468# a_15165_n2672# a_13896_n2837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3889 gnd a_4399_4361# a_4191_4361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3890 a_22095_8105# a_21882_8105# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3891 a_3063_7637# a_3158_8044# a_3109_8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3892 a_24692_n9470# a_24945_n9674# a_24642_n9050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3893 a_36272_8032# a_36529_7842# a_35260_8213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3894 a_37651_n7362# a_38137_n7347# a_38345_n7347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3895 a_39250_1592# a_39136_1473# a_39344_1473# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3896 a_11154_n7812# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3897 gnd d1 a_30263_n2795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3898 a_11303_1284# a_11090_1284# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3899 a_133_5375# a_133_5093# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3900 a_22396_n8339# a_21975_n8339# a_21709_n8153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3901 a_5520_n4244# a_5518_n3847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3902 a_29697_2819# a_29954_2629# a_29602_4811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3903 a_24420_2663# a_24618_3678# a_24569_3868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3904 a_6199_n6387# a_5778_n6387# a_5508_n6021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3905 a_33932_n5084# a_33719_n5084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3906 a_14795_6516# a_14798_5924# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3907 a_28514_n2675# a_28301_n2675# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3908 a_22981_1486# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3909 a_150_2058# a_636_1842# a_844_1842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3910 a_33773_6951# a_33560_6951# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3911 gnd a_41911_n7520# a_41703_n7520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3912 gnd d2 a_40768_3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3913 vdd d2 a_19270_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3914 a_8376_1739# a_8471_2146# a_8422_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3915 a_16579_2244# a_16366_2244# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3916 a_12278_7961# a_12065_7961# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3917 vdd a_4415_1005# a_4207_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3918 gnd d0 a_4487_n5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3919 a_227_n6042# a_710_n6408# a_918_n6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3920 a_27615_1792# a_27194_1792# a_26921_2008# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3921 gnd a_31155_7247# a_30947_7247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3922 a_16448_n4853# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3923 a_23392_n2939# a_23020_n2696# a_22429_n2877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3924 a_37664_n4424# a_38150_n4409# a_38358_n4409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3925 a_28262_1465# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3926 a_21643_1429# a_21643_1147# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3927 a_33567_5972# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3928 gnd d1 a_3475_n5786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3929 a_13591_2700# a_13789_3715# a_13740_3905# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3930 a_38262_5151# a_37841_5151# a_37565_5333# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3931 a_33664_n5645# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3932 gnd a_19379_n3393# a_19171_n3393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3933 a_641_861# a_428_861# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3934 a_12543_n6893# a_12171_n6650# a_11580_n6831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3935 a_6925_2522# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3936 gnd a_30157_4077# a_29949_4077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3937 a_39585_338# a_39476_338# a_37394_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3938 a_1617_7953# a_1404_7953# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3939 a_28924_330# a_29651_4621# a_29606_4634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3940 vdd a_40837_n9241# a_40629_n9241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3941 a_36393_n3608# a_36650_n3624# a_35381_n3789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3942 a_17740_5538# a_17626_5419# a_17834_5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3943 a_28497_n5616# a_28284_n5616# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3944 a_24670_n3361# a_24774_n2816# a_24725_n2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3945 a_12474_1523# a_12365_1523# a_12573_1523# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3946 a_642_1276# a_429_1276# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3947 a_22007_n2462# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3948 a_16085_3024# a_16092_2640# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3949 a_27264_n7754# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3950 a_22195_n7360# a_21982_n7360# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3951 a_3235_n2829# a_4296_n2664# a_4251_n2460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3952 a_10888_n5455# a_11374_n5440# a_11582_n5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3953 a_14909_n3071# a_14912_n2468# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3954 a_1902_n2968# a_1793_n3145# a_2001_n3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3955 a_7213_4447# a_7000_4447# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3956 a_2907_n10402# a_2857_n10418# a_2808_n10402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3957 a_17433_1502# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3958 a_32287_4378# a_32776_4196# a_32984_4196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3959 vdd d0 a_31243_n8491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3960 a_6106_6153# a_5685_6153# a_5409_6335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3961 a_21620_5946# a_22106_5730# a_22314_5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3962 a_25722_n6763# a_25718_n6951# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3963 a_23390_3446# a_23347_2514# a_23531_4439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3964 a_6930_2055# a_6717_2055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3965 a_14782_8061# a_15039_7871# a_13770_8242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3966 a_16161_n7391# a_16166_n7005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3967 a_22919_3026# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3968 a_5903_5172# a_5690_5172# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3969 a_17923_n7049# a_17868_n8077# a_18076_n8077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3970 a_40578_1334# a_41639_963# a_41590_1153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3971 vdd d4 a_19030_4658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3972 a_38365_n3430# a_37944_n3430# a_37671_n3445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3973 a_35071_n6293# a_35328_n6309# a_34959_n10381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3974 a_22208_n4422# a_21995_n4422# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3975 a_38903_5390# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3976 a_6215_n3866# a_5794_n3866# a_5518_n3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3977 a_11563_n9772# a_11142_n9772# a_10866_n9753# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3978 gnd d0 a_4410_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3979 a_818_7153# a_1622_6972# a_1781_7392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3980 a_5098_n10469# a_10656_n10500# a_10498_n10484# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3981 a_24585_1731# a_24838_1718# a_24416_2840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3982 vdd d1 a_30137_7994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3983 a_5417_4096# a_5419_3997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3984 a_23251_n8993# a_23038_n8993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3985 a_27684_n7339# a_27263_n7339# a_26995_n6968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3986 a_29917_1326# a_30978_955# a_30933_968# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3987 a_32989_3215# a_32568_3215# a_32292_3115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3988 a_29998_n4551# a_30251_n4755# a_29939_n5300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3989 a_825_6174# a_404_6174# a_128_6074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3990 a_33944_5411# a_33572_4991# a_32981_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3991 a_11498_2829# a_12303_3063# a_12462_3483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3992 a_3172_n5162# a_3267_n5786# a_3222_n5582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3993 a_21729_n4236# a_21727_n3839# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3994 a_24693_n8677# a_25754_n8512# a_25709_n8308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3995 vdd d0 a_20421_n7549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3996 a_21720_n4536# a_21722_n4437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3997 a_21906_2792# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3998 a_24642_n9050# a_24895_n9254# a_24489_n8022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3999 a_8407_5272# a_8664_5082# a_8352_5833# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4000 a_27603_3752# a_28408_3986# a_28577_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4001 a_33857_n9562# a_33644_n9562# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4002 vdd d0 a_31149_7813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4003 gnd d1 a_40919_n3784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4004 a_35210_7793# a_35314_7042# a_35269_7055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4005 a_33052_n9328# a_32631_n9328# a_32363_n8957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4006 a_39307_n8980# a_38925_n9541# a_38333_n9307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4007 a_40570_3117# a_40823_3104# a_40511_3855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4008 a_13791_5124# a_14044_5111# a_13732_5862# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4009 a_26907_4349# a_26907_4067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4010 a_2907_n10402# a_5256_n10485# a_5098_n10469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4011 gnd d0 a_9774_n5018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4012 a_26892_7285# a_27381_7103# a_27589_7103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4013 gnd d3 a_29934_6546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4014 vdd d2 a_35487_3686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4015 a_32845_n9743# a_32632_n9743# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4016 a_1798_5551# a_1416_5993# a_825_6174# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4017 gnd d0 a_20337_4909# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4018 a_32287_4378# a_32287_4096# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4019 a_39170_n3664# a_38957_n3664# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4020 a_40495_7595# a_40590_8002# a_40545_8015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4021 a_23038_n8993# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4022 vdd d3 a_35403_n8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4023 a_5917_1821# a_5704_1821# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4024 vdd d0 a_15044_6890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4025 a_39312_7350# a_39269_6418# a_39477_6418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4026 a_9517_n5002# a_9774_n5018# a_8508_n4580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4027 a_24720_n3781# a_25781_n3616# a_25736_n3412# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4028 a_26894_6904# a_26901_6520# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4029 a_27469_n8318# a_27256_n8318# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4030 vdd d0 a_25983_n5010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4031 vdd d1 a_35638_n3805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4032 a_19088_1363# a_20149_992# a_20100_1182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4033 vdd a_4399_4361# a_4191_4361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4034 a_21695_n9716# a_21695_n9434# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4035 a_36365_n9297# a_36618_n9501# a_35349_n9666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4036 a_29786_n4272# a_30000_n3356# a_29955_n3152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4037 a_3063_7637# a_3158_8044# a_3113_8057# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4038 a_31006_n4558# a_31018_n3806# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4039 a_13871_n7735# a_14932_n7570# a_14887_n7366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4040 a_24505_n4293# a_24762_n4309# a_24410_n6285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4041 vdd a_15051_5911# a_14843_5911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4042 a_17413_5419# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4043 a_39076_2501# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4044 gnd d0 a_20447_n3066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4045 a_1525_n3706# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4046 a_13656_n8247# a_13913_n8263# a_13585_n6134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4047 a_26909_3968# a_27395_3752# a_27603_3752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4048 a_9501_n8731# a_9754_n8935# a_8488_n8497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4049 a_8433_n9058# a_8528_n9682# a_8483_n9478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4050 a_24700_n7698# a_25761_n7533# a_25712_n7517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4051 vdd a_41836_3338# a_41628_3338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4052 a_3138_3159# a_3391_3146# a_3079_3897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4053 a_28443_7342# a_28230_7342# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4054 a_11499_3244# a_11078_3244# a_10802_3144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4055 a_35335_n3181# a_35430_n3805# a_35381_n3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4056 a_17844_n2955# a_17472_n2712# a_16881_n2893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4057 vdd a_36554_2944# a_36346_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4058 vdd d2 a_40768_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4059 a_32663_n3451# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4060 a_8376_1739# a_8471_2146# a_8426_2159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4061 a_40592_n7265# a_40849_n7281# a_40427_n8197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4062 a_24489_n8022# a_24742_n8226# a_24414_n6097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4063 a_21640_2624# a_22119_2792# a_22327_2792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4064 a_3109_8234# a_4170_7863# a_4125_7876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4065 vdd a_9765_n6560# a_9557_n6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4066 a_20193_n2447# a_20446_n2651# a_19177_n2816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4067 a_27496_n3422# a_27283_n3422# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4068 a_39081_2034# a_38868_2034# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4069 vdd d0 a_41899_n9480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4070 a_26588_n10440# a_32146_n10471# a_21397_n10599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4071 a_37828_6696# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4072 a_20152_n9493# a_20162_n8739# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4073 vdd d0 a_9659_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4074 a_13591_2700# a_13789_3715# a_13744_3728# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4075 a_12705_388# a_12492_388# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4076 gnd d8 a_21654_n10615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4077 a_16863_n5419# a_16442_n5419# a_16169_n5434# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4078 a_27251_n9299# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4079 gnd d0 a_9685_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4080 gnd d0 a_36535_7276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4081 a_37553_7011# a_38042_7111# a_38250_7111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4082 gnd a_41830_3904# a_41622_3904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4083 a_513_n3887# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4084 a_7193_1494# a_6772_1494# a_7099_1613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4085 a_17822_7379# a_17779_6447# a_17987_6447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4086 gnd d0 a_4505_n3079# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4087 gnd d1 a_35537_4106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4088 a_23201_n8573# a_22988_n8573# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4089 a_22983_n9554# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4090 a_838_3236# a_417_3236# a_141_3418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4091 gnd a_15141_n7985# a_14933_n7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4092 a_19090_n9254# a_19194_n8709# a_19149_n8505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4093 a_19094_n9066# a_19347_n9270# a_18941_n8038# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4094 a_41565_6051# a_41822_5861# a_40553_6232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4095 a_19080_3146# a_19333_3133# a_19021_3884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4096 a_35349_n9666# a_36410_n9501# a_36365_n9297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4097 gnd d3 a_35423_n4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4098 vdd d0 a_15166_n3087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4099 a_12310_2084# a_12097_2084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4100 a_4146_3155# a_4158_2414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4101 a_41674_n3587# a_41931_n3603# a_40662_n3768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4102 a_7007_n5645# a_6794_n5645# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4103 a_6202_n5411# a_5781_n5411# a_5513_n5040# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4104 a_24608_7047# a_25666_7268# a_25617_7458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4105 a_27168_7103# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4106 a_11283_5201# a_11070_5201# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4107 a_731_n2906# a_518_n2906# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4108 vdd a_15064_2973# a_14856_2973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4109 a_16058_8021# a_16547_8121# a_16755_8121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4110 gnd d2 a_40869_n3364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4111 a_1798_5551# a_1684_5432# a_1892_5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4112 a_30010_n2591# a_31068_n3029# a_31019_n3013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4113 a_1718_n7623# a_1505_n7623# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4114 a_39322_n4886# a_38950_n4643# a_38359_n4824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4115 a_12394_n4181# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4116 a_24573_3691# a_24668_4098# a_24619_4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4117 a_32870_n4845# a_32657_n4845# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4118 a_39136_1473# a_38923_1473# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4119 a_39056_6418# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4120 a_1895_n5105# a_1513_n5666# a_922_n5847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4121 a_933_n3472# a_512_n3472# a_244_n3101# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4122 a_32856_n7368# a_32643_n7368# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4123 a_38068_1800# a_37855_1800# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4124 a_22111_4749# a_21898_4749# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4125 a_26894_7499# a_27375_7669# a_27583_7669# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4126 vdd d1 a_14136_n5794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4127 a_20182_n4822# a_20435_n5026# a_19169_n4588# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4128 a_9515_n5380# a_9768_n5584# a_8499_n5749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4129 vdd d3 a_40615_2637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4130 a_4133_6093# a_4390_5903# a_3121_6274# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4131 a_32383_n5040# a_32381_n4826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4132 a_32580_1255# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4133 gnd d0 a_20434_n4611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4134 a_5992_n6802# a_5779_n6802# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4135 a_40352_n6272# a_40609_n6288# a_40240_n10360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4136 a_37929_n6366# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4137 gnd d0 a_15045_7305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4138 a_27182_3752# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4139 a_17743_3462# a_17371_3042# a_16780_3223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4140 a_27387_5709# a_27174_5709# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4141 a_21717_n5418# a_22203_n5403# a_22411_n5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4142 vdd d1 a_24982_n2816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4143 a_13787_5301# a_14044_5111# a_13732_5862# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4144 a_8280_n8030# a_8478_n9262# a_8433_n9058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4145 a_6199_n6387# a_7004_n6621# a_7163_n6864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4146 a_2920_n6314# a_3064_n4338# a_3019_n4134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4147 a_13492_4869# a_13636_2687# a_13591_2700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4148 vdd d3 a_29934_6546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4149 a_622_5193# a_409_5193# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4150 a_37856_2215# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4151 a_35166_n4301# a_35380_n3385# a_35331_n3369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4152 a_33555_7932# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4153 a_32267_8295# a_32756_8113# a_32964_8113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4154 a_14884_n7969# a_15141_n7985# a_13875_n7547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4155 a_21720_n4818# a_21720_n4536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4156 a_8500_n6537# a_8753_n6741# a_8441_n7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4157 gnd d2 a_19290_1734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4158 a_17655_n8077# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4159 vdd a_36639_n5999# a_36431_n5999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4160 vdd d0 a_36644_n5018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4161 vdd a_9664_6861# a_9456_6861# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4162 a_37674_n2845# a_38163_n2864# a_38371_n2864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4163 vdd d0 a_4395_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4164 a_30921_2928# a_31174_2915# a_29905_3286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4165 a_19067_6084# a_20125_6305# a_20080_6318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4166 a_5493_n8957# a_5974_n9328# a_6182_n9328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4167 a_25648_2385# a_25901_2372# a_24635_2151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4168 a_39334_n2926# a_39225_n3103# a_39433_n3103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4169 a_23347_2514# a_23134_2514# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4170 a_29981_n7677# a_31042_n7512# a_30993_n7496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4171 a_3134_3336# a_3391_3146# a_3079_3897# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4172 a_9512_n5983# a_9515_n5380# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4173 a_7176_n5084# a_7062_n5084# a_7270_n5084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4174 gnd d0 a_36624_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4175 a_16423_n9751# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4176 a_14897_n5031# a_15154_n5047# a_13888_n4609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4177 a_5979_n8347# a_5766_n8347# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4178 a_29770_n8001# a_30023_n8205# a_29695_n6076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4179 a_33058_n8762# a_33862_n8581# a_34021_n8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4180 a_21734_n2477# a_21123_n2239# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4181 a_11090_1284# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4182 a_24635_2151# a_24888_2138# a_24585_1731# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4183 a_16572_3223# a_16359_3223# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4184 a_5397_8295# a_5397_8013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4185 a_8499_n5749# a_9560_n5584# a_9515_n5380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4186 a_8410_4296# a_8667_4106# a_8364_3699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4187 a_16172_n4834# a_16172_n4552# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4188 a_30916_3909# a_30912_4086# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4189 a_40634_n9457# a_40887_n9661# a_40584_n9037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4190 a_33090_n2885# a_32669_n2885# a_32393_n2584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4191 a_33560_6951# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4192 vdd d0 a_9761_n7956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4193 a_500_n5432# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4194 a_40616_n3160# a_40711_n3784# a_40662_n3768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4195 a_28351_n3095# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4196 a_16366_2244# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4197 a_12065_7961# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4198 a_30929_2364# a_31182_2351# a_29916_2130# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4199 vdd d0 a_36535_7276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4200 a_40550_7034# a_40803_7021# a_40491_7772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4201 a_16791_848# a_17596_1082# a_17755_1502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4202 a_19145_n8693# a_20206_n8528# a_20157_n8512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4203 a_6006_n3451# a_5793_n3451# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4204 a_8211_2671# a_8464_2658# a_8112_4840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4205 a_35289_3138# a_36347_3359# a_36302_3372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4206 a_33644_n9562# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4207 a_10903_n2895# a_10903_n2613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4208 a_1404_7953# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4209 a_9439_2393# a_9435_2570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4210 a_19076_3323# a_19333_3133# a_19021_3884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4211 gnd a_24907_n7294# a_24699_n7294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4212 a_10816_1680# a_11297_1850# a_11505_1850# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4213 a_26921_2603# a_26919_2389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4214 gnd a_31271_n4010# a_31063_n4010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4215 a_39165_n4131# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4216 gnd d0 a_31187_1370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4217 vdd a_35611_n8701# a_35403_n8701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4218 a_5690_5172# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4219 a_22392_n9735# a_23196_n9554# a_23365_n8993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4220 a_13794_4148# a_14852_4369# a_14807_4382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4221 a_9431_2957# a_9427_3134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4222 vdd d0 a_9748_n9501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4223 a_21714_n6989# a_21712_n6775# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4224 vdd d0 a_20447_n3066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4225 a_20095_2163# a_20105_1420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4226 a_38037_8092# a_37824_8092# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4227 a_22307_6709# a_21886_6709# a_21620_6541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4228 gnd d0 a_36638_n5584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4229 a_11154_n7812# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4230 a_38346_n7762# a_39150_n7581# a_39319_n7020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4231 a_7089_n6077# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4232 vdd a_30137_7994# a_29929_7994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4233 a_16552_7140# a_16339_7140# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4234 a_38061_2779# a_37848_2779# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4235 a_10883_n6530# a_11372_n6831# a_11580_n6831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4236 a_693_n9349# a_480_n9349# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4237 a_14881_n8760# a_14877_n8948# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4238 gnd a_41810_7821# a_41602_7821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4239 a_11493_3810# a_11072_3810# a_10804_3640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4240 a_41680_n3021# a_41683_n2418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4241 gnd a_8597_7603# a_8389_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4242 a_9533_n2854# a_9786_n3058# a_8520_n2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4243 vdd d0 a_4504_n2664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4244 gnd d1 a_35517_8023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4245 gnd d0 a_25995_n3050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4246 a_39661_n6056# a_39240_n6056# a_39562_n5879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4247 a_36361_n9485# a_36371_n8731# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4248 a_40635_n8664# a_41696_n8499# a_41651_n8295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4249 vdd d2 a_19290_1734# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4250 a_217_n7785# a_217_n7503# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4251 vdd a_20320_7850# a_20112_7850# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4252 vdd d0 a_41912_n7935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4253 gnd d1 a_30246_n5736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4254 a_32393_n2866# a_32393_n2584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4255 a_13900_n2649# a_14958_n3087# a_14913_n2883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4256 a_36310_1589# a_36567_1399# a_35301_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4257 gnd a_35618_n7722# a_35410_n7722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4258 gnd d1 a_35623_n6741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4259 gnd a_29934_6546# a_29726_6546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4260 a_32963_7698# a_32542_7698# a_32269_7914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4261 gnd a_20337_4909# a_20129_4909# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4262 a_12650_n5113# a_12607_n4181# a_12791_n5929# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4263 a_25644_2562# a_25901_2372# a_24635_2151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4264 a_28497_n5616# a_28284_n5616# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4265 a_5704_1821# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4266 vdd a_15044_6890# a_14836_6890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4267 a_40447_n4280# a_40661_n3364# a_40612_n3348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4268 a_31014_n3994# a_31271_n4010# a_30005_n3572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4269 a_27264_n7754# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4270 a_17750_n6085# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4271 a_7302_n6077# a_7089_n6077# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4272 a_10888_n6050# a_10886_n5836# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4273 a_24553_7608# a_24648_8015# a_24599_8205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4274 a_39358_n8048# a_39145_n8048# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4275 gnd a_41900_n9895# a_41692_n9895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4276 a_20165_n7948# a_20422_n7964# a_19156_n7526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4277 a_832_3802# a_411_3802# a_138_4018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4278 a_26993_n6472# a_27482_n6773# a_27690_n6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4279 a_23385_n5076# a_23003_n5637# a_22412_n5818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4280 a_16547_8121# a_16334_8121# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4281 a_13752_1945# a_13856_1194# a_13807_1384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4282 a_5419_4592# a_5902_4757# a_6110_4757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4283 a_212_n8383# a_219_n8182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4284 a_13833_n5170# a_13928_n5794# a_13883_n5590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4285 vdd d0 a_41925_n4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4286 a_23308_1605# a_23194_1486# a_23402_1486# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4287 a_10811_2066# a_10816_1680# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4288 a_28230_7342# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4289 a_23174_5403# a_22961_5403# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4290 a_29866_1710# a_29961_2117# a_29912_2307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4291 a_15842_n2260# a_16672_n2478# a_16880_n2478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4292 a_22208_n4422# a_21995_n4422# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4293 gnd a_25885_4893# a_25677_4893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4294 a_32361_n8461# a_32850_n8762# a_33058_n8762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4295 a_16844_n9751# a_17648_n9570# a_17817_n9009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4296 a_6215_n3866# a_5794_n3866# a_5518_n3565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4297 a_30925_2541# a_31182_2351# a_29916_2130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4298 a_11510_869# a_11089_869# a_10816_1085# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4299 a_40546_7211# a_40803_7021# a_40491_7772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4300 a_11563_n9772# a_11142_n9772# a_10866_n9471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4301 a_6791_n6621# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4302 vdd a_8761_n4784# a_8553_n4784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4303 a_16058_8303# a_16058_8021# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4304 gnd d1 a_14027_8052# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4305 a_23719_n6069# a_23298_n6069# a_23624_n8061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4306 a_37844_4175# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4307 a_12241_n3153# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4308 a_32788_2236# a_32575_2236# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4309 gnd a_31170_4311# a_30962_4311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4310 a_19157_n6733# a_19414_n6749# a_19102_n7294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4311 a_32559_4757# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4312 a_7250_n9001# a_7207_n8069# a_7415_n8069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4313 a_135_4994# a_621_4778# a_829_4778# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4314 a_29943_n5112# a_30038_n5736# a_29993_n5532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4315 vdd a_19422_n4792# a_19214_n4792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4316 a_237_n3586# a_726_n3887# a_934_n3887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4317 a_14820_1618# a_15077_1428# a_13811_1207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4318 a_22320_5164# a_21899_5164# a_21623_5346# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4319 a_11473_7727# a_11052_7727# a_10779_7943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4320 gnd a_36535_7276# a_36327_7276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4321 a_35378_n4580# a_36436_n5018# a_36391_n4814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4322 a_4921_292# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4323 a_21709_n7375# a_22195_n7360# a_22403_n7360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4324 gnd d1 a_19340_2154# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4325 a_28703_4418# a_28490_4418# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4326 a_5761_n9328# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4327 gnd a_14116_n9711# a_13908_n9711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4328 a_39012_n3103# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4329 a_30914_5300# a_30910_5477# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4330 gnd a_35537_4106# a_35329_4106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4331 a_27596_6124# a_27175_6124# a_26899_6306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4332 a_28792_n6048# a_28579_n6048# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4333 a_11386_n3480# a_11173_n3480# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4334 a_35081_2671# a_35279_3686# a_35230_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4335 vdd d0 a_31187_1370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4336 a_35358_n8497# a_36416_n8935# a_36367_n8919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4337 a_9521_n4814# a_9517_n5002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4338 a_33642_1494# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4339 gnd a_4379_8278# a_4171_8278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4340 a_11070_5201# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4341 a_36378_n6544# a_36635_n6560# a_35366_n6725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4342 a_34403_359# a_33982_359# a_34291_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4343 vdd d0 a_20410_n9924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4344 a_29986_n6696# a_30243_n6712# a_29931_n7257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4345 gnd d1 a_8773_n2824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4346 a_37562_5933# a_38048_5717# a_38256_5717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4347 a_7062_n5084# a_6849_n5084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4348 a_4228_n6980# a_4485_n6996# a_3219_n6558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4349 gnd d1 a_14121_n8730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4350 vdd a_36643_n4603# a_36435_n4603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4351 a_18072_n5908# a_17675_n4160# a_17931_n5092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4352 a_26978_n9909# a_31239_n9887# a_29973_n9449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4353 a_1525_n3706# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4354 a_28425_1045# a_28212_1045# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4355 a_22396_n8339# a_21975_n8339# a_21702_n8354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4356 vdd d0 a_20358_1407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4357 a_7168_n7041# a_7054_n7041# a_7262_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4358 a_25721_n5975# a_25724_n5372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4359 a_17844_n2955# a_17472_n2712# a_16880_n2478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4360 vdd a_8706_n5345# a_8498_n5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4361 a_11298_2265# a_11085_2265# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4362 a_11069_4786# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4363 a_40582_1157# a_41640_1378# a_41595_1391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4364 a_11375_n5855# a_11162_n5855# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4365 a_5431_2632# a_5429_2418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4366 vdd d1 a_35517_8023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4367 vdd d0 a_25888_3917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4368 a_28463_3425# a_28250_3425# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4369 a_27496_n3422# a_27283_n3422# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4370 a_37649_n7461# a_38138_n7762# a_38346_n7762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4371 gnd a_4473_n8956# a_4265_n8956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4372 a_12434_n7070# a_12221_n7070# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4373 gnd a_15045_7305# a_14837_7305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4374 a_3198_n9687# a_3455_n9703# a_3152_n9079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4375 a_27174_5709# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4376 a_19114_n5149# a_19209_n5773# a_19160_n5757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4377 a_13680_n4142# a_13878_n5374# a_13833_n5170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4378 gnd a_36651_n4039# a_36443_n4039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4379 gnd d0 a_36656_n3058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4380 a_11599_n2499# a_12404_n2733# a_12563_n2976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4381 gnd d0 a_25905_976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4382 vdd d1 a_19402_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4383 a_6849_n5084# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4384 a_5491_n8461# a_5493_n8362# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4385 a_37671_n4223# a_38150_n4409# a_38358_n4409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4386 gnd a_40899_n7701# a_40691_n7701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4387 a_23479_n5076# a_23058_n5076# a_23385_n5076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4388 vdd d2 a_3425_n5366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4389 vdd a_29934_6546# a_29726_6546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4390 a_34051_3454# a_34008_2522# a_34192_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4391 a_5511_n4544# a_6000_n4845# a_6208_n4845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4392 a_22423_n3443# a_22002_n3443# a_21729_n3458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4393 a_4226_n7358# a_4222_n7546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4394 vdd d0 a_9679_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4395 a_32306_1056# a_32792_840# a_33000_840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4396 vdd d0 a_36529_7842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4397 a_17812_n8832# a_17703_n9009# a_17911_n9009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4398 a_17510_n5092# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4399 a_26983_n8333# a_27469_n8318# a_27677_n8318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4400 a_30910_5477# a_30913_4885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4401 gnd d3 a_35314_6575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4402 a_24553_7608# a_24648_8015# a_24603_8028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4403 a_23201_n8573# a_22988_n8573# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4404 a_22983_n9554# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4405 a_19161_n6545# a_20219_n6983# a_20170_n6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4406 a_10893_n5069# a_11374_n5440# a_11582_n5440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4407 a_23370_7363# a_22949_7363# a_23271_7363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4408 a_408_4778# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4409 a_36294_5329# a_36290_5506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4410 gnd d0 a_15076_1013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4411 vdd a_9754_n8935# a_9546_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4412 vdd a_4395_4922# a_4187_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4413 a_27010_n3437# a_27015_n3051# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4414 a_35246_1739# a_35499_1726# a_35077_2848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4415 a_27485_n5797# a_27272_n5797# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4416 gnd d1 a_40904_n6720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4417 a_23134_2514# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4418 a_10789_6364# a_10789_6082# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4419 a_24628_3130# a_24881_3117# a_24569_3868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4420 a_3184_n3202# a_3437_n3406# a_3015_n4322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4421 a_32984_4196# a_32563_4196# a_32287_4096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4422 a_29973_n9449# a_31031_n9887# a_26978_n9909# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4423 a_39155_n6600# a_38942_n6600# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4424 a_27709_n2441# a_28514_n2675# a_28673_n2918# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4425 a_5898_6153# a_5685_6153# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4426 a_731_n2906# a_518_n2906# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4427 a_24599_8205# a_25660_7834# a_25615_7847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4428 a_14807_4382# a_15060_4369# a_13794_4148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4429 gnd a_14066_n9291# a_13858_n9291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4430 a_39322_n4886# a_38950_n4643# a_38358_n4409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4431 a_1718_n7623# a_1505_n7623# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4432 a_12541_7400# a_12120_7400# a_12442_7400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4433 a_38143_n6781# a_37930_n6781# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4434 gnd d0 a_4488_n6020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4435 a_24325_4655# a_24445_6567# a_24396_6757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4436 a_10898_n3876# a_10898_n3594# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4437 gnd a_31275_n2614# a_31067_n2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4438 a_32870_n4845# a_32657_n4845# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4439 gnd d1 a_19409_n7730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4440 vdd d1 a_14027_8052# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4441 a_1895_n5105# a_1513_n5666# a_921_n5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4442 a_16583_848# a_16370_848# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4443 vdd a_31170_4311# a_30962_4311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4444 a_34033_n6864# a_33661_n6621# a_33070_n6802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4445 a_9528_n2627# a_9785_n2643# a_8516_n2808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4446 a_27684_n7339# a_27263_n7339# a_26990_n7354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4447 gnd d0 a_41836_3338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4448 a_26887_8266# a_27376_8084# a_27584_8084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4449 a_40646_n7497# a_41704_n7935# a_41659_n7731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4450 vdd a_36535_7276# a_36327_7276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4451 a_37553_7011# a_37555_6912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4452 a_35311_n7286# a_35415_n6741# a_35366_n6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4453 vdd d1 a_19340_2154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4454 a_35058_n10381# a_35008_n10397# a_34959_n10381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4455 a_4226_n7358# a_4479_n7562# a_3210_n7727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4456 a_8191_6588# a_8389_7603# a_8340_7793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4457 vdd d0 a_15039_7871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4458 a_21611_7024# a_22100_7124# a_22308_7124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4459 a_35378_n4580# a_35631_n4784# a_35319_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4460 gnd a_4487_n5605# a_4279_n5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4461 gnd d3 a_13824_6604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4462 a_10893_n4474# a_10900_n4273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4463 gnd d1 a_40815_5061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4464 a_6200_n6802# a_7004_n6621# a_7163_n6864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4465 a_33052_n9328# a_32631_n9328# a_32358_n9343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4466 a_21709_n8153# a_21707_n7756# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4467 a_14887_n7366# a_15140_n7570# a_13871_n7735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4468 a_4126_7072# a_4138_6331# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4469 a_34043_5411# a_33988_6439# a_34196_6439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4470 a_33912_n9001# a_33699_n9001# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4471 a_39230_5509# a_38848_5951# a_38257_6132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4472 a_35081_2671# a_35279_3686# a_35234_3699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4473 a_21700_n8453# a_21702_n8354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4474 a_27697_n4401# a_27276_n4401# a_27003_n4416# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4475 a_21652_847# a_22131_832# a_22339_832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4476 gnd d0 a_20341_4348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4477 gnd a_13913_n8263# a_13705_n8263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4478 vdd d4 a_3177_n6330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4479 a_16085_3619# a_16566_3789# a_16774_3789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4480 a_40659_n4559# a_41717_n4997# a_41672_n4793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4481 a_13732_5862# a_13836_5111# a_13787_5301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4482 gnd d0 a_15154_n5047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4483 a_18961_n4121# a_19159_n5353# a_19110_n5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4484 a_23288_5522# a_23174_5403# a_23382_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4485 a_9407_8270# a_9660_8257# a_8394_8036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4486 a_604_7719# a_391_7719# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4487 gnd a_25888_3917# a_25680_3917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4488 a_498_n6823# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4489 a_39238_3552# a_38856_3994# a_38264_3760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4490 gnd a_40849_n7281# a_40641_n7281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4491 a_39476_338# a_39263_338# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4492 a_21633_3603# a_22114_3773# a_22322_3773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4493 a_838_3236# a_1642_3055# a_1801_3475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4494 a_16459_n2478# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4495 gnd a_3472_n6762# a_3264_n6762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4496 vdd d1 a_24957_n7714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4497 a_22126_1813# a_21913_1813# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4498 a_16423_n9751# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4499 a_1672_7392# a_1459_7392# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4500 gnd d6 a_5256_n10485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4501 a_37824_8092# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4502 a_22323_4188# a_21902_4188# a_21626_4370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4503 a_41659_n6523# a_41916_n6539# a_40647_n6704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4504 a_6994_n8069# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4505 a_41579_3528# a_41836_3338# a_40570_3117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4506 a_28740_n8972# a_28697_n8040# a_28905_n8040# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4507 a_16881_n2893# a_16460_n2893# a_16184_n2874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4508 a_21982_n7360# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4509 a_3210_n7727# a_4271_n7562# a_4226_n7358# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4510 a_17653_n8589# a_17440_n8589# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4511 a_1870_n8845# a_1498_n8602# a_907_n8783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4512 a_37555_6912# a_37562_6528# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4513 a_918_n6408# a_497_n6408# a_227_n6042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4514 a_32304_1437# a_32793_1255# a_33001_1255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4515 a_21914_2228# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4516 gnd a_35517_8023# a_35309_8023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4517 a_2995_n8239# a_3252_n8255# a_2924_n6126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4518 a_40358_2827# a_40572_1705# a_40523_1895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4519 a_18862_n6301# a_19006_n4325# a_18957_n4309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4520 a_10802_3426# a_10802_3144# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4521 a_7183_n2947# a_6811_n2704# a_6220_n2885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4522 vdd d3 a_35314_6575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4523 a_27608_2771# a_27187_2771# a_26921_2603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4524 vdd d0 a_15076_1013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4525 gnd d0 a_41937_n3037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4526 a_33644_n9562# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4527 a_38370_n2449# a_37949_n2449# a_37332_n2231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4528 a_35242_1916# a_35499_1726# a_35077_2848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4529 a_39061_5951# a_38848_5951# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4530 a_12229_n5113# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4531 a_6985_1494# a_6772_1494# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4532 a_33944_5411# a_33835_5411# a_34043_5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4533 a_8461_n3369# a_8565_n2824# a_8516_n2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4534 a_34982_4840# a_35126_2658# a_35081_2671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4535 a_17987_6447# a_17566_6447# a_17834_5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4536 a_13809_n9275# a_13913_n8730# a_13864_n8714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4537 a_27621_1226# a_28425_1045# a_28584_1465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4538 gnd d7 a_32146_n10471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4539 a_10809_2447# a_11298_2265# a_11506_2265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4540 a_36301_2957# a_36554_2944# a_35285_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4541 a_1719_4468# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4542 vdd a_25983_n5010# a_25775_n5010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4543 a_907_n8783# a_486_n8783# a_210_n8764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4544 a_16334_8121# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4545 a_11278_6182# a_11065_6182# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4546 a_26733_263# a_28602_330# a_28924_330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4547 a_9504_n7940# a_9507_n7337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4548 a_32284_5072# a_32286_4973# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4549 vdd a_15134_n8964# a_14926_n8964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4550 a_20089_3557# a_20346_3367# a_19080_3146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4551 a_9496_n8504# a_9508_n7752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4552 a_28602_330# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4553 a_14812_3401# a_14808_3578# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4554 a_32856_n7368# a_32643_n7368# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4555 a_32781_3215# a_32568_3215# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4556 a_1892_5432# a_1471_5432# a_1793_5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4557 a_20157_n8512# a_20414_n8528# a_19145_n8693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4558 a_35390_n2620# a_36448_n3058# a_36399_n3042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4559 vdd a_13749_4679# a_13541_4679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4560 a_23296_3565# a_22914_4007# a_22322_3773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4561 a_38345_n7347# a_37924_n7347# a_37651_n7362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4562 a_28641_n8795# a_28269_n8552# a_27678_n8733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4563 a_4145_3959# a_4398_3946# a_3129_4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4564 a_39473_4426# a_39364_4426# a_39572_4426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4565 vdd d0 a_36655_n2643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4566 a_22106_5730# a_21893_5730# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4567 a_8116_4663# a_8369_4650# a_7434_359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4568 a_16164_n6791# a_16164_n6509# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4569 gnd d1 a_8672_3125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4570 a_32292_3115# a_32294_3016# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4571 gnd a_14027_8052# a_13819_8052# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4572 a_40604_n5120# a_40699_n5744# a_40650_n5728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4573 a_28339_n5055# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4574 a_40558_5251# a_41619_4880# a_41574_4893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4575 a_5787_n4845# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4576 a_30990_n8287# a_31243_n8491# a_29974_n8656# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4577 vdd d2 a_24915_n5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4578 a_32575_2236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4579 a_14888_n6573# a_14896_n5824# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4580 a_29701_2642# a_29954_2629# a_29602_4811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4581 a_10883_n6812# a_11372_n6831# a_11580_n6831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4582 a_38062_3194# a_37849_3194# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4583 vdd d1 a_40815_5061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4584 a_14892_n6012# a_14895_n5409# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4585 a_32968_6717# a_33773_6951# a_33932_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4586 a_22894_7924# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4587 a_19164_n5569# a_20222_n6007# a_20173_n5991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4588 a_36309_2393# a_36562_2380# a_35296_2159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4589 a_7151_n8824# a_7042_n9001# a_7250_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4590 a_40553_6232# a_41614_5861# a_41565_6051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4591 a_13656_n8247# a_13870_n7331# a_13825_n7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4592 a_28490_4418# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4593 a_13732_5862# a_13836_5111# a_13791_5124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4594 a_1479_3475# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4595 a_18868_2856# a_19082_1734# a_19033_1924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4596 a_25628_6302# a_25881_6289# a_24615_6068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4597 a_38281_819# a_39086_1053# a_39245_1473# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4598 a_14811_2986# a_15064_2973# a_13795_3344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4599 gnd d4 a_19119_n6317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4600 a_40659_n4559# a_40912_n4763# a_40600_n5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4601 a_27199_811# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4602 a_32964_8113# a_32543_8113# a_32267_8013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4603 a_3126_5293# a_4187_4922# a_4142_4935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4604 a_225_n5546# a_227_n5447# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4605 a_32299_2418# a_32299_2136# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4606 a_11473_7727# a_12278_7961# a_12447_7519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4607 a_20168_n7345# a_20421_n7549# a_19152_n7714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4608 gnd a_30043_n4288# a_29835_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4609 vdd a_41917_n6954# a_41709_n6954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4610 vdd d0 a_25963_n8927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4611 a_23208_n7594# a_22995_n7594# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4612 a_21881_7690# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4613 a_29905_3286# a_30966_2915# a_30917_3105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4614 vdd d0 a_9676_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4615 a_26906_4944# a_26909_4563# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4616 a_11291_3244# a_11078_3244# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4617 a_26993_n6754# a_27482_n6773# a_27690_n6773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4618 a_23385_n5076# a_23003_n5637# a_22411_n5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4619 a_6125_1821# a_6930_2055# a_7099_1613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4620 a_17983_4455# a_17874_4455# a_18082_4455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4621 a_12913_388# a_15795_300# a_10504_285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4622 a_12568_n3153# a_12454_n3153# a_12662_n3153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4623 a_32286_4973# a_32289_4592# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4624 a_5414_5354# a_5903_5172# a_6111_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4625 a_28212_1045# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4626 vdd a_20358_1407# a_20150_1407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4627 a_14808_3578# a_14811_2986# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4628 a_34285_n8069# a_33864_n8069# a_34132_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4629 a_16567_4204# a_16354_4204# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4630 a_11085_2265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4631 vdd a_15148_n5613# a_14940_n5613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4632 a_16075_5362# a_16564_5180# a_16772_5180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4633 a_33793_3034# a_33580_3034# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4634 a_22949_7363# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4635 gnd d4 a_19030_4658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4636 vdd d1 a_30238_n7693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4637 a_32643_n7368# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4638 a_32361_n8743# a_32850_n8762# a_33058_n8762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4639 vdd a_35517_8023# a_35309_8023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4640 a_28250_3425# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4641 a_6791_n6621# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4642 a_19063_6261# a_20124_5890# a_20075_6080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4643 gnd a_25977_n5576# a_25769_n5576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4644 a_26489_n10440# a_26746_n10456# a_26588_n10440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4645 gnd d0 a_20345_2952# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4646 a_6111_5172# a_6915_4991# a_7074_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4647 a_33587_2055# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4648 gnd a_25905_976# a_25697_976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4649 a_5431_2037# a_5436_1651# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4650 a_35061_6588# a_35259_7603# a_35214_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4651 a_38282_1234# a_37861_1234# a_37585_1134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4652 a_36309_2393# a_36305_2570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4653 a_40515_3678# a_40768_3665# a_40362_2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4654 a_12374_n8098# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4655 a_41574_4893# a_41570_5070# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4656 a_2808_n10402# a_2969_n6330# a_2924_n6126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4657 a_1637_4036# a_1424_4036# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4658 a_29916_2130# a_30974_2351# a_30925_2541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4659 a_9411_6874# a_9664_6861# a_8395_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4660 vdd a_24555_n10389# a_24347_n10389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4661 a_13888_n4609# a_14946_n5047# a_14897_n5031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4662 vdd a_24982_n2816# a_24774_n2816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4663 a_16843_n9336# a_16422_n9336# a_16149_n9351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4664 vdd d4 a_24667_n6301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4665 a_11474_8142# a_11053_8142# a_10777_8042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4666 gnd d0 a_25970_n7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4667 vdd a_14133_n6770# a_13925_n6770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4668 a_39218_7469# a_38836_7911# a_38244_7677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4669 gnd a_35314_6575# a_35106_6575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4670 gnd d0 a_31167_5287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4671 a_17743_3462# a_17634_3462# a_17842_3462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4672 gnd a_15076_1013# a_14868_1013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4673 a_6126_2236# a_5705_2236# a_5429_2136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4674 a_24654_n7090# a_24749_n7714# a_24704_n7510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4675 a_26909_4563# a_27392_4728# a_27600_4728# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4676 a_5891_7132# a_5678_7132# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4677 gnd a_24962_n6733# a_24754_n6733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4678 a_40634_n9457# a_41692_n9895# a_41643_n9879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4679 a_36301_2957# a_36297_3134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4680 a_31672_256# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4681 a_10871_n8490# a_10873_n8391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4682 gnd d0 a_20409_n9509# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4683 a_18937_n8226# a_19151_n7310# a_19102_n7294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4684 a_5685_6153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4685 a_17735_5419# a_17363_4999# a_16771_4765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4686 a_8415_3315# a_9476_2944# a_9431_2957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4687 a_11511_1284# a_11090_1284# a_10814_1466# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4688 a_9412_7289# a_9408_7466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4689 a_12303_3063# a_12090_3063# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4690 a_28484_n8040# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4691 a_205_n9463# a_207_n9364# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4692 a_33862_n8581# a_33649_n8581# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4693 vdd a_41931_n3603# a_41723_n3603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4694 a_8112_4840# a_8369_4650# a_7434_359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4695 vdd a_40684_n8213# a_40476_n8213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4696 a_30999_n6930# a_31256_n6946# a_29990_n6508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4697 vdd d1 a_8672_3125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4698 vdd a_14027_8052# a_13819_8052# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4699 vdd a_31264_n4989# a_31056_n4989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4700 a_813_8134# a_392_8134# a_116_8316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4701 a_29854_3670# a_29949_4077# a_29904_4090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4702 a_28671_3425# a_28628_2493# a_28812_4418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4703 vdd d0 a_15128_n9530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4704 a_8410_4296# a_9471_3925# a_9422_4115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4705 gnd d0 a_9780_n3624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4706 a_30893_8418# a_30896_7826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4707 a_17579_4023# a_17366_4023# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4708 a_41659_n7731# a_41655_n7919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4709 a_12097_2084# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4710 a_40338_6744# a_40552_5622# a_40503_5812# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4711 a_37840_4736# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4712 a_33078_n4845# a_32657_n4845# a_32381_n4826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4713 gnd a_41836_3338# a_41628_3338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4714 vdd a_20415_n8943# a_20207_n8943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4715 a_693_n9349# a_480_n9349# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4716 a_11375_n5855# a_11162_n5855# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4717 a_36305_2570# a_36562_2380# a_35296_2159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4718 a_36277_8270# a_36273_8447# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4719 gnd d0 a_25957_n9493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4720 vdd d0 a_36619_n9916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4721 a_40671_n2599# a_41729_n3037# a_41680_n3021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4722 a_37649_n7743# a_38138_n7762# a_38346_n7762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4723 gnd a_36550_4340# a_36342_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4724 a_29969_n9637# a_30226_n9653# a_29923_n9029# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4725 a_11600_n2914# a_12404_n2733# a_12563_n2976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4726 a_4211_n9921# a_4468_n9937# a_3202_n9499# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4727 a_7411_n5900# a_7014_n4152# a_7282_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4728 a_36367_n8919# a_36624_n8935# a_35358_n8497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4729 gnd a_13824_6604# a_13616_6604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4730 vdd a_21654_n10615# a_21446_n10615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4731 a_18868_2856# a_19082_1734# a_19037_1747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4732 gnd a_40815_5061# a_40607_5061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4733 a_5511_n4826# a_6000_n4845# a_6208_n4845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4734 a_22423_n3443# a_22002_n3443# a_21734_n3072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4735 a_32301_2037# a_32787_1821# a_32995_1821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4736 a_13883_n5590# a_14136_n5794# a_13833_n5170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4737 a_33982_359# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4738 vdd a_20442_n4047# a_20234_n4047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4739 a_11574_n7397# a_11153_n7397# a_10885_n7026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4740 a_222_n6522# a_711_n6823# a_919_n6823# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4741 a_23303_1486# a_22931_1066# a_22339_832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4742 a_7067_7490# a_6685_7932# a_6094_8113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4743 a_4162_1018# a_4415_1005# a_3146_1376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4744 vref a_116_8316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4745 a_391_7719# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4746 a_409_5193# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4747 a_32361_n8461# a_32363_n8362# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4748 a_25736_n3412# a_25989_n3616# a_24720_n3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4749 a_35386_n2808# a_36447_n2643# a_36402_n2439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4750 gnd a_30119_1697# a_29911_1697# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4751 a_29955_n3152# a_30208_n3356# a_29786_n4272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4752 a_29951_n3340# a_30055_n2795# a_30010_n2591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4753 a_24636_1347# a_24893_1157# a_24581_1908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4754 a_9408_7466# a_9411_6874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4755 a_1969_n9022# a_1548_n9022# a_1870_n8845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4756 a_37932_n5390# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4757 a_3239_n2641# a_4297_n3079# a_4252_n2875# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4758 a_27710_n2856# a_28514_n2675# a_28673_n2918# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4759 a_22196_n7775# a_21983_n7775# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4760 a_26981_n8714# a_26981_n8432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4761 a_12474_1523# a_12102_1103# a_11510_869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4762 a_30897_7022# a_31154_6832# a_29885_7203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4763 a_225_n5828# a_225_n5546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4764 a_24509_n4105# a_24707_n5337# a_24662_n5133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4765 a_27277_n4816# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4766 a_12283_6980# a_12070_6980# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4767 a_25713_n7932# a_25716_n7329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4768 vdd d0 a_31244_n8906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4769 a_24485_n8210# a_24699_n7294# a_24654_n7090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4770 a_16843_n9336# a_17648_n9570# a_17817_n9009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4771 a_7282_n3124# a_6861_n3124# a_7183_n2947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4772 a_36378_n7752# a_36631_n7956# a_35365_n7518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4773 a_25705_n8496# a_25717_n7744# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4774 a_34033_n6864# a_33661_n6621# a_33069_n6387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4775 a_5409_6335# a_5409_6053# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4776 a_40511_3855# a_40768_3665# a_40362_2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4777 vdd d0 a_31270_n3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4778 a_36273_8447# a_36276_7855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4779 a_32579_840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4780 a_25632_4906# a_25885_4893# a_24616_5264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4781 vdd d0 a_41830_3904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4782 vdd d0 a_41848_1378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4783 a_17559_7940# a_17346_7940# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4784 a_29916_2130# a_30974_2351# a_30929_2364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4785 a_7012_n4664# a_6799_n4664# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4786 a_38366_n3845# a_37945_n3845# a_37669_n3826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4787 a_25652_989# a_25648_1166# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4788 vdd a_20429_n5592# a_20221_n5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4789 a_1459_7392# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4790 a_135_5589# a_133_5375# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4791 a_629_2821# a_416_2821# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4792 a_40596_n7077# a_40691_n7701# a_40642_n7685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4793 gnd d3 a_40615_2637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4794 a_27692_n5382# a_28497_n5616# a_28666_n5055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4795 a_18750_n10389# a_18911_n6317# a_18862_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4796 a_14782_8061# a_14792_7318# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4797 a_21714_n6989# a_22195_n7360# a_22403_n7360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4798 vdd a_35314_6575# a_35106_6575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4799 a_13811_1207# a_14869_1428# a_14824_1441# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4800 gnd a_31258_n5555# a_31050_n5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4801 vdd a_15076_1013# a_14868_1013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4802 gnd d0 a_36561_1965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4803 a_8211_2671# a_8409_3686# a_8360_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4804 a_24697_n8489# a_25755_n8927# a_25710_n8723# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4805 a_21717_n5418# a_21722_n5032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4806 a_23397_n3116# a_23283_n3116# a_23491_n3116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4807 a_6772_1494# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4808 a_16159_n7772# a_16159_n7490# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4809 a_27697_n4401# a_27276_n4401# a_27010_n4215# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4810 a_8500_n6537# a_9558_n6975# a_9513_n6771# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4811 a_32286_5568# a_32767_5738# a_32975_5738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4812 vdd d4 a_29948_n6280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4813 a_16078_4386# a_16567_4204# a_16775_4204# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4814 gnd d0 a_31251_n7927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4815 a_32980_4757# a_32559_4757# a_32289_4592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4816 a_39124_3433# a_38911_3433# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4817 a_498_n6823# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4818 a_21729_n4236# a_22208_n4422# a_22416_n4422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4819 a_31011_n4785# a_31007_n4973# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4820 a_11065_6182# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4821 a_39145_n8048# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4822 a_24631_2328# a_25692_1957# a_25643_2147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4823 a_35264_8036# a_36322_8257# a_36277_8270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4824 vdd d0 a_4479_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4825 gnd d5 a_29836_n10368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4826 a_13833_n5170# a_14086_n5374# a_13680_n4142# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4827 a_1654_1095# a_1441_1095# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4828 gnd d2 a_30196_n5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4829 a_40338_6744# a_40552_5622# a_40507_5635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4830 a_16154_n8370# a_16161_n8169# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4831 vdd d0 a_25868_7834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4832 a_28281_n6592# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4833 gnd d2 a_35576_n5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4834 vdd a_3475_n5786# a_3267_n5786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4835 a_12454_5440# a_12082_5020# a_11491_5201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4836 a_29681_6559# a_29879_7574# a_29830_7764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4837 vdd a_36550_4340# a_36342_4340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4838 a_21626_4370# a_21626_4088# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4839 a_24298_n10373# a_24459_n6301# a_24414_n6097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4840 vdd a_40780_1705# a_40572_1705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4841 a_7181_3454# a_7138_2522# a_7322_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4842 vdd a_40815_5061# a_40607_5061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4843 a_24704_n7510# a_25762_n7948# a_25713_n7932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4844 a_12551_n4936# a_12442_n5113# a_12650_n5113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4845 a_40358_2827# a_40615_2637# a_40263_4819# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4846 a_1870_n8845# a_1498_n8602# a_906_n8368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4847 gnd d0 a_15071_1994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4848 a_19021_3884# a_19278_3694# a_18872_2679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4849 a_10885_n6431# a_10888_n6050# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4850 a_23288_5522# a_22906_5964# a_22315_6145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4851 gnd d0 a_31238_n9472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4852 a_7183_n2947# a_6811_n2704# a_6219_n2470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4853 a_26990_n8132# a_27469_n8318# a_27677_n8318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4854 a_12531_n8853# a_12159_n8610# a_11567_n8376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4855 a_9444_1412# a_9697_1399# a_8431_1178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4856 a_8376_1739# a_8629_1726# a_8207_2848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4857 a_11490_4786# a_11069_4786# a_10799_4621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4858 a_35289_3138# a_36347_3359# a_36298_3549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4859 a_41648_n8898# a_41905_n8914# a_40639_n8476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4860 vdd a_40892_n8680# a_40684_n8680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4861 a_16864_n5834# a_16443_n5834# a_16167_n5815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4862 a_16166_n7005# a_16647_n7376# a_16855_n7376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4863 a_22183_n9320# a_21970_n9320# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4864 a_39585_338# a_40312_4629# a_40267_4642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4865 a_17923_n7049# a_17502_n7049# a_17824_n6872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4866 vdd a_8736_n9682# a_8528_n9682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4867 vdd d1 a_8741_n8701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4868 a_4251_n2460# a_4504_n2664# a_3235_n2829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4869 a_16766_5746# a_16345_5746# a_16077_5576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4870 a_41659_n6523# a_41667_n5774# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4871 a_28651_7342# a_28608_6410# a_28816_6410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4872 a_32289_4592# a_32287_4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4873 a_37575_3590# a_38056_3760# a_38264_3760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4874 a_37651_n8140# a_37649_n7743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4875 gnd a_15133_n8549# a_14925_n8549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4876 a_28661_n4878# a_28552_n5055# a_28760_n5055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4877 a_16077_5576# a_16075_5362# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4878 a_35222_5833# a_35326_5082# a_35277_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4879 a_3239_n2641# a_3492_n2845# a_3180_n3390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4880 a_12077_6001# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4881 a_27015_n3051# a_27496_n3422# a_27704_n3422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4882 a_36285_6487# a_36542_6297# a_35276_6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4883 gnd d0 a_4404_3380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4884 a_22429_n2877# a_23233_n2696# a_23392_n2939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4885 vdd a_15060_4369# a_14852_4369# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4886 a_24688_n9658# a_25749_n9493# a_25700_n9477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4887 a_35353_n9478# a_36411_n9916# a_32358_n9938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4888 a_148_2157# a_150_2058# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4889 a_15660_n10477# a_18799_n10405# a_18750_n10389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4890 a_38353_n5390# a_37932_n5390# a_37664_n5019# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4891 a_16354_4204# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4892 a_2001_n3145# a_1946_n4173# a_2130_n5921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4893 a_13794_4148# a_14852_4369# a_14803_4559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4894 a_41675_n4002# a_41932_n4018# a_40666_n3580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4895 a_849_861# a_428_861# a_155_1077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4896 a_33580_3034# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4897 a_18957_n4309# a_19214_n4325# a_18862_n6301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4898 a_38345_n7347# a_37924_n7347# a_37656_n6976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4899 a_33869_n7602# a_33656_n7602# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4900 a_28641_n8795# a_28269_n8552# a_27677_n8318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4901 a_12174_n5674# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4902 a_428_861# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4903 gnd a_4411_2401# a_4203_2401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4904 a_22107_6145# a_21894_6145# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4905 a_5787_n4845# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4906 a_5523_n2584# a_5525_n2485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4907 gnd a_20345_2952# a_20137_2952# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4908 a_32383_n5040# a_32864_n5411# a_33072_n5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4909 a_10866_n9471# a_10868_n9372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4910 a_13736_5685# a_13831_6092# a_13782_6282# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4911 a_41659_n7731# a_41912_n7935# a_40646_n7497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4912 gnd a_8718_n3385# a_8510_n3385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4913 a_8516_n2808# a_8773_n2824# a_8461_n3369# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4914 a_12702_4476# a_12305_2551# a_12573_1523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4915 a_1424_4036# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4916 a_8211_2671# a_8409_3686# a_8364_3699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4917 a_9516_n5795# a_9769_n5999# a_8503_n5561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4918 a_32869_n4430# a_32656_n4430# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4919 a_26926_1027# a_26933_826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4920 a_32269_7914# a_32274_7528# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4921 a_24697_n8489# a_24950_n8693# a_24638_n9238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4922 gnd d1 a_30162_3096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4923 a_20073_7297# a_20069_7474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4924 gnd a_31167_5287# a_30959_5287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4925 a_4215_n8525# a_4472_n8541# a_3203_n8706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4926 gnd a_30099_5614# a_29891_5614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4927 gnd a_31276_n3029# a_31068_n3029# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4928 a_31994_256# a_37072_271# a_34403_359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4929 a_6829_n9001# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4930 gnd a_41916_n6539# a_41708_n6539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4931 a_23459_n8993# a_23038_n8993# a_23360_n8816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4932 a_116_8034# a_118_7935# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4933 a_37072_271# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4934 vdd a_9660_8257# a_9452_8257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4935 gnd a_9760_n7541# a_9552_n7541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4936 a_719_n4866# a_506_n4866# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4937 a_25635_3930# a_25888_3917# a_24619_4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4938 a_12090_3063# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4939 a_8089_n10381# a_8346_n10397# a_4999_n10469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4940 a_41557_7834# a_41553_8011# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4941 a_29606_4634# a_29859_4621# a_28924_330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4942 a_17490_n9009# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4943 a_32567_2800# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4944 a_12587_n8098# a_12374_n8098# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4945 a_29681_6559# a_29879_7574# a_29834_7587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4946 a_143_3037# a_629_2821# a_837_2821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4947 a_12702_4476# a_12593_4476# a_12801_4476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4948 a_5486_n9442# a_5975_n9743# a_6183_n9743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4949 gnd a_4488_n6020# a_4280_n6020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4950 a_19165_n4776# a_20226_n4611# a_20181_n4407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4951 vdd d0 a_36546_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4952 a_17366_4023# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4953 a_28502_n4635# a_28289_n4635# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4954 a_16095_1163# a_16097_1064# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4955 a_12367_n9591# a_12154_n9591# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4956 vdd a_8686_n9262# a_8478_n9262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4957 vdd a_3272_n4338# a_3064_n4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4958 a_16779_2808# a_16358_2808# a_16085_3024# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4959 a_21886_6709# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4960 a_23534_351# a_23321_351# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4961 a_21982_n7360# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4962 a_22200_n6379# a_21987_n6379# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4963 a_40647_n6704# a_40904_n6720# a_40592_n7265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4964 a_29994_n4739# a_31055_n4574# a_31006_n4558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4965 a_8399_7055# a_9457_7276# a_9408_7466# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4966 a_918_n6408# a_497_n6408# a_224_n6423# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4967 a_22969_3446# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4968 a_7042_n9001# a_6829_n9001# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4969 a_8503_n5561# a_9561_n5999# a_9516_n5795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4970 a_19094_n9066# a_19189_n9690# a_19140_n9674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4971 vdd d0 a_9696_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4972 a_8364_3699# a_8459_4106# a_8410_4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4973 a_27396_4167# a_27183_4167# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4974 a_6187_n8347# a_6992_n8581# a_7151_n8824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4975 a_33085_n3866# a_33889_n3685# a_34058_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4976 a_133_5093# a_135_4994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4977 a_37651_n8140# a_38130_n8326# a_38338_n8326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4978 a_5511_n4544# a_5513_n4445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4979 a_8372_1916# a_8629_1726# a_8207_2848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4980 a_28400_5943# a_28187_5943# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4981 a_12706_6468# a_12285_6468# a_12541_7400# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4982 a_39238_3552# a_39124_3433# a_39332_3433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4983 a_24616_5264# a_25677_4893# a_25632_4906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4984 a_16843_n9336# a_16422_n9336# a_16154_n8965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4985 a_14824_1441# a_15077_1428# a_13811_1207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4986 a_4246_n3441# a_4242_n3629# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4987 a_38370_n2449# a_37949_n2449# a_37676_n2464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4988 a_10504_285# a_15582_300# a_12913_388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4989 a_21995_n4422# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4990 a_20069_7474# a_20072_6882# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4991 a_10784_6962# a_11270_6746# a_11478_6746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4992 a_28812_4418# a_28703_4418# a_28911_4418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4993 gnd d3 a_40704_n4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4994 a_25700_n9477# a_25710_n8723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4995 a_6220_n2885# a_5799_n2885# a_5523_n2866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4996 a_15582_300# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4997 a_9512_n6356# a_9508_n6544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4998 a_27615_1792# a_28420_2026# a_28589_1584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4999 vdd d0 a_31161_5853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5000 a_35222_5833# a_35326_5082# a_35281_5095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5001 a_9503_n7525# a_9760_n7541# a_8491_n7706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5002 a_26904_5325# a_27393_5143# a_27601_5143# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5003 a_19149_n8505# a_19402_n8709# a_19090_n9254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5004 a_19172_n3797# a_20233_n3632# a_20184_n3616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5005 gnd d0 a_25880_5874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5006 a_39322_n4886# a_39213_n5063# a_39421_n5063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5007 vdd d0 a_4404_3380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5008 a_25721_n5975# a_25978_n5991# a_24712_n5553# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5009 vdd a_25969_n7533# a_25761_n7533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5010 vdd a_24965_n5757# a_24757_n5757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5011 a_41570_6289# a_41566_6466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5012 vdd d0 a_15056_4930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5013 a_12070_6980# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5014 a_4163_1433# a_4159_1610# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5015 a_14900_n4428# a_14896_n4616# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5016 a_5411_5954# a_5416_5568# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5017 a_27601_5143# a_28405_4962# a_28564_5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5018 a_3148_n9267# a_3252_n8722# a_3203_n8706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5019 a_34097_n4152# a_33884_n4152# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5020 gnd a_20414_n8528# a_20206_n8528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5021 a_21732_n2576# a_22221_n2877# a_22429_n2877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5022 gnd d0 a_15051_5911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5023 gnd a_41932_n4018# a_41724_n4018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5024 a_130_6570# a_609_6738# a_817_6738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5025 a_37642_n8722# a_37642_n8440# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5026 a_33078_n4845# a_32657_n4845# a_32381_n4544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5027 a_26921_2008# a_27407_1792# a_27615_1792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5028 vdd a_41848_1378# a_41640_1378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5029 a_7138_2522# a_6925_2522# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5030 a_37841_5151# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5031 vdd d0 a_25974_n6552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5032 a_22340_1247# a_21919_1247# a_21643_1147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5033 vdd a_35638_n3805# a_35430_n3805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5034 vdd d1 a_35643_n2824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5035 a_40582_1157# a_41640_1378# a_41591_1568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5036 a_38057_4175# a_37844_4175# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5037 a_416_2821# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5038 a_9424_5329# a_9677_5316# a_8411_5095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5039 a_17440_n8589# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5040 a_5910_2800# a_5697_2800# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5041 a_27616_2207# a_27195_2207# a_26919_2107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5042 a_1530_n2725# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5043 a_8426_2159# a_8679_2146# a_8376_1739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5044 a_29884_8007# a_30137_7994# a_29834_7587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5045 a_23276_7482# a_22894_7924# a_22302_7690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5046 a_14872_n9929# a_14875_n9326# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5047 a_29900_4267# a_30961_3896# a_30912_4086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5048 a_8429_n9246# a_8533_n8701# a_8488_n8497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5049 vdd a_30099_5614# a_29891_5614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5050 vdd d0 a_9671_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5051 a_13896_n2837# a_14153_n2853# a_13841_n3398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5052 a_32375_n6402# a_32861_n6387# a_33069_n6387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5053 gnd d0 a_41811_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5054 a_39213_7350# a_39104_7350# a_39312_7350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5055 gnd d4 a_8369_4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5056 vdd d0 a_4505_n3079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5057 gnd d0 a_9697_1399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5058 a_222_n6804# a_711_n6823# a_919_n6823# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5059 a_27501_n2441# a_27288_n2441# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5060 a_13795_3344# a_14856_2973# a_14807_3163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5061 a_29602_4811# a_29859_4621# a_28924_330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5062 a_37587_1630# a_37585_1416# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5063 a_25635_3930# a_25631_4107# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5064 a_11057_6746# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5065 a_25648_1166# a_25905_976# a_24636_1347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5066 a_37573_3376# a_37573_3094# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5067 a_26907_4067# a_26909_3968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5068 a_39453_n6056# a_39240_n6056# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5069 a_16439_n6395# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5070 a_14803_4943# a_14799_5120# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5071 a_19092_1186# a_19345_1173# a_19033_1924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5072 a_22196_n7775# a_21983_n7775# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5073 a_32287_4096# a_32289_3997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5074 a_12682_n6106# a_12469_n6106# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5075 vdd a_25868_7834# a_25660_7834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5076 a_38945_n5624# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5077 a_32651_n5411# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5078 a_1900_3475# a_1479_3475# a_1806_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5079 a_26832_263# a_31885_256# a_20996_141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5080 a_4159_1610# a_4162_1018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5081 a_27277_n4816# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5082 a_24620_5087# a_25678_5308# a_25629_5498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5083 a_32272_7314# a_32272_7032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5084 a_16070_6061# a_16559_6161# a_16767_6161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5085 a_33788_4015# a_33575_4015# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5086 a_32643_n7368# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5087 a_19092_1186# a_20150_1407# a_20101_1597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5088 a_21606_8005# a_21608_7906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5089 a_8399_7055# a_9457_7276# a_9412_7289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5090 gnd a_15146_n7004# a_14938_n7004# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5091 a_20174_n6779# a_20170_n6967# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5092 a_8445_n7098# a_8540_n7722# a_8491_n7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5093 a_23271_7363# a_22899_6943# a_22308_7124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5094 gnd a_13726_n10426# a_13518_n10426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5095 a_9439_1174# a_5443_855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5096 a_25648_1166# a_21652_847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5097 a_7012_n4664# a_6799_n4664# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5098 a_27400_2771# a_27187_2771# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5099 a_38366_n3845# a_37945_n3845# a_37669_n3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5100 gnd d1 a_30142_7013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5101 a_38277_2215# a_37856_2215# a_37580_2397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5102 a_16184_n2592# a_16673_n2893# a_16881_n2893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5103 a_7118_6439# a_6905_6439# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5104 a_27693_n5797# a_28497_n5616# a_28666_n5055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5105 a_37860_819# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5106 a_28557_7461# a_28175_7903# a_27584_8084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5107 a_24720_n3781# a_24977_n3797# a_24674_n3173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5108 a_25652_989# a_25905_976# a_24636_1347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5109 a_1723_n6642# a_1510_n6642# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5110 gnd d2 a_24927_n3377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5111 a_6098_6717# a_5677_6717# a_5411_6549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5112 a_33773_6951# a_33560_6951# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5113 a_41583_3351# a_41579_3528# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5114 gnd a_30149_6034# a_29941_6034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5115 a_39401_n8980# a_39358_n8048# a_39566_n8048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5116 a_32388_n3565# a_32877_n3866# a_33085_n3866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5117 a_8496_n6725# a_9557_n6560# a_9508_n6544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5118 a_32775_3781# a_32562_3781# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5119 vdd d1 a_14141_n4813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5120 a_9520_n4399# a_9773_n4603# a_8504_n4768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5121 vdd a_35588_n3385# a_35380_n3385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5122 a_849_861# a_1654_1095# a_1813_1515# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5123 a_33567_5972# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5124 vdd d0 a_36630_n7541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5125 gnd d0 a_25982_n4595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5126 a_34291_4447# a_33870_4447# a_34192_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5127 a_5518_n3565# a_5520_n3466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5128 a_22408_n6379# a_21987_n6379# a_21717_n6013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5129 a_5918_2236# a_5705_2236# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5130 a_32279_6335# a_32768_6153# a_32976_6153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5131 a_5762_n9743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5132 a_1617_7953# a_1404_7953# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5133 gnd d1 a_24970_n4776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5134 a_3227_n4601# a_4285_n5039# a_4236_n5023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5135 a_33944_n3124# a_33731_n3124# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5136 a_40541_8192# a_40798_8002# a_40495_7595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5137 a_21722_n4437# a_22208_n4422# a_22416_n4422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5138 a_4235_n4608# a_4247_n3856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5139 a_12298_4044# a_12085_4044# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5140 gnd a_4404_3380# a_4196_3380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5141 a_30933_968# a_31186_955# a_29917_1326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5142 a_921_n5432# a_500_n5432# a_227_n5447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5143 a_3059_7814# a_3163_7063# a_3114_7253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5144 a_22100_7124# a_21887_7124# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5145 a_9524_n4023# a_9527_n3420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5146 a_36277_7051# a_36534_6861# a_35265_7232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5147 gnd d2 a_3336_3707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5148 a_25636_4345# a_25632_4522# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5149 a_9516_n4587# a_9528_n3835# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5150 a_1786_7511# a_1672_7392# a_1880_7392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5151 vdd a_31250_n7512# a_31042_n7512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5152 vdd a_30246_n5736# a_30038_n5736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5153 a_2252_380# a_1831_380# a_2153_380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5154 a_14824_1441# a_14820_1618# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5155 a_6779_n8581# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5156 a_9420_5506# a_9677_5316# a_8411_5095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5157 a_37917_n8326# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5158 vdd a_36644_n5018# a_36436_n5018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5159 a_33676_n3685# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5160 a_8344_7616# a_8439_8023# a_8390_8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5161 gnd a_3391_3146# a_3183_3146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5162 a_21631_3389# a_22120_3207# a_22328_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5163 a_40342_6567# a_40595_6554# a_40267_4642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5164 a_22319_4749# a_23124_4983# a_23283_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5165 a_16584_1263# a_16371_1263# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5166 a_41583_3351# a_41836_3338# a_40570_3117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5167 a_22397_n8754# a_21976_n8754# a_21700_n8735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5168 a_8422_2336# a_8679_2146# a_8376_1739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5169 a_12283_6980# a_12070_6980# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5170 a_14908_n2656# a_15842_n2260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5171 a_7099_1613# a_6985_1494# a_7193_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5172 a_4121_8053# a_4378_7863# a_3109_8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5173 a_35234_3699# a_35329_4106# a_35284_4119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5174 a_10900_n3495# a_11386_n3480# a_11594_n3480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5175 a_39250_1592# a_38868_2034# a_38276_1800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5176 a_34051_3454# a_33630_3454# a_33952_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5177 a_14787_8299# a_16058_8303# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5178 gnd a_36624_n8935# a_36416_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5179 a_35349_n9666# a_35606_n9682# a_35303_n9058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5180 vdd d0 a_41811_8236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5181 vdd d4 a_8369_4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5182 vdd d1 a_40924_n2803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5183 a_17559_7940# a_17346_7940# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5184 a_41579_3528# a_41582_2936# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5185 gnd a_30162_3096# a_29954_3096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5186 a_13571_6617# a_13824_6604# a_13496_4692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5187 a_40562_5074# a_40815_5061# a_40503_5812# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5188 a_1622_6972# a_1409_6972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5189 a_7262_n7041# a_6841_n7041# a_7168_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5190 a_41651_n8295# a_41904_n8499# a_40635_n8664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5191 a_13821_n7315# a_14078_n7331# a_13656_n8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5192 a_5488_n9343# a_5493_n8957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5193 a_9434_2155# a_9691_1965# a_8422_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5194 vdd d0 a_4384_7297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5195 a_37662_n4523# a_38151_n4824# a_38359_n4824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5196 vdd d2 a_35568_n7302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5197 a_40639_n8476# a_40892_n8680# a_40580_n9225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5198 a_32995_1821# a_32574_1821# a_32306_1651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5199 a_35280_4296# a_36341_3925# a_36296_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5200 a_16864_n5834# a_16443_n5834# a_16167_n5533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5201 a_19001_7801# a_19105_7050# a_19056_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5202 gnd d0 a_15165_n2672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5203 a_16161_n7391# a_16647_n7376# a_16855_n7376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5204 a_28552_n5055# a_28339_n5055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5205 vdd d1 a_3386_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5206 a_6898_7932# a_6685_7932# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5207 vdd d1 a_19429_n3813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5208 a_34982_4840# a_35126_2658# a_35077_2848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5209 a_6111_5172# a_5690_5172# a_5414_5354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5210 a_25721_n6348# a_25717_n6536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5211 a_19088_1363# a_19345_1173# a_19033_1924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5212 a_31003_n6742# a_30999_n6930# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5213 a_11575_n7812# a_11154_n7812# a_10878_n7793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5214 a_22008_n2877# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5215 a_38856_3994# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5216 a_21727_n3557# a_21729_n3458# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5217 a_10886_n5554# a_11375_n5855# a_11583_n5855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5218 a_6011_n2470# a_5798_n2470# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5219 a_37568_4357# a_38057_4175# a_38265_4175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5220 a_19156_n7526# a_19409_n7730# a_19106_n7106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5221 a_8515_n3601# a_9573_n4039# a_9524_n4023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5222 a_27010_n3437# a_27496_n3422# a_27704_n3422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5223 a_12479_1642# a_12097_2084# a_11506_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5224 a_24705_n6717# a_25766_n6552# a_25721_n6348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5225 a_35331_n3369# a_35435_n2824# a_35390_n2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5226 a_23372_n6856# a_23263_n7033# a_23471_n7033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5227 gnd a_19417_n5773# a_19209_n5773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5228 vdd a_36546_4901# a_36338_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5229 gnd d5 a_40497_n10376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5230 a_29885_7203# a_30946_6832# a_30901_6845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5231 a_20093_3380# a_20346_3367# a_19080_3146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5232 a_25725_n4579# a_25982_n4595# a_24713_n4760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5233 a_16174_n4453# a_16660_n4438# a_16868_n4438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5234 a_32292_3115# a_32781_3215# a_32989_3215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5235 a_21902_4188# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5236 a_14820_1618# a_14823_1026# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5237 a_33869_n7602# a_33656_n7602# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5238 a_12174_n5674# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5239 vdd d1 a_30142_7013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5240 gnd a_13749_4679# a_13541_4679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5241 a_40527_1718# a_40622_2125# a_40573_2315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5242 a_25633_5321# a_25629_5498# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5243 a_38049_6132# a_37836_6132# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5244 a_830_5193# a_409_5193# a_133_5093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5245 gnd d0 a_41815_6840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5246 a_11587_n4459# a_12392_n4693# a_12551_n4936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5247 a_29880_8184# a_30941_7813# a_30892_8003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5248 a_22319_4749# a_21898_4749# a_21628_4584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5249 a_32378_n5426# a_32864_n5411# a_33072_n5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5250 a_5994_n5411# a_5781_n5411# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5251 vdd a_4390_5903# a_4182_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5252 vdd a_30149_6034# a_29941_6034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5253 a_27183_4167# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5254 a_16169_n6029# a_16167_n5815# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5255 a_1733_n4173# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5256 a_16564_5180# a_16351_5180# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5257 gnd a_20427_n6983# a_20219_n6983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5258 a_27685_n7754# a_27264_n7754# a_26988_n7735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5259 a_9529_n3042# a_9786_n3058# a_8520_n2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5260 vdd d0 a_9753_n8520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5261 vdd d0 a_25995_n3050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5262 a_26996_n5496# a_27485_n5797# a_27693_n5797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5263 a_11505_1850# a_11084_1850# a_10816_1680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5264 vdd d0 a_20325_6869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5265 a_10797_4125# a_11286_4225# a_11494_4225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5266 a_29985_n7489# a_30238_n7693# a_29935_n7069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5267 a_12392_n4693# a_12179_n4693# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5268 a_1793_5432# a_1421_5012# a_830_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5269 gnd a_36638_n5584# a_36430_n5584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5270 gnd d0 a_36643_n4603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5271 a_25710_n8723# a_25963_n8927# a_24697_n8489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5272 a_38351_n6781# a_39155_n6600# a_39314_n6843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5273 gnd d0 a_20320_7850# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5274 a_33053_n9743# a_32632_n9743# a_32356_n9724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5275 a_17735_n3132# a_17522_n3132# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5276 a_21697_n9335# a_21702_n8949# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5277 a_8499_n5749# a_8756_n5765# a_8453_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5278 gnd d2 a_8706_n5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5279 a_32975_5738# a_32554_5738# a_32281_5954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5280 vdd a_4404_3380# a_4196_3380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5281 vdd d4 a_35328_n6309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5282 a_1880_7392# a_1459_7392# a_1786_7511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5283 a_3059_7814# a_3163_7063# a_3118_7076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5284 a_35299_n9246# a_35556_n9262# a_35150_n8030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5285 a_20105_1420# a_20101_1597# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5286 a_19072_5103# a_20130_5324# a_20081_5514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5287 vdd a_15056_4930# a_14848_4930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5288 a_14900_n4428# a_15153_n4632# a_13884_n4797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5289 a_719_n4866# a_506_n4866# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5290 a_30991_n8702# a_30987_n8890# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5291 gnd d1 a_30251_n4755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5292 gnd d1 a_19397_n9690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5293 a_8344_7616# a_8439_8023# a_8394_8036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5294 a_7161_7371# a_7118_6439# a_7326_6439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5295 gnd a_35623_n6741# a_35415_n6741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5296 a_844_1842# a_423_1842# a_150_2058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5297 a_1912_1515# a_1857_2543# a_2041_4468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5298 a_10791_6578# a_10789_6364# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5299 vdd a_3391_3146# a_3183_3146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5300 a_5486_n9724# a_5975_n9743# a_6183_n9743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5301 a_7161_7371# a_6740_7371# a_7062_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5302 a_40338_6744# a_40595_6554# a_40267_4642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5303 a_1580_n3145# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5304 a_13581_n6322# a_13838_n6338# a_13469_n10410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5305 a_28502_n4635# a_28289_n4635# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5306 gnd d0 a_9760_n7541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5307 a_32989_3215# a_33793_3034# a_33952_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5308 a_22914_4007# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5309 a_24505_n4293# a_24719_n3377# a_24670_n3361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5310 a_8419_3138# a_8672_3125# a_8360_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5311 a_25629_5498# a_25632_4906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5312 gnd d0 a_31175_3330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5313 a_23213_n6613# a_23000_n6613# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5314 gnd a_41905_n8914# a_41697_n8914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5315 a_32664_n3866# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5316 a_36383_n6771# a_36379_n6959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5317 a_8390_8213# a_9451_7842# a_9406_7855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5318 a_33823_7371# a_33610_7371# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5319 a_40558_5251# a_40815_5061# a_40503_5812# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5320 gnd a_9749_n9916# a_9541_n9916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5321 a_13829_n5358# a_13933_n4813# a_13888_n4609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5322 a_8116_4663# a_8236_6575# a_8187_6765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5323 a_35361_n7706# a_36422_n7541# a_36377_n7337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5324 gnd a_19367_n5353# a_19159_n5353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5325 a_12531_n8853# a_12159_n8610# a_11568_n8791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5326 a_37644_n8341# a_38130_n8326# a_38338_n8326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5327 a_29935_n7069# a_30030_n7693# a_29985_n7489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5328 a_10498_n10484# a_10448_n10500# a_10399_n10484# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5329 a_7019_n3685# a_6806_n3685# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5330 a_3214_n7539# a_4272_n7977# a_4227_n7773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5331 vdd a_9696_984# a_9488_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5332 a_19001_7801# a_19105_7050# a_19060_7063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5333 a_24658_n5321# a_24762_n4776# a_24713_n4760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5334 a_4146_4374# a_4142_4551# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5335 vdd a_9679_3925# a_9471_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5336 a_11494_4225# a_12298_4044# a_12467_3602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5337 a_27252_n9714# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5338 a_41671_n4378# a_41667_n4566# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5339 a_21995_n4422# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5340 a_11485_5767# a_11064_5767# a_10791_5983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5341 a_22183_n9320# a_21970_n9320# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5342 a_23382_5403# a_23327_6431# a_23535_6431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5343 a_39213_n5063# a_39000_n5063# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5344 a_1890_n4928# a_1781_n5105# a_1989_n5105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5345 a_17680_n3693# a_17467_n3693# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5346 a_29691_n6264# a_29948_n6280# a_29579_n10352# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5347 a_1907_n3145# a_1525_n3706# a_934_n3887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5348 a_5402_7032# a_5891_7132# a_6099_7132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5349 a_4220_n8752# a_4216_n8940# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5350 a_32390_n4244# a_32388_n3847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5351 gnd d2 a_3316_7624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5352 a_20848_n805# a_20739_n805# vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5353 a_29986_n6696# a_31047_n6531# a_31002_n6327# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5354 a_32381_n4544# a_32383_n4445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5355 a_5098_n10469# a_5048_n10485# a_4999_n10469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5356 a_3126_5293# a_3383_5103# a_3071_5854# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5357 a_20101_1597# a_20104_1005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5358 vdd d0 a_31181_1936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5359 a_40562_5074# a_41620_5295# a_41575_5308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5360 gnd d0 a_20446_n2651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5361 a_3138_3159# a_4196_3380# a_4147_3570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5362 a_29935_n7069# a_30188_n7273# a_29766_n8189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5363 a_28269_n8552# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5364 a_27412_811# a_27199_811# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5365 vdd d3 a_3183_2679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5366 a_27001_n4797# a_27001_n4515# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5367 a_6203_n5826# a_5782_n5826# a_5506_n5807# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5368 a_40527_1718# a_40622_2125# a_40577_2138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5369 a_33575_4015# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5370 a_1773_n7062# a_1560_n7062# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5371 a_13845_n3210# a_13940_n3834# a_13891_n3818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5372 a_25733_n4015# a_25736_n3412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5373 a_17773_367# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5374 a_38270_3194# a_37849_3194# a_37573_3376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5375 a_7079_5530# a_6965_5411# a_7173_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5376 gnd a_19214_n4325# a_19006_n4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5377 a_21727_n3839# a_21727_n3557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5378 a_21732_n2858# a_22221_n2877# a_22429_n2877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5379 a_11391_n2499# a_11178_n2499# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5380 a_27672_n9299# a_27251_n9299# a_26983_n8928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5381 a_29854_3670# a_29949_4077# a_29900_4267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5382 a_39319_n7020# a_38937_n7581# a_38346_n7762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5383 a_3198_n9687# a_4259_n9522# a_4214_n9318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5384 a_121_7335# a_610_7153# a_818_7153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5385 a_40612_n3348# a_40716_n2803# a_40671_n2599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5386 a_934_n3887# a_513_n3887# a_237_n3868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5387 a_27392_4728# a_27179_4728# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5388 a_32857_n7783# a_32644_n7783# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5389 gnd a_30142_7013# a_29934_7013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5390 a_38346_n7762# a_37925_n7762# a_37649_n7743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5391 vdd a_36651_n4039# a_36443_n4039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5392 vdd d0 a_36656_n3058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5393 gnd a_8773_n2824# a_8565_n2824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5394 a_38269_2779# a_37848_2779# a_37575_2995# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5395 a_34043_5411# a_33622_5411# a_33944_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5396 a_32869_n4430# a_32656_n4430# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5397 gnd d2 a_19347_n9270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5398 a_5503_n6501# a_5505_n6402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5399 a_37861_1234# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5400 a_6114_4196# a_5693_4196# a_5417_4378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5401 a_28475_1465# a_28262_1465# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5402 a_33560_6951# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5403 a_20184_n3616# a_20441_n3632# a_19172_n3797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5404 a_13896_n2837# a_14957_n2672# a_14908_n2656# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5405 a_1530_n2725# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5406 a_18866_n6113# a_19119_n6317# a_18750_n10389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5407 a_5911_3215# a_5698_3215# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5408 a_3141_2357# a_4202_1986# a_4157_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5409 a_4142_4551# a_4145_3959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5410 a_39401_n8980# a_38980_n8980# a_39307_n8980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5411 a_19068_5280# a_19325_5090# a_19013_5841# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5412 a_32562_3781# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5413 a_31017_n3391# a_31270_n3595# a_30001_n3760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5414 a_10804_3640# a_10802_3426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5415 a_11380_n4874# a_11167_n4874# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5416 a_16179_n3855# a_16179_n3573# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5417 vdd d1 a_35626_n5765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5418 vdd d0 a_9691_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5419 a_21631_3107# a_21633_3008# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5420 a_32547_6717# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5421 a_12791_n5929# a_12394_n4181# a_12650_n5113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5422 a_19072_5103# a_20130_5324# a_20085_5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5423 a_27501_n2441# a_27288_n2441# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5424 a_5705_2236# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5425 vdd d0 a_36541_5882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5426 a_3203_n8706# a_3460_n8722# a_3148_n9267# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5427 a_1404_7953# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5428 gnd a_3405_n9283# a_3197_n9283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5429 a_19110_n5337# a_19214_n4792# a_19165_n4776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5430 a_17646_1502# a_17433_1502# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5431 gnd a_36656_n3058# a_36448_n3058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5432 gnd d0 a_41924_n4582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5433 a_16652_n6395# a_16439_n6395# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5434 gnd d0 a_20435_n5026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5435 a_833_4217# a_412_4217# a_136_4117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5436 a_12085_4044# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5437 a_128_6356# a_128_6074# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5438 a_153_1176# a_642_1276# a_850_1276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5439 a_11058_7161# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5440 gnd a_3336_3707# a_3128_3707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5441 a_24640_1170# a_24893_1157# a_24581_1908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5442 a_32651_n5411# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5443 a_38945_n5624# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5444 a_8415_3315# a_8672_3125# a_8360_3876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5445 a_40580_n9225# a_40837_n9241# a_40431_n8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5446 a_16174_n4453# a_16181_n4252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5447 a_20996_141# a_20887_141# a_20853_n686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5448 vdd d0 a_31175_3330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5449 gnd d3 a_19194_n8242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5450 a_24611_6245# a_25672_5874# a_25627_5887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5451 a_34380_n6077# a_33959_n6077# a_34285_n8069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5452 a_14819_2422# a_15072_2409# a_13806_2188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5453 a_39233_3433# a_38861_3013# a_38269_2779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5454 a_38053_4736# a_37840_4736# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5455 a_23223_n4144# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5456 a_16371_1263# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5457 a_8116_4663# a_8236_6575# a_8191_6588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5458 a_12070_6980# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5459 vdd a_25994_n2635# a_25786_n2635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5460 a_21638_2410# a_21638_2128# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5461 a_32294_3611# a_32775_3781# a_32983_3781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5462 vdd d0 a_15141_n7985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5463 vdd a_15149_n6028# a_14941_n6028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5464 vdd d5 a_8346_n10397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5465 a_35374_n4768# a_36435_n4603# a_36386_n4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5466 gnd d0 a_41848_1378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5467 a_12662_n3153# a_12241_n3153# a_12568_n3153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5468 a_20084_4922# a_20080_5099# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5469 a_501_n5847# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5470 a_7087_3573# a_6705_4015# a_6113_3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5471 a_1723_n6642# a_1510_n6642# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5472 a_10905_n2514# a_10462_n2231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5473 a_37930_n6781# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5474 gnd a_25978_n5991# a_25770_n5991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5475 gnd d0 a_4493_n5039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5476 a_397_7153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5477 a_5488_n9938# a_9492_n9900# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5478 a_22404_n7775# a_23208_n7594# a_23377_n7033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5479 a_1831_380# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5480 a_21613_7520# a_22094_7690# a_22302_7690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5481 a_21623_5064# a_22112_5164# a_22320_5164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5482 a_32388_n3847# a_32877_n3866# a_33085_n3866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5483 a_13811_1207# a_14869_1428# a_14820_1618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5484 gnd a_15129_n9945# a_14921_n9945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5485 a_21712_n6493# a_21714_n6394# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5486 a_6007_n3866# a_5794_n3866# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5487 vdd d2 a_3316_7624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5488 a_16844_n9751# a_16423_n9751# a_16147_n9732# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5489 a_20156_n9305# a_20409_n9509# a_19140_n9674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5490 vdd d0 a_15154_n5047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5491 a_6685_7932# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5492 gnd d3 a_30023_n8205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5493 a_28532_n8972# a_28319_n8972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5494 a_23298_n6069# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5495 a_3138_3159# a_4196_3380# a_4151_3393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5496 a_14888_n7781# a_14884_n7969# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5497 a_5762_n9743# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5498 gnd d0 a_20353_2388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5499 a_2930_2692# a_3128_3707# a_3083_3720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5500 a_4231_n6377# a_4484_n6581# a_3215_n6746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5501 a_16097_1659# a_16578_1829# a_16786_1829# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5502 a_41679_n2606# a_41558_8249# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5503 a_39289_2501# a_39076_2501# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5504 a_705_n7389# a_492_n7389# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5505 a_23070_n3116# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5506 a_30913_4885# a_30909_5062# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5507 a_32301_2632# a_32299_2418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5508 a_9419_6310# a_9672_6297# a_8406_6076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5509 a_616_5759# a_403_5759# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5510 a_921_n5432# a_500_n5432# a_232_n5061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5511 a_28772_n3095# a_28351_n3095# a_28678_n3095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5512 a_38042_7111# a_37829_7111# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5513 a_35264_8036# a_36322_8257# a_36273_8447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5514 vdd a_30142_7013# a_29934_7013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5515 a_28608_6410# a_28395_6410# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5516 a_23416_n8061# a_23203_n8061# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5517 a_37917_n8326# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5518 a_22335_2228# a_21914_2228# a_21638_2410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5519 gnd a_41815_6840# a_41607_6840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5520 a_37836_6132# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5521 a_39213_7350# a_38841_6930# a_38250_7111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5522 a_22397_n8754# a_21976_n8754# a_21700_n8453# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5523 a_41573_4094# a_41830_3904# a_40561_4275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5524 a_10886_n5554# a_10888_n5455# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5525 a_41591_1568# a_41848_1378# a_40582_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5526 gnd d1 a_35522_7042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5527 a_16351_5180# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5528 a_4228_n6980# a_4231_n6377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5529 a_17842_3462# a_17421_3462# a_17743_3462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5530 vdd d1 a_24962_n6733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5531 a_20173_n5991# a_20176_n5388# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5532 a_40362_2650# a_40615_2637# a_40263_4819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5533 a_1568_n5105# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5534 a_694_n9764# a_481_n9764# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5535 vdd a_20325_6869# a_20117_6869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5536 gnd d0 a_25958_n9908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5537 vdd a_14121_n8730# a_13913_n8730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5538 a_39562_n5879# a_39165_n4131# a_39433_n3103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5539 gnd a_35529_6063# a_35321_6063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5540 a_32792_840# a_32579_840# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5541 a_141_3418# a_141_3136# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5542 vdd d0 a_41937_n3037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5543 a_5419_3997# a_5424_3611# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5544 a_19140_n9674# a_20201_n9509# a_20156_n9305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5545 a_37944_n3430# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5546 gnd a_24950_n8693# a_24742_n8693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5547 a_37662_n4805# a_38151_n4824# a_38359_n4824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5548 gnd d1 a_3366_8044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5549 a_20085_5337# a_20081_5514# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5550 a_12221_n7070# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5551 gnd a_8346_n10397# a_8138_n10397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5552 a_22424_n3858# a_22003_n3858# a_21727_n3557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5553 a_24549_7785# a_24653_7034# a_24604_7224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5554 a_25616_8262# a_25612_8439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5555 a_29969_n9637# a_31030_n9472# a_30981_n9456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5556 a_16856_n7791# a_17660_n7610# a_17829_n7049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5557 a_32373_n6501# a_32862_n6802# a_33070_n6802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5558 a_39585_338# a_40312_4629# a_40263_4819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5559 a_7227_n4152# a_7014_n4152# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5560 a_24636_1347# a_25697_976# a_25652_989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5561 a_23276_7482# a_23162_7363# a_23370_7363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5562 a_11575_n7812# a_11154_n7812# a_10878_n7511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5563 a_22008_n2877# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5564 a_23263_n7033# a_23050_n7033# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5565 vdd d1 a_40907_n5744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5566 a_10886_n5836# a_11375_n5855# a_11583_n5855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5567 a_36313_997# a_36566_984# a_35297_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5568 a_32358_n9343# a_32363_n8957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5569 a_16346_6161# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5570 gnd a_24977_n3797# a_24769_n3797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5571 gnd a_15060_4369# a_14852_4369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5572 a_35390_n2620# a_36448_n3058# a_36403_n2854# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5573 a_28589_1584# a_28475_1465# a_28683_1465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5574 a_6093_7698# a_5672_7698# a_5404_7528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5575 a_25611_8024# a_25868_7834# a_24599_8205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5576 a_20083_4123# a_20340_3933# a_19071_4304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5577 a_39307_n8980# a_39193_n8980# a_39401_n8980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5578 a_12447_7519# a_12333_7400# a_12541_7400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5579 gnd d1 a_14032_7071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5580 gnd a_14128_n7751# a_13920_n7751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5581 a_28455_5382# a_28242_5382# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5582 gnd a_31175_3330# a_30967_3330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5583 a_32793_1255# a_32580_1255# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5584 a_9528_n3835# a_9524_n4023# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5585 a_22209_n4837# a_21996_n4837# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5586 a_23308_1605# a_22926_2047# a_22334_1813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5587 a_33610_7371# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5588 a_5994_n5411# a_5781_n5411# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5589 gnd d1 a_19308_8031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5590 gnd a_14039_6092# a_13831_6092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5591 a_517_n2491# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5592 a_27685_n7754# a_27264_n7754# a_26988_n7453# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5593 vdd d0 a_31271_n4010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5594 a_850_1276# a_429_1276# a_153_1176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5595 a_35323_n5141# a_35418_n5765# a_35373_n5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5596 a_32861_n6387# a_32648_n6387# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5597 gnd a_8458_n6309# a_8250_n6309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5598 a_17822_7379# a_17401_7379# a_17728_7498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5599 a_22906_5964# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5600 vdd d0 a_20422_n7964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5601 vdd a_20430_n6007# a_20222_n6007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5602 a_7074_n3124# a_6861_n3124# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5603 a_27601_5143# a_27180_5143# a_26904_5325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5604 a_40655_n4747# a_41716_n4582# a_41667_n4566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5605 a_16754_7706# a_16333_7706# a_16060_7922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5606 gnd a_24895_n9254# a_24687_n9254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5607 vdd a_36655_n2643# a_36447_n2643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5608 vdd a_30263_n2795# a_30055_n2795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5609 vdd a_19409_n7730# a_19201_n7730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5610 a_4141_4136# a_4151_3393# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5611 a_21707_n7474# a_22196_n7775# a_22404_n7775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5612 a_20081_5514# a_20084_4922# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5613 a_9532_n2439# a_9528_n2627# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5614 gnd a_31259_n5970# a_31051_n5970# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5615 gnd a_4384_7297# a_4176_7297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5616 a_33053_n9743# a_32632_n9743# a_32356_n9442# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5617 a_29691_n6264# a_29835_n4288# a_29786_n4272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5618 a_1813_1515# a_1441_1095# a_850_1276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5619 gnd a_3316_7624# a_3108_7624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5620 a_25612_8439# a_25615_7847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5621 a_16186_n3088# a_16184_n2874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5622 gnd a_20410_n9924# a_20202_n9924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5623 a_21626_4370# a_22115_4188# a_22323_4188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5624 a_32976_6153# a_32555_6153# a_32279_6053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5625 a_14799_6339# a_15052_6326# a_13786_6105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5626 gnd a_9660_8257# a_9452_8257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5627 vdd d6 a_15917_n10493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5628 a_3210_n7727# a_3467_n7743# a_3164_n7119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5629 a_39240_n6056# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5630 a_22095_8105# a_21882_8105# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5631 a_24724_n3593# a_25782_n4031# a_25737_n3827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5632 a_39245_1473# a_39136_1473# a_39344_1473# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5633 vdd d1 a_19414_n6749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5634 a_31002_n5954# a_31005_n5351# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5635 a_29917_1326# a_30978_955# a_30929_1145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5636 a_32358_n9938# a_36619_n9916# a_35353_n9478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5637 a_13875_n7547# a_14933_n7985# a_14888_n7781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5638 a_40578_1334# a_41639_963# a_41594_976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5639 a_5411_5954# a_5897_5738# a_6105_5738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5640 vdd d0 a_4480_n7977# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5641 a_155_1672# a_636_1842# a_844_1842# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5642 a_5709_840# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5643 vdd d1 a_35522_7042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5644 a_9495_n9297# a_9491_n9485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5645 a_17522_n3132# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5646 a_37662_n4805# a_37662_n4523# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5647 vdd d0 a_4379_8278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5648 a_16579_2244# a_16366_2244# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5649 a_33805_1074# a_33592_1074# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5650 a_22995_n7594# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5651 a_23213_n6613# a_23000_n6613# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5652 a_9521_n4814# a_9774_n5018# a_8508_n4580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5653 a_32664_n3866# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5654 a_36394_n4023# a_36397_n3420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5655 vdd d2 a_8698_n7302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5656 vdd a_9766_n6975# a_9558_n6975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5657 a_5411_6549# a_5409_6335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5658 vdd a_35529_6063# a_35321_6063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5659 a_12159_n8610# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5660 a_27497_n3837# a_27284_n3837# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5661 a_28262_1465# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5662 vdd a_25900_1957# a_25692_1957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5663 vdd d0 a_41900_n9895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5664 a_13888_n4609# a_14946_n5047# a_14901_n4843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5665 gnd d0 a_20357_992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5666 a_14888_n6573# a_15145_n6589# a_13876_n6754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5667 a_641_861# a_428_861# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5668 a_11147_n8791# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5669 vdd d1 a_3366_8044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5670 vdd a_24653_6567# a_24445_6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5671 a_3118_7076# a_4176_7297# a_4131_7310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5672 vdd a_15153_n4632# a_14945_n4632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5673 a_39332_3433# a_39289_2501# a_39473_4426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5674 a_17735_5419# a_17626_5419# a_17834_5419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5675 a_24549_7785# a_24653_7034# a_24608_7047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5676 gnd a_14078_n7331# a_13870_n7331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5677 a_12593_4476# a_12380_4476# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5678 vdd d1 a_30243_n6712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5679 a_1649_2076# a_1436_2076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5680 a_9423_4914# a_9676_4901# a_8407_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5681 a_27252_n9714# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5682 a_39334_n2926# a_38962_n2683# a_38370_n2449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5683 a_11486_6182# a_11065_6182# a_10789_6082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5684 a_3083_3720# a_3178_4127# a_3133_4140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5685 gnd d0 a_9749_n9916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5686 a_32882_n2885# a_32669_n2885# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5687 a_35265_7232# a_36326_6861# a_36277_7051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5688 gnd a_25982_n4595# a_25774_n4595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5689 a_1907_n3145# a_1525_n3706# a_933_n3472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5690 a_26981_n8432# a_27470_n8733# a_27678_n8733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5691 a_17433_1502# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5692 a_39230_5509# a_38848_5951# a_38256_5717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5693 a_10804_3045# a_10811_2661# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5694 a_29834_7587# a_29929_7994# a_29884_8007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5695 a_23402_1486# a_23347_2514# a_23531_4439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5696 a_28651_7342# a_28230_7342# a_28552_7342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5697 a_35170_n4113# a_35368_n5345# a_35323_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5698 a_6011_n2470# a_5798_n2470# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5699 a_33089_n2470# a_33894_n2704# a_34053_n2947# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5700 a_5903_5172# a_5690_5172# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5701 gnd a_30231_n8672# a_30023_n8672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5702 gnd d3 a_3163_6596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5703 a_16159_n7490# a_16648_n7791# a_16856_n7791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5704 vdd a_24667_n6301# a_24459_n6301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5705 gnd a_15161_n4068# a_14953_n4068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5706 a_37585_1416# a_37585_1134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5707 a_28269_n8552# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5708 vdd d1 a_3455_n9703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5709 vdd d1 a_14032_7071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5710 vdd a_19359_n7310# a_19151_n7310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5711 a_16181_n4252# a_16660_n4438# a_16868_n4438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5712 a_35390_n2620# a_35643_n2824# a_35331_n3369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5713 a_21707_n7474# a_21709_n7375# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5714 a_6203_n5826# a_5782_n5826# a_5506_n5525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5715 vdd a_31175_3330# a_30967_3330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5716 a_13770_8242# a_14831_7871# a_14782_8061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5717 a_24654_n7090# a_24907_n7294# a_24485_n8210# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5718 a_24650_n7278# a_24754_n6733# a_24709_n6529# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5719 a_29606_4634# a_29726_6546# a_29677_6736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5720 a_20182_n4822# a_20178_n5010# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5721 a_32989_3215# a_32568_3215# a_32292_3397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5722 gnd d1 a_3383_5103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5723 vdd d1 a_19308_8031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5724 a_825_6174# a_404_6174# a_128_6356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5725 gnd d0 a_9786_n3058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5726 a_17931_n5092# a_17510_n5092# a_17837_n5092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5727 a_28420_2026# a_28207_2026# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5728 a_225_n5546# a_714_n5847# a_922_n5847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5729 a_8422_2336# a_9483_1965# a_9434_2155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5730 a_40671_n2599# a_41729_n3037# a_41684_n2833# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5731 gnd a_41848_1378# a_41640_1378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5732 a_12353_3483# a_12140_3483# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5733 gnd a_15917_n10493# a_15709_n10493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5734 a_38346_n7762# a_37925_n7762# a_37649_n7461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5735 a_19067_6084# a_19320_6071# a_19017_5664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5736 a_17842_3462# a_17799_2530# a_17983_4455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5737 vdd a_41936_n2622# a_41728_n2622# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5738 a_5431_2632# a_5910_2800# a_6118_2800# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5739 vdd a_9780_n3624# a_9572_n3624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5740 a_26892_7003# a_27381_7103# a_27589_7103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5741 a_36382_n5983# a_36385_n5380# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5742 vdd a_30196_n5316# a_29988_n5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5743 a_1560_n7062# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5744 gnd a_31169_3896# a_30961_3896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5745 gnd d2 a_3437_n3406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5746 gnd d3 a_19105_6583# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5747 vdd a_3316_7624# a_3108_7624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5748 a_16435_n7791# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5749 a_230_n4847# a_230_n4565# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5750 a_926_n4451# a_1731_n4685# a_1890_n4928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5751 a_11380_n4874# a_11167_n4874# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5752 a_39324_5390# a_39269_6418# a_39477_6418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5753 a_24628_3130# a_25686_3351# a_25637_3541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5754 gnd d0 a_25962_n8512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5755 a_16149_n9946# a_20153_n9908# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5756 a_14795_6516# a_15052_6326# a_13786_6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5757 gnd a_13838_n6338# a_13630_n6338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5758 gnd a_20353_2388# a_20145_2388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5759 a_29974_n8656# a_30231_n8672# a_29919_n9217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5760 a_32373_n6501# a_32375_n6402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5761 a_7079_5530# a_6697_5972# a_6106_6153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5762 a_4216_n8940# a_4473_n8956# a_3207_n8518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5763 a_23479_n5076# a_23436_n4144# a_23620_n5892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5764 a_39076_2501# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5765 a_403_5759# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5766 a_9435_2570# a_9438_1978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5767 a_26914_3582# a_27395_3752# a_27603_3752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5768 vdd d0 a_41828_5295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5769 a_11499_3244# a_11078_3244# a_10802_3426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5770 a_12814_388# a_12705_388# a_12913_388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5771 vdd d1 a_40899_n7701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5772 a_13888_n4609# a_14141_n4813# a_13829_n5358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5773 a_32301_2037# a_32306_1651# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5774 a_28395_6410# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5775 a_20168_n7345# a_20164_n7533# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5776 a_30909_5062# a_31166_4872# a_29897_5243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5777 a_6953_7371# a_6740_7371# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5778 a_12422_n9030# a_12209_n9030# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5779 a_27484_n5382# a_27271_n5382# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5780 a_39081_2034# a_38868_2034# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5781 vdd a_19119_n6317# a_18911_n6317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5782 gnd d0 a_36644_n5018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5783 a_38054_5151# a_37841_5151# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5784 gnd d0 a_15140_n7570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5785 vdd d3 a_29954_2629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5786 a_19169_n4588# a_20227_n5026# a_20182_n4822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5787 gnd a_35522_7042# a_35314_7042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5788 a_41558_7030# a_41570_6289# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5789 a_30908_5866# a_31161_5853# a_29892_6224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5790 a_18082_4455# a_17986_367# a_15904_300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5791 a_40356_n6084# a_40476_n8213# a_40427_n8197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5792 a_22411_n5403# a_21990_n5403# a_21717_n5418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5793 a_12573_1523# a_12152_1523# a_12474_1523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5794 a_21983_n7775# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5795 gnd d1 a_8736_n9682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5796 a_22201_n6794# a_21988_n6794# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5797 vdd d0 a_20333_6305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5798 a_3015_n4322# a_3229_n3406# a_3184_n3202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5799 vdd d0 a_41842_1944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5800 a_30896_7826# a_30892_8003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5801 a_501_n5847# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5802 a_29998_n4551# a_31056_n4989# a_31007_n4973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5803 a_9439_1174# a_9696_984# a_8427_1355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5804 a_9503_n7525# a_9513_n6771# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5805 a_919_n6823# a_498_n6823# a_222_n6804# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5806 a_17834_5419# a_17779_6447# a_17987_6447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5807 a_22894_7924# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5808 a_32969_7132# a_33773_6951# a_33932_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5809 a_14803_4943# a_15056_4930# a_13787_5301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5810 a_35315_n7098# a_35410_n7722# a_35365_n7518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5811 a_19149_n8505# a_20207_n8943# a_20158_n8927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5812 a_19087_2167# a_20145_2388# a_20100_2401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5813 a_17817_n9009# a_17435_n9570# a_16843_n9336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5814 a_27268_n6358# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5815 a_6007_n3866# a_5794_n3866# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5816 a_21606_8287# a_22095_8105# a_22303_8105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5817 a_5508_n5426# a_5513_n5040# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5818 gnd a_3366_8044# a_3158_8044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5819 a_12642_n7070# a_12587_n8098# a_12795_n8098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5820 a_37642_n8440# a_38131_n8741# a_38339_n8741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5821 a_41558_8249# a_41811_8236# a_40545_8015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5822 a_2995_n8239# a_3209_n7323# a_3160_n7307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5823 a_11173_n3480# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5824 a_20169_n6552# a_20426_n6568# a_19157_n6733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5825 a_11077_2829# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5826 a_16844_n9751# a_16423_n9751# a_16147_n9450# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5827 a_3168_n5350# a_3272_n4805# a_3227_n4601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5828 a_38371_n2864# a_37950_n2864# a_37674_n2845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5829 a_28532_n8972# a_28319_n8972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5830 a_3172_n5162# a_3425_n5366# a_3019_n4134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5831 a_23742_351# a_26624_263# a_26832_263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5832 vdd a_20434_n4611# a_20226_n4611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5833 a_6214_n3451# a_7019_n3685# a_7188_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5834 a_210_n8764# a_210_n8482# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5835 a_25741_n2431# a_25737_n2619# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5836 a_11283_5201# a_11070_5201# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5837 a_11562_n9357# a_12367_n9591# a_12536_n9030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5838 a_31002_n6327# a_31255_n6531# a_29986_n6696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5839 a_25611_8024# a_25621_7281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5840 a_14891_n5597# a_14901_n4843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5841 a_1793_5432# a_1684_5432# a_1892_5432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5842 a_1706_n9583# a_1493_n9583# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5843 a_16090_2426# a_16579_2244# a_16787_2244# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5844 gnd a_31263_n4574# a_31055_n4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5845 a_11474_8142# a_12278_7961# a_12447_7519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5846 a_14799_5120# a_14807_4382# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5847 a_9504_n7940# a_9761_n7956# a_8495_n7518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5848 a_8515_n3601# a_8768_n3805# a_8465_n3181# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5849 a_39136_1473# a_38923_1473# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5850 a_29606_4634# a_29726_6546# a_29681_6559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5851 a_16166_n6410# a_16169_n6029# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5852 a_6219_n2470# a_5798_n2470# a_5181_n2252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5853 a_35315_n7098# a_35568_n7302# a_35146_n8218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5854 a_23291_3446# a_22919_3026# a_22327_2792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5855 a_22111_4749# a_21898_4749# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5856 a_10814_1184# a_11303_1284# a_11511_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5857 vdd d3 a_3252_n8255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5858 gnd a_14032_7071# a_13824_7071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5859 vdd d0 a_36555_3359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5860 a_26978_n9909# a_26976_n9695# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5861 a_812_7719# a_1617_7953# a_1786_7511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5862 a_32580_1255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5863 a_14792_7318# a_14788_7495# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5864 a_9411_6874# a_9407_7051# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5865 a_19063_6261# a_19320_6071# a_19017_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5866 a_4214_n9318# a_4467_n9522# a_3198_n9687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5867 gnd a_730_n2491# a_938_n2491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5868 a_27387_5709# a_27174_5709# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5869 a_9426_3938# a_9679_3925# a_8410_4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5870 a_25704_n9289# a_25700_n9477# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5871 gnd a_3065_n10418# a_2857_n10418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5872 gnd a_19308_8031# a_19100_8031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5873 a_32542_7698# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5874 a_12543_n6893# a_12434_n7070# a_12642_n7070# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5875 a_37856_2215# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5876 a_4137_5916# a_4133_6093# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5877 a_17888_n4160# a_17675_n4160# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5878 a_30909_6281# a_30905_6458# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5879 vdd d2 a_40849_n7281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5880 a_21734_n3072# a_21732_n2858# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5881 vdd d3 a_19105_6583# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5882 a_694_n9764# a_481_n9764# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5883 vdd d0 a_25975_n6967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5884 a_20068_8278# a_20321_8265# a_19055_8044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5885 a_5409_6053# a_5411_5954# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5886 a_12553_5440# a_12132_5440# a_12459_5559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5887 a_5906_4196# a_5693_4196# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5888 a_32267_8013# a_32756_8113# a_32964_8113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5889 a_5677_6717# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5890 a_36276_7855# a_36272_8032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5891 a_24628_3130# a_25686_3351# a_25641_3364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5892 a_17668_n5653# a_17455_n5653# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5893 a_16880_n2478# a_16459_n2478# a_15842_n2260# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5894 a_33681_n2704# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5895 a_23203_n8061# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5896 a_40639_n8476# a_41697_n8914# a_41652_n8710# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5897 a_11366_n7397# a_11153_n7397# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5898 a_9491_n9485# a_9748_n9501# a_8479_n9666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5899 gnd a_40837_n9241# a_40629_n9241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5900 vdd a_15160_n3653# a_14952_n3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5901 a_33870_4447# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5902 vdd d0 a_20414_n8528# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5903 a_34140_n5084# a_34097_n4152# a_34281_n5900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5904 a_23347_2514# a_23134_2514# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5905 a_35301_1178# a_36359_1399# a_36310_1589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5906 vdd d1 a_24945_n9674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5907 a_32373_n6783# a_32862_n6802# a_33070_n6802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5908 a_3235_n2829# a_4296_n2664# a_4247_n2648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5909 gnd d1 a_3386_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5910 a_8407_5272# a_9468_4901# a_9423_4914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5911 a_12295_5020# a_12082_5020# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5912 a_16147_n9450# a_16149_n9351# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5913 a_8465_n3181# a_8560_n3805# a_8515_n3601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5914 a_20193_n2447# a_20189_n2635# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5915 gnd d0 a_31243_n8491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5916 a_5508_n6021# a_5991_n6387# a_6199_n6387# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5917 a_35146_n8218# a_35360_n7302# a_35315_n7098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5918 a_16572_3223# a_16359_3223# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5919 vdd d0 a_9785_n2643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5920 a_38145_n5390# a_37932_n5390# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5921 a_39238_3552# a_38856_3994# a_38265_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5922 vdd a_35522_7042# a_35314_7042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5923 a_21970_n9320# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5924 a_35075_n6105# a_35328_n6309# a_34959_n10381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5925 vdd d2 a_14098_n3414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5926 a_16366_2244# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5927 a_13806_2188# a_14864_2409# a_14815_2599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5928 a_33592_1074# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5929 gnd a_40830_2125# a_40622_2125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5930 a_10878_n7511# a_10880_n7412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5931 a_36391_n4814# a_36387_n5002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5932 a_22209_n4837# a_21996_n4837# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5933 a_32644_n7783# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5934 gnd a_31149_7813# a_30941_7813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5935 a_26926_1622# a_26924_1408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5936 a_1642_3055# a_1429_3055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5937 a_20165_n7948# a_20168_n7345# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5938 a_23050_n7033# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5939 a_1518_n4685# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5940 a_32983_3781# a_32562_3781# a_32289_3997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5941 a_20157_n8512# a_20169_n7760# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5942 gnd a_20357_992# a_20149_992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5943 a_150_2653# a_148_2439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5944 a_24693_n8677# a_25754_n8512# a_25705_n8496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5945 a_38868_2034# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5946 gnd d0 a_20421_n7549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5947 a_34058_n3124# a_33944_n3124# a_34152_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5948 vdd a_3366_8044# a_3158_8044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5949 a_36289_6310# a_36285_6487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5950 a_41554_8426# a_41811_8236# a_40545_8015# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5951 a_39213_7350# a_38841_6930# a_38249_6696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5952 a_21626_4088# a_21628_3989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5953 a_12380_4476# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5954 a_6918_4015# a_6705_4015# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5955 a_1436_2076# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5956 a_33874_n6621# a_33661_n6621# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5957 vdd d4 a_40609_n6288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5958 a_6131_1255# a_5710_1255# a_5434_1155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5959 a_16755_8121# a_16334_8121# a_16058_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5960 a_38264_3760# a_37843_3760# a_37575_3590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5961 a_21707_n7756# a_22196_n7775# a_22404_n7775# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5962 a_30912_4086# a_31169_3896# a_29900_4267# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5963 a_7415_n8069# a_6994_n8069# a_7250_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5964 a_5690_5172# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5965 a_7067_7490# a_6685_7932# a_6093_7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5966 a_11387_n3895# a_11174_n3895# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5967 gnd a_3163_6596# a_2955_6596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5968 a_32358_n9938# a_36362_n9900# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5969 a_27583_7669# a_27162_7669# a_26894_7499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5970 vdd d0 a_36631_n7956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5971 gnd d0 a_25983_n5010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5972 gnd d1 a_35638_n3805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5973 a_7156_n9001# a_6774_n9562# a_6183_n9743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5974 a_35378_n4580# a_36436_n5018# a_36387_n5002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5975 vdd a_14032_7071# a_13824_7071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5976 a_38333_n9307# a_37912_n9307# a_37639_n9322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5977 a_13871_n7735# a_14932_n7570# a_14883_n7554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5978 a_24509_n4105# a_24762_n4309# a_24410_n6285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5979 a_22307_6709# a_21886_6709# a_21613_6925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5980 a_30922_3343# a_30918_3520# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5981 a_36379_n6959# a_36636_n6975# a_35370_n6537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5982 a_12795_n8098# a_12374_n8098# a_12642_n7070# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5983 a_9434_2155# a_9444_1412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5984 a_17584_3042# a_17371_3042# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5985 a_37575_3590# a_37573_3376# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5986 a_13660_n8059# a_13913_n8263# a_13585_n6134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5987 a_34959_n10381# a_35120_n6309# a_35075_n6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5988 a_5523_n2866# a_6012_n2885# a_6220_n2885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5989 a_8433_n9058# a_8528_n9682# a_8479_n9666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5990 a_10871_n8772# a_11360_n8791# a_11568_n8791# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5991 vdd a_19308_8031# a_19100_8031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5992 a_13895_n3630# a_14148_n3834# a_13845_n3210# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5993 a_40596_n7077# a_40849_n7281# a_40427_n8197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5994 a_40592_n7265# a_40696_n6720# a_40651_n6516# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5995 a_17378_2063# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5996 gnd a_9765_n6560# a_9557_n6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5997 a_32274_7528# a_32272_7314# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5998 vdd a_31251_n7927# a_31043_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5999 a_41562_6853# a_41815_6840# a_40546_7211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6000 a_21898_4749# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6001 a_20064_8455# a_20321_8265# a_19055_8044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6002 a_4121_8053# a_4131_7310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6003 gnd d0 a_41899_n9480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6004 a_33937_7490# a_33823_7371# a_34031_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6005 a_37918_n8741# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6006 a_32849_n8347# a_32636_n8347# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6007 a_27497_n3837# a_27284_n3837# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6008 a_26988_n7735# a_26988_n7453# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6009 a_10782_7061# a_10784_6962# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6010 a_26588_n10440# a_26538_n10456# a_24397_n10373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6011 a_6806_n3685# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6012 gnd a_19105_6583# a_18897_6583# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6013 a_37944_n3430# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6014 a_7062_7371# a_6690_6951# a_6099_7132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6015 vdd d0 a_36618_n9501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6016 a_25712_n7517# a_25722_n6763# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6017 a_19172_n3797# a_19429_n3813# a_19126_n3189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6018 a_28905_n8040# a_28484_n8040# a_28752_n7012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6019 a_22424_n3858# a_22003_n3858# a_21727_n3839# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6020 vdd d0 a_31256_n6946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6021 a_24298_n10373# a_24555_n10389# a_24397_n10373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6022 a_37582_2016# a_38068_1800# a_38276_1800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6023 a_16855_n7376# a_17660_n7610# a_17829_n7049# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6024 a_5243_292# a_7112_359# a_7434_359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6025 a_10796_5002# a_11282_4786# a_11490_4786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6026 a_26981_n8714# a_27470_n8733# a_27678_n8733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6027 a_40566_3294# a_41627_2923# a_41582_2936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6028 a_19090_n9254# a_19194_n8709# a_19145_n8693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6029 a_7112_359# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6030 a_26983_n8333# a_26990_n8132# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6031 gnd d2 a_8609_5643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6032 a_33090_n2885# a_33894_n2704# a_34053_n2947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6033 vdd d1 a_40823_3104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6034 a_35349_n9666# a_36410_n9501# a_36361_n9485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6035 a_7024_n2704# a_6811_n2704# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6036 a_26901_5925# a_27387_5709# a_27595_5709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6037 a_41678_n3399# a_41931_n3603# a_40662_n3768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6038 vdd a_41828_5295# a_41620_5295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6039 a_30994_n7911# a_30997_n7308# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6040 vdd d1 a_30226_n9653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6041 gnd a_40704_n4296# a_40496_n4296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6042 a_30918_3520# a_30921_2928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6043 a_39049_7911# a_38836_7911# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6044 gnd d3 a_3183_2679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6045 a_32631_n9328# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6046 gnd a_26746_n10456# a_26538_n10456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6047 vdd d0 a_4468_n9937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6048 vdd a_40830_2125# a_40622_2125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6049 a_40427_n8197# a_40641_n7281# a_40596_n7077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6050 a_17564_6959# a_17351_6959# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6051 a_5885_7698# a_5672_7698# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6052 a_24709_n6529# a_25767_n6967# a_25722_n6763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6053 vdd a_29954_2629# a_29746_2629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6054 a_32559_4757# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6055 gnd d1 a_14136_n5794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6056 a_10797_4407# a_10797_4125# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6057 a_225_n5828# a_714_n5847# a_922_n5847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6058 a_25726_n4994# a_25983_n5010# a_24717_n4572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6059 a_41589_1957# a_41585_2134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6060 a_138_4613# a_621_4778# a_829_4778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6061 a_31018_n3806# a_31014_n3994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6062 a_28752_n7012# a_28331_n7012# a_28653_n6835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6063 vdd a_20333_6305# a_20125_6305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6064 vdd a_41842_1944# a_41634_1944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6065 a_17358_5980# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6066 a_40356_n6084# a_40609_n6288# a_40240_n10360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6067 a_24573_3691# a_24668_4098# a_24623_4111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6068 a_10784_6962# a_10791_6578# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6069 a_33884_n4152# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6070 vdd d0 a_31150_8228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6071 a_8280_n8030# a_8478_n9262# a_8429_n9246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6072 a_2920_n6314# a_3064_n4338# a_3015_n4322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6073 a_5422_3397# a_5911_3215# a_6119_3215# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6074 a_24642_n9050# a_24737_n9674# a_24692_n9470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6075 a_35281_5095# a_36339_5316# a_36290_5506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6076 a_36398_n3835# a_36394_n4023# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6077 gnd d2 a_30208_n3356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6078 a_19076_3323# a_20137_2952# a_20092_2965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6079 a_6110_4757# a_6915_4991# a_7074_5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6080 a_23288_5522# a_22906_5964# a_22314_5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6081 a_21397_n10599# a_21654_n10615# a_20848_n805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6082 a_5778_n6387# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6083 vdd a_35643_n2824# a_35435_n2824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6084 a_14888_n7781# a_15141_n7985# a_13875_n7547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6085 a_27698_n4816# a_27277_n4816# a_27001_n4797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6086 a_31010_n4370# a_31006_n4558# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6087 a_24619_4288# a_25680_3917# a_25635_3930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6088 gnd d0 a_41823_6276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6089 a_11070_5201# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6090 gnd a_36639_n5999# a_36431_n5999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6091 a_37567_5547# a_38048_5717# a_38256_5717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6092 a_19071_4304# a_20132_3933# a_20083_4123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6093 a_24321_4832# a_24465_2650# a_24416_2840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6094 vdd a_41919_n5563# a_41711_n5563# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6095 a_10504_285# a_10395_285# a_10603_285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6096 a_38073_819# a_37860_819# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6097 a_5416_5568# a_5414_5354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6098 a_37676_n3059# a_37674_n2845# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6099 vdd d0 a_25873_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6100 a_8201_n6293# a_8345_n4317# a_8300_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6101 a_13786_6105# a_14844_6326# a_14795_6516# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6102 a_27380_6688# a_27167_6688# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6103 a_19122_n3377# a_19379_n3393# a_18957_n4309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6104 a_36402_n2439# a_36398_n2627# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6105 vdd a_36555_3359# a_36347_3359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6106 a_3113_8057# a_4171_8278# a_4126_8291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6107 vdd a_25880_5874# a_25672_5874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6108 a_30982_n9871# a_30985_n9268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6109 a_8499_n5749# a_9560_n5584# a_9511_n5568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6110 a_27174_5709# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6111 a_17735_5419# a_17363_4999# a_16772_5180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6112 a_8205_n6105# a_8325_n8234# a_8276_n8218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6113 a_41660_n6938# a_41917_n6954# a_40651_n6516# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6114 a_5243_292# a_5134_292# a_5342_292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6115 a_12159_n8610# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6116 a_40240_n10360# a_40401_n6288# a_40356_n6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6117 a_34063_1494# a_34008_2522# a_34192_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6118 vdd d0 a_9660_8257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6119 a_21606_8287# a_21606_8005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6120 a_39312_7350# a_38891_7350# a_39213_7350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6121 vdd d1 a_8753_n6741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6122 vdd a_19105_6583# a_18897_6583# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6123 a_22411_n5403# a_21990_n5403# a_21722_n5032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6124 a_4248_n3063# a_4251_n2460# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6125 a_21983_n7775# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6126 vdd d1 a_3480_n4805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6127 a_1548_n9022# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6128 a_2021_n6098# a_1808_n6098# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6129 a_34058_n3124# a_33676_n3685# a_33085_n3866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6130 a_5693_4196# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6131 gnd d1 a_30154_5053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6132 a_36374_n7940# a_36377_n7337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6133 a_919_n6823# a_498_n6823# a_222_n6522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6134 a_36366_n8504# a_36378_n7752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6135 a_30929_1145# a_31186_955# a_29917_1326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6136 a_9427_4353# a_9680_4340# a_8414_4119# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6137 a_38339_n8741# a_39143_n8560# a_39302_n8803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6138 a_624_3802# a_411_3802# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6139 a_28569_5501# a_28187_5943# a_27596_6124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6140 a_222_n6804# a_222_n6522# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6141 a_23370_7363# a_22949_7363# a_23276_7482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6142 a_35365_n7518# a_36423_n7956# a_36378_n7752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6143 a_33785_4991# a_33572_4991# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6144 a_37642_n8722# a_38131_n8741# a_38339_n8741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6145 a_25724_n5372# a_25977_n5576# a_24708_n5741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6146 vdd d2 a_8609_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6147 a_23134_2514# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6148 a_16771_4765# a_16350_4765# a_16080_4600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6149 a_28653_n6835# a_28281_n6592# a_27689_n6358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6150 a_12186_n3714# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6151 a_38371_n2864# a_37950_n2864# a_37674_n2563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6152 a_32281_5954# a_32286_5568# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6153 a_29939_n5300# a_30043_n4755# a_29998_n4551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6154 a_10462_n2231# a_11391_n2499# a_11599_n2499# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6155 a_12082_5020# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6156 a_28577_3544# a_28195_3986# a_27603_3752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6157 a_22184_n9735# a_21971_n9735# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6158 a_3227_n4601# a_4285_n5039# a_4240_n4835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6159 a_10893_n5069# a_10891_n4855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6160 a_5799_n2885# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6161 a_24725_n2800# a_24982_n2816# a_24670_n3361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6162 a_4211_n9921# a_4214_n9318# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6163 a_24489_n8022# a_24687_n9254# a_24642_n9050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6164 a_1629_5993# a_1416_5993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6165 gnd a_35611_n8701# a_35403_n8701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6166 a_7270_n5084# a_6849_n5084# a_7171_n4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6167 a_32378_n5426# a_32383_n5040# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6168 a_34021_n8824# a_33649_n8581# a_33057_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6169 a_16460_n2893# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6170 a_5434_1155# a_5436_1056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6171 gnd d0 a_9748_n9501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6172 a_22112_5164# a_21899_5164# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6173 a_3071_5854# a_3175_5103# a_3126_5293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6174 a_24709_n6529# a_24962_n6733# a_24650_n7278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6175 a_11265_7727# a_11052_7727# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6176 a_38354_n5805# a_37933_n5805# a_37657_n5786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6177 a_37573_3094# a_37575_2995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6178 a_38861_3013# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6179 a_4134_6508# a_4391_6318# a_3125_6097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6180 a_39413_n7020# a_38992_n7020# a_39314_n6843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6181 a_41672_n4793# a_41668_n4981# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6182 vdd d3 a_35334_2658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6183 a_26892_7003# a_26894_6904# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6184 a_417_3236# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6185 a_27388_6124# a_27175_6124# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6186 a_3160_n7307# a_3417_n7323# a_2995_n8239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6187 a_28296_n3656# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6188 gnd d3 a_13933_n4346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6189 a_21643_1429# a_22132_1247# a_22340_1247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6190 a_36288_5895# a_36541_5882# a_35272_6253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6191 a_30991_n8702# a_31244_n8906# a_29978_n8468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6192 a_35281_5095# a_36339_5316# a_36294_5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6193 vdd d5 a_13726_n10426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6194 a_41595_1391# a_41848_1378# a_40582_1157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6195 a_35303_n9058# a_35398_n9682# a_35353_n9478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6196 gnd d0 a_4504_n2664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6197 a_17983_4455# a_17586_2530# a_17854_1502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6198 a_6705_4015# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6199 vdd a_31255_n6531# a_31047_n6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6200 a_18076_n8077# a_17963_n6085# a_18171_n6085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6201 a_40635_n8664# a_41696_n8499# a_41647_n8483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6202 a_34063_1494# a_33642_1494# a_33964_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6203 a_5500_n7383# a_5505_n6997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6204 a_17668_n5653# a_17455_n5653# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6205 gnd d2 a_24806_7595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6206 vdd d0 a_41823_6276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6207 a_33069_n6387# a_32648_n6387# a_32375_n6402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6208 a_33681_n2704# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6209 a_28400_5943# a_28187_5943# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6210 a_16097_1064# a_16583_848# a_16791_848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6211 a_23283_5403# a_23174_5403# a_23382_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6212 a_232_n5061# a_713_n5432# a_921_n5432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6213 a_24321_4832# a_24465_2650# a_24420_2663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6214 a_486_n8783# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6215 a_19177_n2816# a_20238_n2651# a_20193_n2447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6216 a_604_7719# a_391_7719# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6217 a_36305_2570# a_36308_1978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6218 gnd d1 a_8659_6063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6219 a_837_2821# a_1642_3055# a_1801_3475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6220 a_12379_n7631# a_12166_n7631# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6221 vdd d0 a_4396_5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6222 gnd a_24861_7034# a_24653_7034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6223 vdd d3 a_19214_n4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6224 a_25640_2949# a_25893_2936# a_24624_3307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6225 a_12556_n5113# a_12174_n5674# a_11583_n5855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6226 a_31018_n3806# a_31271_n4010# a_30005_n3572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6227 a_13786_6105# a_14844_6326# a_14799_6339# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6228 a_19013_5841# a_19117_5090# a_19068_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6229 a_35292_2336# a_36353_1965# a_36308_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6230 a_2045_6460# a_1624_6460# a_1880_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6231 a_35354_n8685# a_35611_n8701# a_35299_n9246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6232 vdd d1 a_3398_2167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6233 a_22126_1813# a_21913_1813# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6234 a_20169_n7760# a_20422_n7964# a_19156_n7526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6235 vdd a_4467_n9522# a_4259_n9522# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6236 a_11158_n6416# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6237 gnd d2 a_13977_7632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6238 a_8515_n3601# a_9573_n4039# a_9528_n3835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6239 a_13833_n5170# a_13928_n5794# a_13879_n5778# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6240 gnd d0 a_41925_n4997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6241 a_17371_3042# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6242 a_16653_n6810# a_16440_n6810# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6243 a_11379_n4459# a_11166_n4459# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6244 a_25726_n4994# a_25729_n4391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6245 a_18941_n8038# a_19139_n9270# a_19094_n9066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6246 a_37575_2995# a_37582_2611# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6247 a_29897_5243# a_30958_4872# a_30913_4885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6248 a_9515_n5380# a_9511_n5568# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6249 a_20105_1420# a_20358_1407# a_19092_1186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6250 a_12531_n8853# a_12422_n9030# a_12630_n9030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6251 a_32304_1155# a_32793_1255# a_33001_1255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6252 a_11580_n6831# a_11159_n6831# a_10883_n6812# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6253 a_21914_2228# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6254 gnd a_8761_n4784# a_8553_n4784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6255 gnd a_35487_3686# a_35279_3686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6256 vdd d0 a_4472_n8541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6257 vdd d1 a_30154_5053# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6258 a_28489_n7573# a_28276_n7573# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6259 a_27401_3186# a_27188_3186# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6260 a_22307_6709# a_23112_6943# a_23271_7363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6261 a_19161_n6545# a_19414_n6749# a_19102_n7294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6262 a_9423_4530# a_9680_4340# a_8414_4119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6263 a_27608_2771# a_27187_2771# a_26914_2987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6264 gnd d0 a_41827_4880# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6265 a_29892_6224# a_30953_5853# a_30904_6043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6266 a_34077_n8069# a_33864_n8069# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6267 gnd a_19422_n4792# a_19214_n4792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6268 a_27268_n6358# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6269 a_17817_n9009# a_17435_n9570# a_16844_n9751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6270 a_16154_n8965# a_16635_n9336# a_16843_n9336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6271 a_17987_6447# a_17566_6447# a_17822_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6272 a_33874_n6621# a_33661_n6621# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6273 a_17911_n9009# a_17490_n9009# a_17812_n8832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6274 a_27620_811# a_28425_1045# a_28584_1465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6275 a_13787_5301# a_14848_4930# a_14799_5120# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6276 a_37649_n7743# a_37649_n7461# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6277 a_10809_2165# a_11298_2265# a_11506_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6278 a_16065_6941# a_16551_6725# a_16759_6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6279 a_34196_6439# a_34083_4447# a_34291_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6280 vdd a_40823_3104# a_40615_3104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6281 a_27690_n6773# a_27269_n6773# a_26993_n6754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6282 gnd d0 a_20332_5890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6283 a_25742_n2846# a_25995_n3050# a_24729_n2612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6284 a_41663_n5962# a_41920_n5978# a_40654_n5540# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6285 a_6219_n2470# a_5798_n2470# a_5525_n2485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6286 a_36382_n6356# a_36635_n6560# a_35366_n6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6287 vdd d2 a_35467_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6288 a_1892_5432# a_1471_5432# a_1798_5551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6289 a_7156_n9001# a_6774_n9562# a_6182_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6290 a_11567_n8376# a_11146_n8376# a_10873_n8391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6291 a_29990_n6508# a_30243_n6712# a_29931_n7257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6292 a_38333_n9307# a_37912_n9307# a_37644_n8936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6293 a_38836_7911# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6294 a_23296_3565# a_22914_4007# a_22323_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6295 a_1981_n7062# a_1926_n8090# a_2134_n8090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6296 a_14871_n9514# a_14881_n8760# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6297 gnd a_36643_n4603# a_36435_n4603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6298 a_37644_n8341# a_37651_n8140# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6299 a_22308_7124# a_21887_7124# a_21611_7024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6300 a_8441_n7286# a_8545_n6741# a_8500_n6537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6301 a_17351_6959# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6302 a_130_6570# a_128_6356# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6303 a_40550_7034# a_41608_7255# a_41559_7445# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6304 a_4999_n10469# a_8138_n10397# a_7510_n6077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6305 a_5672_7698# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6306 a_901_n9349# a_1706_n9583# a_1875_n9022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6307 a_8504_n4768# a_8761_n4784# a_8449_n5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6308 a_16667_n3459# a_16454_n3459# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6309 gnd a_8706_n5345# a_8498_n5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6310 a_23209_4439# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6311 a_34196_6439# a_33775_6439# a_34043_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6312 a_23511_n6069# a_23298_n6069# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6313 a_22926_2047# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6314 gnd d0 a_4379_8278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6315 gnd a_36529_7842# a_36321_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6316 a_24400_6580# a_24598_7595# a_24553_7608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6317 a_34046_n5084# a_33932_n5084# a_34140_n5084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6318 a_27621_1226# a_27200_1226# a_26924_1126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6319 a_8431_1178# a_8684_1165# a_8372_1916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6320 a_3202_n9499# a_3455_n9703# a_3152_n9079# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6321 a_17832_n4915# a_17723_n5092# a_17931_n5092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6322 a_23271_7363# a_22899_6943# a_22307_6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6323 a_13680_n4142# a_13878_n5374# a_13829_n5358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6324 a_37918_n8741# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6325 a_32849_n8347# a_32636_n8347# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6326 a_35230_3876# a_35334_3125# a_35285_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6327 gnd d1 a_19402_n8709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6328 a_8402_6253# a_9463_5882# a_9418_5895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6329 a_22322_3773# a_21901_3773# a_21633_3603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6330 a_33957_3573# a_33843_3454# a_34051_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6331 vdd d1 a_8659_6063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6332 a_32964_8113# a_32543_8113# a_32267_8295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6333 a_28557_7461# a_28175_7903# a_27583_7669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6334 vdd a_24861_7034# a_24653_7034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6335 gnd a_24653_6567# a_24445_6567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6336 gnd d0 a_9680_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6337 a_40584_n9037# a_40679_n9661# a_40634_n9457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6338 a_23000_n6613# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6339 vdd a_9691_1965# a_9483_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6340 gnd a_41823_6276# a_41615_6276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6341 a_9414_6072# a_9424_5329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6342 a_11506_2265# a_12310_2084# a_12479_1642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6343 vdd d2 a_13977_7632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6344 a_3083_3720# a_3178_4127# a_3129_4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6345 a_5402_7032# a_5404_6933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6346 a_36292_4115# a_36549_3925# a_35280_4296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6347 a_23058_n5076# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6348 a_32393_n2584# a_32395_n2485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6349 vdd a_14148_n3834# a_13940_n3834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6350 a_23459_n8993# a_23416_n8061# a_23624_n8061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6351 a_5404_7528# a_5885_7698# a_6093_7698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6352 a_20887_141# a_20674_141# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6353 a_5414_5072# a_5903_5172# a_6111_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6354 vdd a_25873_6853# a_25665_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6355 a_7024_n2704# a_6811_n2704# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6356 a_19060_7063# a_20118_7284# a_20069_7474# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6357 a_26624_263# a_26411_263# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6358 gnd d2 a_3328_5664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6359 a_39378_n4131# a_39165_n4131# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6360 a_29973_n9449# a_31031_n9887# a_30982_n9871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6361 a_29790_n4084# a_29988_n5316# a_29939_n5300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6362 a_33793_3034# a_33580_3034# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6363 a_21970_n9320# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6364 a_39000_n5063# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6365 a_16855_n7376# a_16434_n7376# a_16161_n7391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6366 a_13581_n6322# a_13725_n4346# a_13676_n4330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6367 vdd a_35487_3686# a_35279_3686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6368 gnd a_15039_7871# a_14831_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6369 a_33587_2055# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6370 vdd d1 a_14153_n2853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6371 a_38282_1234# a_37861_1234# a_37585_1416# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6372 a_9532_n2439# a_9785_n2643# a_8516_n2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6373 gnd d0 a_25994_n2635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6374 a_4242_n3629# a_4252_n2875# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6375 a_25648_2385# a_25644_2562# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6376 a_28552_7342# a_28180_6922# a_27589_7103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6377 a_1637_4036# a_1424_4036# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6378 a_36398_n3835# a_36651_n4039# a_35385_n3601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6379 a_118_7935# a_604_7719# a_812_7719# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6380 a_133_5375# a_622_5193# a_830_5193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6381 a_41643_n9879# a_41646_n9276# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6382 a_23271_n5076# a_23058_n5076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6383 a_11474_8142# a_11053_8142# a_10777_8324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6384 a_38244_7677# a_37823_7677# a_37555_7507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6385 gnd a_30154_5053# a_29946_5053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6386 a_5922_840# a_5709_840# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6387 a_7282_n3124# a_7227_n4152# a_7411_n5900# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6388 a_411_3802# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6389 a_6194_n7368# a_5773_n7368# a_5505_n6997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6390 a_21640_2029# a_22126_1813# a_22334_1813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6391 a_6126_2236# a_5705_2236# a_5429_2418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6392 a_33572_4991# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6393 a_14802_4144# a_15059_3954# a_13790_4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6394 a_28717_n4123# a_28504_n4123# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6395 a_5923_1255# a_5710_1255# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6396 gnd d4 a_3088_4671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6397 a_1622_6972# a_1409_6972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6398 vdd a_25957_n9493# a_25749_n9493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6399 a_143_3632# a_141_3418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6400 a_27698_n4816# a_27277_n4816# a_27001_n4515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6401 a_40659_n4559# a_41717_n4997# a_41668_n4981# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6402 vdd a_36656_n3058# a_36448_n3058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6403 a_5404_6933# a_5411_6549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6404 a_36304_2155# a_36314_1412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6405 a_39572_4426# a_39151_4426# a_39473_4426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6406 a_12303_3063# a_12090_3063# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6407 a_37560_6314# a_38049_6132# a_38257_6132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6408 a_6898_7932# a_6685_7932# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6409 a_1416_5993# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6410 a_2140_4468# a_1719_4468# a_2041_4468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6411 a_21720_n4536# a_22209_n4837# a_22417_n4837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6412 a_40550_7034# a_41608_7255# a_41563_7268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6413 a_20085_5337# a_20338_5324# a_19072_5103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6414 gnd d1 a_24957_n7714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6415 a_17579_4023# a_17366_4023# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6416 a_16186_n2493# a_15842_n2260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6417 a_845_2257# a_424_2257# a_148_2157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6418 a_27381_7103# a_27168_7103# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6419 a_8340_7793# a_8444_7042# a_8395_7232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6420 a_11052_7727# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6421 a_21633_3603# a_21631_3389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6422 vdd a_35626_n5765# a_35418_n5765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6423 vdd d1 a_35631_n4784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6424 vdd d0 a_25893_2936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6425 a_41663_n6335# a_41916_n6539# a_40647_n6704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6426 a_7067_7490# a_6953_7371# a_7161_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6427 a_26998_n5992# a_26996_n5778# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6428 a_27271_n5382# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6429 a_8427_1355# a_8684_1165# a_8372_1916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6430 a_7183_n2947# a_7074_n3124# a_7282_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6431 vdd a_35334_2658# a_35126_2658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6432 a_4126_7072# a_4383_6882# a_3114_7253# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6433 vdd d0 a_31169_3896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6434 a_27175_6124# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6435 a_39245_1473# a_38873_1053# a_38281_819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6436 a_35230_3876# a_35334_3125# a_35289_3138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6437 a_28564_n3095# a_28351_n3095# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6438 gnd d3 a_29954_2629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6439 a_3210_n7727# a_4271_n7562# a_4222_n7546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6440 a_20068_8278# a_20064_8455# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6441 a_2134_n8090# a_1713_n8090# a_1981_n7062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6442 a_9402_8032# a_9659_7842# a_8390_8213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6443 a_10789_6082# a_11278_6182# a_11486_6182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6444 a_32306_1651# a_32787_1821# a_32995_1821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6445 a_2999_n8051# a_3252_n8255# a_2924_n6126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6446 a_12890_n6106# a_13726_n10426# a_13568_n10410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6447 vdd d0 a_4493_n5039# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6448 a_33982_359# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6449 vdd d0 a_9680_4340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6450 a_210_n8764# a_699_n8783# a_907_n8783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6451 vdd d0 a_36530_8257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6452 a_23303_1486# a_22931_1066# a_22340_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6453 gnd a_24806_7595# a_24598_7595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6454 vdd a_41823_6276# a_41615_6276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6455 a_17358_5980# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6456 a_7099_1613# a_6717_2055# a_6125_1821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6457 a_18082_4455# a_17661_4455# a_17983_4455# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6458 a_391_7719# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6459 a_6903_6951# a_6690_6951# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6460 a_21625_5560# a_22106_5730# a_22314_5730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6461 a_31002_n6327# a_30998_n6515# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6462 a_16186_n2493# a_16672_n2478# a_16880_n2478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6463 vdd a_4396_5337# a_4188_5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6464 a_41594_976# a_41590_1153# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6465 a_1713_n8090# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6466 a_12186_n3714# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6467 a_16427_n8355# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6468 a_19060_7063# a_20118_7284# a_20073_7297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6469 vdd d2 a_3328_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6470 a_22184_n9735# a_21971_n9735# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6471 a_6697_5972# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6472 vdd a_3398_2167# a_3190_2167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6473 a_12474_1523# a_12102_1103# a_11511_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6474 gnd a_13977_7632# a_13769_7632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6475 a_16090_2144# a_16092_2045# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6476 a_3129_4317# a_4190_3946# a_4145_3959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6477 a_8276_n8218# a_8533_n8234# a_8205_n6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6478 a_16167_n5533# a_16169_n5434# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6479 a_1493_n9583# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6480 gnd a_25983_n5010# a_25775_n5010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6481 a_24603_8028# a_25661_8249# a_25616_8262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6482 a_32631_n9328# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6483 gnd d0 a_4383_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6484 a_41571_5485# a_41828_5295# a_40562_5074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6485 gnd a_15134_n8964# a_14926_n8964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6486 a_13859_n9695# a_14116_n9711# a_13813_n9087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6487 a_6012_n2885# a_5799_n2885# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6488 vdd d0 a_9765_n6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6489 a_37848_2779# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6490 a_12561_3483# a_12140_3483# a_12467_3602# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6491 vdd d5 a_24555_n10389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6492 a_33719_n5084# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6493 a_27008_n3536# a_27497_n3837# a_27705_n3837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6494 a_17715_n7049# a_17502_n7049# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6495 a_118_7935# a_123_7549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6496 a_35276_6076# a_36334_6297# a_36285_6487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6497 a_5417_4378# a_5906_4196# a_6114_4196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6498 a_38354_n5805# a_37933_n5805# a_37657_n5504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6499 gnd a_36650_n3624# a_36442_n3624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6500 gnd d0 a_36655_n2643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6501 a_16172_n4552# a_16661_n4853# a_16869_n4853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6502 gnd a_30258_n3776# a_30050_n3776# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6503 a_37573_3094# a_38062_3194# a_38270_3194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6504 gnd d0 a_36555_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6505 a_128_6074# a_130_5975# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6506 vdd d2 a_14078_n7331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6507 vdd a_30154_5053# a_29946_5053# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6508 a_25712_n7517# a_25969_n7533# a_24700_n7698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6509 a_1711_n8602# a_1498_n8602# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6510 a_24708_n5741# a_24965_n5757# a_24662_n5133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6511 gnd d2 a_24915_n5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6512 a_10898_n3594# a_10900_n3495# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6513 vdd d4 a_40520_4629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6514 a_710_n6408# a_497_n6408# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6515 a_28296_n3656# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6516 gnd a_41827_4880# a_41619_4880# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6517 a_20185_n4031# a_20188_n3428# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6518 a_4154_2591# a_4411_2401# a_3145_2180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6519 a_32376_n5525# a_32865_n5826# a_33073_n5826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6520 a_10603_285# a_10182_285# a_10504_285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6521 a_39225_5390# a_38853_4970# a_38262_5151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6522 a_8484_n8685# a_9545_n8520# a_9496_n8504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6523 a_20177_n4595# a_20189_n3843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6524 a_41585_2134# a_41842_1944# a_40573_2315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6525 a_26924_1408# a_26924_1126# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6526 a_34038_n7041# a_33924_n7041# a_34132_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6527 gnd d1 a_35534_5082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6528 a_10182_285# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6529 a_11486_6182# a_12290_6001# a_12459_5559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6530 vdd d4 a_3088_4671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6531 vdd a_35576_n5345# a_35368_n5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6532 a_41679_n3814# a_41932_n4018# a_40666_n3580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6533 a_27188_3186# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6534 a_16078_4104# a_16567_4204# a_16775_4204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6535 a_5498_n7764# a_5987_n7783# a_6195_n7783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6536 a_227_n5447# a_713_n5432# a_921_n5432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6537 a_32980_4757# a_32559_4757# a_32286_4973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6538 a_1818_1634# a_1704_1515# a_1912_1515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6539 a_12379_n7631# a_12166_n7631# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6540 a_605_8134# a_392_8134# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6541 a_33077_n4430# a_33882_n4664# a_34041_n4907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6542 a_4158_2414# a_4154_2591# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6543 gnd d1 a_3378_6084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6544 gnd a_20332_5890# a_20124_5890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6545 a_12556_n5113# a_12174_n5674# a_11582_n5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6546 a_20081_5514# a_20338_5324# a_19072_5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6547 gnd a_41917_n6954# a_41709_n6954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6548 gnd d1 a_8679_2146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6549 a_24561_5825# a_24665_5074# a_24616_5264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6550 vdd a_35467_7603# a_35259_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6551 a_11158_n6416# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6552 a_8340_7793# a_8444_7042# a_8399_7055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6553 vdd a_31238_n9472# a_31030_n9472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6554 gnd a_9761_n7956# a_9553_n7956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6555 a_32370_n7383# a_32375_n6997# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6556 a_25624_6479# a_25881_6289# a_24615_6068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6557 a_8300_n4113# a_8553_n4317# a_8201_n6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6558 a_13841_n3398# a_13945_n2853# a_13900_n2649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6559 gnd d0 a_15065_3388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6560 gnd d2 a_13997_3715# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6561 a_7193_1494# a_7138_2522# a_7322_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6562 a_13807_1384# a_14064_1194# a_13752_1945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6563 a_36382_n6356# a_36378_n6544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6564 gnd a_15148_n5613# a_14940_n5613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6565 a_41566_6466# a_41569_5874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6566 a_4150_2978# a_4146_3155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6567 gnd d1 a_30238_n7693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6568 a_41664_n6750# a_41660_n6938# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6569 a_16861_n6810# a_17665_n6629# a_17824_n6872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6570 a_5342_292# a_4921_292# a_2252_380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6571 a_39225_n3103# a_39012_n3103# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6572 a_7014_n4152# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6573 a_11580_n6831# a_11159_n6831# a_10883_n6530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6574 a_20095_2163# a_20352_1973# a_19083_2344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6575 a_32388_n3565# a_32390_n3466# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6576 a_28489_n7573# a_28276_n7573# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6577 vdd d1 a_40912_n4763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6578 a_28772_n3095# a_28717_n4123# a_28901_n5871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6579 gnd a_31187_1370# a_30979_1370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6580 a_20075_6080# a_20085_5337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6581 a_7250_n9001# a_6829_n9001# a_7156_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6582 a_17760_1621# a_17646_1502# a_17854_1502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6583 a_13809_n9275# a_14066_n9291# a_13660_n8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6584 vdd a_9684_2944# a_9476_2944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6585 a_38338_n8326# a_39143_n8560# a_39302_n8803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6586 vdd d2 a_35556_n9262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6587 gnd a_24555_n10389# a_24347_n10389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6588 a_31018_n2598# a_31275_n2614# a_30006_n2779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6589 gnd d4 a_24667_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6590 a_23377_n7033# a_22995_n7594# a_22404_n7775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6591 a_16149_n9351# a_16635_n9336# a_16843_n9336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6592 gnd d0 a_15153_n4632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6593 gnd a_14133_n6770# a_13925_n6770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6594 a_37568_4357# a_37568_4075# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6595 a_16775_4204# a_17579_4023# a_17748_3581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6596 a_21996_n4837# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6597 vdd a_13977_7632# a_13769_7632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6598 a_16766_5746# a_16345_5746# a_16072_5962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6599 a_24654_n7090# a_24749_n7714# a_24700_n7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6600 a_2001_n3145# a_1580_n3145# a_1902_n2968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6601 a_29701_2642# a_29899_3657# a_29854_3670# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6602 a_12077_6001# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6603 a_26998_n5397# a_27484_n5382# a_27692_n5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6604 a_27690_n6773# a_27269_n6773# a_26993_n6472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6605 a_35319_n5329# a_35423_n4784# a_35378_n4580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6606 a_27003_n4416# a_27010_n4215# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6607 a_11174_n3895# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6608 a_38365_n3430# a_39170_n3664# a_39339_n3103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6609 a_4230_n5589# a_4487_n5605# a_3218_n5770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6610 gnd a_3328_5664# a_3120_5664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6611 a_16166_n7005# a_16164_n6791# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6612 a_38068_1800# a_37855_1800# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6613 a_33580_3034# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6614 vdd a_20435_n5026# a_20227_n5026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6615 a_6861_n3124# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6616 a_11089_869# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6617 a_11567_n8376# a_11146_n8376# a_10880_n8190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6618 a_10395_285# a_10182_285# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6619 gnd a_41931_n3603# a_41723_n3603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6620 vdd d0 a_31167_5287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6621 gnd a_40684_n8213# a_40476_n8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6622 a_29850_3847# a_29954_3096# a_29905_3286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6623 vdd a_3437_n3406# a_3229_n3406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6624 a_22107_6145# a_21894_6145# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6625 gnd a_31264_n4989# a_31056_n4989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6626 a_38856_3994# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6627 a_40541_8192# a_41602_7821# a_41557_7834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6628 a_29850_3847# a_30107_3657# a_29701_2642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6629 a_12702_4476# a_12305_2551# a_12561_3483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6630 a_26909_3968# a_26914_3582# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6631 gnd a_20415_n8943# a_20207_n8943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6632 a_11392_n2914# a_11179_n2914# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6633 a_27673_n9714# a_27252_n9714# a_26976_n9695# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6634 a_1424_4036# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6635 a_32289_3997# a_32294_3611# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6636 vdd a_4492_n4624# a_4284_n4624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6637 vdd d1 a_35534_5082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6638 gnd a_3417_n7323# a_3209_n7323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6639 a_3215_n6746# a_3472_n6762# a_3160_n7307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6640 vdd a_40857_n5324# a_40649_n5324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6641 a_19122_n3377# a_19226_n2832# a_19177_n2816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6642 a_29973_n9449# a_30226_n9653# a_29923_n9029# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6643 gnd d0 a_41936_n2622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6644 a_207_n9959# a_4468_n9937# a_3202_n9499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6645 a_16459_n2478# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6646 a_21608_7906# a_21613_7520# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6647 vdd a_36566_984# a_36358_984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6648 gnd a_21654_n10615# a_21446_n10615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6649 a_212_n8978# a_210_n8764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6650 a_16181_n3474# a_16186_n3088# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6651 a_17723_n5092# a_17510_n5092# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6652 a_5710_1255# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6653 vdd d1 a_3378_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6654 a_33855_1494# a_33642_1494# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6655 a_3130_5116# a_4188_5337# a_4143_5350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6656 gnd a_4500_n4060# a_4292_n4060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6657 a_23000_n6613# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6658 a_24561_5825# a_24665_5074# a_24620_5087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6659 vdd d1 a_8679_2146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6660 a_12090_3063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6661 vdd a_8698_n7302# a_8490_n7302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6662 a_16754_7706# a_17559_7940# a_17728_7498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6663 a_35277_5272# a_36338_4901# a_36289_5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6664 a_27502_n2856# a_27289_n2856# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6665 a_143_3037# a_150_2653# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6666 a_6685_7932# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6667 a_9492_n9900# a_9749_n9916# a_8483_n9478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6668 a_37555_6912# a_38041_6696# a_38249_6696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6669 a_150_2653# a_629_2821# a_837_2821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6670 vdd a_15161_n4068# a_14953_n4068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6671 vdd d2 a_13997_3715# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6672 a_35386_n2808# a_36447_n2643# a_36398_n2627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6673 a_16653_n6810# a_16440_n6810# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6674 a_5397_8295# a_5886_8113# a_6094_8113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6675 a_21697_n9930# a_25701_n9892# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6676 a_11379_n4459# a_11166_n4459# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6677 a_29951_n3340# a_30055_n2795# a_30006_n2779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6678 a_28663_5382# a_28242_5382# a_28564_5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6679 a_19051_8221# a_20112_7850# a_20067_7863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6680 a_17366_4023# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6681 a_25615_7847# a_25611_8024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6682 a_21886_6709# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6683 a_24509_n4105# a_24707_n5337# a_24658_n5321# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6684 a_20100_1182# a_16104_863# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6685 a_37659_n6000# a_38142_n6366# a_38350_n6366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6686 a_23534_351# a_23321_351# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6687 vdd a_25893_2936# a_25685_2936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6688 gnd a_8617_3686# a_8409_3686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6689 a_16855_n7376# a_16434_n7376# a_16166_n7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6690 vdd d0 a_20441_n3632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6691 a_24485_n8210# a_24699_n7294# a_24650_n7278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6692 a_14819_1203# a_10823_884# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6693 a_32652_n5826# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6694 a_28911_4418# a_28815_330# a_26733_263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6695 a_34281_n5900# a_33884_n4152# a_34140_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6696 vdd a_31187_1370# a_30979_1370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6697 vdd a_20340_3933# a_20132_3933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6698 a_33711_n7041# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6699 a_34285_n8069# a_34172_n6077# a_34380_n6077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6700 vdd d0 a_9786_n3058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6701 vdd a_30119_1697# a_29911_1697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6702 a_27396_4167# a_27183_4167# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6703 gnd d0 a_31270_n3595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6704 gnd a_29954_2629# a_29746_2629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6705 a_27167_6688# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6706 a_3202_n9499# a_4260_n9937# a_207_n9959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6707 a_10885_n7026# a_11366_n7397# a_11574_n7397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6708 a_7082_3454# a_6710_3034# a_6118_2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6709 a_3172_n5162# a_3267_n5786# a_3218_n5770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6710 gnd a_15166_n3087# a_14958_n3087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6711 a_39233_3433# a_39124_3433# a_39332_3433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6712 gnd a_20429_n5592# a_20221_n5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6713 a_5774_n7783# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6714 a_37659_n6000# a_37657_n5786# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6715 vdd d1 a_3460_n8722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6716 a_10791_6578# a_11270_6746# a_11478_6746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6717 a_16868_n4438# a_16447_n4438# a_16181_n4252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6718 a_33669_n4664# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6719 a_2229_n6098# a_1808_n6098# a_2134_n8090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6720 a_29939_n5300# a_30196_n5316# a_29790_n4084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6721 a_36386_n4587# a_36398_n3835# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6722 gnd d0 a_31150_8228# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6723 a_6690_6951# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6724 a_11161_n5440# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6725 a_242_n2887# a_242_n2605# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6726 a_16338_6725# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6727 a_26904_5043# a_27393_5143# a_27601_5143# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6728 a_29974_n8656# a_31035_n8491# a_30990_n8287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6729 a_8500_n6537# a_9558_n6975# a_9509_n6959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6730 vdd a_3328_5664# a_3120_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6731 vdd a_25888_3917# a_25680_3917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6732 gnd d4 a_29948_n6280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6733 a_23194_1486# a_22981_1486# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6734 a_34021_n8824# a_33912_n9001# a_34120_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6735 a_29923_n9029# a_30176_n9233# a_29770_n8001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6736 a_24720_n3781# a_25781_n3616# a_25732_n3600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6737 a_24640_1170# a_25698_1391# a_25649_1581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6738 a_621_4778# a_408_4778# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6739 a_23620_n5892# a_23223_n4144# a_23491_n3116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6740 a_8419_3138# a_9477_3359# a_9432_3372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6741 a_39566_n8048# a_39145_n8048# a_39401_n8980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6742 a_22409_n6794# a_21988_n6794# a_21712_n6493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6743 a_29786_n4272# a_30000_n3356# a_29951_n3340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6744 a_34152_n3124# a_33731_n3124# a_34058_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6745 a_20172_n5576# a_20182_n4822# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6746 a_40566_3294# a_40823_3104# a_40511_3855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6747 a_1761_n9022# a_1548_n9022# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6748 gnd d1 a_14047_4135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6749 a_4231_n6004# a_4234_n5401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6750 a_17452_n6629# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6751 a_21720_n4818# a_22209_n4837# a_22417_n4837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6752 a_706_n7804# a_493_n7804# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6753 gnd d0 a_4479_n7562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6754 a_25628_6302# a_25624_6479# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6755 a_20075_6080# a_20332_5890# a_19063_6261# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6756 vdd d3 a_40684_n8213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6757 a_9497_n8919# a_9500_n8316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6758 a_16440_n6810# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6759 a_28504_n4123# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6760 a_922_n5847# a_501_n5847# a_225_n5828# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6761 a_40600_n5308# a_40704_n4763# a_40659_n4559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6762 a_16667_n3459# a_16454_n3459# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6763 a_12890_n6106# a_12469_n6106# a_12795_n8098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6764 a_7138_2522# a_6925_2522# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6765 a_37841_5151# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6766 a_22340_1247# a_21919_1247# a_21643_1429# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6767 a_11493_3810# a_11072_3810# a_10799_4026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6768 a_19088_1363# a_20149_992# a_20104_1005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6769 a_148_2439# a_637_2257# a_845_2257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6770 a_38334_n9722# a_37913_n9722# a_37637_n9703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6771 gnd a_36555_3359# a_36347_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6772 a_5525_n3080# a_5523_n2866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6773 a_19152_n7714# a_20213_n7549# a_20168_n7345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6774 a_29786_n4272# a_30043_n4288# a_29691_n6264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6775 a_6118_2800# a_5697_2800# a_5431_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6776 a_3113_8057# a_4171_8278# a_4122_8468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6777 a_24298_n10373# a_24459_n6301# a_24410_n6285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6778 a_13884_n4797# a_14945_n4632# a_14896_n4616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6779 a_27616_2207# a_27195_2207# a_26919_2389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6780 a_33988_6439# a_33775_6439# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6781 a_4146_3155# a_4403_2965# a_3134_3336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6782 a_23719_n6069# a_23298_n6069# a_23620_n5892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6783 gnd d0 a_9660_8257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6784 gnd a_35534_5082# a_35326_5082# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6785 a_10898_n3876# a_11387_n3895# a_11595_n3895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6786 gnd d1 a_3371_7063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6787 a_23491_n3116# a_23070_n3116# a_23392_n2939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6788 a_17648_n9570# a_17435_n9570# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6789 gnd a_36644_n5018# a_36436_n5018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6790 a_38957_n3664# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6791 a_39175_n2683# a_38962_n2683# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6792 a_20100_2401# a_20096_2578# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6793 a_22906_5964# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6794 a_39116_5390# a_38903_5390# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6795 a_23630_4439# a_23209_4439# a_23531_4439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6796 a_41652_n8710# a_41905_n8914# a_40639_n8476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6797 a_29000_n6048# a_28579_n6048# a_28905_n8040# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6798 gnd a_40892_n8680# a_40684_n8680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6799 a_392_8134# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6800 a_37945_n3845# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6801 gnd a_3378_6084# a_3170_6084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6802 a_21618_6327# a_22107_6145# a_22315_6145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6803 a_16427_n8355# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6804 a_41570_6289# a_41823_6276# a_40557_6055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6805 a_227_n6042# a_225_n5828# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6806 gnd d1 a_8741_n8701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6807 gnd a_8736_n9682# a_8528_n9682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6808 a_19181_n2628# a_20239_n3066# a_20190_n3050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6809 a_29830_7764# a_29934_7013# a_29885_7203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6810 vdd a_24927_n3377# a_24719_n3377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6811 a_31994_256# a_31885_256# a_20996_141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6812 a_9440_1589# a_9697_1399# a_8431_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6813 a_28557_7461# a_28443_7342# a_28651_7342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6814 vdd a_8617_3686# a_8409_3686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6815 a_30898_7437# a_31155_7247# a_29889_7026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6816 vdd d1 a_35537_4106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6817 a_22119_2792# a_21906_2792# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6818 a_25616_7043# a_25873_6853# a_24604_7224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6819 a_13567_6794# a_13781_5672# a_13732_5862# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6820 gnd a_15065_3388# a_14857_3388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6821 a_20092_2965# a_20088_3142# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6822 gnd a_13997_3715# a_13789_3715# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6823 a_20072_6882# a_20325_6869# a_19056_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6824 a_1989_n5105# a_1568_n5105# a_1895_n5105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6825 a_29900_4267# a_30157_4077# a_29854_3670# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6826 a_18072_n5908# a_17675_n4160# a_17943_n3132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6827 a_27008_n3818# a_27497_n3837# a_27705_n3837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6828 a_12498_6468# a_12285_6468# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6829 a_4247_n3856# a_4243_n4044# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6830 a_40667_n2787# a_41728_n2622# a_41679_n2606# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6831 vdd d0 a_15129_n9945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6832 vdd d0 a_41831_4319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6833 a_16172_n4834# a_16661_n4853# a_16869_n4853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6834 a_155_1077# a_162_876# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6835 gnd d1 a_19313_7050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6836 vdd d0 a_36549_3925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6837 a_12650_n5113# a_12229_n5113# a_12556_n5113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6838 a_4138_6331# a_4391_6318# a_3125_6097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6839 a_1711_n8602# a_1498_n8602# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6840 a_33065_n7783# a_32644_n7783# a_32368_n7482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6841 a_6098_6717# a_5677_6717# a_5404_6933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6842 a_12642_n7070# a_12221_n7070# a_12548_n7070# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6843 gnd d3 a_35334_2658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6844 a_28589_1584# a_28207_2026# a_27615_1792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6845 a_38891_7350# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6846 a_23390_3446# a_22969_3446# a_23291_3446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6847 a_32376_n5807# a_32865_n5826# a_33073_n5826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6848 gnd d1 a_24982_n2816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6849 a_5995_n5826# a_5782_n5826# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6850 a_6194_n7368# a_5773_n7368# a_5500_n7383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6851 gnd a_19320_6071# a_19112_6071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6852 vdd a_4499_n3645# a_4291_n3645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6853 a_38036_7677# a_37823_7677# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6854 vdd d0 a_9754_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6855 a_34291_4447# a_33870_4447# a_34196_6439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6856 a_20080_6318# a_20333_6305# a_19067_6084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6857 a_25641_3364# a_25637_3541# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6858 vdd d0 a_15045_7305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6859 a_14901_n4843# a_14897_n5031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6860 a_5918_2236# a_5705_2236# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6861 a_32279_6053# a_32768_6153# a_32976_6153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6862 a_5689_4757# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6863 a_4219_n8337# a_4472_n8541# a_3203_n8706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6864 a_35071_n6293# a_35215_n4317# a_35166_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6865 a_37669_n3826# a_37669_n3544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6866 a_17817_n9009# a_17703_n9009# a_17911_n9009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6867 a_34291_4447# a_34195_359# a_34403_359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6868 a_32981_5172# a_32560_5172# a_32284_5072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6869 vdd d1 a_14047_4135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6870 a_33078_n4845# a_33882_n4664# a_34041_n4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6871 a_30928_1949# a_30924_2126# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6872 gnd a_9665_7276# a_9457_7276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6873 a_817_6738# a_396_6738# a_130_6570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6874 a_22100_7124# a_21887_7124# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6875 gnd d0 a_4396_5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6876 a_28760_n5055# a_28339_n5055# a_28666_n5055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6877 a_16159_n7490# a_16161_n7391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6878 a_26907_4349# a_27396_4167# a_27604_4167# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6879 gnd a_8667_4106# a_8459_4106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6880 a_7510_n6077# a_8346_n10397# a_4999_n10469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6881 a_23392_n2939# a_23020_n2696# a_22428_n2462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6882 a_33959_n6077# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6883 gnd d1 a_3398_2167# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6884 vdd a_31167_5287# a_30959_5287# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6885 a_207_n9959# a_205_n9745# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6886 a_17673_n4672# a_17460_n4672# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6887 a_3150_1199# a_4208_1420# a_4159_1610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6888 a_1932_4468# a_1719_4468# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6889 vdd a_41920_n5978# a_41712_n5978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6890 a_27376_8084# a_27163_8084# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6891 a_938_n2491# a_517_n2491# a_244_n2506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6892 vdd d0 a_15059_3954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6893 a_21631_3107# a_22120_3207# a_22328_3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6894 a_37664_n4424# a_37671_n4223# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6895 a_9496_n8504# a_9753_n8520# a_8484_n8685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6896 a_19165_n4776# a_20226_n4611# a_20177_n4595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6897 vdd a_30169_2117# a_29961_2117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6898 vdd a_15165_n2672# a_14957_n2672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6899 a_16584_1263# a_16371_1263# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6900 gnd d1 a_40835_1144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6901 gnd d3 a_13844_2687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6902 gnd a_8686_n9262# a_8478_n9262# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6903 gnd a_3272_n4338# a_3064_n4338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6904 vdd d1 a_24950_n8693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6905 gnd d0 a_31154_6832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6906 gnd d0 a_9761_n7956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6907 a_39250_1592# a_38868_2034# a_38277_2215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6908 vdd a_35534_5082# a_35326_5082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6909 a_34051_3454# a_33630_3454# a_33957_3573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6910 a_32313_855# a_32792_840# a_33000_840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6911 a_8503_n5561# a_9561_n5999# a_9512_n5983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6912 vdd d1 a_3371_7063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6913 a_10799_4621# a_10797_4407# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6914 gnd a_31161_5853# a_30953_5853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6915 a_23360_n8816# a_23251_n8993# a_23459_n8993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6916 a_37932_n5390# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6917 a_33699_n9001# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6918 a_32995_1821# a_32574_1821# a_32301_2037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6919 vdd d0 a_25989_n3616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6920 vdd d1 a_3467_n7743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6921 a_22412_n5818# a_21991_n5818# a_21715_n5517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6922 a_9443_997# a_9439_1174# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6923 vdd a_3378_6084# a_3170_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6924 a_24553_7608# a_24806_7595# a_24400_6580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6925 vdd a_8553_n4317# a_8345_n4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6926 a_20189_n3843# a_20185_n4031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6927 a_25637_3541# a_25640_2949# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6928 a_41566_6466# a_41823_6276# a_40557_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6929 a_39225_5390# a_38853_4970# a_38261_4736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6930 a_29830_7764# a_29934_7013# a_29889_7026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6931 a_17874_4455# a_17661_4455# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6932 a_1692_3475# a_1479_3475# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6933 a_21996_n4837# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6934 a_23251_n8993# a_23038_n8993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6935 a_933_n3472# a_1738_n3706# a_1907_n3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6936 a_16767_6161# a_16346_6161# a_16070_6061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6937 a_9507_n7337# a_9760_n7541# a_8491_n7706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6938 a_13567_6794# a_13781_5672# a_13736_5685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6939 a_37568_4075# a_38057_4175# a_38265_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6940 a_12541_7400# a_12120_7400# a_12447_7519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6941 a_17943_n3132# a_17522_n3132# a_17849_n3132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6942 a_492_n7389# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6943 vdd a_13997_3715# a_13789_3715# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6944 a_25725_n5787# a_25978_n5991# a_24712_n5553# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6945 a_38366_n3845# a_39170_n3664# a_39339_n3103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6946 a_3114_7253# a_4175_6882# a_4126_7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6947 gnd a_8533_n8234# a_8325_n8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6948 a_31001_n5539# a_31258_n5555# a_29989_n5720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6949 gnd a_24965_n5757# a_24757_n5757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6950 a_13724_7645# a_13977_7632# a_13571_6617# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6951 a_7079_5530# a_6697_5972# a_6105_5738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6952 gnd d3 a_8444_6575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6953 a_16791_848# a_16370_848# a_16104_863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6954 a_38069_2215# a_37856_2215# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6955 gnd d0 a_9664_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6956 a_16370_848# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6957 vdd d1 a_19313_7050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6958 vdd a_30208_n3356# a_30000_n3356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6959 vdd d0 a_15145_n6589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6960 a_22328_3207# a_23132_3026# a_23291_3446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6961 a_29834_7587# a_30087_7574# a_29681_6559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6962 a_22319_4749# a_21898_4749# a_21625_4965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6963 a_23038_n8993# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6964 a_17596_1082# a_17383_1082# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6965 a_27183_4167# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6966 a_710_n6408# a_497_n6408# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6967 a_505_n4451# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6968 a_11392_n2914# a_11179_n2914# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6969 vdd d0 a_31259_n5970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6970 a_27673_n9714# a_27252_n9714# a_26976_n9413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6971 gnd d0 a_25974_n6552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6972 vdd a_19320_6071# a_19112_6071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6973 gnd a_35638_n3805# a_35430_n3805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6974 a_33964_1494# a_33855_1494# a_34063_1494# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6975 a_7151_n8824# a_6779_n8581# a_6188_n8762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6976 a_32395_n2485# a_32881_n2470# a_33089_n2470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6977 a_41663_n5962# a_41666_n5359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6978 a_41574_4893# a_41827_4880# a_40558_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6979 vdd a_19397_n9690# a_19189_n9690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6980 a_232_n4466# a_239_n4265# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6981 a_21695_n9434# a_22184_n9735# a_22392_n9735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6982 a_20068_8278# a_21606_8287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6983 a_12814_388# a_13541_4679# a_13496_4692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6984 a_23228_n3677# a_23015_n3677# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6985 a_8429_n9246# a_8533_n8701# a_8484_n8685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6986 gnd a_20321_8265# a_20113_8265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6987 a_13900_n2649# a_14153_n2853# a_13841_n3398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6988 vdd a_9665_7276# a_9457_7276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6989 a_37394_271# a_39263_338# a_39585_338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6990 vdd a_8597_7603# a_8389_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6991 a_39421_n5063# a_39000_n5063# a_39327_n5063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6992 a_39263_338# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6993 a_1912_1515# a_1491_1515# a_1813_1515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6994 a_5134_292# a_4921_292# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6995 a_16070_6343# a_16070_6061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6996 a_24712_n5553# a_25770_n5991# a_25725_n5787# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6997 a_20739_n805# a_20526_n805# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6998 a_27502_n2856# a_27289_n2856# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6999 a_3150_1199# a_4208_1420# a_4163_1433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7000 a_22396_n8339# a_23201_n8573# a_23360_n8816# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7001 a_19181_n2628# a_20239_n3066# a_20194_n2862# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7002 a_7173_5411# a_7118_6439# a_7326_6439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7003 gnd a_14047_4135# a_13839_4135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7004 a_13863_n9507# a_14921_n9945# a_10868_n9967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7005 a_7161_7371# a_6740_7371# a_7067_7490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7006 a_4142_4935# a_4395_4922# a_3126_5293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7007 gnd d1 a_8748_n7722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7008 vdd d1 a_40835_1144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7009 vdd d0 a_9697_1399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7010 vdd d0 a_36623_n8520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7011 vdd a_36618_n9501# a_36410_n9501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7012 a_32988_2800# a_33793_3034# a_33952_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7013 a_22914_4007# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7014 a_513_n3887# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7015 a_19177_n2816# a_19434_n2832# a_19122_n3377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7016 a_37656_n6381# a_38142_n6366# a_38350_n6366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7017 a_11159_n6831# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7018 vdd d0 a_4410_1986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7019 a_4131_7310# a_4127_7487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7020 a_21887_7124# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7021 a_16860_n6395# a_17665_n6629# a_17824_n6872# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7022 a_40573_2315# a_41634_1944# a_41585_2134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7023 a_32652_n5826# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7024 a_17829_n7049# a_17447_n7610# a_16855_n7376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7025 a_1981_n7062# a_1560_n7062# a_1887_n7062# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7026 vdd d2 a_8686_n9262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7027 a_33823_7371# a_33610_7371# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7028 a_13752_1945# a_13856_1194# a_13811_1207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7029 a_33775_6439# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7030 a_14876_n8533# a_15133_n8549# a_13864_n8714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7031 a_813_8134# a_1617_7953# a_1786_7511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7032 a_28544_n7012# a_28331_n7012# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7033 a_3180_n3390# a_3284_n2845# a_3239_n2641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7034 vdd a_20446_n2651# a_20238_n2651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7035 a_29943_n5112# a_30038_n5736# a_29989_n5720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7036 a_11574_n7397# a_12379_n7631# a_12548_n7070# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7037 a_24620_5087# a_25678_5308# a_25633_5321# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7038 vdd d1 a_30231_n8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7039 a_11493_3810# a_12298_4044# a_12467_3602# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7040 a_17854_1502# a_17433_1502# a_17755_1502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7041 vdd d0 a_4473_n8956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7042 a_19092_1186# a_20150_1407# a_20105_1420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7043 a_12394_n4181# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7044 a_24724_n3593# a_24977_n3797# a_24674_n3173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7045 a_33669_n4664# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7046 a_10782_7343# a_11271_7161# a_11479_7161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7047 a_123_6954# a_130_6570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7048 a_21901_3773# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7049 vdd d0 a_31162_6268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7050 gnd d1 a_14141_n4813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7051 a_26976_n9413# a_26978_n9314# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7052 a_27269_n6773# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7053 a_5434_1437# a_5923_1255# a_6131_1255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7054 a_26914_2987# a_26921_2603# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7055 gnd a_35588_n3385# a_35380_n3385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7056 a_31022_n2410# a_31018_n2598# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7057 gnd a_8647_8023# a_8439_8023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7058 gnd d0 a_36630_n7541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7059 a_16147_n9450# a_16636_n9751# a_16844_n9751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7060 a_10893_n4474# a_11379_n4459# a_11587_n4459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7061 a_26733_263# a_28602_330# a_28911_4418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7062 a_8461_n3369# a_8718_n3385# a_8296_n4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7063 gnd a_15149_n6028# a_14941_n6028# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7064 a_16358_2808# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7065 a_13720_7822# a_13977_7632# a_13571_6617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7066 a_16095_1445# a_16584_1263# a_16792_1263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7067 a_28602_330# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7068 vdd d3 a_8444_6575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7069 vdd a_19347_n9270# a_19139_n9270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7070 a_9516_n5795# a_9512_n5983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7071 vdd a_13933_n4346# a_13725_n4346# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7072 a_24631_2328# a_25692_1957# a_25647_1970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7073 a_21613_6925# a_21620_6541# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7074 gnd a_29859_4621# a_29651_4621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7075 vdd a_35537_4106# a_35329_4106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7076 gnd d2 a_8597_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7077 a_4232_n6792# a_4485_n6996# a_3219_n6558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7078 a_21732_n2576# a_21734_n2477# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7079 a_19083_2344# a_20144_1973# a_20095_2163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7080 a_24638_n9238# a_24742_n8693# a_24697_n8489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7081 a_29830_7764# a_30087_7574# a_29681_6559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7082 a_7074_5411# a_6965_5411# a_7173_5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7083 a_8112_4840# a_8256_2658# a_8211_2671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7084 a_27684_n7339# a_28489_n7573# a_28658_n7012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7085 a_706_n7804# a_493_n7804# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7086 a_16755_8121# a_17559_7940# a_17728_7498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7087 a_121_7053# a_610_7153# a_818_7153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7088 a_922_n5847# a_501_n5847# a_225_n5546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7089 a_12285_6468# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7090 gnd a_31250_n7512# a_31042_n7512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7091 a_34132_n7041# a_34077_n8069# a_34285_n8069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7092 a_4127_7487# a_4130_6895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7093 a_9431_2957# a_9684_2944# a_8415_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7094 a_28572_3425# a_28200_3005# a_27608_2771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7095 a_27392_4728# a_27179_4728# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7096 a_11568_n8791# a_11147_n8791# a_10871_n8772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7097 a_38334_n9722# a_37913_n9722# a_37637_n9421# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7098 a_11494_4225# a_11073_4225# a_10797_4125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7099 gnd a_19313_7050# a_19105_7050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7100 a_27689_n6358# a_27268_n6358# a_26998_n5992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7101 a_1634_5012# a_1421_5012# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7102 a_34043_5411# a_33622_5411# a_33949_5530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7103 vdd a_41924_n4582# a_41716_n4582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7104 a_37861_1234# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7105 a_33052_n9328# a_33857_n9562# a_34026_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7106 gnd a_35334_2658# a_35126_2658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7107 vdd a_9768_n5584# a_9560_n5584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7108 a_11594_n3480# a_11173_n3480# a_10900_n3495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7109 vdd d0 a_20426_n6568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7110 a_5911_3215# a_5698_3215# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7111 vdd d2 a_3336_3707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7112 gnd d2 a_3425_n5366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7113 a_16174_n5048# a_16172_n4834# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7114 vdd a_20321_8265# a_20113_8265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7115 a_16083_3405# a_16083_3123# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7116 a_26926_1027# a_27412_811# a_27620_811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7117 a_37823_7677# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7118 vdd a_30176_n9233# a_29968_n9233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7119 a_32767_5738# a_32554_5738# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7120 a_35353_n9478# a_35606_n9682# a_35303_n9058# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7121 a_39324_5390# a_38903_5390# a_39225_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7122 gnd d0 a_31255_n6531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7123 a_13825_n7127# a_13920_n7751# a_13875_n7547# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7124 gnd d1 a_40924_n2803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7125 vdd d7 a_10656_n10500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7126 vdd a_19194_n8242# a_18986_n8242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7127 a_32547_6717# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7128 vdd a_15045_7305# a_14837_7305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7129 a_5705_2236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7130 gnd d0 a_36530_8257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7131 a_37548_7992# a_38037_8092# a_38245_8092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7132 a_38957_n3664# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7133 a_6098_6717# a_6903_6951# a_7062_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7134 gnd d2 a_35568_n7302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7135 a_636_1842# a_423_1842# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7136 a_9439_2393# a_9692_2380# a_8426_2159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7137 a_2041_4468# a_1644_2543# a_1912_1515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7138 gnd d1 a_3391_3146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7139 a_22200_n6379# a_21987_n6379# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7140 a_17346_7940# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7141 vdd a_14047_4135# a_13839_4135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7142 a_19144_n9486# a_20202_n9924# a_16149_n9946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7143 a_37945_n3845# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7144 a_15904_300# a_15795_300# a_10504_285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7145 a_833_4217# a_412_4217# a_136_4399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7146 a_35284_4119# a_36342_4340# a_36293_4530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7147 gnd a_4396_5337# a_4188_5337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7148 vdd a_8753_n6741# a_8545_n6741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7149 gnd d1 a_19429_n3813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7150 a_11058_7161# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7151 a_20164_n7533# a_20174_n6779# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7152 a_28628_2493# a_28415_2493# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7153 a_13876_n6754# a_14937_n6589# a_14892_n6385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7154 gnd d0 a_4467_n9522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7155 a_16075_5080# a_16564_5180# a_16772_5180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7156 a_37565_5051# a_37567_4952# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7157 gnd a_3398_2167# a_3190_2167# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7158 gnd d2 a_40780_1705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7159 vdd a_25869_8249# a_25661_8249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7160 a_24603_8028# a_25661_8249# a_25612_8439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7161 a_27163_8084# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7162 a_24705_n6717# a_25766_n6552# a_25717_n6536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7163 a_39233_3433# a_38861_3013# a_38270_3194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7164 a_30993_n7496# a_31250_n7512# a_29981_n7677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7165 a_39158_n5624# a_38945_n5624# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7166 a_16371_1263# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7167 a_25729_n4391# a_25982_n4595# a_24713_n4760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7168 a_32668_n2470# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7169 gnd a_13844_2687# a_13636_2687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7170 gnd a_40835_1144# a_40627_1144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7171 vdd a_30023_n8205# a_29815_n8205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7172 a_38146_n5805# a_37933_n5805# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7173 a_12191_n2733# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7174 a_13587_2877# a_13801_1755# a_13752_1945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7175 gnd a_31154_6832# a_30946_6832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7176 vdd d0 a_41904_n8499# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7177 a_21971_n9735# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7178 a_3019_n4134# a_3217_n5366# a_3172_n5162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7179 a_4162_1018# a_4158_1195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7180 a_11277_5767# a_11064_5767# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7181 a_16856_n7791# a_16435_n7791# a_16159_n7772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7182 a_23624_n8061# a_23203_n8061# a_23459_n8993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7183 a_23535_6431# a_23114_6431# a_23382_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7184 a_38873_1053# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7185 a_7087_3573# a_6705_4015# a_6114_4196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7186 gnd d4 a_40520_4629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7187 a_16868_n4438# a_16447_n4438# a_16174_n4453# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7188 a_6099_7132# a_5678_7132# a_5402_7032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7189 a_27256_n8318# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7190 gnd d0 a_15040_8286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7191 a_6923_3034# a_6710_3034# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7192 a_1441_1095# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7193 a_26906_5539# a_26904_5325# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7194 a_5995_n5826# a_5782_n5826# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7195 a_429_1276# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7196 a_11161_n5440# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7197 a_7168_n7041# a_6786_n7602# a_6195_n7783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7198 a_16760_7140# a_16339_7140# a_16063_7040# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7199 a_26892_7285# a_26892_7003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7200 a_32286_5568# a_32284_5354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7201 a_2229_n6098# a_3065_n10418# a_2907_n10402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7202 vdd a_8647_8023# a_8439_8023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7203 a_39314_n6843# a_38942_n6600# a_38351_n6781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7204 a_22988_n8573# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7205 a_6202_n5411# a_7007_n5645# a_7176_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7206 a_35297_1355# a_36358_984# a_36313_997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7207 a_39433_n3103# a_39378_n4131# a_39562_n5879# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7208 a_6717_2055# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7209 a_17661_4455# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7210 a_30917_3105# a_31174_2915# a_29905_3286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7211 a_8191_6588# a_8389_7603# a_8344_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7212 a_224_n7018# a_705_n7389# a_913_n7389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7213 a_36365_n9297# a_36361_n9485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7214 vdd d2 a_35588_n3385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7215 a_7062_7371# a_6690_6951# a_6098_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7216 vdd a_29859_4621# a_29651_4621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7217 a_219_n8182# a_217_n7785# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7218 a_28301_n2675# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7219 vdd d3 a_13824_6604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7220 a_35354_n8685# a_36415_n8520# a_36370_n8316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7221 a_8503_n5561# a_8756_n5765# a_8453_n5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7222 a_41679_n2606# a_41936_n2622# a_40667_n2787# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7223 a_616_5759# a_403_5759# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7224 a_25631_4107# a_25888_3917# a_24619_4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7225 a_1907_n3145# a_1793_n3145# a_2001_n3145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7226 a_6113_3781# a_5692_3781# a_5424_3611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7227 gnd d4 a_35328_n6309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7228 a_17452_n6629# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7229 a_6207_n4430# a_5786_n4430# a_5520_n4244# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7230 vdd d0 a_4390_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7231 a_35303_n9058# a_35556_n9262# a_35150_n8030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7232 a_19106_n7106# a_19201_n7730# a_19152_n7714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7233 vdd a_25958_n9908# a_25750_n9908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7234 a_37567_4952# a_37570_4571# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7235 gnd a_8444_6575# a_8236_6575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7236 gnd d0 a_41911_n7520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7237 a_6841_n7041# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7238 a_16440_n6810# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7239 a_7411_n5900# a_7302_n6077# a_7510_n6077# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7240 a_23471_n7033# a_23050_n7033# a_23377_n7033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7241 a_17673_n4672# a_17460_n4672# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7242 a_17911_n9009# a_17868_n8077# a_18076_n8077# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7243 a_1890_n4928# a_1518_n4685# a_927_n4866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7244 a_10814_1466# a_10814_1184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7245 vdd a_19313_7050# a_19105_7050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7246 a_9426_3938# a_9422_4115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7247 a_239_n4265# a_718_n4451# a_926_n4451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7248 vdd a_25905_976# a_25697_976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7249 a_27588_6688# a_27167_6688# a_26894_6904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7250 a_13585_n6134# a_13838_n6338# a_13469_n10410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7251 a_17383_1082# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7252 a_21732_n2858# a_21732_n2576# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7253 a_39049_7911# a_38836_7911# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7254 a_12551_n4936# a_12179_n4693# a_11588_n4874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7255 a_17842_3462# a_17421_3462# a_17748_3581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7256 a_4122_8468# a_4379_8278# a_3113_8057# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7257 a_35166_n4301# a_35423_n4317# a_35071_n6293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7258 a_17564_6959# a_17351_6959# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7259 a_13829_n5358# a_13933_n4813# a_13884_n4797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7260 a_24724_n3593# a_25782_n4031# a_25733_n4015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7261 a_38853_4970# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7262 a_16566_3789# a_16353_3789# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7263 a_35361_n7706# a_36422_n7541# a_36373_n7525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7264 a_33000_840# a_32579_840# a_32313_855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7265 a_19068_5280# a_20129_4909# a_20084_4922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7266 a_29935_n7069# a_30030_n7693# a_29981_n7677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7267 a_11354_n9357# a_11141_n9357# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7268 a_17648_n9570# a_17435_n9570# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7269 a_30993_n7496# a_31003_n6742# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7270 a_29766_n8189# a_29980_n7273# a_29935_n7069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7271 a_3214_n7539# a_4272_n7977# a_4223_n7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7272 a_9435_2570# a_9692_2380# a_8426_2159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7273 vdd d1 a_3391_3146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7274 a_35150_n8030# a_35403_n8234# a_35075_n6105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7275 a_14889_n6988# a_15146_n7004# a_13880_n6566# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7276 a_1837_6460# a_1624_6460# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7277 a_35284_4119# a_36342_4340# a_36297_4353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7278 a_3223_n4789# a_4284_n4624# a_4235_n4608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7279 a_15795_300# a_15582_300# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7280 gnd a_9680_4340# a_9472_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7281 a_16184_n2874# a_16184_n2592# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7282 a_40358_2827# a_40572_1705# a_40527_1718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7283 a_23271_7363# a_23162_7363# a_23370_7363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7284 a_28494_n6592# a_28281_n6592# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7285 a_29695_n6076# a_29948_n6280# a_29579_n10352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7286 a_32304_1155# a_32306_1056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7287 a_934_n3887# a_1738_n3706# a_1907_n3145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7288 a_20526_n805# d9 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7289 a_5500_n8161# a_5979_n8347# a_6187_n8347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7290 a_16077_4981# a_16563_4765# a_16771_4765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7291 a_29701_2642# a_29899_3657# a_29850_3847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7292 gnd d1 a_14148_n3834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7293 a_33864_n8069# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7294 a_237_n3868# a_726_n3887# a_934_n3887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7295 a_25738_n3034# a_25995_n3050# a_24729_n2612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7296 a_5431_2037# a_5917_1821# a_6125_1821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7297 a_17812_n8832# a_17440_n8589# a_16849_n8770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7298 vdd a_40835_1144# a_40627_1144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7299 a_28584_1465# a_28475_1465# a_28683_1465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7300 gnd d0 a_31182_2351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7301 a_25725_n5787# a_25721_n5975# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7302 a_28678_n3095# a_28564_n3095# a_28772_n3095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7303 a_13587_2877# a_13801_1755# a_13756_1768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7304 a_29889_7026# a_30947_7247# a_30902_7260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7305 a_37656_n6381# a_37659_n6000# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7306 a_13469_n10410# a_13630_n6338# a_13585_n6134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7307 vdd d2 a_14086_n5374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7308 a_8504_n4768# a_9565_n4603# a_9520_n4399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7309 a_27464_n9299# a_27251_n9299# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7310 a_7171_n4907# a_7062_n5084# a_7270_n5084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7311 a_38848_5951# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7312 a_32632_n9743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7313 a_23308_1605# a_22926_2047# a_22335_2228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7314 a_33610_7371# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7315 vdd a_41810_7821# a_41602_7821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7316 a_5525_n3080# a_6006_n3451# a_6214_n3451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7317 gnd d0 a_9684_2944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7318 gnd d2 a_19278_3694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7319 gnd d0 a_36534_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7320 a_505_n4451# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7321 a_40612_n3348# a_40716_n2803# a_40667_n2787# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7322 vdd d0 a_15040_8286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7323 a_850_1276# a_429_1276# a_153_1458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7324 vdd a_4391_6318# a_4183_6318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7325 a_29854_3670# a_30107_3657# a_29701_2642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7326 a_24569_3868# a_24673_3117# a_24628_3130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7327 vdd d0 a_25977_n5576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7328 gnd a_36541_5882# a_36333_5882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7329 a_33649_n8581# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7330 a_21695_n9716# a_22184_n9735# a_22392_n9735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7331 a_16786_1829# a_16365_1829# a_16097_1659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7332 a_23283_5403# a_22911_4983# a_22319_4749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7333 a_23228_n3677# a_23015_n3677# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7334 a_35242_1916# a_35346_1165# a_35297_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7335 gnd d0 a_4378_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7336 vdd a_31162_6268# a_30954_6268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7337 a_3145_2180# a_4203_2401# a_4154_2591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7338 a_29579_n10352# a_29740_n6280# a_29695_n6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7339 a_24604_7224# a_25665_6853# a_25616_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7340 a_30981_n9456# a_30991_n8702# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7341 a_32976_6153# a_32555_6153# a_32279_6335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7342 a_28569_5501# a_28187_5943# a_27595_5709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7343 gnd d1 a_35626_n5765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7344 a_3130_5116# a_4188_5337# a_4139_5527# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7345 vdd a_8444_6575# a_8236_6575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7346 a_8511_n3789# a_9572_n3624# a_9523_n3608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7347 gnd d0 a_9692_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7348 a_13859_n9695# a_14920_n9530# a_14871_n9514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7349 a_14893_n6800# a_14889_n6988# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7350 a_22397_n8754# a_23201_n8573# a_23360_n8816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7351 a_24397_n10373# a_24347_n10389# a_23719_n6069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7352 a_37637_n9421# a_37639_n9322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7353 a_22127_2228# a_21914_2228# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7354 a_34132_n7041# a_33711_n7041# a_34038_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7355 gnd d0 a_9677_5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7356 a_36373_n7525# a_36383_n6771# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7357 vdd d1 a_3492_n2845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7358 a_13756_1768# a_13851_2175# a_13802_2365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7359 a_5416_5568# a_5897_5738# a_6105_5738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7360 a_9517_n5002# a_9520_n4399# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7361 gnd d0 a_15044_6890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7362 a_40580_n9225# a_40684_n8680# a_40639_n8476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7363 a_40584_n9037# a_40837_n9241# a_40431_n8009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7364 gnd a_9753_n8520# a_9545_n8520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7365 a_16647_n7376# a_16434_n7376# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7366 a_11159_n6831# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7367 vdd a_31239_n9887# a_31031_n9887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7368 a_33805_1074# a_33592_1074# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7369 a_35214_7616# a_35467_7603# a_35061_6588# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7370 a_39150_n7581# a_38937_n7581# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7371 a_32760_6717# a_32547_6717# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7372 a_12791_n5929# a_12682_n6106# a_12890_n6106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7373 a_1421_5012# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7374 a_698_n8368# a_485_n8368# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7375 a_11302_869# a_11089_869# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7376 a_24397_n10373# a_26746_n10456# a_26588_n10440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7377 a_8394_8036# a_9452_8257# a_9407_8270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7378 a_5486_n9724# a_5486_n9442# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7379 a_27485_n5797# a_27272_n5797# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7380 a_36394_n4023# a_36651_n4039# a_35385_n3601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7381 a_36313_997# a_36309_1174# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7382 vdd a_3336_3707# a_3128_3707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7383 gnd d0 a_15141_n7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7384 a_6794_n5645# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7385 a_10891_n4573# a_10893_n4474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7386 a_41655_n7919# a_41658_n7316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7387 gnd d5 a_8346_n10397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7388 a_27609_3186# a_27188_3186# a_26912_3086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7389 a_32554_5738# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7390 a_41647_n8483# a_41659_n7731# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7391 a_4210_n9506# a_4220_n8752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7392 a_11575_n7812# a_12379_n7631# a_12548_n7070# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7393 a_39344_1473# a_39289_2501# a_39473_4426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7394 a_224_n6423# a_227_n6042# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7395 gnd a_24982_n2816# a_24774_n2816# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7396 a_19160_n5757# a_19417_n5773# a_19114_n5149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7397 a_1649_2076# a_1436_2076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7398 a_28564_5382# a_28192_4962# a_27601_5143# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7399 a_12593_4476# a_12380_4476# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7400 a_1946_n4173# a_1733_n4173# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7401 a_25632_4906# a_25628_5083# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7402 a_22412_n5818# a_21991_n5818# a_21715_n5799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7403 a_14815_2599# a_15072_2409# a_13806_2188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7404 a_130_5975# a_616_5759# a_824_5759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7405 a_9424_5329# a_9420_5506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7406 vdd a_9680_4340# a_9472_4340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7407 a_16860_n6395# a_16439_n6395# a_16166_n6410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7408 a_40447_n4280# a_40704_n4296# a_40352_n6272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7409 a_28663_5382# a_28608_6410# a_28816_6410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7410 a_38937_n7581# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7411 a_423_1842# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7412 a_40642_n7685# a_41703_n7520# a_41654_n7504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7413 a_28651_7342# a_28230_7342# a_28557_7461# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7414 a_27269_n6773# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7415 a_31019_n3013# a_31276_n3029# a_30010_n2591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7416 a_30905_6458# a_30908_5866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7417 a_16147_n9732# a_16636_n9751# a_16844_n9751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7418 a_17655_n8077# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7419 a_28331_n7012# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7420 a_28901_n5871# a_28792_n6048# a_29000_n6048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7421 a_20170_n6967# a_20427_n6983# a_19161_n6545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7422 vdd d0 a_31182_2351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7423 a_28415_2493# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7424 a_23380_n4899# a_23008_n4656# a_22417_n4837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7425 a_23107_7924# a_22894_7924# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7426 a_20848_n805# a_21446_n10615# a_10498_n10484# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7427 a_17750_n6085# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7428 a_39339_n3103# a_39225_n3103# a_39433_n3103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7429 a_34195_359# a_33982_359# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7430 a_8419_3138# a_9477_3359# a_9428_3549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7431 a_31003_n6742# a_31256_n6946# a_29990_n6508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7432 a_27685_n7754# a_28489_n7573# a_28658_n7012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7433 a_36381_n5568# a_36638_n5584# a_35369_n5749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7434 a_11270_6746# a_11057_6746# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7435 a_4231_n6004# a_4488_n6020# a_3222_n5582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7436 a_20104_1005# a_20100_1182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7437 a_28420_2026# a_28207_2026# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7438 vdd a_25962_n8512# a_25754_n8512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7439 vdd d0 a_20353_2388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7440 a_1793_n3145# a_1580_n3145# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7441 a_17614_7379# a_17401_7379# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7442 gnd a_35479_5643# a_35271_5643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7443 a_27393_5143# a_27180_5143# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7444 a_11064_5767# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7445 a_8352_5833# a_8456_5082# a_8407_5272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7446 gnd d0 a_36619_n9916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7447 a_10804_3045# a_11290_2829# a_11498_2829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7448 a_9533_n2854# a_9529_n3042# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7449 a_31952_n2202# a_32881_n2470# a_33089_n2470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7450 a_9415_6487# a_9672_6297# a_8406_6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7451 a_33053_n9743# a_33857_n9562# a_34026_n9001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7452 a_6987_n9562# a_6774_n9562# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7453 a_22094_7690# a_21881_7690# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7454 a_6710_3034# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7455 a_12568_n3153# a_12186_n3714# a_11595_n3895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7456 a_35242_1916# a_35346_1165# a_35301_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7457 a_26924_1408# a_27413_1226# a_27621_1226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7458 a_35366_n6725# a_35623_n6741# a_35311_n7286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7459 gnd d0 a_25900_1957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7460 a_22308_7124# a_23112_6943# a_23271_7363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7461 vdd a_4479_n7562# a_4271_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7462 a_9420_5506# a_9423_4914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7463 a_5766_n8347# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7464 vdd a_19007_n10405# a_18799_n10405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7465 a_34403_359# a_37285_271# a_31994_256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7466 a_4137_5916# a_4390_5903# a_3121_6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7467 vdd d0 a_9692_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7468 a_32548_7132# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7469 a_19140_n9674# a_20201_n9509# a_20152_n9493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7470 a_16881_n2893# a_16460_n2893# a_16184_n2592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7471 vdd a_13824_6604# a_13616_6604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7472 a_28564_5382# a_28455_5382# a_28663_5382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7473 a_20087_3946# a_20083_4123# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7474 a_32567_2800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7475 a_29602_4811# a_29746_2629# a_29701_2642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7476 vdd d0 a_9677_5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7477 a_403_5759# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7478 a_36285_6487# a_36288_5895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7479 a_37570_4571# a_37568_4357# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7480 a_21628_3989# a_21633_3603# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7481 a_13756_1768# a_13851_2175# a_13806_2188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7482 a_19110_n5337# a_19367_n5353# a_18961_n4121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7483 gnd a_35239_4650# a_35031_4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7484 gnd d1 a_40907_n5744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7485 a_4158_1195# a_4415_1005# a_3146_1376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7486 a_5793_n3451# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7487 a_28678_n3095# a_28296_n3656# a_27705_n3837# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7488 vdd d2 a_3417_n7323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7489 a_27407_1792# a_27194_1792# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7490 a_6953_7371# a_6740_7371# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7491 gnd d2 a_19258_7611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7492 a_30902_7260# a_31155_7247# a_29889_7026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7493 gnd a_13989_5672# a_13781_5672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7494 gnd d0 a_31244_n8906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7495 a_30897_8241# a_32267_8295# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7496 a_39158_n5624# a_38945_n5624# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7497 gnd a_19434_n2832# a_19226_n2832# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7498 a_17829_n7049# a_17447_n7610# a_16856_n7791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7499 a_38054_5151# a_37841_5151# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7500 a_16063_7322# a_16063_7040# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7501 a_38836_7911# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7502 a_29904_4090# a_30157_4077# a_29854_3670# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7503 a_38146_n5805# a_37933_n5805# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7504 a_12191_n2733# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7505 a_24708_n5741# a_25769_n5576# a_25724_n5372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7506 a_18095_367# a_17986_367# a_15904_300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7507 a_10777_8042# a_10779_7943# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7508 a_17834_5419# a_17413_5419# a_17735_5419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7509 a_12573_1523# a_12152_1523# a_12479_1642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7510 a_21971_n9735# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7511 a_37654_n6480# a_38143_n6781# a_38351_n6781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7512 a_5697_2800# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7513 a_17351_6959# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7514 gnd d0 a_41831_4319# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7515 a_34046_n5084# a_33664_n5645# a_33073_n5826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7516 a_907_n8783# a_486_n8783# a_210_n8482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7517 gnd d0 a_36567_1399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7518 a_22314_5730# a_21893_5730# a_21625_5560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7519 a_16353_3789# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7520 a_27588_6688# a_28393_6922# a_28552_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7521 a_13864_n8714# a_14121_n8730# a_13809_n9275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7522 gnd d0 a_31271_n4010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7523 a_22428_n2462# a_22007_n2462# a_21734_n2477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7524 a_23531_4439# a_23134_2514# a_23402_1486# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7525 a_35323_n5141# a_35418_n5765# a_35369_n5749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7526 a_21606_8005# a_22095_8105# a_22303_8105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7527 a_37651_n7362# a_37656_n6976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7528 a_7168_n7041# a_6786_n7602# a_6194_n7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7529 a_11579_n6416# a_11158_n6416# a_10885_n6431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7530 a_11077_2829# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7531 a_1624_6460# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7532 gnd d1 a_40810_6042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7533 gnd d0 a_20422_n7964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7534 gnd a_20430_n6007# a_20222_n6007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7535 gnd a_36655_n2643# a_36447_n2643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7536 a_22988_n8573# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7537 a_6203_n5826# a_7007_n5645# a_7176_n5084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7538 a_26733_263# a_26624_263# a_26832_263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7539 a_10900_n4273# a_11379_n4459# a_11587_n4459# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7540 gnd a_30263_n2795# a_30055_n2795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7541 a_22339_832# a_21918_832# a_21652_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7542 a_3230_n3810# a_3487_n3826# a_3184_n3202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7543 a_24713_n4760# a_24970_n4776# a_24658_n5321# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7544 a_33070_n6802# a_32649_n6802# a_32373_n6783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7545 a_913_n7389# a_1718_n7623# a_1887_n7062# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7546 a_28301_n2675# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7547 a_16090_2144# a_16579_2244# a_16787_2244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7548 a_7302_n6077# a_7089_n6077# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7549 a_29978_n8468# a_31036_n8906# a_30991_n8702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7550 a_23291_3446# a_22919_3026# a_22328_3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7551 a_617_6174# a_404_6174# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7552 a_32370_n7383# a_32856_n7368# a_33064_n7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7553 a_33785_4991# a_33572_4991# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7554 a_833_4217# a_1637_4036# a_1806_3594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7555 a_12469_n6106# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7556 a_3214_n7539# a_3467_n7743# a_3164_n7119# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7557 a_17346_7940# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7558 gnd d6 a_15917_n10493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7559 a_2045_6460# a_1932_4468# a_2140_4468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7560 vdd a_35479_5643# a_35271_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7561 gnd d1 a_19414_n6749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7562 gnd a_3475_n5786# a_3267_n5786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7563 a_30001_n3760# a_31062_n3595# a_31017_n3391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7564 a_20088_3142# a_20100_2401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7565 vdd a_4384_7297# a_4176_7297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7566 a_8352_5833# a_8456_5082# a_8411_5095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7567 a_39401_n8980# a_38980_n8980# a_39302_n8803# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7568 a_232_n4466# a_718_n4451# a_926_n4451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7569 a_28577_3544# a_28195_3986# a_27604_4167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7570 a_13875_n7547# a_14933_n7985# a_14884_n7969# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7571 a_14807_4382# a_14803_4559# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7572 a_27689_n6358# a_27268_n6358# a_26995_n6373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7573 a_12384_n6650# a_12171_n6650# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7574 a_40511_3855# a_40615_3104# a_40566_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7575 a_3148_n9267# a_3405_n9283# a_2999_n8051# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7576 a_28284_n5616# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7577 a_27589_7103# a_27168_7103# a_26892_7003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7578 vdd a_3386_4127# a_3178_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7579 gnd a_19278_3694# a_19070_3694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7580 gnd d0 a_4480_n7977# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7581 a_22931_1066# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7582 gnd a_30169_2117# a_29961_2117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7583 gnd a_36534_6861# a_36326_6861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7584 a_1629_5993# a_1416_5993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7585 a_41662_n5547# a_41919_n5563# a_40650_n5728# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7586 a_41574_4509# a_41831_4319# a_40565_4098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7587 a_23436_n4144# a_23223_n4144# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7588 a_16668_n3874# a_16455_n3874# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7589 gnd d0 a_4492_n4624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7590 gnd d2 a_40857_n5324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7591 a_39477_6418# a_39056_6418# a_39324_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7592 vdd a_31243_n8491# a_31035_n8491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7593 a_5677_6717# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7594 a_8491_n7706# a_8748_n7722# a_8445_n7098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7595 gnd d2 a_8698_n7302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7596 gnd a_9766_n6975# a_9558_n6975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7597 a_33057_n8347# a_32636_n8347# a_32363_n8362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7598 a_32299_2418# a_32788_2236# a_32996_2236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7599 gnd d0 a_41900_n9895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7600 a_28552_7342# a_28180_6922# a_27588_6688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7601 a_10868_n9372# a_10873_n8986# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7602 a_20173_n5991# a_20430_n6007# a_19164_n5569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7603 a_11354_n9357# a_11141_n9357# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7604 a_14892_n6385# a_15145_n6589# a_13876_n6754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7605 a_28579_n6048# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7606 gnd a_4378_7863# a_4170_7863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7607 a_29985_n7489# a_31043_n7927# a_30994_n7911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7608 a_4231_n6377# a_4227_n6565# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7609 a_33870_4447# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7610 a_27603_3752# a_27182_3752# a_26914_3582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7611 a_20176_n5388# a_20172_n5576# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7612 gnd d1 a_30243_n6712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7613 vdd d0 a_15071_1994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7614 a_3079_3897# a_3183_3146# a_3134_3336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7615 a_39012_n3103# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7616 a_22120_3207# a_21907_3207# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7617 a_38157_n3430# a_37944_n3430# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7618 a_36297_3134# a_36554_2944# a_35285_3315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7619 a_1806_3594# a_1692_3475# a_1900_3475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7620 a_22327_2792# a_21906_2792# a_21633_3008# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7621 vdd a_35239_4650# a_35031_4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7622 a_16149_n9946# a_20410_n9924# a_19144_n9486# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7623 a_1857_2543# a_1644_2543# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7624 a_5493_n8362# a_5979_n8347# a_6187_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7625 a_16787_2244# a_17591_2063# a_17760_1621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7626 a_33889_n3685# a_33676_n3685# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7627 vdd d2 a_19258_7611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7628 vdd a_13989_5672# a_13781_5672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7629 a_35170_n4113# a_35368_n5345# a_35319_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7630 a_33084_n3451# a_32663_n3451# a_32390_n3466# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7631 a_41642_n9464# a_41652_n8710# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7632 a_16428_n8770# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7633 gnd a_24667_n6301# a_24459_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7634 a_28697_n8040# a_28484_n8040# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7635 a_23283_n3116# a_23070_n3116# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7636 a_4141_4136# a_4398_3946# a_3129_4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7637 a_35353_n9478# a_36411_n9916# a_36362_n9900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7638 a_19017_5664# a_19270_5651# a_18848_6773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7639 gnd d1 a_3455_n9703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7640 a_14872_n9929# a_15129_n9945# a_13863_n9507# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7641 vdd d0 a_25885_4893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7642 a_32668_n2470# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7643 a_25612_8439# a_25869_8249# a_24603_8028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7644 gnd a_15044_6890# a_14836_6890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7645 gnd a_19359_n7310# a_19151_n7310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7646 a_20084_4538# a_20341_4348# a_19075_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7647 a_33592_1074# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7648 a_14803_4559# a_14806_3967# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7649 a_32632_n9743# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7650 a_28477_n9533# a_28264_n9533# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7651 a_4143_5350# a_4139_5527# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7652 a_12462_3483# a_12353_3483# a_12561_3483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7653 a_40582_1157# a_40835_1144# a_40523_1895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7654 a_13591_2700# a_13844_2687# a_13492_4869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7655 a_1642_3055# a_1429_3055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7656 a_5520_n3466# a_6006_n3451# a_6214_n3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7657 vdd a_35403_n8234# a_35195_n8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7658 a_3215_n6746# a_4276_n6581# a_4231_n6377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7659 a_1882_n6885# a_1773_n7062# a_1981_n7062# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7660 a_40553_6232# a_41614_5861# a_41569_5874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7661 a_4235_n4608# a_4492_n4624# a_3223_n4789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7662 a_38370_n2449# a_39175_n2683# a_39334_n2926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7663 a_38868_2034# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7664 a_27256_n8318# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7665 a_19021_3884# a_19125_3133# a_19076_3323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7666 a_25742_n2846# a_25738_n3034# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7667 vdd d1 a_40810_6042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7668 a_1436_2076# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7669 a_32963_7698# a_33768_7932# a_33937_7490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7670 a_12380_4476# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7671 a_6918_4015# a_6705_4015# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7672 a_33862_n8581# a_33649_n8581# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7673 a_6131_1255# a_5710_1255# a_5434_1437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7674 a_41569_5874# a_41565_6051# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7675 a_23479_n5076# a_23058_n5076# a_23380_n4899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7676 vdd a_4411_2401# a_4203_2401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7677 gnd a_20447_n3066# a_20239_n3066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7678 a_16755_8121# a_16334_8121# a_16058_8303# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7679 a_14807_3163# a_15064_2973# a_13795_3344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7680 a_13736_5685# a_13831_6092# a_13786_6105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7681 a_38249_6696# a_37828_6696# a_37555_6912# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7682 a_12814_388# a_13541_4679# a_13492_4869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7683 a_6195_n7783# a_5774_n7783# a_5498_n7764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7684 a_38853_4970# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7685 a_37664_n5019# a_38145_n5390# a_38353_n5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7686 vdd a_4500_n4060# a_4292_n4060# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7687 a_26996_n5496# a_26998_n5397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7688 a_27583_7669# a_27162_7669# a_26889_7885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7689 gnd d0 a_4398_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7690 a_29905_3286# a_30966_2915# a_30921_2928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7691 gnd a_40748_7582# a_40540_7582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7692 a_37565_5333# a_38054_5151# a_38262_5151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7693 a_8441_n7286# a_8698_n7302# a_8276_n8218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7694 a_6207_n4430# a_5786_n4430# a_5513_n4445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7695 a_27283_n3422# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7696 a_6903_6951# a_6690_6951# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7697 a_36370_n8316# a_36623_n8520# a_35354_n8685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7698 a_3121_6274# a_4182_5903# a_4137_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7699 vdd d2 a_24907_n7294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7700 a_5429_2136# a_5431_2037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7701 a_29978_n8468# a_30231_n8672# a_29919_n9217# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7702 a_14904_n4052# a_14907_n3449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7703 vdd d1 a_30162_3096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7704 a_36296_3938# a_36292_4115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7705 a_14896_n4616# a_14908_n3864# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7706 a_14908_n3864# a_15161_n4068# a_13895_n3630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7707 a_2252_380# a_1831_380# a_2140_4468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7708 a_37568_4075# a_37570_3976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7709 a_17584_3042# a_17371_3042# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7710 a_5905_3781# a_5692_3781# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7711 a_25717_n7744# a_25713_n7932# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7712 gnd d0 a_41835_2923# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7713 a_16766_5746# a_17571_5980# a_17740_5538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7714 gnd d5 a_3065_n10418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7715 a_6697_5972# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7716 a_9407_8270# a_9403_8447# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7717 a_7421_4447# a_7000_4447# a_7322_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7718 a_16655_n5419# a_16442_n5419# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7719 gnd d1 a_40899_n7701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7720 a_5409_6335# a_5898_6153# a_6106_6153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7721 vdd a_20353_2388# a_20145_2388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7722 gnd d0 a_36547_5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7723 a_16647_n7376# a_16434_n7376# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7724 gnd a_4505_n3079# a_4297_n3079# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7725 a_17378_2063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7726 a_32267_8013# a_32269_7914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7727 a_17401_7379# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7728 a_27180_5143# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7729 vdd d0 a_20345_2952# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7730 a_21898_4749# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7731 a_4139_5527# a_4142_4935# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7732 a_26983_n8928# a_26981_n8714# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7733 a_33932_7371# a_33823_7371# a_34031_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7734 vdd d1 a_35618_n7722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7735 a_9407_7051# a_9664_6861# a_8395_7232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7736 gnd a_35423_n4317# a_35215_n4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7737 vdd a_15166_n3087# a_14958_n3087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7738 a_25709_n8308# a_25705_n8496# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7739 gnd d0 a_20340_3933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7740 a_6794_n5645# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7741 a_24485_n8210# a_24742_n8226# a_24414_n6097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7742 vdd a_3183_2679# a_2975_2679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7743 a_28653_n6835# a_28544_n7012# a_28752_n7012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7744 a_30917_3105# a_30929_2364# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7745 a_9523_n3608# a_9780_n3624# a_8511_n3789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7746 a_3079_3897# a_3183_3146# a_3138_3159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7747 a_1505_n7623# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7748 a_2924_n6126# a_3177_n6330# a_2808_n10402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7749 a_7094_1494# a_6722_1074# a_6130_840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7750 a_2044_380# a_1831_380# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7751 a_13871_n7735# a_14128_n7751# a_13825_n7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7752 a_5243_292# a_7112_359# a_7421_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7753 a_155_1077# a_641_861# a_849_861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7754 gnd d0 a_25886_5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7755 a_2134_n8090# a_2021_n6098# a_2229_n6098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7756 a_32356_n9724# a_32356_n9442# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7757 vdd a_14136_n5794# a_13928_n5794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7758 a_7112_359# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7759 a_8364_3699# a_8459_4106# a_8414_4119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7760 a_20173_n6364# a_20426_n6568# a_19157_n6733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7761 gnd d0 a_31162_6268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7762 a_7181_3454# a_6760_3454# a_7082_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7763 a_31885_256# a_31672_256# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7764 a_26906_5539# a_27387_5709# a_27595_5709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7765 a_3168_n5350# a_3272_n4805# a_3223_n4789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7766 gnd a_20434_n4611# a_20226_n4611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7767 a_27692_n5382# a_27271_n5382# a_26998_n5397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7768 a_19013_5841# a_19270_5651# a_18848_6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7769 a_23380_n4899# a_23008_n4656# a_22416_n4422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7770 a_32306_1056# a_32313_855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7771 a_20184_n3616# a_20194_n2862# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7772 a_16152_n8469# a_16154_n8370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7773 a_8201_n6293# a_8458_n6309# a_8089_n10381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7774 gnd d0 a_15057_5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7775 a_27194_1792# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7776 a_17755_1502# a_17383_1082# a_16792_1263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7777 gnd a_19258_7611# a_19050_7611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7778 a_8410_4296# a_9471_3925# a_9426_3938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7779 a_33843_3454# a_33630_3454# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7780 a_9403_8447# a_9406_7855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7781 a_40578_1334# a_40835_1144# a_40523_1895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7782 a_39138_n9541# a_38925_n9541# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7783 a_40451_n4092# a_40649_n5324# a_40600_n5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7784 a_8112_4840# a_8256_2658# a_8207_2848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7785 gnd d3 a_3252_n8255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7786 a_31002_n5954# a_31259_n5970# a_29993_n5532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7787 a_19021_3884# a_19125_3133# a_19080_3146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7788 vdd d0 a_41847_963# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7789 a_11505_1850# a_11084_1850# a_10811_2066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7790 a_5436_1056# a_5922_840# a_6130_840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7791 a_10883_n6530# a_10885_n6431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7792 gnd a_36567_1399# a_36359_1399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7793 a_41654_n7504# a_41911_n7520# a_40642_n7685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7794 vdd a_9676_4901# a_9468_4901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7795 a_6987_n9562# a_6774_n9562# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7796 gnd a_35499_1726# a_35291_1726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7797 a_11491_5201# a_12295_5020# a_12454_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7798 a_6182_n9328# a_5761_n9328# a_5493_n8957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7799 a_25647_1970# a_25643_2147# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7800 a_5422_3115# a_5911_3215# a_6119_3215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7801 a_16848_n8355# a_16427_n8355# a_16154_n8370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7802 a_12568_n3153# a_12186_n3714# a_11594_n3480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7803 a_711_n6823# a_498_n6823# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7804 gnd d2 a_40849_n7281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7805 gnd d0 a_25975_n6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7806 a_16672_n2478# a_16459_n2478# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7807 a_5766_n8347# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7808 a_11141_n9357# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7809 vdd d3 a_8533_n8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7810 a_32850_n8762# a_32637_n8762# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7811 vdd a_40919_n3784# a_40711_n3784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7812 gnd d0 a_9672_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7813 a_18773_4848# a_19030_4658# a_18095_367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7814 a_1875_n9022# a_1493_n9583# a_902_n9764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7815 a_26904_5325# a_26904_5043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7816 a_39205_n7020# a_38992_n7020# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7817 vdd a_40748_7582# a_40540_7582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7818 vdd d1 a_8768_n3805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7819 a_610_7153# a_397_7153# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7820 a_22099_6709# a_21886_6709# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7821 a_32284_5354# a_32284_5072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7822 a_40639_n8476# a_41697_n8914# a_41648_n8898# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7823 vdd d1 a_14116_n9711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7824 a_13568_n10410# a_13518_n10426# a_13469_n10410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7825 a_12229_n5113# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7826 a_38073_819# a_37860_819# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7827 a_9495_n9297# a_9748_n9501# a_8479_n9666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7828 a_36385_n5380# a_36381_n5568# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7829 a_4157_1999# a_4410_1986# a_3141_2357# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7830 gnd a_15160_n3653# a_14952_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7831 a_29880_8184# a_30137_7994# a_29834_7587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7832 a_32568_3215# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7833 gnd d1 a_24945_n9674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7834 a_404_6174# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7835 a_33572_4991# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7836 a_11285_3810# a_11072_3810# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7837 a_141_3418# a_630_3236# a_838_3236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7838 a_21697_n9335# a_22183_n9320# a_22391_n9320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7839 a_8465_n3181# a_8560_n3805# a_8511_n3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7840 a_5520_n3466# a_5525_n3080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7841 a_26996_n5778# a_26996_n5496# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7842 vdd d0 a_36547_5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7843 a_5793_n3451# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7844 a_29842_5804# a_29946_5053# a_29897_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7845 a_35146_n8218# a_35360_n7302# a_35311_n7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7846 a_28678_n3095# a_28296_n3656# a_27704_n3422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7847 vdd d2 a_30188_n7273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7848 gnd a_25869_8249# a_25661_8249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7849 a_38962_n2683# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7850 gnd d0 a_9785_n2643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7851 a_41595_1391# a_41591_1568# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7852 vdd a_14086_n5374# a_13878_n5374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7853 a_20189_n3843# a_20442_n4047# a_19176_n3609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7854 a_35301_1178# a_36359_1399# a_36314_1412# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7855 a_698_n8368# a_485_n8368# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7856 gnd a_14009_1755# a_13801_1755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7857 a_32755_7698# a_32542_7698# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7858 a_1416_5993# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7859 a_20084_4922# a_20337_4909# a_19068_5280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7860 vdd a_36619_n9916# a_36411_n9916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7861 a_22423_n3443# a_23228_n3677# a_23397_n3116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7862 a_14802_4144# a_14812_3401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7863 a_28339_n5055# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7864 a_12442_n5113# a_12229_n5113# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7865 gnd d2 a_14098_n3414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7866 a_14787_7080# a_15044_6890# a_13775_7261# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7867 a_34046_n5084# a_33664_n5645# a_33072_n5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7868 a_25627_5887# a_25880_5874# a_24611_6245# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7869 vdd d0 a_41843_2359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7870 vdd d0 a_36650_n3624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7871 a_36387_n5002# a_36390_n4399# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7872 vdd d0 a_36561_1965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7873 gnd d1 a_19325_5090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7874 a_25713_n7932# a_25970_n7948# a_24704_n7510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7875 a_624_3802# a_411_3802# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7876 a_22428_n2462# a_22007_n2462# a_21123_n2239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7877 a_6119_3215# a_6923_3034# a_7082_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7878 a_7156_n9001# a_7042_n9001# a_7250_n9001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7879 a_26993_n6754# a_26993_n6472# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7880 a_4242_n3629# a_4499_n3645# a_3230_n3810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7881 a_38903_5390# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7882 a_23402_1486# a_22981_1486# a_23303_1486# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7883 a_5493_n8957# a_5491_n8743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7884 vdd a_20447_n3066# a_20239_n3066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7885 a_13806_2188# a_14864_2409# a_14819_2422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7886 a_11579_n6416# a_11158_n6416# a_10888_n6050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7887 a_725_n3472# a_512_n3472# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7888 a_16780_3223# a_17584_3042# a_17743_3462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7889 a_16771_4765# a_16350_4765# a_16077_4981# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7890 a_11078_3244# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7891 a_8479_n9666# a_9540_n9501# a_9495_n9297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7892 gnd d4 a_40609_n6288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7893 a_25717_n6536# a_25725_n5787# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7894 gnd d3 a_8553_n4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7895 a_14903_n3637# a_15160_n3653# a_13891_n3818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7896 a_30001_n3760# a_30258_n3776# a_29955_n3152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7897 a_33070_n6802# a_32649_n6802# a_32373_n6501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7898 a_914_n7804# a_1718_n7623# a_1887_n7062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7899 vdd d0 a_15057_5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7900 a_480_n9349# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7901 a_27620_811# a_27199_811# a_26933_826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7902 vdd a_19258_7611# a_19050_7611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7903 a_6000_n4845# a_5787_n4845# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7904 vdd a_4504_n2664# a_4296_n2664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7905 vdd a_40869_n3364# a_40661_n3364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7906 gnd a_25995_n3050# a_25787_n3050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7907 a_17703_n9009# a_17490_n9009# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7908 a_5986_n7368# a_5773_n7368# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7909 a_829_4778# a_408_4778# a_138_4613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7910 a_16072_6557# a_16070_6343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7911 a_22112_5164# a_21899_5164# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7912 a_11265_7727# a_11052_7727# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7913 gnd a_8609_5643# a_8401_5643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7914 a_36282_7289# a_36535_7276# a_35269_7055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7915 a_210_n8482# a_212_n8383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7916 a_16848_n8355# a_17653_n8589# a_17812_n8832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7917 a_36383_n6771# a_36636_n6975# a_35370_n6537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7918 a_38861_3013# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7919 vdd a_41912_n7935# a_41704_n7935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7920 vdd d2 a_14066_n9291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7921 gnd a_30246_n5736# a_30038_n5736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7922 a_21729_n3458# a_21734_n3072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7923 a_25700_n9477# a_25957_n9493# a_24688_n9658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7924 a_34959_n10381# a_35120_n6309# a_35071_n6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7925 a_35284_4119# a_35537_4106# a_35234_3699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7926 vdd d0 a_31275_n2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7927 a_417_3236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7928 a_28284_n5616# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7929 a_27388_6124# a_27175_6124# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7930 vdd a_35499_1726# a_35291_1726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7931 a_21397_n10599# a_31938_n10471# a_26588_n10440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7932 a_21643_1147# a_22132_1247# a_22340_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7933 a_36290_5506# a_36293_4914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7934 a_27697_n4401# a_28502_n4635# a_28661_n4878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7935 a_16668_n3874# a_16455_n3874# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7936 a_1808_n6098# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7937 a_4126_8291# a_4379_8278# a_3113_8057# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7938 a_6705_4015# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7939 a_21717_n6013# a_22200_n6379# a_22408_n6379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7940 gnd d0 a_31166_4872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7941 vout a_20526_n805# a_20853_n686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7942 a_5678_7132# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7943 vdd a_41925_n4997# a_41717_n4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7944 a_33057_n8347# a_32636_n8347# a_32370_n8161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7945 a_16875_n3459# a_17680_n3693# a_17849_n3132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7946 a_38256_5717# a_37835_5717# a_37567_5547# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7947 a_16104_863# a_16583_848# a_16791_848# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7948 a_11595_n3895# a_11174_n3895# a_10898_n3876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7949 vdd a_9769_n5999# a_9561_n5999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7950 a_12367_n9591# a_12154_n9591# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7951 a_36403_n2854# a_36399_n3042# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7952 gnd d0 a_36618_n9501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7953 a_19176_n3609# a_19429_n3813# a_19126_n3189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7954 a_28242_5382# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7955 vdd d3 a_24762_n4309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7956 a_24725_n2800# a_25786_n2635# a_25741_n2431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7957 a_16759_6725# a_17564_6959# a_17723_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7958 gnd a_4398_3946# a_4190_3946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7959 a_23719_n6069# a_24555_n10389# a_24397_n10373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7960 a_6690_6951# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7961 a_23535_6431# a_23422_4439# a_23630_4439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7962 vdd d3 a_13913_n8263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7963 a_1926_n8090# a_1713_n8090# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7964 vdd a_30162_3096# a_29954_3096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7965 a_13567_6794# a_13824_6604# a_13496_4692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7966 a_29842_5804# a_29946_5053# a_29901_5066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7967 a_14792_7318# a_15045_7305# a_13779_7084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7968 a_6188_n8762# a_6992_n8581# a_7151_n8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7969 a_17371_3042# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7970 a_5692_3781# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7971 vdd d0 a_4484_n6581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7972 a_33084_n3451# a_32663_n3451# a_32395_n3080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7973 gnd a_41835_2923# a_41627_2923# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7974 a_37657_n5504# a_37659_n5405# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7975 gnd d3 a_24742_n8226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7976 a_14875_n9326# a_15128_n9530# a_13859_n9695# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7977 a_3184_n3202# a_3279_n3826# a_3230_n3810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7978 a_35226_5656# a_35321_6063# a_35272_6253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7979 gnd a_20441_n3632# a_20233_n3632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7980 vdd d1 a_3472_n6762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7981 a_34192_4447# a_33795_2522# a_34063_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7982 gnd d1 a_35542_3125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7983 vdd a_14009_1755# a_13801_1755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7984 gnd d1 a_30226_n9653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7985 gnd d0 a_4399_4361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7986 a_6220_n2885# a_5799_n2885# a_5523_n2584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7987 gnd a_36547_5316# a_36339_5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7988 a_13736_5685# a_13989_5672# a_13567_6794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7989 gnd d0 a_4468_n9937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7990 a_29889_7026# a_30947_7247# a_30898_7437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7991 vdd a_20345_2952# a_20137_2952# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7992 vdd d2 a_24826_3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7993 a_28477_n9533# a_28264_n9533# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7994 a_20161_n8324# a_20157_n8512# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7995 a_11173_n3480# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7996 gnd d0 a_9676_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7997 a_40427_n8197# a_40641_n7281# a_40592_n7265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7998 gnd a_35549_2146# a_35341_2146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7999 a_30994_n7911# a_31251_n7927# a_29985_n7489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8000 a_24709_n6529# a_25767_n6967# a_25718_n6951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8001 a_23162_7363# a_22949_7363# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8002 gnd a_3460_n8722# a_3252_n8722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8003 a_5506_n5807# a_5506_n5525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8004 a_25730_n4806# a_25983_n5010# a_24717_n4572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8005 a_31006_n4558# a_31263_n4574# a_29994_n4739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8006 gnd a_24673_2650# a_24465_2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8007 vdd a_24881_3117# a_24673_3117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8008 a_10868_n9967# a_14872_n9929# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8009 a_23365_n8993# a_22983_n9554# a_22392_n9735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8010 a_41675_n4002# a_41678_n3399# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8011 gnd a_4391_6318# a_4183_6318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8012 a_24569_3868# a_24673_3117# a_24624_3307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8013 a_13813_n9087# a_13908_n9711# a_13863_n9507# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8014 a_244_n2506# gnd SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8015 a_32776_4196# a_32563_4196# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8016 a_19140_n9674# a_19397_n9690# a_19094_n9066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8017 a_23296_3565# a_23182_3446# a_23390_3446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8018 gnd d0 a_20326_7284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8019 a_33780_5972# a_33567_5972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8020 a_19126_n3189# a_19221_n3813# a_19176_n3609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8021 a_16072_6557# a_16551_6725# a_16759_6725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8022 a_24642_n9050# a_24737_n9674# a_24688_n9658# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8023 a_16085_3619# a_16083_3405# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8024 vdd d0 a_41931_n3603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8025 a_12333_7400# a_12120_7400# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8026 a_16869_n4853# a_16448_n4853# a_16172_n4834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8027 a_5424_3611# a_5905_3781# a_6113_3781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8028 a_16169_n6029# a_16652_n6395# a_16860_n6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8029 a_22188_n8339# a_21975_n8339# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8030 a_34192_4447# a_34083_4447# a_34291_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8031 a_20064_8455# a_20067_7863# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8032 gnd a_31162_6268# a_30954_6268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8033 vdd a_8741_n8701# a_8533_n8701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8034 a_10498_n10484# a_21654_n10615# a_20848_n805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8035 a_11162_n5855# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8036 a_38353_n5390# a_39158_n5624# a_39327_n5063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8037 a_37285_271# a_37072_271# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8038 a_12221_n7070# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8039 a_27283_n3422# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8040 a_27584_8084# a_27163_8084# a_26887_7984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8041 gnd d1 a_14052_3154# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8042 a_32375_n6997# a_32856_n7368# a_33064_n7368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8043 vdd a_8609_5643# a_8401_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8044 gnd a_41919_n5563# a_41711_n5563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8045 a_36278_7466# a_36535_7276# a_35269_7055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8046 vdd a_19402_n8709# a_19194_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8047 gnd a_15057_5345# a_14849_5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8048 a_26671_n2223# a_27501_n2441# a_27709_n2441# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8049 vdd a_3425_n5366# a_3217_n5366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8050 a_4216_n8940# a_4219_n8337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8051 a_22308_7124# a_21887_7124# a_21611_7306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8052 a_23015_n3677# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8053 a_23233_n2696# a_23020_n2696# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8054 a_33630_3454# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8055 a_38358_n4409# a_37937_n4409# a_37671_n4223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8056 gnd d1 a_19328_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8057 a_19126_n3189# a_19379_n3393# a_18957_n4309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8058 gnd a_14059_2175# a_13851_2175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8059 a_23209_4439# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8060 a_12384_n6650# a_12171_n6650# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8061 a_12179_n4693# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8062 a_138_4018# a_624_3802# a_832_3802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8063 a_39562_n5879# a_39453_n6056# a_39661_n6056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8064 a_34196_6439# a_33775_6439# a_34031_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8065 a_35381_n3789# a_36442_n3624# a_36397_n3420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8066 a_22926_2047# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8067 a_27621_1226# a_27200_1226# a_26924_1408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8068 a_32274_6933# a_32760_6717# a_32968_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8069 a_16774_3789# a_16353_3789# a_16080_4005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8070 a_21899_5164# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8071 a_11582_n5440# a_11161_n5440# a_10893_n5069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8072 a_41664_n6750# a_41917_n6954# a_40651_n6516# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8073 a_23382_5403# a_22961_5403# a_23283_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8074 a_27272_n5797# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8075 gnd a_40904_n6720# a_40696_n6720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8076 a_8394_8036# a_9452_8257# a_9403_8447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8077 a_40240_n10360# a_40401_n6288# a_40352_n6272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8078 a_39069_3994# a_38856_3994# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8079 a_16439_n6395# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8080 a_22322_3773# a_21901_3773# a_21628_3989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8081 a_33952_3454# a_33843_3454# a_34051_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8082 gnd a_8748_n7722# a_8540_n7722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8083 gnd d1 a_8753_n6741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8084 gnd d1 a_3480_n4805# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8085 vdd a_36623_n8520# a_36415_n8520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8086 gnd d2 a_30176_n9233# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8087 a_18076_n8077# a_17655_n8077# a_17911_n9009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8088 a_825_6174# a_1629_5993# a_1798_5551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8089 a_1505_n7623# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8090 a_32996_2236# a_32575_2236# a_32299_2136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8091 a_130_5975# a_135_5589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8092 a_22911_4983# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8093 a_38157_n3430# a_37944_n3430# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8094 a_17824_n6872# a_17452_n6629# a_16860_n6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8095 a_22115_4188# a_21902_4188# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8096 a_37548_7992# a_37550_7893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8097 gnd a_3383_5103# a_3175_5103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8098 a_10779_7943# a_11265_7727# a_11473_7727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8099 vdd d0 a_25880_5874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8100 a_27490_n4816# a_27277_n4816# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8101 a_26894_7499# a_26892_7285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8102 a_11355_n9772# a_11142_n9772# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8103 a_40570_3117# a_41628_3338# a_41583_3351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8104 a_28901_n5871# a_28504_n4123# a_28760_n5055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8105 a_20887_141# a_20674_141# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8106 a_27476_n7339# a_27263_n7339# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8107 a_28911_4418# a_28490_4418# a_28812_4418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8108 a_12140_3483# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8109 a_16184_n2874# a_16673_n2893# a_16881_n2893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8110 a_26624_263# a_26411_263# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8111 a_13660_n8059# a_13858_n9291# a_13813_n9087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8112 a_29939_n5300# a_30043_n4755# a_29994_n4739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8113 a_35226_5656# a_35321_6063# a_35276_6076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8114 a_11072_3810# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8115 a_26899_6306# a_27388_6124# a_27596_6124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8116 vdd d1 a_35542_3125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8117 gnd a_8659_6063# a_8451_6063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8118 a_16428_n8770# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8119 vdd d3 a_30043_n4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8120 a_21640_2029# a_21645_1643# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8121 a_37582_2611# a_37580_2397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8122 vdd d0 a_4399_4361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8123 vdd a_36547_5316# a_36339_5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8124 a_35264_8036# a_35517_8023# a_35214_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8125 a_13732_5862# a_13989_5672# a_13567_6794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8126 vdd d0 a_20429_n5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8127 a_12442_7400# a_12333_7400# a_12541_7400# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8128 a_18957_n4309# a_19171_n3393# a_19126_n3189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8129 a_5491_n8461# a_5980_n8762# a_6188_n8762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8130 a_24489_n8022# a_24687_n9254# a_24638_n9238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8131 vdd d0 a_15051_5911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8132 a_14798_5924# a_14794_6101# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8133 vdd a_35549_2146# a_35341_2146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8134 a_39138_n9541# a_38925_n9541# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8135 a_2153_380# a_2880_4671# a_2831_4861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8136 a_14908_n3864# a_14904_n4052# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8137 a_4154_2591# a_4157_1999# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8138 a_30897_7022# a_30909_6281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8139 a_21987_n6379# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8140 vdd d0 a_9766_n6975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8141 vdd a_3177_n6330# a_2969_n6330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8142 a_16767_6161# a_17571_5980# a_17740_5538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8143 a_10873_n8986# a_11354_n9357# a_11562_n9357# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8144 vdd a_24673_2650# a_24465_2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8145 gnd a_15154_n5047# a_14946_n5047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8146 a_17467_n3693# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8147 a_123_7549# a_604_7719# a_812_7719# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8148 a_17779_6447# a_17566_6447# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8149 a_28584_1465# a_28212_1045# a_27620_811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8150 a_21643_1147# a_21645_1048# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8151 a_38244_7677# a_37823_7677# a_37550_7893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8152 a_8508_n4580# a_9566_n5018# a_9521_n4814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8153 a_9443_997# a_9696_984# a_8427_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8154 vdd a_41843_2359# a_41635_2359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8155 a_12556_n5113# a_12442_n5113# a_12650_n5113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8156 a_11506_2265# a_11085_2265# a_10809_2165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8157 vdd d0 a_20326_7284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8158 gnd a_19325_5090# a_19117_5090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8159 a_35285_3315# a_36346_2944# a_36297_3134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8160 a_38041_6696# a_37828_6696# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8161 a_411_3802# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8162 a_29770_n8001# a_29968_n9233# a_29923_n9029# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8163 a_27689_n6358# a_28494_n6592# a_28653_n6835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8164 a_24410_n6285# a_24554_n4309# a_24509_n4105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8165 vdd a_24957_n7714# a_24749_n7714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8166 a_16848_n8355# a_16427_n8355# a_16161_n8169# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8167 a_20158_n8927# a_20161_n8324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8168 a_21645_1643# a_22126_1813# a_22334_1813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8169 a_711_n6823# a_498_n6823# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8170 a_13879_n5778# a_14940_n5613# a_14895_n5409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8171 a_39302_n8803# a_38930_n8560# a_38338_n8326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8172 a_35303_n9058# a_35398_n9682# a_35349_n9666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8173 a_28671_3425# a_28250_3425# a_28572_3425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8174 a_33937_7490# a_33555_7932# a_32964_8113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8175 a_13585_n6134# a_13705_n8263# a_13660_n8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8176 a_19080_3146# a_20138_3367# a_20093_3380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8177 a_37671_n3445# a_37676_n3059# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8178 a_14912_n2468# a_14908_n2656# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8179 a_5923_1255# a_5710_1255# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8180 vdd d2 a_3348_1747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8181 a_8488_n8497# a_9546_n8935# a_9497_n8919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8182 a_11141_n9357# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8183 a_18937_n8226# a_19194_n8242# a_18866_n6113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8184 a_32850_n8762# a_32637_n8762# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8185 gnd d0 a_41830_3904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8186 a_13795_3344# a_14856_2973# a_14811_2986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8187 a_17685_n2712# a_17472_n2712# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8188 a_6740_7371# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8189 a_6779_n8581# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8190 a_1684_5432# a_1471_5432# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8191 a_13492_4869# a_13749_4679# a_12814_388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8192 a_39572_4426# a_39151_4426# a_39477_6418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8193 a_23127_4007# a_22914_4007# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8194 vdd d1 a_14052_3154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8195 a_24414_n6097# a_24534_n8226# a_24485_n8210# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8196 a_37654_n6762# a_37654_n6480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8197 a_9508_n6544# a_9765_n6560# a_8496_n6725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8198 a_19177_n2816# a_20238_n2651# a_20189_n2635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8199 a_37560_6032# a_38049_6132# a_38257_6132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8200 vdd a_15057_5345# a_14849_5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8201 a_40600_n5308# a_40857_n5324# a_40451_n4092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8202 gnd d0 a_36542_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8203 vdd a_9773_n4603# a_9565_n4603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8204 a_13774_8065# a_14027_8052# a_13724_7645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8205 a_26983_n8928# a_27464_n9299# a_27672_n9299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8206 a_2140_4468# a_1719_4468# a_2045_6460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8207 a_13790_4325# a_14851_3954# a_14802_4144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8208 vdd a_24970_n4776# a_24762_n4776# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8209 a_29602_4811# a_29746_2629# a_29697_2819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8210 gnd d1 a_3403_1186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8211 vdd d1 a_19328_4114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8212 vdd a_14059_2175# a_13851_2175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8213 vdd d0 a_25874_7268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8214 a_845_2257# a_424_2257# a_148_2439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8215 a_35358_n8497# a_35611_n8701# a_35299_n9246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8216 a_4158_1195# a_162_876# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8217 a_28666_n5055# a_28552_n5055# a_28760_n5055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8218 a_35296_2159# a_36354_2380# a_36305_2570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8219 a_27381_7103# a_27168_7103# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8220 a_16655_n5419# a_16442_n5419# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8221 a_11052_7727# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8222 a_10873_n8986# a_10871_n8772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8223 a_5709_840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8224 a_14884_n7969# a_14887_n7366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8225 a_19087_2167# a_19340_2154# a_19037_1747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8226 a_7062_7371# a_6953_7371# a_7161_7371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8227 a_14876_n8533# a_14888_n7781# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8228 gnd a_41937_n3037# a_41729_n3037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8229 a_1989_n5105# a_1946_n4173# a_2130_n5921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8230 a_29695_n6076# a_29815_n8205# a_29770_n8001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8231 gnd a_9781_n4039# a_9573_n4039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8232 a_24615_6068# a_25673_6289# a_25624_6479# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8233 a_27175_6124# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8234 a_39245_1473# a_38873_1053# a_38282_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8235 a_26912_3086# a_27401_3186# a_27609_3186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8236 a_36277_7051# a_36289_6310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8237 a_18941_n8038# a_19139_n9270# a_19090_n9254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8238 a_22424_n3858# a_23228_n3677# a_23397_n3116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8239 a_41642_n9464# a_41899_n9480# a_40630_n9645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8240 a_32756_8113# a_32543_8113# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8241 gnd d3 a_19125_2666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8242 a_16648_n7791# a_16435_n7791# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8243 gnd d0 a_4472_n8541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8244 a_12447_7519# a_12065_7961# a_11474_8142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8245 a_40662_n3768# a_41723_n3603# a_41678_n3399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8246 gnd a_31166_4872# a_30958_4872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8247 a_4130_6895# a_4126_7072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8248 a_7099_1613# a_6717_2055# a_6126_2236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8249 a_18082_4455# a_17661_4455# a_17987_6447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8250 a_18171_n6085# a_17750_n6085# a_18072_n5908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8251 a_39163_n4643# a_38950_n4643# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8252 a_25647_1970# a_25900_1957# a_24631_2328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8253 a_10888_n5455# a_10893_n5069# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8254 a_1726_n5666# a_1513_n5666# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8255 a_20101_1597# a_20358_1407# a_19092_1186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8256 a_37933_n5805# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8257 a_6935_1074# a_6722_1074# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8258 a_725_n3472# a_512_n3472# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8259 a_21695_n9434# a_21697_n9335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8260 a_16772_5180# a_16351_5180# a_16075_5080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8261 a_19169_n4588# a_20227_n5026# a_20178_n5010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8262 vdd a_8659_6063# a_8451_6063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8263 a_11588_n4874# a_12392_n4693# a_12551_n4936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8264 vdd a_24915_n5337# a_24707_n5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8265 a_32395_n3080# a_32393_n2866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8266 a_20083_4123# a_20093_3380# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8267 a_35260_8213# a_35517_8023# a_35214_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8268 a_6973_3454# a_6760_3454# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8269 a_7074_5411# a_6702_4991# a_6110_4757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8270 a_6000_n4845# a_5787_n4845# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8271 a_38074_1234# a_37861_1234# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8272 a_37848_2779# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8273 a_41662_n5547# a_41672_n4793# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8274 a_32363_n8957# a_32361_n8743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8275 a_2153_380# a_2880_4671# a_2835_4684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8276 a_7163_n6864# a_6791_n6621# a_6200_n6802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8277 a_41667_n5774# a_41920_n5978# a_40654_n5540# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8278 a_26996_n5778# a_27485_n5797# a_27693_n5797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8279 gnd a_35542_3125# a_35334_3125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8280 a_8395_7232# a_9456_6861# a_9407_7051# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8281 a_30928_1949# a_31181_1936# a_29912_2307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8282 a_32648_n6387# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8283 a_16442_n5419# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8284 a_11266_8142# a_11053_8142# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8285 gnd a_9697_1399# a_9489_1399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8286 vdd a_24826_3678# a_24618_3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8287 a_153_1458# a_153_1176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8288 a_8441_n7286# a_8545_n6741# a_8496_n6725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8289 a_35061_6588# a_35314_6575# a_34986_4663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8290 a_4999_n10469# a_8138_n10397# a_8089_n10381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8291 a_17854_1502# a_17799_2530# a_17983_4455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8292 a_12630_n9030# a_12209_n9030# a_12536_n9030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8293 a_36382_n5983# a_36639_n5999# a_35373_n5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8294 a_14823_1026# a_15076_1013# a_13807_1384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8295 a_8508_n4580# a_8761_n4784# a_8449_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8296 a_27609_3186# a_28413_3005# a_28572_3425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8297 gnd a_3386_4127# a_3178_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8298 a_6182_n9328# a_5761_n9328# a_5488_n9343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8299 a_27698_n4816# a_28502_n4635# a_28661_n4878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8300 a_41578_4332# a_41831_4319# a_40565_4098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8301 vdd a_25963_n8927# a_25755_n8927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8302 a_4247_n2648# a_5181_n2252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8303 a_39433_n3103# a_39012_n3103# a_39339_n3103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8304 a_11485_5767# a_12290_6001# a_12459_5559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8305 a_7042_n9001# a_6829_n9001# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8306 a_32563_4196# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8307 a_22408_n6379# a_23213_n6613# a_23372_n6856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8308 a_21893_5730# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8309 a_17576_4999# a_17363_4999# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8310 gnd a_20326_7284# a_20118_7284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8311 a_32393_n2584# a_32882_n2885# a_33090_n2885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8312 a_11303_1284# a_11090_1284# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8313 a_913_n7389# a_492_n7389# a_219_n7404# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8314 gnd d0 a_31186_955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8315 a_1813_1515# a_1704_1515# a_1912_1515# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8316 a_12120_7400# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8317 a_35075_n6105# a_35195_n8234# a_35146_n8218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8318 vdd d0 a_31258_n5555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8319 a_40557_6055# a_40810_6042# a_40507_5635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8320 gnd d1 a_3487_n3826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8321 a_13770_8242# a_14027_8052# a_13724_7645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8322 vdd a_36630_n7541# a_36422_n7541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8323 vdd d0 a_36635_n6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8324 a_605_8134# a_392_8134# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8325 a_28812_4418# a_28415_2493# a_28683_1465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8326 a_18095_367# a_18822_4658# a_18777_4671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8327 vdd a_30238_n7693# a_30030_n7693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8328 vdd a_4480_n7977# a_4272_n7977# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8329 a_40584_n9037# a_40679_n9661# a_40630_n9645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8330 vdd d1 a_3403_1186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8331 a_5767_n8762# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8332 a_19005_7624# a_19100_8031# a_19051_8221# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8333 a_35296_2159# a_36354_2380# a_36309_2393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8334 gnd a_14052_3154# a_13844_3154# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8335 a_21702_n8949# a_22183_n9320# a_22391_n9320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8336 a_39327_n5063# a_39213_n5063# a_39421_n5063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8337 vdd d0 a_9769_n5999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8338 a_19083_2344# a_19340_2154# a_19037_1747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8339 a_926_n4451# a_505_n4451# a_232_n4466# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8340 gnd a_19328_4114# a_19120_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8341 a_22131_832# a_21918_832# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8342 vdd a_37407_n10464# a_37199_n10464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8343 a_12913_388# a_12492_388# a_12814_388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8344 vdd d3 a_19125_2666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8345 a_25616_8262# a_25869_8249# a_24603_8028# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8346 vdd d0 a_41815_6840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8347 a_20088_4361# a_20341_4348# a_19075_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8348 a_29880_8184# a_30941_7813# a_30896_7826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8349 a_32287_4096# a_32776_4196# a_32984_4196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8350 a_12492_388# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8351 a_3146_1376# a_4207_1005# a_4158_1195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8352 a_4153_2176# a_4163_1433# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8353 a_27003_n5011# a_27001_n4797# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8354 a_17755_1502# a_17646_1502# a_17854_1502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8355 gnd d1 a_14153_n2853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8356 a_24670_n3361# a_24927_n3377# a_24505_n4293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8357 a_34140_n5084# a_33719_n5084# a_34041_n4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8358 a_25624_6479# a_25627_5887# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8359 a_10905_n2514# a_11391_n2499# a_11599_n2499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8360 gnd d0 a_41810_7821# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8361 a_13775_7261# a_14836_6890# a_14791_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8362 a_25729_n4391# a_25725_n4579# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8363 gnd d0 a_9696_984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8364 gnd d0 a_36546_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8365 a_23365_n8993# a_22983_n9554# a_22391_n9320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8366 a_12548_n7070# a_12434_n7070# a_12642_n7070# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8367 a_29866_1710# a_30119_1697# a_29697_2819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8368 a_24581_1908# a_24685_1157# a_24640_1170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8369 vdd d0 a_25969_n7533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8370 a_17888_n4160# a_17675_n4160# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8371 a_12315_1103# a_12102_1103# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8372 a_36367_n8919# a_36370_n8316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8373 a_29579_n10352# a_29836_n10368# a_26489_n10440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8374 a_16774_3789# a_17579_4023# a_17748_3581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8375 vdd d0 a_20320_7850# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8376 vdd a_15128_n9530# a_14920_n9530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8377 gnd a_8652_7042# a_8444_7042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8378 a_16869_n4853# a_16448_n4853# a_16172_n4552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8379 a_16063_7322# a_16552_7140# a_16760_7140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8380 vdd a_14039_6092# a_13831_6092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8381 a_39319_n7020# a_38937_n7581# a_38345_n7347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8382 a_32376_n5807# a_32376_n5525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8383 a_934_n3887# a_513_n3887# a_237_n3586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8384 vdd d1 a_19434_n2832# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8385 a_480_n9349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8386 a_32857_n7783# a_32644_n7783# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8387 a_11162_n5855# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8388 gnd a_25957_n9493# a_25749_n9493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8389 a_38354_n5805# a_39158_n5624# a_39327_n5063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8390 a_21906_2792# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8391 a_24616_5264# a_25677_4893# a_25628_5083# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8392 vdd a_35542_3125# a_35334_3125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8393 a_6099_7132# a_6903_6951# a_7062_7371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8394 a_38841_6930# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8395 a_11089_869# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8396 a_10891_n4573# a_11380_n4874# a_11588_n4874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8397 a_26894_6904# a_27380_6688# a_27588_6688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8398 a_5986_n7368# a_5773_n7368# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8399 a_16181_n4252# a_16179_n3855# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8400 a_33064_n7368# a_33869_n7602# a_34038_n7041# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8401 a_8520_n2620# a_9578_n3058# a_9529_n3042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8402 a_27015_n2456# a_27501_n2441# a_27709_n2441# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8403 a_16172_n4552# a_16174_n4453# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8404 a_39453_n6056# a_39240_n6056# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8405 a_20096_2578# a_20099_1986# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8406 vdd d0 a_15133_n8549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8407 a_23015_n3677# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8408 a_37582_2016# a_37587_1630# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8409 a_35057_6765# a_35314_6575# a_34986_4663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8410 vdd a_30188_n7273# a_29980_n7273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8411 a_27187_2771# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8412 a_14819_1203# a_15076_1013# a_13807_1384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8413 a_35365_n7518# a_35618_n7722# a_35315_n7098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8414 a_10816_1085# a_10823_884# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8415 gnd a_35626_n5765# a_35418_n5765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8416 gnd d1 a_35631_n4784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8417 a_12791_n5929# a_12394_n4181# a_12662_n3153# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8418 a_17566_6447# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8419 gnd d0 a_25894_3351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8420 a_32383_n4445# a_32869_n4430# a_33077_n4430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8421 a_30005_n3572# a_31063_n4010# a_31018_n3806# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8422 a_32984_4196# a_33788_4015# a_33957_3573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8423 a_21709_n7375# a_21714_n6989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8424 a_10900_n4273# a_10898_n3876# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8425 a_16775_4204# a_16354_4204# a_16078_4104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8426 vdd a_20326_7284# a_20118_7284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8427 gnd d0 a_31170_4311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8428 a_19156_n7526# a_20214_n7964# a_20169_n7760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8429 a_10903_n2613# a_10905_n2514# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8430 a_32772_4757# a_32559_4757# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8431 a_23216_n5637# a_23003_n5637# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8432 a_10868_n9967# a_10866_n9753# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8433 gnd a_25901_2372# a_25693_2372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8434 a_31889_n10455# a_37199_n10464# a_35058_n10381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8435 a_40553_6232# a_40810_6042# a_40507_5635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8436 vdd a_41911_n7520# a_41703_n7520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8437 a_5710_1255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8438 vdd a_3348_1747# a_3140_1747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8439 gnd a_3183_2679# a_2975_2679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8440 a_40352_n6272# a_40496_n4296# a_40451_n4092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8441 vdd a_31244_n8906# a_31036_n8906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8442 a_1471_5432# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8443 a_19005_7624# a_19100_8031# a_19055_8044# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8444 vdd d2 a_19379_n3393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8445 vdd a_14052_3154# a_13844_3154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8446 a_12295_5020# a_12082_5020# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8447 a_33058_n8762# a_32637_n8762# a_32361_n8743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8448 a_41679_n3814# a_41675_n4002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8449 a_37828_6696# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8450 a_41573_4094# a_41583_3351# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8451 a_11355_n9772# a_11142_n9772# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8452 a_27490_n4816# a_27277_n4816# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8453 a_25741_n2431# a_25994_n2635# a_24725_n2800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8454 a_12705_388# a_12492_388# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8455 gnd a_36542_6297# a_36334_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8456 vdd d0 a_20357_992# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8457 a_19102_n7294# a_19206_n6749# a_19161_n6545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8458 gnd a_3403_1186# a_3195_1186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8459 a_5397_8013# a_5886_8113# a_6094_8113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8460 vdd a_19328_4114# a_19120_4114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8461 vdd d0 a_41916_n6539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8462 a_40263_4819# a_40407_2637# a_40362_2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8463 vdd a_25874_7268# a_25666_7268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8464 a_11580_n6831# a_12384_n6650# a_12543_n6893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8465 a_7415_n8069# a_6994_n8069# a_7262_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8466 a_33944_n3124# a_33731_n3124# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8467 a_19165_n4776# a_19422_n4792# a_19110_n5337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8468 a_28641_n8795# a_28532_n8972# a_28740_n8972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8469 a_13779_7084# a_14837_7305# a_14788_7495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8470 a_2907_n10402# a_2857_n10418# a_2229_n6098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8471 a_5491_n8743# a_5980_n8762# a_6188_n8762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8472 a_41582_2936# a_41835_2923# a_40566_3294# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8473 a_3133_4140# a_4191_4361# a_4142_4551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8474 a_22403_n7360# a_21982_n7360# a_21714_n6989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8475 a_23119_5964# a_22906_5964# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8476 a_17986_367# a_17773_367# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8477 a_7000_4447# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8478 a_13863_n9507# a_14116_n9711# a_13813_n9087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8479 a_34008_2522# a_33795_2522# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8480 gnd d0 a_9765_n6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8481 a_41683_n2418# a_41679_n2606# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8482 a_8431_1178# a_9489_1399# a_9440_1589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8483 gnd d5 a_24555_n10389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8484 vdd d3 a_3163_6596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8485 a_11282_4786# a_11069_4786# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8486 a_10868_n9372# a_11354_n9357# a_11562_n9357# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8487 vdd a_29948_n6280# a_29740_n6280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8488 a_32669_n2885# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8489 gnd a_19125_2666# a_18917_2666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8490 a_7082_3454# a_6710_3034# a_6119_3215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8491 a_40240_n10360# a_40497_n10376# a_37150_n10448# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8492 a_4232_n6792# a_4228_n6980# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8493 a_20177_n5803# a_20173_n5991# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8494 a_217_n7503# a_219_n7404# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8495 a_116_8316# a_605_8134# a_813_8134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8496 a_24712_n5553# a_24965_n5757# a_24662_n5133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8497 a_38245_8092# a_37824_8092# a_37548_7992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8498 a_37671_n3445# a_38157_n3430# a_38365_n3430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8499 a_35366_n6725# a_36427_n6560# a_36382_n6356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8500 a_16558_5746# a_16345_5746# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8501 a_28816_6410# a_28395_6410# a_28663_5382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8502 a_29931_n7257# a_30035_n6712# a_29990_n6508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8503 a_38264_3760# a_37843_3760# a_37570_3976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8504 a_3219_n6558# a_4277_n6996# a_4232_n6792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8505 a_36386_n4587# a_36643_n4603# a_35374_n4768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8506 a_31018_n2598# a_31952_n2202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8507 vdd a_8652_7042# a_8444_7042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8508 vdd d1 a_3383_5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8509 gnd a_30196_n5316# a_29988_n5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8510 a_16338_6725# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8511 a_27013_n2837# a_27013_n2555# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8512 vdd a_25970_n7948# a_25762_n7948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8513 a_27257_n8733# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8514 gnd d2 a_8629_1726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8515 a_35276_6076# a_36334_6297# a_36289_6310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8516 a_22188_n8339# a_21975_n8339# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8517 a_6722_1074# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8518 gnd a_35576_n5345# a_35368_n5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8519 a_7262_n7041# a_6841_n7041# a_7163_n6864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8520 a_17685_n2712# a_17472_n2712# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8521 a_41646_n9276# a_41642_n9464# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8522 a_8449_n5329# a_8706_n5345# a_8300_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8523 a_18777_4671# a_19030_4658# a_18095_367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8524 vdd d0 a_31250_n7512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8525 a_621_4778# a_408_4778# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8526 a_6760_3454# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8527 a_6992_n8581# a_6779_n8581# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8528 a_4220_n8752# a_4473_n8956# a_3207_n8518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8529 a_3152_n9079# a_3247_n9703# a_3202_n9499# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8530 a_20092_2965# a_20345_2952# a_19076_3323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8531 vdd a_20409_n9509# a_20201_n9509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8532 a_12563_n2976# a_12191_n2733# a_11600_n2914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8533 a_27672_n9299# a_28477_n9533# a_28646_n8972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8534 a_32269_7914# a_32755_7698# a_32963_7698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8535 a_41570_5070# a_41578_4332# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8536 a_38358_n4409# a_37937_n4409# a_37664_n4424# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8537 a_12518_2551# a_12305_2551# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8538 vdd a_4484_n6581# a_4276_n6581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8539 gnd a_31238_n9472# a_31030_n9472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8540 a_6208_n4845# a_5787_n4845# a_5511_n4826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8541 a_22215_n3443# a_22002_n3443# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8542 a_30908_5866# a_30904_6043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8543 a_13841_n3398# a_13945_n2853# a_13896_n2837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8544 vdd d3 a_24653_6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8545 a_148_2157# a_637_2257# a_845_2257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8546 a_11053_8142# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8547 vdd d0 a_25894_3351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8548 a_23377_n7033# a_23263_n7033# a_23471_n7033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8549 a_20853_n686# a_20674_141# a_20996_141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8550 a_27677_n8318# a_27256_n8318# a_26990_n8132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8551 a_36397_n3420# a_36650_n3624# a_35381_n3789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8552 a_30914_5300# a_31167_5287# a_29901_5066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8553 a_11582_n5440# a_11161_n5440# a_10888_n5455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8554 vdd d0 a_31170_4311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8555 a_33988_6439# a_33775_6439# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8556 a_9497_n8919# a_9754_n8935# a_8488_n8497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8557 a_24700_n7698# a_25761_n7533# a_25716_n7329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8558 vdd a_25901_2372# a_25693_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8559 a_38848_5951# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8560 a_32968_6717# a_32547_6717# a_32281_6549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8561 a_3015_n4322# a_3229_n3406# a_3180_n3390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8562 gnd d1 a_40912_n4763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8563 vdd d0 a_15065_3388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8564 a_28673_n2918# a_28301_n2675# a_27710_n2856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8565 a_17363_4999# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8566 a_25623_6064# a_25633_5321# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8567 a_11090_1284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8568 gnd d0 a_41843_2359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8569 a_13813_n9087# a_14066_n9291# a_13660_n8059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8570 a_37587_1630# a_38068_1800# a_38276_1800# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8571 a_39163_n4643# a_38950_n4643# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8572 a_17824_n6872# a_17452_n6629# a_16861_n6810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8573 gnd d2 a_35556_n9262# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8574 a_31022_n2410# a_31275_n2614# a_30006_n2779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8575 a_23630_4439# a_23209_4439# a_23535_6431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8576 a_837_2821# a_416_2821# a_150_2653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8577 gnd d0 a_4416_1420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8578 a_392_8134# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8579 a_1726_n5666# a_1513_n5666# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8580 a_37933_n5805# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8581 a_21618_6045# a_22107_6145# a_22315_6145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8582 a_33656_n7602# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8583 vdd a_3403_1186# a_3195_1186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8584 vdd d0 a_25990_n4031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8585 a_8516_n2808# a_9577_n2643# a_9532_n2439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8586 a_6130_840# a_5709_840# a_5443_855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8587 a_27476_n7339# a_27263_n7339# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8588 a_13864_n8714# a_14925_n8549# a_14880_n8345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8589 a_34041_n4907# a_33669_n4664# a_33078_n4845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8590 gnd a_40595_6554# a_40387_6554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8591 a_28552_7342# a_28443_7342# a_28651_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8592 a_3133_4140# a_4191_4361# a_4146_4374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8593 a_25724_n5372# a_25720_n5560# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8594 a_517_n2491# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8595 a_31006_n5766# a_31002_n5954# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8596 a_35319_n5329# a_35423_n4784# a_35374_n4768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8597 a_9508_n7752# a_9761_n7956# a_8495_n7518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8598 a_17844_n2955# a_17735_n3132# a_17943_n3132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8599 a_4234_n5401# a_4487_n5605# a_3218_n5770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8600 a_32861_n6387# a_32648_n6387# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8601 a_7163_n6864# a_6791_n6621# a_6199_n6387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8602 a_32656_n4430# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8603 vdd d3 a_35423_n4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8604 a_37849_3194# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8605 a_12498_6468# a_12285_6468# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8606 a_39332_3433# a_38911_3433# a_39233_3433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8607 vdd a_19125_2666# a_18917_2666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8608 a_16149_n9351# a_16154_n8965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8609 a_27489_n4401# a_27276_n4401# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8610 a_36288_5895# a_36284_6072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8611 a_845_2257# a_1649_2076# a_1818_1634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8612 vdd a_41815_6840# a_41607_6840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8613 a_11478_6746# a_11057_6746# a_10791_6578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8614 gnd d1 a_30174_1136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8615 a_2999_n8051# a_3197_n9283# a_3152_n9079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8616 a_37555_7507# a_37553_7293# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8617 gnd d3 a_35403_n8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8618 vdd d0 a_15146_n7004# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8619 a_28589_1584# a_28207_2026# a_27616_2207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8620 a_23390_3446# a_22969_3446# a_23296_3565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8621 a_13676_n4330# a_13933_n4346# a_13581_n6322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8622 a_38036_7677# a_37823_7677# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8623 gnd a_36546_4901# a_36338_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8624 a_506_n4866# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8625 vdd d2 a_8629_1726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8626 a_3219_n6558# a_3472_n6762# a_3160_n7307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8627 a_41586_2549# a_41843_2359# a_40577_2138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8628 a_16063_7040# a_16065_6941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8629 a_39302_n8803# a_38930_n8560# a_38339_n8741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8630 a_12374_n8098# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8631 a_37664_n5019# a_37662_n4805# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8632 a_22409_n6794# a_23213_n6613# a_23372_n6856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8633 a_10880_n7412# a_10885_n7026# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8634 a_12102_1103# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8635 a_5689_4757# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8636 a_22981_1486# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8637 a_40647_n6704# a_41708_n6539# a_41663_n6335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8638 a_34304_359# a_34195_359# a_34403_359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8639 a_32981_5172# a_32560_5172# a_32284_5354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8640 a_28564_5382# a_28192_4962# a_27600_4728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8641 a_12154_n9591# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8642 gnd d1 a_40798_8002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8643 a_41667_n4566# a_41924_n4582# a_40655_n4747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8644 gnd a_4390_5903# a_4182_5903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8645 a_817_6738# a_396_6738# a_123_6954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8646 a_1895_n5105# a_1781_n5105# a_1989_n5105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8647 a_11142_n9772# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8648 a_16673_n2893# a_16460_n2893# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8649 a_5767_n8762# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8650 a_30929_1145# a_26933_826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8651 a_27615_1792# a_27194_1792# a_26926_1622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8652 a_22132_1247# a_21919_1247# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8653 a_3091_1937# a_3195_1186# a_3146_1376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8654 a_26907_4067# a_27396_4167# a_27604_4167# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8655 gnd a_8698_n7302# a_8490_n7302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8656 a_13724_7645# a_13819_8052# a_13770_8242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8657 a_8411_5095# a_9469_5316# a_9420_5506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8658 a_1932_4468# a_1719_4468# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8659 a_41654_n7504# a_41664_n6750# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8660 a_2924_n6126# a_3044_n8255# a_2999_n8051# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8661 a_926_n4451# a_505_n4451# a_239_n4265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8662 a_4236_n5023# a_4239_n4420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8663 a_27408_2207# a_27195_2207# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8664 a_23107_7924# a_22894_7924# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8665 a_36308_1978# a_36561_1965# a_35292_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8666 a_25636_3126# a_25648_2385# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8667 a_38162_n2449# a_37949_n2449# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8668 vdd d0 a_36624_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8669 a_39312_7350# a_38891_7350# a_39218_7469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8670 gnd a_25894_3351# a_25686_3351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8671 a_27015_n2456# a_26671_n2223# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8672 a_21623_5346# a_21623_5064# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8673 gnd d2 a_24826_3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8674 a_39314_n6843# a_39205_n7020# a_39413_n7020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8675 a_23303_1486# a_23194_1486# a_23402_1486# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8676 a_699_n8783# a_486_n8783# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8677 a_16159_n7772# a_16648_n7791# a_16856_n7791# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8678 a_36386_n5795# a_36382_n5983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8679 vdd a_9685_3359# a_9477_3359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8680 a_3202_n9499# a_4260_n9937# a_4211_n9921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8681 a_16065_6941# a_16072_6557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8682 vdd d0 a_4416_1420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8683 a_14877_n8948# a_15134_n8964# a_13868_n8526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8684 gnd a_24881_3117# a_24673_3117# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8685 a_19033_1924# a_19137_1173# a_19088_1363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8686 a_19145_n8693# a_20206_n8528# a_20161_n8324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8687 a_37949_n2449# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8688 a_32975_5738# a_33780_5972# a_33949_5530# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8689 a_17874_4455# a_17661_4455# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8690 a_1692_3475# a_1479_3475# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8691 a_38137_n7347# a_37924_n7347# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8692 a_28482_n8552# a_28269_n8552# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8693 a_30934_1383# a_30930_1560# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8694 vdd a_40595_6554# a_40387_6554# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8695 a_12082_5020# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8696 a_16767_6161# a_16346_6161# a_16070_6343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8697 a_4247_n3856# a_4500_n4060# a_3234_n3622# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8698 a_37560_6032# a_37562_5933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8699 vdd a_20357_992# a_20149_992# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8700 a_29974_n8656# a_31035_n8491# a_30986_n8475# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8701 vdd a_25974_n6552# a_25766_n6552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8702 a_23112_6943# a_22899_6943# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8703 a_4921_292# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8704 a_8483_n9478# a_9541_n9916# a_5488_n9938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8705 a_10799_4026# a_10804_3640# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8706 gnd d0 a_36631_n7956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8707 a_232_n5061# a_230_n4847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8708 a_10891_n4855# a_11380_n4874# a_11588_n4874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8709 a_14818_2007# a_15071_1994# a_13802_2365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8710 a_14904_n4052# a_15161_n4068# a_13895_n3630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8711 a_16791_848# a_16370_848# a_16097_1064# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8712 a_38069_2215# a_37856_2215# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8713 a_33065_n7783# a_33869_n7602# a_34038_n7041# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8714 a_4133_6093# a_4143_5350# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8715 a_6915_4991# a_6702_4991# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8716 a_6999_n7602# a_6786_n7602# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8717 a_16370_848# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8718 a_28388_7903# a_28175_7903# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8719 a_16442_n5419# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8720 vdd d1 a_30174_1136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8721 a_38350_n6366# a_37929_n6366# a_37656_n6381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8722 a_22327_2792# a_23132_3026# a_23291_3446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8723 a_10794_5101# a_10796_5002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8724 a_33795_2522# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8725 a_5513_n5040# a_5994_n5411# a_6202_n5411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8726 a_29896_6047# a_30149_6034# a_29846_5627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8727 gnd d3 a_40684_n8213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8728 a_927_n4866# a_1731_n4685# a_1890_n4928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8729 gnd d0 a_41847_963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8730 vdd a_4505_n3079# a_4297_n3079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8731 a_29912_2307# a_30973_1936# a_30924_2126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8732 vdd a_3163_6596# a_2955_6596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8733 vdd d1 a_19417_n5773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8734 a_40600_n5308# a_40704_n4763# a_40655_n4747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8735 a_16551_6725# a_16338_6725# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8736 a_34380_n6077# a_33959_n6077# a_34281_n5900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8737 a_39225_5390# a_39116_5390# a_39324_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8738 a_24569_3868# a_24826_3678# a_24420_2663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8739 a_10802_3144# a_10804_3045# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8740 a_34083_4447# a_33870_4447# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8741 a_19152_n7714# a_20213_n7549# a_20164_n7533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8742 a_17983_4455# a_17586_2530# a_17842_3462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8743 a_29790_n4084# a_30043_n4288# a_29691_n6264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8744 a_5999_n4430# a_5786_n4430# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8745 a_26887_8266# a_26887_7984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8746 a_13807_1384# a_14868_1013# a_14819_1203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8747 a_25701_n9892# a_25958_n9908# a_24692_n9470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8748 a_12536_n9030# a_12422_n9030# a_12630_n9030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8749 a_33800_2055# a_33587_2055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8750 vdd d0 a_31276_n3029# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8751 a_16085_3024# a_16571_2808# a_16779_2808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8752 a_32267_8295# a_32267_8013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8753 a_23216_n5637# a_23003_n5637# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8754 a_12662_n3153# a_12241_n3153# a_12563_n2976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8755 a_20178_n5010# a_20181_n4407# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8756 a_16660_n4438# a_16447_n4438# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8757 a_11069_4786# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8758 vdd d0 a_20427_n6983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8759 a_4151_3393# a_4404_3380# a_3138_3159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8760 a_26588_n10440# a_26538_n10456# a_26489_n10440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8761 a_31014_n3994# a_31017_n3391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8762 gnd d0 a_20352_1973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8763 a_21633_3008# a_22119_2792# a_22327_2792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8764 a_37394_271# a_39263_338# a_39572_4426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8765 a_35265_7232# a_36326_6861# a_36281_6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8766 a_34077_n8069# a_33864_n8069# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8767 vdd d3 a_8464_2658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8768 a_27589_7103# a_28393_6922# a_28552_7342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8769 a_21712_n6493# a_22201_n6794# a_22409_n6794# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8770 a_14891_n5597# a_15148_n5613# a_13879_n5778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8771 a_30930_1560# a_30933_968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8772 gnd d0 a_31256_n6946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8773 a_1912_1515# a_1491_1515# a_1818_1634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8774 a_39263_338# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8775 a_3091_1937# a_3195_1186# a_3150_1199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8776 a_33058_n8762# a_32637_n8762# a_32361_n8461# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8777 a_13724_7645# a_13819_8052# a_13774_8065# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8778 a_12541_7400# a_12498_6468# a_12706_6468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8779 a_9418_5895# a_9671_5882# a_8402_6253# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8780 a_37562_5933# a_37567_5547# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8781 a_8411_5095# a_9469_5316# a_9424_5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8782 a_9507_n7337# a_9503_n7525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8783 a_37674_n2845# a_37674_n2563# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8784 a_37829_7111# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8785 vdd a_35618_n7722# a_35410_n7722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8786 a_34120_n9001# a_33699_n9001# a_34026_n9001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8787 a_22328_3207# a_21907_3207# a_21631_3107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8788 a_35260_8213# a_36321_7842# a_36272_8032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8789 a_40267_4642# a_40387_6554# a_40338_6744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8790 a_41578_4332# a_41574_4509# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8791 a_40570_3117# a_41628_3338# a_41579_3528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8792 a_23283_5403# a_22911_4983# a_22320_5164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8793 a_10809_2447# a_10809_2165# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8794 a_22201_n6794# a_21988_n6794# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8795 a_12305_2551# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8796 a_7193_1494# a_6772_1494# a_7094_1494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8797 a_16164_n6509# a_16166_n6410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8798 a_28646_n8972# a_28532_n8972# a_28740_n8972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8799 a_1510_n6642# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8800 vdd d0 a_15149_n6028# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8801 vdd a_3480_n4805# a_3272_n4805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8802 gnd a_24927_n3377# a_24719_n3377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8803 a_16635_n9336# a_16422_n9336# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8804 a_23630_4439# a_23534_351# a_23742_351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8805 a_13770_8242# a_14831_7871# a_14786_7884# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8806 a_21887_7124# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8807 gnd a_36549_3925# a_36341_3925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8808 a_13880_n6566# a_14938_n7004# a_14893_n6800# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8809 vdd a_25894_3351# a_25686_3351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8810 a_10796_5002# a_10799_4621# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8811 a_13876_n6754# a_14133_n6770# a_13821_n7315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8812 a_38841_6930# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8813 a_29909_3109# a_30162_3096# a_29850_3847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8814 a_13496_4692# a_13616_6604# a_13567_6794# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8815 a_40503_5812# a_40607_5061# a_40558_5251# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8816 vdd d0 a_4485_n6996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8817 a_14895_n5409# a_14891_n5597# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8818 gnd a_19270_5651# a_19062_5651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8819 gnd a_3088_4671# a_2880_4671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8820 a_8422_2336# a_9483_1965# a_9438_1978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8821 a_33775_6439# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8822 vdd a_20341_4348# a_20133_4348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8823 a_12310_2084# a_12097_2084# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8824 a_37843_3760# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8825 a_32787_1821# a_32574_1821# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8826 gnd d0 a_15129_n9945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8827 a_6215_n3866# a_7019_n3685# a_7188_n3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8828 a_32984_4196# a_32563_4196# a_32287_4378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8829 a_11563_n9772# a_12367_n9591# a_12536_n9030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8830 a_33731_n3124# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8831 a_17854_1502# a_17433_1502# a_17760_1621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8832 a_22961_5403# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8833 vdd a_15065_3388# a_14857_3388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8834 a_23511_n6069# a_23298_n6069# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8835 a_19033_1924# a_19137_1173# a_19092_1186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8836 gnd d0 a_36550_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8837 vdd d0 a_41905_n8914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8838 a_41553_8011# a_41563_7268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8839 gnd a_41843_2359# a_41635_2359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8840 a_10782_7061# a_11271_7161# a_11479_7161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8841 a_14819_2422# a_14815_2599# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8842 a_21901_3773# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8843 a_1568_n5105# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8844 vdd a_13726_n10426# a_13518_n10426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8845 a_40427_n8197# a_40684_n8213# a_40356_n6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8846 a_29990_n6508# a_31048_n6946# a_31003_n6742# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8847 a_38925_n9541# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8848 a_38265_4175# a_37844_4175# a_37568_4075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8849 vdd d2 a_19367_n5353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8850 a_32299_2136# a_32301_2037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8851 gnd a_4499_n3645# a_4291_n3645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8852 gnd a_4416_1420# a_4208_1420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8853 a_27257_n8733# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8854 a_31007_n4973# a_31264_n4989# a_29998_n4551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8855 a_5434_1155# a_5923_1255# a_6131_1255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8856 a_16339_7140# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8857 a_26887_7984# a_27376_8084# a_27584_8084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8858 a_36289_5091# a_36546_4901# a_35277_5272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8859 a_19080_3146# a_20138_3367# a_20089_3557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8860 gnd d2 a_3348_1747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8861 gnd a_3487_n3826# a_3279_n3826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8862 a_20158_n8927# a_20415_n8943# a_19149_n8505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8863 a_21715_n5517# a_21717_n5418# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8864 a_20194_n2862# a_20190_n3050# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8865 a_16095_1163# a_16584_1263# a_16792_1263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8866 a_16358_2808# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8867 a_244_n2506# a_730_n2491# a_938_n2491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8868 a_13496_4692# a_13749_4679# a_12814_388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8869 a_18750_n10389# a_19007_n10405# a_15660_n10477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8870 a_12459_5559# a_12345_5440# a_12553_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8871 a_24623_4111# a_25681_4332# a_25632_4522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8872 a_622_5193# a_409_5193# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8873 vdd d0 a_41932_n4018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8874 a_29923_n9029# a_30018_n9653# a_29973_n9449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8875 a_14811_2986# a_14807_3163# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8876 gnd a_15059_3954# a_14851_3954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8877 a_12563_n2976# a_12191_n2733# a_11599_n2499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8878 a_27673_n9714# a_28477_n9533# a_28646_n8972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8879 a_7227_n4152# a_7014_n4152# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8880 a_35358_n8497# a_36416_n8935# a_36371_n8731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8881 gnd d2 a_30119_1697# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8882 a_29892_6224# a_30149_6034# a_29846_5627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8883 gnd d0 a_25874_7268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8884 a_12285_6468# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8885 a_6208_n4845# a_5787_n4845# a_5511_n4544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8886 vdd a_40924_n2803# a_40716_n2803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8887 a_22215_n3443# a_22002_n3443# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8888 a_28572_3425# a_28200_3005# a_27609_3186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8889 a_32368_n7482# a_32857_n7783# a_33065_n7783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8890 a_14794_6101# a_14804_5358# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8891 a_38992_n7020# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8892 a_1781_n5105# a_1568_n5105# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8893 a_11297_1850# a_11084_1850# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8894 gnd d0 a_41912_n7935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8895 gnd a_41920_n5978# a_41712_n5978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8896 vdd a_8768_n3805# a_8560_n3805# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8897 vdd d1 a_8773_n2824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8898 a_11494_4225# a_11073_4225# a_10797_4407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8899 a_20185_n4031# a_20442_n4047# a_19176_n3609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8900 gnd a_30174_1136# a_29966_1136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8901 gnd d1 a_24876_4098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8902 vdd d1 a_14121_n8730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8903 a_11366_n7397# a_11153_n7397# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8904 a_1634_5012# a_1421_5012# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8905 a_7326_6439# a_7213_4447# a_7421_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8906 a_32390_n4244# a_32869_n4430# a_33077_n4430# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8907 vdd a_35568_n7302# a_35360_n7302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8908 a_13807_1384# a_14868_1013# a_14823_1026# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8909 gnd a_25881_6289# a_25673_6289# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8910 gnd a_15165_n2672# a_14957_n2672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8911 a_230_n4565# a_719_n4866# a_927_n4866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8912 a_30904_6043# a_31161_5853# a_29892_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8913 gnd d1 a_24950_n8693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8914 a_14787_8299# a_14783_8476# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8915 a_26933_826# a_27412_811# a_27620_811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8916 a_9406_7855# a_9402_8032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8917 a_37823_7677# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8918 a_33957_3573# a_33575_4015# a_32983_3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8919 a_33924_n7041# a_33711_n7041# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8920 a_32767_5738# a_32554_5738# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8921 a_4147_3570# a_4404_3380# a_3138_3159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8922 a_21702_n8354# a_22188_n8339# a_22396_n8339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8923 a_1672_7392# a_1459_7392# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8924 a_5505_n6402# a_5991_n6387# a_6199_n6387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8925 a_14799_5120# a_15056_4930# a_13787_5301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8926 a_28673_n2918# a_28301_n2675# a_27709_n2441# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8927 gnd a_4383_6882# a_4175_6882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8928 vdd a_35216_n10397# a_35008_n10397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8929 vdd d3 a_13844_2687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8930 a_5505_n6997# a_5503_n6783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8931 a_37580_2397# a_38069_2215# a_38277_2215# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8932 a_7326_6439# a_6905_6439# a_7173_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8933 a_7074_n3124# a_6861_n3124# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8934 a_636_1842# a_423_1842# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8935 a_2041_4468# a_1644_2543# a_1900_3475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8936 gnd a_40798_8002# a_40590_8002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8937 a_32964_8113# a_33768_7932# a_33937_7490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8938 a_35365_n7518# a_36423_n7956# a_36374_n7940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8939 a_40267_4642# a_40387_6554# a_40342_6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8940 a_41577_3917# a_41830_3904# a_40561_4275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8941 gnd d1 a_3467_n7743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8942 a_14798_5924# a_15051_5911# a_13782_6282# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8943 gnd a_9659_7842# a_9451_7842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8944 a_33656_n7602# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8945 a_16792_1263# a_17596_1082# a_17755_1502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8946 a_34041_n4907# a_33669_n4664# a_33077_n4430# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8947 a_8360_3876# a_8464_3125# a_8415_3315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8948 a_32644_n7783# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8949 a_11579_n6416# a_12384_n6650# a_12543_n6893# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8950 a_38158_n3845# a_37945_n3845# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8951 a_20172_n5576# a_20429_n5592# a_19160_n5757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8952 a_5781_n5411# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8953 a_7087_3573# a_6973_3454# a_7181_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8954 vdd d2 a_3405_n9283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8955 a_28666_n5055# a_28284_n5616# a_27693_n5797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8956 a_1518_n4685# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8957 a_24729_n2612# a_24982_n2816# a_24670_n3361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8958 a_26904_5043# a_26906_4944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8959 a_40503_5812# a_40607_5061# a_40562_5074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8960 a_22403_n7360# a_21982_n7360# a_21709_n7375# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8961 vdd a_25995_n3050# a_25787_n3050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8962 a_25617_7458# a_25874_7268# a_24608_7047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8963 gnd d4 a_24578_4642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8964 vdd d1 a_40904_n6720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8965 a_27195_2207# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8966 vdd a_19270_5651# a_19062_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8967 vdd a_3088_4671# a_2880_4671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8968 a_39240_n6056# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8969 a_31005_n5351# a_31258_n5555# a_29989_n5720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8970 a_730_n2491# a_517_n2491# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8971 vdd d0 a_20337_4909# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8972 a_27489_n4401# a_27276_n4401# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8973 a_9422_4115# a_9679_3925# a_8410_4296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8974 a_12467_3602# a_12085_4044# a_11493_3810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8975 a_11277_5767# a_11064_5767# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8976 vdd d0 a_20430_n6007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8977 a_23535_6431# a_23114_6431# a_23370_7363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8978 gnd d0 a_15145_n6589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8979 vdd d0 a_36550_4340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8980 a_38873_1053# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8981 gnd a_24826_3678# a_24618_3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8982 vdd d1 a_19409_n7730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8983 a_17522_n3132# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8984 a_5922_840# a_5709_840# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8985 a_9419_6310# a_9415_6487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8986 a_37676_n3059# a_38157_n3430# a_38365_n3430# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8987 a_6099_7132# a_5678_7132# a_5402_7314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8988 a_14783_8476# a_14786_7884# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8989 vdd a_35328_n6309# a_35120_n6309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8990 a_22416_n4422# a_21995_n4422# a_21722_n4437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8991 a_31023_n2825# a_31019_n3013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8992 a_6923_3034# a_6710_3034# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8993 gnd d0 a_31259_n5970# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8994 a_429_1276# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8995 a_21988_n6794# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8996 a_5518_n3565# a_6007_n3866# a_6215_n3866# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8997 a_14903_n3637# a_14913_n2883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8998 vdd a_4416_1420# a_4208_1420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8999 a_10866_n9471# a_11355_n9772# a_11563_n9772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9000 a_506_n4866# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9001 a_3071_5854# a_3175_5103# a_3130_5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9002 gnd d0 a_20410_n9924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9003 a_38037_8092# a_37824_8092# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9004 a_26990_n7354# a_27476_n7339# a_27684_n7339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9005 gnd a_19397_n9690# a_19189_n9690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9006 a_6717_2055# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9007 a_38244_7677# a_39049_7911# a_39218_7469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9008 a_17661_4455# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9009 a_3218_n5770# a_3475_n5786# a_3172_n5162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9010 a_25705_n8496# a_25962_n8512# a_24693_n8677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9011 vdd d0 a_25978_n5991# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9012 a_24623_4111# a_25681_4332# a_25636_4345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9013 a_11178_n2499# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9014 a_16849_n8770# a_16428_n8770# a_16152_n8469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9015 a_38062_3194# a_37849_3194# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9016 a_7173_5411# a_6752_5411# a_7074_5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9017 gnd d0 a_4403_2965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9018 a_26990_n8132# a_26988_n7735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9019 vdd a_19030_4658# a_18822_4658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9020 a_13883_n5590# a_14941_n6028# a_14896_n5824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9021 a_26981_n8432# a_26983_n8333# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9022 a_18095_367# a_18822_4658# a_18773_4848# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9023 a_11142_n9772# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9024 a_818_7153# a_397_7153# a_121_7053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9025 a_32358_n9343# a_32844_n9328# a_33052_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9026 a_25716_n7329# a_25712_n7517# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9027 a_29889_7026# a_30142_7013# a_29830_7764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9028 a_24712_n5553# a_25770_n5991# a_25721_n5975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9029 a_22335_2228# a_23139_2047# a_23308_1605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9030 gnd a_4410_1986# a_4202_1986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9031 vdd d2 a_24806_7595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9032 a_29989_n5720# a_31050_n5555# a_31005_n5351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9033 a_6702_4991# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9034 a_21715_n5799# a_21715_n5517# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9035 a_28175_7903# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9036 a_33835_5411# a_33622_5411# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9037 vdd a_30174_1136# a_29966_1136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9038 a_32963_7698# a_32542_7698# a_32274_7528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9039 a_12290_6001# a_12077_6001# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9040 a_13863_n9507# a_14921_n9945# a_14872_n9929# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9041 vdd a_9774_n5018# a_9566_n5018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9042 a_6806_n3685# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9043 a_27677_n8318# a_27256_n8318# a_26983_n8333# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9044 a_12372_n8610# a_12159_n8610# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9045 vdd d0 a_15060_4369# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9046 gnd a_41847_963# a_41639_963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9047 gnd a_36618_n9501# a_36410_n9501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9048 vdd a_24762_n4309# a_24554_n4309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9049 a_19013_5841# a_19117_5090# a_19072_5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9050 a_16656_n5834# a_16443_n5834# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9051 gnd d1 a_35554_1165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9052 vdd a_31149_7813# a_30941_7813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9053 a_17715_n7049# a_17502_n7049# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9054 gnd d0 a_4411_2401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9055 gnd a_9754_n8935# a_9546_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9056 a_8479_n9666# a_8736_n9682# a_8433_n9058# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9057 a_29901_5066# a_30959_5287# a_30910_5477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9058 gnd d2 a_8686_n9262# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9059 gnd a_24742_n8226# a_24534_n8226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9060 a_14880_n8345# a_15133_n8549# a_13864_n8714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9061 a_3180_n3390# a_3284_n2845# a_3235_n2829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9062 gnd a_20446_n2651# a_20238_n2651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9063 a_625_4217# a_412_4217# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9064 a_27704_n3422# a_27283_n3422# a_27010_n3437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9065 gnd d1 a_30231_n8672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9066 gnd a_20352_1973# a_20144_1973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9067 a_2130_n5921# a_1733_n4173# a_1989_n5105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9068 vdd a_8464_2658# a_8256_2658# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9069 a_3083_3720# a_3336_3707# a_2930_2692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9070 a_40666_n3580# a_41724_n4018# a_41679_n3814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9071 a_1560_n7062# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9072 gnd d0 a_15161_n4068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9073 a_24581_1908# a_24685_1157# a_24636_1347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9074 a_18862_n6301# a_19006_n4325# a_18961_n4121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9075 a_8360_3876# a_8464_3125# a_8419_3138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9076 a_38137_n7347# a_37924_n7347# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9077 a_28482_n8552# a_28269_n8552# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9078 vdd d2 a_19359_n7310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9079 gnd d2 a_30099_5614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9080 a_33877_n5645# a_33664_n5645# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9081 a_39074_3013# a_38861_3013# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9082 a_16080_4600# a_16563_4765# a_16771_4765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9083 a_25616_7043# a_25628_6302# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9084 a_12345_5440# a_12132_5440# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9085 a_33072_n5411# a_32651_n5411# a_32378_n5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9086 vdd d4 a_24578_4642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9087 a_5436_1651# a_5917_1821# a_6125_1821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9088 a_40646_n7497# a_41704_n7935# a_41655_n7919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9089 a_8465_n3181# a_8718_n3385# a_8296_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9090 a_8461_n3369# a_8565_n2824# a_8520_n2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9091 a_13809_n9275# a_13913_n8730# a_13868_n8526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9092 a_32656_n4430# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9093 gnd d1 a_24856_8015# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9094 a_9432_3372# a_9428_3549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9095 gnd a_19347_n9270# a_19139_n9270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9096 a_6999_n7602# a_6786_n7602# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9097 a_32780_2800# a_32567_2800# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9098 gnd d1 a_14064_1194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9099 a_24638_n9238# a_24742_n8693# a_24693_n8677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9100 a_38350_n6366# a_37929_n6366# a_37659_n6000# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9101 a_12209_n9030# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9102 a_26978_n9909# a_30982_n9871# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9103 a_21975_n8339# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9104 a_5508_n5426# a_5994_n5411# a_6202_n5411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9105 a_22302_7690# a_21881_7690# a_21608_7906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9106 a_3203_n8706# a_4264_n8541# a_4219_n8337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9107 a_33642_1494# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9108 a_1870_n8845# a_1761_n9022# a_1969_n9022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9109 a_17660_n7610# a_17447_n7610# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9110 a_32862_n6802# a_32649_n6802# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9111 a_5778_n6387# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9112 vdd d1 a_24977_n3797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9113 a_31023_n2825# a_31276_n3029# a_30010_n2591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9114 a_32574_1821# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9115 a_1818_1634# a_1436_2076# a_844_1842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9116 a_41558_7030# a_41815_6840# a_40546_7211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9117 a_1887_n7062# a_1505_n7623# a_914_n7804# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9118 gnd d4 a_3177_n6330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9119 a_36297_4353# a_36293_4530# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9120 a_4240_n4835# a_4236_n5023# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9121 vdd d1 a_14128_n7751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9122 gnd a_41924_n4582# a_41716_n4582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9123 a_237_n3586# a_239_n3487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9124 a_2906_6786# a_3120_5664# a_3071_5854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9125 a_5414_5072# a_5416_4973# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9126 gnd a_20435_n5026# a_20227_n5026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9127 a_16786_1829# a_16365_1829# a_16092_2045# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9128 a_41557_7834# a_41810_7821# a_40541_8192# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9129 a_32286_4973# a_32772_4757# a_32980_4757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9130 gnd d0 a_20426_n6568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9131 gnd a_9768_n5584# a_9560_n5584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9132 a_23020_n2696# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9133 a_28683_1465# a_28628_2493# a_28812_4418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9134 a_12097_2084# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9135 a_8406_6076# a_9464_6297# a_9415_6487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9136 a_6183_n9743# a_5762_n9743# a_5486_n9724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9137 vdd a_40609_n6288# a_40401_n6288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9138 a_10779_7943# a_10784_7557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9139 a_13825_n7127# a_13920_n7751# a_13871_n7735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9140 a_4235_n5816# a_4488_n6020# a_3222_n5582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9141 gnd a_3348_1747# a_3140_1747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9142 gnd a_19194_n8242# a_18986_n8242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9143 gnd d7 a_10656_n10500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9144 vdd d4 a_8458_n6309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9145 a_8429_n9246# a_8686_n9262# a_8280_n8030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9146 a_3015_n4322# a_3272_n4338# a_2920_n6314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9147 vdd d2 a_24895_n9254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9148 a_29885_7203# a_30142_7013# a_29830_7764# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9149 a_8296_n4301# a_8510_n3385# a_8465_n3181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9150 a_22127_2228# a_21914_2228# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9151 a_207_n9959# a_4211_n9921# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9152 vdd d4 a_19119_n6317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9153 a_224_n7018# a_222_n6804# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9154 a_39054_6930# a_38841_6930# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9155 a_10791_5983# a_11277_5767# a_11485_5767# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9156 vdd a_36631_n7956# a_36423_n7956# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9157 gnd a_8753_n6741# a_8545_n6741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9158 a_40561_4275# a_41622_3904# a_41577_3917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9159 a_9428_3549# a_9431_2957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9160 a_34058_n3124# a_33676_n3685# a_33084_n3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9161 a_38338_n8326# a_37917_n8326# a_37644_n8341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9162 a_13876_n6754# a_14937_n6589# a_14888_n6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9163 gnd a_25874_7268# a_25666_7268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9164 a_17634_3462# a_17421_3462# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9165 a_40263_4819# a_40407_2637# a_40358_2827# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9166 a_1510_n6642# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9167 a_20067_7863# a_20063_8040# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9168 a_16635_n9336# a_16422_n9336# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9169 vdd a_30251_n4755# a_30043_n4755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9170 gnd a_4493_n5039# a_4285_n5039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9171 a_11084_1850# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9172 a_20068_7059# a_20325_6869# a_19056_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9173 a_38162_n2449# a_37949_n2449# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9174 vdd d1 a_35554_1165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9175 a_32760_6717# a_32547_6717# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9176 a_1421_5012# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9177 gnd a_24876_4098# a_24668_4098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9178 a_30997_n7308# a_31250_n7512# a_29981_n7677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9179 a_5794_n3866# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9180 a_35276_6076# a_35529_6063# a_35226_5656# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9181 a_409_5193# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9182 a_11302_869# a_11089_869# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9183 a_11360_n8791# a_11147_n8791# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9184 vdd d1 a_35606_n9682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9185 gnd a_30023_n8205# a_29815_n8205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9186 a_27481_n6358# a_27268_n6358# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9187 vdd a_15154_n5047# a_14946_n5047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9188 a_20067_7863# a_20320_7850# a_19051_8221# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9189 a_8491_n7706# a_9552_n7541# a_9507_n7337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9190 a_32554_5738# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9191 gnd d0 a_41904_n8499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9192 a_32876_n3451# a_32663_n3451# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9193 a_155_1672# a_153_1458# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9194 a_26995_n6373# a_26998_n5992# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9195 a_135_5589# a_616_5759# a_824_5759# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9196 a_492_n7389# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9197 a_37949_n2449# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9198 vdd a_13844_2687# a_13636_2687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9199 a_35297_1355# a_36358_984# a_36309_1174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9200 a_39143_n8560# a_38930_n8560# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9201 a_38925_n9541# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9202 vdd d2 a_30099_5614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9203 a_423_1842# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9204 a_37575_2995# a_38061_2779# a_38269_2779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9205 a_20161_n8324# a_20414_n8528# a_19145_n8693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9206 a_22429_n2877# a_22008_n2877# a_21732_n2858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9207 a_28683_1465# a_28262_1465# a_28584_1465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
C0 a_10603_285# a_10504_285# 5.04fF
C1 a_39661_n6056# a_40240_n10360# 3.90fF
C2 a_34304_359# a_34291_4447# 3.90fF
C3 a_29000_n6048# a_29579_n10352# 3.90fF
C4 a_20996_141# a_26832_263# 3.01fF
C5 a_39585_338# a_39572_4426# 3.89fF
C6 d2 vdd 4.27fF
C7 a_7434_359# a_7421_4447# 3.89fF
C8 a_18095_367# a_18082_4455# 3.89fF
C9 a_2229_n6098# a_2808_n10402# 3.89fF
C10 d2 gnd 10.12fF
C11 a_12814_388# a_12801_4476# 3.90fF
C12 a_2153_380# a_2140_4468# 3.90fF
C13 a_7510_n6077# a_8089_n10381# 3.90fF
C14 a_26588_n10440# a_21397_n10599# 5.04fF
C15 d0 vdd 17.09fF
C16 a_23719_n6069# a_24298_n10373# 3.89fF
C17 a_28924_330# a_28911_4418# 3.89fF
C18 d0 gnd 40.52fF
C19 d4 gnd 2.53fF
C20 a_12890_n6106# a_13469_n10410# 3.89fF
C21 a_18171_n6085# a_18750_n10389# 3.90fF
C22 a_10498_n10484# a_10399_n10484# 3.01fF
C23 d1 vdd 8.55fF
C24 vdd gnd 54.11fF
C25 d3 vdd 2.14fF
C26 d1 gnd 20.24fF
C27 d3 gnd 5.06fF
C28 a_34380_n6077# a_34959_n10381# 3.89fF
C29 a_23643_351# a_23630_4439# 3.90fF
C30 gnd SUB 332.75fF
C31 vdd SUB 1368.84fF
C32 a_37150_n10448# SUB 4.48fF
C33 d6 SUB 2.81fF
C34 a_35058_n10381# SUB 3.05fF
C35 a_31889_n10455# SUB 6.47fF
C36 a_21397_n10599# SUB 12.33fF
C37 d5 SUB 5.76fF
C38 a_26489_n10440# SUB 4.48fF
C39 a_26588_n10440# SUB 6.01fF
C40 a_24397_n10373# SUB 3.05fF
C41 a_15660_n10477# SUB 4.48fF
C42 a_13568_n10410# SUB 3.05fF
C43 a_10399_n10484# SUB 6.47fF
C44 a_10498_n10484# SUB 12.03fF
C45 a_4999_n10469# SUB 4.48fF
C46 a_5098_n10469# SUB 6.01fF
C47 a_2907_n10402# SUB 3.05fF
C48 d0 SUB 168.00fF
C49 a_32358_n9938# SUB 6.03fF
C50 a_26978_n9909# SUB 6.03fF
C51 a_21697_n9930# SUB 6.03fF
C52 a_40634_n9457# SUB 2.20fF
C53 a_35353_n9478# SUB 2.20fF
C54 a_16149_n9946# SUB 6.03fF
C55 a_10868_n9967# SUB 6.03fF
C56 d1 SUB 85.83fF
C57 a_40630_n9645# SUB 2.33fF
C58 a_38334_n9722# SUB 2.33fF
C59 a_29973_n9449# SUB 2.20fF
C60 a_24692_n9470# SUB 2.20fF
C61 a_5488_n9938# SUB 6.03fF
C62 a_207_n9959# SUB 6.03fF
C63 a_35349_n9666# SUB 2.33fF
C64 a_38333_n9307# SUB 2.20fF
C65 a_29969_n9637# SUB 2.33fF
C66 a_27673_n9714# SUB 2.33fF
C67 a_19144_n9486# SUB 2.20fF
C68 a_13863_n9507# SUB 2.20fF
C69 a_24688_n9658# SUB 2.33fF
C70 a_22392_n9735# SUB 2.33fF
C71 a_40584_n9037# SUB 2.04fF
C72 a_19140_n9674# SUB 2.33fF
C73 a_16844_n9751# SUB 2.33fF
C74 a_8483_n9478# SUB 2.20fF
C75 a_3202_n9499# SUB 2.20fF
C76 a_35303_n9058# SUB 2.04fF
C77 d2 SUB 43.28fF
C78 a_27672_n9299# SUB 2.20fF
C79 a_13859_n9695# SUB 2.33fF
C80 a_11563_n9772# SUB 2.33fF
C81 a_29923_n9029# SUB 2.04fF
C82 a_22391_n9320# SUB 2.20fF
C83 a_24642_n9050# SUB 2.04fF
C84 a_16843_n9336# SUB 2.20fF
C85 a_8479_n9666# SUB 2.33fF
C86 a_6183_n9743# SUB 2.33fF
C87 a_3198_n9687# SUB 2.33fF
C88 a_19094_n9066# SUB 2.04fF
C89 a_11562_n9357# SUB 2.20fF
C90 a_13813_n9087# SUB 2.04fF
C91 a_6182_n9328# SUB 2.20fF
C92 a_8433_n9058# SUB 2.04fF
C93 a_901_n9349# SUB 2.20fF
C94 a_3152_n9079# SUB 2.04fF
C95 a_40639_n8476# SUB 2.20fF
C96 a_35358_n8497# SUB 2.20fF
C97 a_40635_n8664# SUB 2.33fF
C98 a_38339_n8741# SUB 2.33fF
C99 a_39302_n8803# SUB 2.04fF
C100 a_29978_n8468# SUB 2.20fF
C101 a_24697_n8489# SUB 2.20fF
C102 a_35354_n8685# SUB 2.33fF
C103 a_33058_n8762# SUB 2.33fF
C104 a_34021_n8824# SUB 2.04fF
C105 a_38338_n8326# SUB 2.20fF
C106 a_29974_n8656# SUB 2.33fF
C107 a_27678_n8733# SUB 2.33fF
C108 a_28641_n8795# SUB 2.04fF
C109 a_19149_n8505# SUB 2.20fF
C110 a_13868_n8526# SUB 2.20fF
C111 a_24693_n8677# SUB 2.33fF
C112 a_22397_n8754# SUB 2.33fF
C113 a_23360_n8816# SUB 2.04fF
C114 a_19145_n8693# SUB 2.33fF
C115 a_16849_n8770# SUB 2.33fF
C116 a_17812_n8832# SUB 2.04fF
C117 a_8488_n8497# SUB 2.20fF
C118 a_3207_n8518# SUB 2.20fF
C119 a_13864_n8714# SUB 2.33fF
C120 a_11568_n8791# SUB 2.33fF
C121 a_12531_n8853# SUB 2.04fF
C122 a_40431_n8009# SUB 2.78fF
C123 d3 SUB 20.35fF
C124 a_35150_n8030# SUB 2.78fF
C125 a_27677_n8318# SUB 2.20fF
C126 a_22396_n8339# SUB 2.20fF
C127 a_16848_n8355# SUB 2.20fF
C128 a_8484_n8685# SUB 2.33fF
C129 a_6188_n8762# SUB 2.33fF
C130 a_7151_n8824# SUB 2.04fF
C131 a_3203_n8706# SUB 2.33fF
C132 a_907_n8783# SUB 2.33fF
C133 a_1870_n8845# SUB 2.04fF
C134 a_11567_n8376# SUB 2.20fF
C135 a_39401_n8980# SUB 2.02fF
C136 a_29770_n8001# SUB 2.78fF
C137 a_24489_n8022# SUB 2.78fF
C138 a_18941_n8038# SUB 2.78fF
C139 a_13660_n8059# SUB 2.78fF
C140 a_6187_n8347# SUB 2.20fF
C141 a_34120_n9001# SUB 2.02fF
C142 a_28740_n8972# SUB 2.02fF
C143 a_23459_n8993# SUB 2.02fF
C144 a_17911_n9009# SUB 2.02fF
C145 a_8280_n8030# SUB 2.78fF
C146 a_2999_n8051# SUB 2.78fF
C147 a_12630_n9030# SUB 2.02fF
C148 a_40646_n7497# SUB 2.20fF
C149 a_35365_n7518# SUB 2.20fF
C150 a_40642_n7685# SUB 2.33fF
C151 a_38346_n7762# SUB 2.33fF
C152 a_29985_n7489# SUB 2.20fF
C153 a_24704_n7510# SUB 2.20fF
C154 a_7250_n9001# SUB 2.02fF
C155 a_1969_n9022# SUB 2.02fF
C156 a_35361_n7706# SUB 2.33fF
C157 a_40427_n8197# SUB 2.02fF
C158 a_38345_n7347# SUB 2.20fF
C159 a_29981_n7677# SUB 2.33fF
C160 a_27685_n7754# SUB 2.33fF
C161 a_19156_n7526# SUB 2.20fF
C162 a_13875_n7547# SUB 2.20fF
C163 a_24700_n7698# SUB 2.33fF
C164 a_22404_n7775# SUB 2.33fF
C165 a_40596_n7077# SUB 2.04fF
C166 a_35146_n8218# SUB 2.02fF
C167 a_19152_n7714# SUB 2.33fF
C168 a_16856_n7791# SUB 2.33fF
C169 a_8495_n7518# SUB 2.20fF
C170 a_3214_n7539# SUB 2.20fF
C171 a_35315_n7098# SUB 2.04fF
C172 a_29766_n8189# SUB 2.02fF
C173 a_27684_n7339# SUB 2.20fF
C174 a_13871_n7735# SUB 2.33fF
C175 a_11575_n7812# SUB 2.33fF
C176 a_29935_n7069# SUB 2.04fF
C177 a_24485_n8210# SUB 2.02fF
C178 a_22403_n7360# SUB 2.20fF
C179 a_24654_n7090# SUB 2.04fF
C180 a_18937_n8226# SUB 2.02fF
C181 a_16855_n7376# SUB 2.20fF
C182 a_8491_n7706# SUB 2.33fF
C183 a_6195_n7783# SUB 2.33fF
C184 a_3210_n7727# SUB 2.33fF
C185 a_19106_n7106# SUB 2.04fF
C186 a_13656_n8247# SUB 2.02fF
C187 a_11574_n7397# SUB 2.20fF
C188 a_13825_n7127# SUB 2.04fF
C189 a_39413_n7020# SUB 2.78fF
C190 a_34132_n7041# SUB 2.78fF
C191 a_28752_n7012# SUB 2.78fF
C192 a_23471_n7033# SUB 2.78fF
C193 a_8276_n8218# SUB 2.02fF
C194 a_6194_n7368# SUB 2.20fF
C195 a_8445_n7098# SUB 2.04fF
C196 a_2995_n8239# SUB 2.02fF
C197 a_913_n7389# SUB 2.20fF
C198 a_3164_n7119# SUB 2.04fF
C199 a_40651_n6516# SUB 2.20fF
C200 a_35370_n6537# SUB 2.20fF
C201 a_17923_n7049# SUB 2.78fF
C202 a_12642_n7070# SUB 2.78fF
C203 a_40647_n6704# SUB 2.33fF
C204 a_38351_n6781# SUB 2.33fF
C205 a_39314_n6843# SUB 2.04fF
C206 a_29990_n6508# SUB 2.20fF
C207 a_24709_n6529# SUB 2.20fF
C208 a_7262_n7041# SUB 2.78fF
C209 a_1981_n7062# SUB 2.78fF
C210 a_35366_n6725# SUB 2.33fF
C211 a_34033_n6864# SUB 2.04fF
C212 a_40240_n10360# SUB 4.80fF
C213 a_38350_n6366# SUB 2.20fF
C214 a_29986_n6696# SUB 2.33fF
C215 a_27690_n6773# SUB 2.33fF
C216 a_28653_n6835# SUB 2.04fF
C217 a_19161_n6545# SUB 2.20fF
C218 a_13880_n6566# SUB 2.20fF
C219 a_24705_n6717# SUB 2.33fF
C220 a_22409_n6794# SUB 2.33fF
C221 a_23372_n6856# SUB 2.04fF
C222 a_40356_n6084# SUB 3.86fF
C223 a_34959_n10381# SUB 4.80fF
C224 a_19157_n6733# SUB 2.33fF
C225 a_16861_n6810# SUB 2.33fF
C226 a_17824_n6872# SUB 2.04fF
C227 a_8500_n6537# SUB 2.20fF
C228 a_3219_n6558# SUB 2.20fF
C229 a_35075_n6105# SUB 3.86fF
C230 d4 SUB 10.50fF
C231 a_29579_n10352# SUB 4.80fF
C232 a_27689_n6358# SUB 2.20fF
C233 a_13876_n6754# SUB 2.33fF
C234 a_11580_n6831# SUB 2.33fF
C235 a_12543_n6893# SUB 2.04fF
C236 a_29695_n6076# SUB 3.86fF
C237 a_24298_n10373# SUB 4.80fF
C238 a_22408_n6379# SUB 2.20fF
C239 a_24414_n6097# SUB 3.86fF
C240 a_18750_n10389# SUB 4.80fF
C241 a_16860_n6395# SUB 2.20fF
C242 a_8496_n6725# SUB 2.33fF
C243 a_6200_n6802# SUB 2.33fF
C244 a_7163_n6864# SUB 2.04fF
C245 a_3215_n6746# SUB 2.33fF
C246 a_919_n6823# SUB 2.33fF
C247 a_1882_n6885# SUB 2.04fF
C248 a_18866_n6113# SUB 3.86fF
C249 a_13469_n10410# SUB 4.80fF
C250 a_11579_n6416# SUB 2.20fF
C251 a_13585_n6134# SUB 3.86fF
C252 a_39566_n8048# SUB 2.93fF
C253 a_39661_n6056# SUB 5.58fF
C254 a_34285_n8069# SUB 2.93fF
C255 a_34380_n6077# SUB 5.58fF
C256 a_28905_n8040# SUB 2.93fF
C257 a_29000_n6048# SUB 5.58fF
C258 a_23624_n8061# SUB 2.93fF
C259 a_23719_n6069# SUB 5.58fF
C260 a_8089_n10381# SUB 4.80fF
C261 a_6199_n6387# SUB 2.20fF
C262 a_8205_n6105# SUB 3.86fF
C263 a_2808_n10402# SUB 4.80fF
C264 a_2924_n6126# SUB 3.86fF
C265 a_40654_n5540# SUB 2.20fF
C266 a_35373_n5561# SUB 2.20fF
C267 a_18076_n8077# SUB 2.93fF
C268 a_18171_n6085# SUB 5.58fF
C269 a_12795_n8098# SUB 2.93fF
C270 a_12890_n6106# SUB 5.58fF
C271 a_40650_n5728# SUB 2.33fF
C272 a_38354_n5805# SUB 2.33fF
C273 a_29993_n5532# SUB 2.20fF
C274 a_24712_n5553# SUB 2.20fF
C275 a_7415_n8069# SUB 2.93fF
C276 a_7510_n6077# SUB 5.58fF
C277 a_2134_n8090# SUB 2.93fF
C278 a_2229_n6098# SUB 5.58fF
C279 a_35369_n5749# SUB 2.33fF
C280 a_38353_n5390# SUB 2.20fF
C281 a_29989_n5720# SUB 2.33fF
C282 a_27693_n5797# SUB 2.33fF
C283 a_19164_n5569# SUB 2.20fF
C284 a_13883_n5590# SUB 2.20fF
C285 a_24708_n5741# SUB 2.33fF
C286 a_22412_n5818# SUB 2.33fF
C287 a_40604_n5120# SUB 2.04fF
C288 a_19160_n5757# SUB 2.33fF
C289 a_16864_n5834# SUB 2.33fF
C290 a_8503_n5561# SUB 2.20fF
C291 a_3222_n5582# SUB 2.20fF
C292 a_35323_n5141# SUB 2.04fF
C293 a_27692_n5382# SUB 2.20fF
C294 a_13879_n5778# SUB 2.33fF
C295 a_11583_n5855# SUB 2.33fF
C296 a_29943_n5112# SUB 2.04fF
C297 a_22411_n5403# SUB 2.20fF
C298 a_24662_n5133# SUB 2.04fF
C299 a_16863_n5419# SUB 2.20fF
C300 a_8499_n5749# SUB 2.33fF
C301 a_6203_n5826# SUB 2.33fF
C302 a_3218_n5770# SUB 2.33fF
C303 a_19114_n5149# SUB 2.04fF
C304 a_11582_n5440# SUB 2.20fF
C305 a_13833_n5170# SUB 2.04fF
C306 a_6202_n5411# SUB 2.20fF
C307 a_8453_n5141# SUB 2.04fF
C308 a_921_n5432# SUB 2.20fF
C309 a_3172_n5162# SUB 2.04fF
C310 a_40659_n4559# SUB 2.20fF
C311 a_35378_n4580# SUB 2.20fF
C312 a_40655_n4747# SUB 2.33fF
C313 a_38359_n4824# SUB 2.33fF
C314 a_39322_n4886# SUB 2.04fF
C315 a_29998_n4551# SUB 2.20fF
C316 a_24717_n4572# SUB 2.20fF
C317 a_35374_n4768# SUB 2.33fF
C318 a_34041_n4907# SUB 2.04fF
C319 a_38358_n4409# SUB 2.20fF
C320 a_29994_n4739# SUB 2.33fF
C321 a_27698_n4816# SUB 2.33fF
C322 a_28661_n4878# SUB 2.04fF
C323 a_19169_n4588# SUB 2.20fF
C324 a_13888_n4609# SUB 2.20fF
C325 a_24713_n4760# SUB 2.33fF
C326 a_22417_n4837# SUB 2.33fF
C327 a_23380_n4899# SUB 2.04fF
C328 a_19165_n4776# SUB 2.33fF
C329 a_16869_n4853# SUB 2.33fF
C330 a_17832_n4915# SUB 2.04fF
C331 a_8508_n4580# SUB 2.20fF
C332 a_3227_n4601# SUB 2.20fF
C333 a_13884_n4797# SUB 2.33fF
C334 a_11588_n4874# SUB 2.33fF
C335 a_12551_n4936# SUB 2.04fF
C336 a_40352_n6272# SUB 2.93fF
C337 a_40451_n4092# SUB 2.78fF
C338 a_35071_n6293# SUB 2.93fF
C339 a_35170_n4113# SUB 2.78fF
C340 a_27697_n4401# SUB 2.20fF
C341 a_22416_n4422# SUB 2.20fF
C342 a_16868_n4438# SUB 2.20fF
C343 a_8504_n4768# SUB 2.33fF
C344 a_6208_n4845# SUB 2.33fF
C345 a_7171_n4907# SUB 2.04fF
C346 a_3223_n4789# SUB 2.33fF
C347 a_1890_n4928# SUB 2.04fF
C348 a_11587_n4459# SUB 2.20fF
C349 a_39421_n5063# SUB 2.02fF
C350 a_39562_n5879# SUB 3.86fF
C351 a_29691_n6264# SUB 2.93fF
C352 a_29790_n4084# SUB 2.78fF
C353 a_24410_n6285# SUB 2.93fF
C354 a_24509_n4105# SUB 2.78fF
C355 a_18862_n6301# SUB 2.93fF
C356 a_18961_n4121# SUB 2.78fF
C357 a_13581_n6322# SUB 2.93fF
C358 a_13680_n4142# SUB 2.78fF
C359 a_6207_n4430# SUB 2.20fF
C360 a_926_n4451# SUB 2.20fF
C361 a_34140_n5084# SUB 2.02fF
C362 a_34281_n5900# SUB 3.86fF
C363 a_28760_n5055# SUB 2.02fF
C364 a_28901_n5871# SUB 3.86fF
C365 a_23479_n5076# SUB 2.02fF
C366 a_23620_n5892# SUB 3.86fF
C367 a_17931_n5092# SUB 2.02fF
C368 a_18072_n5908# SUB 3.86fF
C369 a_8201_n6293# SUB 2.93fF
C370 a_8300_n4113# SUB 2.78fF
C371 a_2920_n6314# SUB 2.93fF
C372 a_3019_n4134# SUB 2.78fF
C373 a_12650_n5113# SUB 2.02fF
C374 a_12791_n5929# SUB 3.86fF
C375 a_40666_n3580# SUB 2.20fF
C376 a_35385_n3601# SUB 2.20fF
C377 a_40662_n3768# SUB 2.33fF
C378 a_38366_n3845# SUB 2.33fF
C379 a_30005_n3572# SUB 2.20fF
C380 a_24724_n3593# SUB 2.20fF
C381 a_7270_n5084# SUB 2.02fF
C382 a_7411_n5900# SUB 3.86fF
C383 a_1989_n5105# SUB 2.02fF
C384 a_2130_n5921# SUB 3.86fF
C385 a_35381_n3789# SUB 2.33fF
C386 a_33085_n3866# SUB 2.33fF
C387 a_40447_n4280# SUB 2.02fF
C388 a_38365_n3430# SUB 2.20fF
C389 a_30001_n3760# SUB 2.33fF
C390 a_27705_n3837# SUB 2.33fF
C391 a_19176_n3609# SUB 2.20fF
C392 a_13895_n3630# SUB 2.20fF
C393 a_24720_n3781# SUB 2.33fF
C394 a_22424_n3858# SUB 2.33fF
C395 a_40616_n3160# SUB 2.04fF
C396 a_35166_n4301# SUB 2.02fF
C397 a_19172_n3797# SUB 2.33fF
C398 a_16876_n3874# SUB 2.33fF
C399 a_8515_n3601# SUB 2.20fF
C400 a_3234_n3622# SUB 2.20fF
C401 a_35335_n3181# SUB 2.04fF
C402 a_29786_n4272# SUB 2.02fF
C403 a_27704_n3422# SUB 2.20fF
C404 a_13891_n3818# SUB 2.33fF
C405 a_11595_n3895# SUB 2.33fF
C406 a_29955_n3152# SUB 2.04fF
C407 a_24505_n4293# SUB 2.02fF
C408 a_22423_n3443# SUB 2.20fF
C409 a_24674_n3173# SUB 2.04fF
C410 a_18957_n4309# SUB 2.02fF
C411 a_16875_n3459# SUB 2.20fF
C412 a_8511_n3789# SUB 2.33fF
C413 a_6215_n3866# SUB 2.33fF
C414 a_3230_n3810# SUB 2.33fF
C415 a_934_n3887# SUB 2.33fF
C416 a_19126_n3189# SUB 2.04fF
C417 a_13676_n4330# SUB 2.02fF
C418 a_11594_n3480# SUB 2.20fF
C419 a_13845_n3210# SUB 2.04fF
C420 a_39433_n3103# SUB 2.78fF
C421 a_34152_n3124# SUB 2.78fF
C422 a_28772_n3095# SUB 2.78fF
C423 a_23491_n3116# SUB 2.78fF
C424 a_8296_n4301# SUB 2.02fF
C425 a_6214_n3451# SUB 2.20fF
C426 a_8465_n3181# SUB 2.04fF
C427 a_3015_n4322# SUB 2.02fF
C428 a_3184_n3202# SUB 2.04fF
C429 a_40671_n2599# SUB 2.20fF
C430 a_35390_n2620# SUB 2.20fF
C431 a_17943_n3132# SUB 2.78fF
C432 a_12662_n3153# SUB 2.78fF
C433 a_40667_n2787# SUB 2.33fF
C434 a_38371_n2864# SUB 2.33fF
C435 a_39334_n2926# SUB 2.04fF
C436 a_30010_n2591# SUB 2.20fF
C437 a_24729_n2612# SUB 2.20fF
C438 a_7282_n3124# SUB 2.78fF
C439 a_2001_n3145# SUB 2.78fF
C440 a_35386_n2808# SUB 2.33fF
C441 a_34053_n2947# SUB 2.04fF
C442 a_30006_n2779# SUB 2.33fF
C443 a_27710_n2856# SUB 2.33fF
C444 a_28673_n2918# SUB 2.04fF
C445 a_19181_n2628# SUB 2.20fF
C446 a_13900_n2649# SUB 2.20fF
C447 a_24725_n2800# SUB 2.33fF
C448 a_22429_n2877# SUB 2.33fF
C449 a_23392_n2939# SUB 2.04fF
C450 a_19177_n2816# SUB 2.33fF
C451 a_16881_n2893# SUB 2.33fF
C452 a_17844_n2955# SUB 2.04fF
C453 a_8520_n2620# SUB 2.20fF
C454 a_3239_n2641# SUB 2.20fF
C455 a_13896_n2837# SUB 2.33fF
C456 a_11600_n2914# SUB 2.33fF
C457 a_12563_n2976# SUB 2.04fF
C458 a_38370_n2449# SUB 2.20fF
C459 a_8516_n2808# SUB 2.33fF
C460 a_6220_n2885# SUB 2.33fF
C461 a_7183_n2947# SUB 2.04fF
C462 a_3235_n2829# SUB 2.33fF
C463 a_1902_n2968# SUB 2.04fF
C464 a_37332_n2231# SUB 2.33fF
C465 a_27709_n2441# SUB 2.20fF
C466 a_22428_n2462# SUB 2.20fF
C467 a_16880_n2478# SUB 2.20fF
C468 a_11599_n2499# SUB 2.20fF
C469 a_31952_n2202# SUB 2.47fF
C470 a_26671_n2223# SUB 2.33fF
C471 a_21123_n2239# SUB 2.66fF
C472 a_15842_n2260# SUB 2.33fF
C473 a_6219_n2470# SUB 2.20fF
C474 a_938_n2491# SUB 2.20fF
C475 a_10462_n2231# SUB 2.47fF
C476 a_5181_n2252# SUB 2.33fF
C477 a_20848_n805# SUB 10.76fF
C478 a_37394_271# SUB 3.05fF
C479 a_31994_256# SUB 6.01fF
C480 a_34403_359# SUB 4.48fF
C481 a_26733_263# SUB 3.05fF
C482 a_26832_263# SUB 6.47fF
C483 a_20996_141# SUB 12.03fF
C484 a_23742_351# SUB 4.48fF
C485 a_15904_300# SUB 3.05fF
C486 a_10504_285# SUB 6.01fF
C487 a_10603_285# SUB 12.33fF
C488 a_12913_388# SUB 4.48fF
C489 a_5243_292# SUB 3.05fF
C490 a_5342_292# SUB 6.47fF
C491 a_2252_380# SUB 4.48fF
C492 a_32313_855# SUB 6.03fF
C493 a_38281_819# SUB 2.20fF
C494 a_40578_1334# SUB 2.33fF
C495 a_38282_1234# SUB 2.33fF
C496 a_33000_840# SUB 2.20fF
C497 a_21652_847# SUB 6.03fF
C498 a_27620_811# SUB 2.20fF
C499 a_35297_1355# SUB 2.33fF
C500 a_40582_1157# SUB 2.20fF
C501 a_33001_1255# SUB 2.33fF
C502 a_16104_863# SUB 6.03fF
C503 a_29917_1326# SUB 2.33fF
C504 a_27621_1226# SUB 2.33fF
C505 a_22339_832# SUB 2.20fF
C506 a_10823_884# SUB 6.03fF
C507 a_24636_1347# SUB 2.33fF
C508 a_39245_1473# SUB 2.04fF
C509 a_35301_1178# SUB 2.20fF
C510 a_33964_1494# SUB 2.04fF
C511 a_29921_1149# SUB 2.20fF
C512 a_22340_1247# SUB 2.33fF
C513 a_16791_848# SUB 2.20fF
C514 a_19088_1363# SUB 2.33fF
C515 a_28584_1465# SUB 2.04fF
C516 a_24640_1170# SUB 2.20fF
C517 a_16792_1263# SUB 2.33fF
C518 a_11510_869# SUB 2.20fF
C519 a_162_876# SUB 6.03fF
C520 a_6130_840# SUB 2.20fF
C521 a_13807_1384# SUB 2.33fF
C522 a_23303_1486# SUB 2.04fF
C523 a_19092_1186# SUB 2.20fF
C524 a_11511_1284# SUB 2.33fF
C525 a_8427_1355# SUB 2.33fF
C526 a_6131_1255# SUB 2.33fF
C527 a_849_861# SUB 2.20fF
C528 a_3146_1376# SUB 2.33fF
C529 a_17755_1502# SUB 2.04fF
C530 a_13811_1207# SUB 2.20fF
C531 a_12474_1523# SUB 2.04fF
C532 a_8431_1178# SUB 2.20fF
C533 a_7094_1494# SUB 2.04fF
C534 a_3150_1199# SUB 2.20fF
C535 a_1813_1515# SUB 2.04fF
C536 a_38276_1800# SUB 2.20fF
C537 a_40527_1718# SUB 2.04fF
C538 a_40573_2315# SUB 2.33fF
C539 a_38277_2215# SUB 2.33fF
C540 a_32995_1821# SUB 2.20fF
C541 a_35246_1739# SUB 2.04fF
C542 a_27615_1792# SUB 2.20fF
C543 a_35292_2336# SUB 2.33fF
C544 a_32996_2236# SUB 2.33fF
C545 a_29866_1710# SUB 2.04fF
C546 a_29912_2307# SUB 2.33fF
C547 a_27616_2207# SUB 2.33fF
C548 a_22334_1813# SUB 2.20fF
C549 a_24585_1731# SUB 2.04fF
C550 a_24631_2328# SUB 2.33fF
C551 a_40577_2138# SUB 2.20fF
C552 a_39344_1473# SUB 2.78fF
C553 a_35296_2159# SUB 2.20fF
C554 a_22335_2228# SUB 2.33fF
C555 a_16786_1829# SUB 2.20fF
C556 a_19037_1747# SUB 2.04fF
C557 a_19083_2344# SUB 2.33fF
C558 a_29916_2130# SUB 2.20fF
C559 a_16787_2244# SUB 2.33fF
C560 a_11505_1850# SUB 2.20fF
C561 a_13756_1768# SUB 2.04fF
C562 a_6125_1821# SUB 2.20fF
C563 a_13802_2365# SUB 2.33fF
C564 a_34063_1494# SUB 2.78fF
C565 a_28683_1465# SUB 2.78fF
C566 a_24635_2151# SUB 2.20fF
C567 a_11506_2265# SUB 2.33fF
C568 a_8376_1739# SUB 2.04fF
C569 a_8422_2336# SUB 2.33fF
C570 a_6126_2236# SUB 2.33fF
C571 a_844_1842# SUB 2.20fF
C572 a_3095_1760# SUB 2.04fF
C573 a_3141_2357# SUB 2.33fF
C574 a_40358_2827# SUB 2.02fF
C575 a_35077_2848# SUB 2.02fF
C576 a_23402_1486# SUB 2.78fF
C577 a_19087_2167# SUB 2.20fF
C578 a_29697_2819# SUB 2.02fF
C579 a_17854_1502# SUB 2.78fF
C580 a_13806_2188# SUB 2.20fF
C581 a_8426_2159# SUB 2.20fF
C582 a_38269_2779# SUB 2.20fF
C583 a_24416_2840# SUB 2.02fF
C584 a_12573_1523# SUB 2.78fF
C585 a_7193_1494# SUB 2.78fF
C586 a_3145_2180# SUB 2.20fF
C587 a_40566_3294# SUB 2.33fF
C588 a_38270_3194# SUB 2.33fF
C589 a_32988_2800# SUB 2.20fF
C590 a_18868_2856# SUB 2.02fF
C591 a_27608_2771# SUB 2.20fF
C592 a_35285_3315# SUB 2.33fF
C593 a_40570_3117# SUB 2.20fF
C594 a_32989_3215# SUB 2.33fF
C595 a_13587_2877# SUB 2.02fF
C596 a_1912_1515# SUB 2.78fF
C597 a_8207_2848# SUB 2.02fF
C598 a_29905_3286# SUB 2.33fF
C599 a_27609_3186# SUB 2.33fF
C600 a_22327_2792# SUB 2.20fF
C601 a_24624_3307# SUB 2.33fF
C602 a_39233_3433# SUB 2.04fF
C603 a_39332_3433# SUB 2.02fF
C604 a_35289_3138# SUB 2.20fF
C605 a_33952_3454# SUB 2.04fF
C606 a_34051_3454# SUB 2.02fF
C607 a_29909_3109# SUB 2.20fF
C608 a_22328_3207# SUB 2.33fF
C609 a_16779_2808# SUB 2.20fF
C610 a_2926_2869# SUB 2.02fF
C611 a_19076_3323# SUB 2.33fF
C612 a_28572_3425# SUB 2.04fF
C613 a_28671_3425# SUB 2.02fF
C614 a_24628_3130# SUB 2.20fF
C615 a_16780_3223# SUB 2.33fF
C616 a_11498_2829# SUB 2.20fF
C617 a_6118_2800# SUB 2.20fF
C618 a_13795_3344# SUB 2.33fF
C619 a_23291_3446# SUB 2.04fF
C620 a_23390_3446# SUB 2.02fF
C621 a_19080_3146# SUB 2.20fF
C622 a_11499_3244# SUB 2.33fF
C623 a_8415_3315# SUB 2.33fF
C624 a_6119_3215# SUB 2.33fF
C625 a_837_2821# SUB 2.20fF
C626 a_3134_3336# SUB 2.33fF
C627 a_40362_2650# SUB 2.78fF
C628 a_17743_3462# SUB 2.04fF
C629 a_17842_3462# SUB 2.02fF
C630 a_13799_3167# SUB 2.20fF
C631 a_35081_2671# SUB 2.78fF
C632 a_29701_2642# SUB 2.78fF
C633 a_12462_3483# SUB 2.04fF
C634 a_12561_3483# SUB 2.02fF
C635 a_8419_3138# SUB 2.20fF
C636 a_838_3236# SUB 2.33fF
C637 a_7082_3454# SUB 2.04fF
C638 a_7181_3454# SUB 2.02fF
C639 a_3138_3159# SUB 2.20fF
C640 a_1801_3475# SUB 2.04fF
C641 a_1900_3475# SUB 2.02fF
C642 a_38264_3760# SUB 2.20fF
C643 a_24420_2663# SUB 2.78fF
C644 a_40515_3678# SUB 2.04fF
C645 a_40561_4275# SUB 2.33fF
C646 a_38265_4175# SUB 2.33fF
C647 a_32983_3781# SUB 2.20fF
C648 a_18872_2679# SUB 2.78fF
C649 a_35234_3699# SUB 2.04fF
C650 a_27603_3752# SUB 2.20fF
C651 a_35280_4296# SUB 2.33fF
C652 a_32984_4196# SUB 2.33fF
C653 a_29854_3670# SUB 2.04fF
C654 a_13591_2700# SUB 2.78fF
C655 a_8211_2671# SUB 2.78fF
C656 a_29900_4267# SUB 2.33fF
C657 a_27604_4167# SUB 2.33fF
C658 a_22322_3773# SUB 2.20fF
C659 a_24573_3691# SUB 2.04fF
C660 a_24619_4288# SUB 2.33fF
C661 a_40565_4098# SUB 2.20fF
C662 a_39473_4426# SUB 3.86fF
C663 a_39572_4426# SUB 4.80fF
C664 a_35284_4119# SUB 2.20fF
C665 a_22323_4188# SUB 2.33fF
C666 a_16774_3789# SUB 2.20fF
C667 a_2930_2692# SUB 2.78fF
C668 a_19025_3707# SUB 2.04fF
C669 a_19071_4304# SUB 2.33fF
C670 a_39585_338# SUB 5.58fF
C671 a_40263_4819# SUB 2.93fF
C672 a_34192_4447# SUB 3.86fF
C673 a_34291_4447# SUB 4.80fF
C674 a_29904_4090# SUB 2.20fF
C675 a_28812_4418# SUB 3.86fF
C676 a_28911_4418# SUB 4.80fF
C677 a_16775_4204# SUB 2.33fF
C678 a_11493_3810# SUB 2.20fF
C679 a_13744_3728# SUB 2.04fF
C680 a_6113_3781# SUB 2.20fF
C681 a_13790_4325# SUB 2.33fF
C682 a_24623_4111# SUB 2.20fF
C683 a_34304_359# SUB 5.58fF
C684 a_34982_4840# SUB 2.93fF
C685 a_28924_330# SUB 5.58fF
C686 a_29602_4811# SUB 2.93fF
C687 a_23531_4439# SUB 3.86fF
C688 a_23630_4439# SUB 4.80fF
C689 a_11494_4225# SUB 2.33fF
C690 a_8364_3699# SUB 2.04fF
C691 a_8410_4296# SUB 2.33fF
C692 a_6114_4196# SUB 2.33fF
C693 a_832_3802# SUB 2.20fF
C694 a_3083_3720# SUB 2.04fF
C695 a_3129_4317# SUB 2.33fF
C696 a_19075_4127# SUB 2.20fF
C697 a_38261_4736# SUB 2.20fF
C698 a_23643_351# SUB 5.58fF
C699 a_24321_4832# SUB 2.93fF
C700 a_17983_4455# SUB 3.86fF
C701 a_18082_4455# SUB 4.80fF
C702 a_13794_4148# SUB 2.20fF
C703 a_40558_5251# SUB 2.33fF
C704 a_38262_5151# SUB 2.33fF
C705 a_32980_4757# SUB 2.20fF
C706 a_18095_367# SUB 5.58fF
C707 a_18773_4848# SUB 2.93fF
C708 a_12702_4476# SUB 3.86fF
C709 a_12801_4476# SUB 4.80fF
C710 a_8414_4119# SUB 2.20fF
C711 a_7322_4447# SUB 3.86fF
C712 a_7421_4447# SUB 4.80fF
C713 a_3133_4140# SUB 2.20fF
C714 a_27600_4728# SUB 2.20fF
C715 a_35277_5272# SUB 2.33fF
C716 a_40562_5074# SUB 2.20fF
C717 a_32981_5172# SUB 2.33fF
C718 a_12814_388# SUB 5.58fF
C719 a_13492_4869# SUB 2.93fF
C720 a_7434_359# SUB 5.58fF
C721 a_8112_4840# SUB 2.93fF
C722 a_2041_4468# SUB 3.86fF
C723 a_2140_4468# SUB 4.80fF
C724 a_29897_5243# SUB 2.33fF
C725 a_27601_5143# SUB 2.33fF
C726 a_22319_4749# SUB 2.20fF
C727 a_24616_5264# SUB 2.33fF
C728 a_39225_5390# SUB 2.04fF
C729 a_35281_5095# SUB 2.20fF
C730 a_33944_5411# SUB 2.04fF
C731 a_29901_5066# SUB 2.20fF
C732 a_22320_5164# SUB 2.33fF
C733 a_16771_4765# SUB 2.20fF
C734 a_2153_380# SUB 5.58fF
C735 a_2831_4861# SUB 2.93fF
C736 a_19068_5280# SUB 2.33fF
C737 a_28564_5382# SUB 2.04fF
C738 a_24620_5087# SUB 2.20fF
C739 a_16772_5180# SUB 2.33fF
C740 a_11490_4786# SUB 2.20fF
C741 a_6110_4757# SUB 2.20fF
C742 a_13787_5301# SUB 2.33fF
C743 a_23283_5403# SUB 2.04fF
C744 a_19072_5103# SUB 2.20fF
C745 a_11491_5201# SUB 2.33fF
C746 a_8407_5272# SUB 2.33fF
C747 a_6111_5172# SUB 2.33fF
C748 a_829_4778# SUB 2.20fF
C749 a_3126_5293# SUB 2.33fF
C750 a_17735_5419# SUB 2.04fF
C751 a_13791_5124# SUB 2.20fF
C752 a_12454_5440# SUB 2.04fF
C753 a_8411_5095# SUB 2.20fF
C754 a_7074_5411# SUB 2.04fF
C755 a_3130_5116# SUB 2.20fF
C756 a_1793_5432# SUB 2.04fF
C757 a_38256_5717# SUB 2.20fF
C758 a_40507_5635# SUB 2.04fF
C759 a_40553_6232# SUB 2.33fF
C760 a_38257_6132# SUB 2.33fF
C761 a_32975_5738# SUB 2.20fF
C762 a_35226_5656# SUB 2.04fF
C763 a_27595_5709# SUB 2.20fF
C764 a_35272_6253# SUB 2.33fF
C765 a_32976_6153# SUB 2.33fF
C766 a_29846_5627# SUB 2.04fF
C767 a_29892_6224# SUB 2.33fF
C768 a_27596_6124# SUB 2.33fF
C769 a_22314_5730# SUB 2.20fF
C770 a_24565_5648# SUB 2.04fF
C771 a_24611_6245# SUB 2.33fF
C772 a_40557_6055# SUB 2.20fF
C773 a_39324_5390# SUB 2.78fF
C774 a_39477_6418# SUB 2.93fF
C775 a_35276_6076# SUB 2.20fF
C776 a_22315_6145# SUB 2.33fF
C777 a_16766_5746# SUB 2.20fF
C778 a_19017_5664# SUB 2.04fF
C779 a_19063_6261# SUB 2.33fF
C780 a_29896_6047# SUB 2.20fF
C781 a_16767_6161# SUB 2.33fF
C782 a_11485_5767# SUB 2.20fF
C783 a_13736_5685# SUB 2.04fF
C784 a_6105_5738# SUB 2.20fF
C785 a_13782_6282# SUB 2.33fF
C786 a_34043_5411# SUB 2.78fF
C787 a_34196_6439# SUB 2.93fF
C788 a_28663_5382# SUB 2.78fF
C789 a_28816_6410# SUB 2.93fF
C790 a_24615_6068# SUB 2.20fF
C791 a_11486_6182# SUB 2.33fF
C792 a_8356_5656# SUB 2.04fF
C793 a_8402_6253# SUB 2.33fF
C794 a_6106_6153# SUB 2.33fF
C795 a_3075_5677# SUB 2.04fF
C796 a_3121_6274# SUB 2.33fF
C797 a_40267_4642# SUB 3.86fF
C798 a_40338_6744# SUB 2.02fF
C799 a_34986_4663# SUB 3.86fF
C800 a_35057_6765# SUB 2.02fF
C801 a_23382_5403# SUB 2.78fF
C802 a_23535_6431# SUB 2.93fF
C803 a_19067_6084# SUB 2.20fF
C804 a_29606_4634# SUB 3.86fF
C805 a_29677_6736# SUB 2.02fF
C806 a_17834_5419# SUB 2.78fF
C807 a_17987_6447# SUB 2.93fF
C808 a_13786_6105# SUB 2.20fF
C809 a_8406_6076# SUB 2.20fF
C810 a_38249_6696# SUB 2.20fF
C811 a_24325_4655# SUB 3.86fF
C812 a_24396_6757# SUB 2.02fF
C813 a_12553_5440# SUB 2.78fF
C814 a_12706_6468# SUB 2.93fF
C815 a_7173_5411# SUB 2.78fF
C816 a_7326_6439# SUB 2.93fF
C817 a_3125_6097# SUB 2.20fF
C818 a_40546_7211# SUB 2.33fF
C819 a_38250_7111# SUB 2.33fF
C820 a_32968_6717# SUB 2.20fF
C821 a_18777_4671# SUB 3.86fF
C822 a_18848_6773# SUB 2.02fF
C823 a_27588_6688# SUB 2.20fF
C824 a_35265_7232# SUB 2.33fF
C825 a_40550_7034# SUB 2.20fF
C826 a_32969_7132# SUB 2.33fF
C827 a_13496_4692# SUB 3.86fF
C828 a_13567_6794# SUB 2.02fF
C829 a_1892_5432# SUB 2.78fF
C830 a_2045_6460# SUB 2.93fF
C831 a_8116_4663# SUB 3.86fF
C832 a_8187_6765# SUB 2.02fF
C833 a_29885_7203# SUB 2.33fF
C834 a_27589_7103# SUB 2.33fF
C835 a_22307_6709# SUB 2.20fF
C836 a_24604_7224# SUB 2.33fF
C837 a_39213_7350# SUB 2.04fF
C838 a_39312_7350# SUB 2.02fF
C839 a_35269_7055# SUB 2.20fF
C840 a_33932_7371# SUB 2.04fF
C841 a_34031_7371# SUB 2.02fF
C842 a_29889_7026# SUB 2.20fF
C843 a_22308_7124# SUB 2.33fF
C844 a_16759_6725# SUB 2.20fF
C845 a_2835_4684# SUB 3.86fF
C846 a_2906_6786# SUB 2.02fF
C847 a_19056_7240# SUB 2.33fF
C848 a_28552_7342# SUB 2.04fF
C849 a_28651_7342# SUB 2.02fF
C850 a_24608_7047# SUB 2.20fF
C851 a_16760_7140# SUB 2.33fF
C852 a_11478_6746# SUB 2.20fF
C853 a_6098_6717# SUB 2.20fF
C854 a_13775_7261# SUB 2.33fF
C855 a_23271_7363# SUB 2.04fF
C856 a_23370_7363# SUB 2.02fF
C857 a_19060_7063# SUB 2.20fF
C858 a_11479_7161# SUB 2.33fF
C859 a_8395_7232# SUB 2.33fF
C860 a_6099_7132# SUB 2.33fF
C861 a_817_6738# SUB 2.20fF
C862 a_3114_7253# SUB 2.33fF
C863 a_40342_6567# SUB 2.78fF
C864 a_17723_7379# SUB 2.04fF
C865 a_17822_7379# SUB 2.02fF
C866 a_13779_7084# SUB 2.20fF
C867 a_35061_6588# SUB 2.78fF
C868 a_29681_6559# SUB 2.78fF
C869 a_12442_7400# SUB 2.04fF
C870 a_12541_7400# SUB 2.02fF
C871 a_8399_7055# SUB 2.20fF
C872 a_818_7153# SUB 2.33fF
C873 a_7062_7371# SUB 2.04fF
C874 a_7161_7371# SUB 2.02fF
C875 a_3118_7076# SUB 2.20fF
C876 a_1781_7392# SUB 2.04fF
C877 a_1880_7392# SUB 2.02fF
C878 a_38244_7677# SUB 2.20fF
C879 a_24400_6580# SUB 2.78fF
C880 a_40495_7595# SUB 2.04fF
C881 a_40541_8192# SUB 2.33fF
C882 a_38245_8092# SUB 2.33fF
C883 a_32963_7698# SUB 2.20fF
C884 a_18852_6596# SUB 2.78fF
C885 a_35214_7616# SUB 2.04fF
C886 a_27583_7669# SUB 2.20fF
C887 a_35260_8213# SUB 2.33fF
C888 a_32964_8113# SUB 2.33fF
C889 a_29834_7587# SUB 2.04fF
C890 a_13571_6617# SUB 2.78fF
C891 a_8191_6588# SUB 2.78fF
C892 a_29880_8184# SUB 2.33fF
C893 a_27584_8084# SUB 2.33fF
C894 a_22302_7690# SUB 2.20fF
C895 a_24553_7608# SUB 2.04fF
C896 a_24599_8205# SUB 2.33fF
C897 a_40545_8015# SUB 2.20fF
C898 a_36277_8270# SUB 2.33fF
C899 a_35264_8036# SUB 2.20fF
C900 a_22303_8105# SUB 2.33fF
C901 a_16754_7706# SUB 2.20fF
C902 a_2910_6609# SUB 2.78fF
C903 a_19005_7624# SUB 2.04fF
C904 a_19051_8221# SUB 2.33fF
C905 a_29884_8007# SUB 2.20fF
C906 a_30897_8241# SUB 2.47fF
C907 a_16755_8121# SUB 2.33fF
C908 a_11473_7727# SUB 2.20fF
C909 a_13724_7645# SUB 2.04fF
C910 a_6093_7698# SUB 2.20fF
C911 a_13770_8242# SUB 2.33fF
C912 a_25616_8262# SUB 2.33fF
C913 a_24603_8028# SUB 2.20fF
C914 a_11474_8142# SUB 2.33fF
C915 a_8344_7616# SUB 2.04fF
C916 a_8390_8213# SUB 2.33fF
C917 a_6094_8113# SUB 2.33fF
C918 a_812_7719# SUB 2.20fF
C919 a_3063_7637# SUB 2.04fF
C920 a_3109_8234# SUB 2.33fF
C921 a_20068_8278# SUB 2.66fF
C922 a_19055_8044# SUB 2.20fF
C923 a_14787_8299# SUB 2.33fF
C924 a_13774_8065# SUB 2.20fF
C925 a_813_8134# SUB 2.33fF
C926 a_8394_8036# SUB 2.20fF
C927 a_4126_8291# SUB 2.33fF
C928 a_3113_8057# SUB 2.20fF
C929 vout gnd 50fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0 0.1ps 0.1ps 5us 10us)
Vd1 d1 0 pulse(0 1.8 0 0.1ps 0.1ps 10us 20us)
Vd2 d2 0 pulse(0 1.8 0 0.1ps 0.1ps 20us 40us)
Vd3 d3 0 pulse(0 1.8 0 0.1ps 0.1ps 40us 80us)
Vd4 d4 0 pulse(0 1.8 0 0.1ps 0.1ps 80us 160us)
Vd5 d5 0 pulse(0 1.8 0 0.1ps 0.1ps 160us 320us)
Vd6 d6 0 pulse(0 1.8 0 0.1ps 0.1ps 320us 640us)
Vd7 d7 0 pulse(0 1.8 0 0.1ps 0.1ps 640us 1280us)
Vd8 d8 0 pulse(0 1.8 0 0.1ps 0.1ps 1280us 2560us)
Vd9 d9 0 pulse(0 1.8 0 0.1ps 0.1ps 2560us 5120us)

.tran 20us 5120us
.control
run
plot V(vout)
.endc
.end
