* SPICE3 file created from 10bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 a_6539_3037# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1 a_37081_7554# a_36784_8525# a_37064_9117# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2 a_39093_6841# a_39099_6115# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3 a_24010_n8233# a_24006_n8421# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4 a_15735_n3462# a_15522_n3462# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5 vdd a_23217_n5945# a_23009_n5945# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6 a_17830_n4910# a_18087_n4926# a_17865_n3606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7 a_35707_n3992# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8 a_36125_n9507# a_35704_n9507# a_35390_n9054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9 a_10149_n6639# a_10678_n6730# a_10886_n6730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X10 a_17972_n9645# a_18956_n10159# a_18907_n10143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X11 a_17975_2515# a_18959_2812# a_18910_3002# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X12 a_20303_n8821# a_20303_n8592# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X13 a_24964_n10698# a_30219_n10835# a_20533_n10895# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X14 gnd a_39352_3342# a_39144_3342# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X15 gnd d0 a_34295_n8996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X16 vdd d1 a_38413_4689# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X17 a_2887_4675# a_3871_4972# a_3826_4985# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X18 a_15205_n6451# a_15205_n6221# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X19 gnd a_29322_n4620# a_29114_n4620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X20 a_25675_8253# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X21 a_117_7425# a_117_7238# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X22 a_3822_6265# a_4079_6075# a_2887_5778# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X23 a_38018_n9115# a_38203_n9830# a_38154_n9814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X24 a_21979_4659# a_21558_4659# a_21041_4903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X25 gnd d0 a_24265_n4025# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X26 a_32991_3211# a_33248_3021# a_32991_5411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X27 a_30651_n5608# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X28 a_3827_n1634# a_3823_n1822# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X29 a_15940_6620# a_16671_6930# a_16879_6930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X30 vdd d0 a_19165_n5193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X31 a_8880_n8293# a_9133_n8497# a_7938_n8725# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X32 a_20305_n4596# a_20305_n4409# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X33 a_25889_n6747# a_25676_n6747# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X34 a_119_n3969# a_647_n3965# a_855_n3965# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X35 a_6859_n5772# a_6539_n3737# a_6861_n3560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X36 a_21558_5762# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X37 a_6640_n8728# a_6427_n8728# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X38 a_5490_n4006# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X39 a_36646_3602# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X40 gnd a_8194_n9844# a_7986_n9844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X41 vdd d0 a_4080_n1838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X42 a_18911_7786# a_19164_7773# a_17969_8207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X43 a_11616_n5383# a_11403_n5383# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X44 a_434_3265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X45 vdd d4 a_38304_n5991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X46 a_34042_7177# a_34295_7164# a_33103_6867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X47 a_16812_6338# a_16599_6338# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X48 a_30335_6121# a_30864_6011# a_31072_6011# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X49 a_30865_n4505# a_30652_n4505# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X50 a_5491_n4560# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X51 a_32020_5194# a_31700_2982# a_32022_2982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X52 vdd d6 a_4936_n10733# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X53 a_21556_9071# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X54 a_35389_9242# a_35389_9012# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X55 a_17973_6927# a_18957_7224# a_18912_7237# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X56 a_36644_6911# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X57 vdd d0 a_14109_4423# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X58 a_11402_n8692# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X59 a_20302_n10111# a_24006_n10078# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X60 a_5913_1654# a_5492_1654# a_5176_1764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X61 gnd d0 a_14108_9389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X62 a_10148_8533# a_10148_8346# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X63 a_2742_n7070# a_2932_n6494# a_2883_n6478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X64 a_10887_n1764# a_10466_n1764# a_9855_n1566# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X65 a_25890_1081# a_25677_1081# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X66 a_35391_n6848# a_35918_n7301# a_36126_n7301# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X67 a_16878_9136# a_16457_9136# a_15940_9380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X68 gnd a_23217_5216# a_23009_5216# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X69 a_37083_3142# a_36786_4113# a_37066_4705# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X70 a_38049_7487# a_38302_7474# a_38051_5275# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X71 a_34896_n10703# a_37895_n10699# a_37846_n10683# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X72 a_855_n5622# a_434_n5622# a_118_n5302# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X73 a_13851_6819# a_13857_6093# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X74 a_11725_5213# a_11512_5213# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X75 a_30864_4908# a_30651_4908# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X76 a_1791_9090# a_1370_9090# a_853_9334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X77 a_11823_6889# a_11756_6297# a_11834_7413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X78 a_18910_n3525# a_19167_n3541# a_17975_n3027# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X79 a_18915_1722# a_18911_1899# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X80 vdd d0 a_24265_6056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X81 a_39096_n4609# a_39099_n3867# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X82 a_36787_n2607# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X83 vdd a_14109_7183# a_13901_7183# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X84 a_3821_7368# a_3824_6637# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X85 a_15944_n2359# a_16674_n2115# a_16882_n2115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X86 a_15207_n2039# a_15207_n1809# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X87 vdd a_28242_n4902# a_28034_n4902# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X88 a_38161_n3008# a_39145_n3522# a_39100_n3318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X89 a_35919_5498# a_35706_5498# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X90 a_35062_466# a_34849_466# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X91 gnd d2 a_2998_n9292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X92 a_34043_n6586# a_34296_n6790# a_33104_n6276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X93 vdd d0 a_19167_n4644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X94 a_1794_2472# a_1373_2472# a_856_2716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X95 a_13858_n3296# a_14111_n3500# a_12919_n2986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X96 a_7832_n8013# a_7846_n9333# a_7797_n9317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X97 a_29067_8316# a_29063_8493# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X98 a_10886_3270# a_11617_3580# a_11825_3580# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X99 gnd a_29322_3891# a_29114_3891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X100 a_29063_n7913# a_29320_n7929# a_28128_n7415# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X101 a_15732_6620# a_15519_6620# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X102 gnd a_8085_7488# a_7877_7488# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X103 gnd d0 a_39351_5548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X104 a_22958_n8141# a_22977_n7067# a_22932_n6863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X105 a_26097_n5644# a_26827_n5400# a_27035_n5400# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X106 vdd a_13172_n4293# a_12964_n4293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X107 a_31074_1599# a_30653_1599# a_30337_1709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X108 a_33098_n9773# a_33355_n9789# a_32962_n9074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X109 vdd a_29319_9406# a_29111_9406# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X110 gnd d0 a_14111_n4603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X111 a_33101_3735# a_33358_3545# a_32960_4327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X112 gnd a_23325_6849# a_23117_6849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X113 a_25360_6157# a_25360_5928# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X114 a_10462_8785# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X115 vdd d0 a_34297_n3481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X116 vdd a_29320_n5169# a_29112_n5169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X117 a_32991_n3734# a_33248_n3750# a_32991_n5934# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X118 a_27987_8598# a_28172_9096# a_28123_9286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X119 vdd d0 a_29320_n9032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X120 a_6850_n4316# a_6429_n4316# a_5911_n4006# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X121 a_6859_5249# a_6539_3037# a_6866_3156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X122 a_18913_3374# a_19166_3361# a_17971_3795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X123 a_1373_n3172# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X124 a_35390_7036# a_35390_6806# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X125 vdd a_8197_3600# a_7989_3600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X126 a_5701_9375# a_5488_9375# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X127 a_30335_5205# a_30863_5457# a_31071_5457# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X128 a_6750_n8149# a_6537_n8149# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X129 vdd a_39352_3342# a_39144_3342# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X130 a_27986_n2680# a_28176_n2104# a_28127_n2088# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X131 a_15519_9380# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X132 gnd a_39351_8308# a_39143_8308# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X133 a_21042_n3397# a_20621_n3397# a_20305_n3077# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X134 a_25675_n7850# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X135 a_4954_480# a_4845_480# a_5053_480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X136 a_18911_n7195# a_18907_n7383# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X137 gnd a_24263_n10094# a_24055_n10094# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X138 a_35921_1086# a_35708_1086# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X139 a_38051_3075# a_38304_3062# a_38047_5452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X140 a_27047_n3541# a_26756_n2602# a_27037_n2091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X141 a_25890_2738# a_25677_2738# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X142 a_32965_1944# a_33150_2442# a_33101_2632# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X143 a_30865_3805# a_30652_3805# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X144 a_20619_7109# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X145 a_35390_8139# a_35919_8258# a_36127_8258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X146 a_10677_n6176# a_10464_n6176# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X147 a_10883_n9485# a_11614_n9795# a_11822_n9795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X148 a_21979_n6462# a_21558_n6462# a_21041_n6706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X149 a_35919_n6198# a_35706_n6198# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X150 a_22930_n2639# a_23187_n2655# a_22960_n3729# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X151 a_6568_6333# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X152 a_32009_n8673# a_31941_n9184# a_32025_n8094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X153 a_35392_n3352# a_35392_n3123# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X154 a_16879_n7630# a_16812_n7038# a_16890_n7977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X155 gnd d1 a_23328_n2063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X156 a_36784_n9225# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X157 a_13856_n8811# a_14109_n9015# a_12917_n8501# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X158 gnd d0 a_9133_9425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X159 a_5910_n8972# a_5489_n8972# a_5173_n8652# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X160 a_25358_9007# a_25886_8802# a_26094_8802# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X161 vdd d1 a_18228_n3231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X162 a_39092_9047# a_39349_8857# a_38154_9291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X163 a_23073_n5168# a_24057_n5682# a_24012_n5478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X164 a_36129_n1786# a_35708_n1786# a_35393_n1790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X165 a_20621_2697# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X166 a_18907_7963# a_19164_7773# a_17969_8207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X167 a_31072_6011# a_31802_5767# a_32010_5767# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X168 a_29063_4630# a_29069_3904# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X169 a_2883_5955# a_3870_5521# a_3821_5711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X170 a_118_5032# a_118_4803# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X171 a_5703_n6766# a_5490_n6766# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X172 a_34038_7354# a_34295_7164# a_33103_6867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X173 a_39095_6292# a_39098_5561# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X174 a_27035_4700# a_26968_4108# a_27052_3137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X175 gnd d0 a_39353_1136# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X176 gnd a_8087_3076# a_7879_3076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X177 vdd a_2999_n7086# a_2791_n7086# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X178 vdd a_24263_n8437# a_24055_n8437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X179 a_6864_n8149# a_6567_n9239# a_6848_n8728# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X180 vdd a_9134_7219# a_8926_7219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X181 vdd a_29321_4994# a_29113_4994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X182 a_31069_n9466# a_30648_n9466# a_30334_n9013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X183 a_31069_8766# a_31800_9076# a_32008_9076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X184 a_4632_480# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X185 a_21989_n7912# a_21880_n8089# a_21994_n5889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X186 a_11834_n7936# a_11543_n6997# a_11823_n7589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X187 a_10465_n6730# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X188 a_649_n2313# a_436_n2313# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X189 gnd a_38271_8590# a_38063_8590# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X190 a_2741_n9276# a_2998_n9292# a_2776_n7972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X191 a_8876_n7378# a_9133_n7394# a_7938_n7622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X192 a_5702_8272# a_5489_8272# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X193 a_25889_6047# a_25676_6047# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X194 vdd a_23217_5216# a_23009_5216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X195 a_26723_n8130# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X196 a_31073_n3402# a_30652_n3402# a_30336_n3082# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X197 a_11841_3120# a_11544_4091# a_11825_3580# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X198 a_8876_n8481# a_8881_n7744# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X199 a_38016_n4891# a_38206_n4315# a_38161_n4111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X200 a_38045_7664# a_38302_7474# a_38051_5275# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X201 a_21042_n1740# a_21773_n2050# a_21981_n2050# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X202 a_17861_n5994# a_18118_n6010# a_17660_n10702# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X203 a_38157_2673# a_39144_2239# a_39095_2429# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X204 gnd d0 a_29321_6097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X205 a_15206_3975# a_15735_3865# a_15943_3865# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X206 a_31728_n9184# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X207 a_36999_n4813# a_36786_n4813# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X208 a_11836_n3524# a_11727_n3701# a_11834_n5736# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X209 gnd d2 a_13032_n2679# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X210 a_23069_5936# a_24056_5502# a_24007_5692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X211 a_31941_8484# a_31728_8484# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X212 a_25360_n6197# a_25888_n6193# a_26096_n6193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X213 a_17861_n3794# a_17880_n2720# a_17831_n2704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X214 a_32009_7973# a_31588_7973# a_31070_7663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X215 a_16672_4724# a_16459_4724# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X216 a_1585_5781# a_1372_5781# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X217 vdd d2 a_28241_n7108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X218 a_12914_n5380# a_13171_n5396# a_12778_n4681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X219 a_5174_n5113# a_5175_n4656# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X220 gnd a_39352_n5728# a_39144_n5728# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X221 a_17970_n5421# a_18957_n5193# a_18912_n4989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X222 a_32020_n5717# a_31700_n3682# a_32027_n3682# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X223 a_28125_5977# a_28382_5787# a_27984_6569# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X224 a_13850_n9548# a_13856_n8811# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X225 a_27050_n8130# a_26753_n9220# a_27034_n8709# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X226 a_648_1059# a_435_1059# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X227 vdd d1 a_8196_5806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X228 a_1584_n8687# a_1371_n8687# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X229 a_8881_5575# a_8877_5752# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X230 gnd a_4078_n7907# a_3870_n7907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X231 a_20304_n6156# a_20832_n6152# a_21040_n6152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X232 gnd d4 a_18118_5281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X233 a_22927_n9257# a_23184_n9273# a_22962_n7953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X234 a_16878_n9836# a_16457_n9836# a_15940_n10080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X235 gnd a_24265_6056# a_24057_6056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X236 vdd d1 a_13171_n6499# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X237 a_15204_n7970# a_15732_n8423# a_15940_n8423# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X238 a_38161_3599# a_38414_3586# a_38016_4368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X239 gnd d0 a_9135_5013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X240 a_35919_n7855# a_35706_n7855# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X241 a_34038_n8980# a_34041_n8238# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X242 a_13852_n6239# a_14109_n6255# a_12914_n6483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X243 a_10147_8990# a_10148_8533# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X244 gnd d0 a_14108_n10118# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X245 gnd a_28382_n6516# a_28174_n6516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X246 gnd a_8198_n2123# a_7990_n2123# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X247 a_37067_n3199# a_37000_n2607# a_37078_n3546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X248 a_26095_7699# a_25674_7699# a_25359_7447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X249 a_26938_n3718# a_26725_n3718# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X250 a_25361_n3347# a_25890_n3438# a_26098_n3438# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X251 gnd d4 a_3031_5235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X252 a_434_4922# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X253 a_1682_500# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X254 a_18909_3551# a_19166_3361# a_17971_3795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X255 a_34039_2388# a_34045_1662# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X256 vdd d1 a_33359_1339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X257 a_35705_n7301# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X258 a_18912_8340# a_18908_8517# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X259 a_13853_6270# a_13856_5539# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X260 a_21700_n2561# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X261 a_8878_n6829# a_9135_n6845# a_7943_n6331# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X262 a_8883_2820# a_8879_2997# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X263 a_3826_n5497# a_3822_n5685# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X264 a_27036_n4297# a_26968_n4808# a_27052_n3718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X265 a_22928_n7051# a_23118_n6475# a_23073_n6271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X266 vdd a_24263_n10094# a_24055_n10094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X267 a_6427_8028# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X268 vdd d0 a_4077_7727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X269 a_38047_3252# a_38304_3062# a_38047_5452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X270 a_39099_n2764# a_39095_n2952# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X271 a_32965_1944# a_33150_2442# a_33105_2455# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X272 a_32961_2121# a_33218_1931# a_32991_3211# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X273 a_16461_n2115# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X274 a_5911_3306# a_5490_3306# a_5175_3054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X275 a_16673_3621# a_16460_3621# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X276 a_30334_n8597# a_30334_n8367# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X277 a_11544_n4791# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X278 vdd a_38413_4689# a_38205_4689# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X279 a_21040_8212# a_20619_8212# a_20303_8322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X280 gnd d2 a_13029_n9297# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X281 a_23071_1524# a_24058_1090# a_24009_1280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X282 a_31943_4072# a_31730_4072# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X283 a_31071_4354# a_30650_4354# a_30335_4559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X284 a_17975_n4130# a_18959_n4644# a_18914_n4440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X285 a_27036_2494# a_26615_2494# a_26097_2184# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X286 a_17970_6001# a_18957_5567# a_18912_5580# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X287 vdd d0 a_9133_9425# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X288 gnd d1 a_3139_6868# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X289 vdd d2 a_8057_1986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X290 a_17834_n4722# a_18019_n5437# a_17974_n5233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X291 a_21041_n5603# a_21771_n5359# a_21979_n5359# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X292 a_16878_9136# a_16811_8544# a_16895_7573# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X293 a_26614_n5400# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X294 gnd a_34297_n1824# a_34089_n1824# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X295 a_39098_7218# a_39351_7205# a_38159_6908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X296 vdd d1 a_8198_1394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X297 gnd a_13170_6873# a_12962_6873# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X298 a_15205_n6680# a_15734_n6771# a_15942_n6771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X299 a_2883_5955# a_3870_5521# a_3825_5534# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X300 a_13855_1858# a_14112_1668# a_12920_1371# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X301 a_25360_4825# a_25360_4595# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X302 a_12919_n4089# a_13903_n4603# a_13854_n4587# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X303 a_5174_n6675# a_5174_n6446# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X304 gnd d5 a_33047_n10658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X305 vdd a_4078_n5147# a_3870_n5147# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X306 a_35392_3497# a_35392_3040# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X307 vdd d0 a_39353_1136# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X308 vdd a_8087_3076# a_7879_3076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X309 a_15733_n6217# a_15520_n6217# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X310 a_27035_n6503# a_26614_n6503# a_26096_n6193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X311 a_30335_n5288# a_30864_n5608# a_31072_n5608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X312 a_37064_n9817# a_36997_n9225# a_37081_n8135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X313 a_26097_3287# a_25676_3287# a_25361_3035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X314 gnd a_19164_n7399# a_18956_n7399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X315 a_2885_n2066# a_3142_n2082# a_2744_n2658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X316 a_6861_n3560# a_6752_n3737# a_6859_n5772# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X317 gnd a_38413_n6521# a_38205_n6521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X318 gnd d0 a_29321_n4066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X319 a_1794_2472# a_1727_1880# a_1805_2996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X320 a_29065_4081# a_29322_3891# a_28130_3594# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X321 a_16781_5254# a_16568_5254# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X322 a_37076_n7958# a_36785_n7019# a_37065_n7611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X323 gnd a_3139_n8700# a_2931_n8700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X324 gnd a_14108_9389# a_13900_9389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X325 a_15735_2762# a_15522_2762# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X326 a_2888_2469# a_3872_2766# a_3823_2956# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X327 a_33098_n9773# a_34085_n9545# a_34040_n9341# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X328 a_27034_8009# a_26613_8009# a_26096_8253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X329 a_645_n10034# a_432_n10034# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X330 vdd d1 a_8196_n6535# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X331 a_15735_n3462# a_15522_n3462# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X332 vdd a_29319_7749# a_29111_7749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X333 a_16599_n7038# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X334 a_10147_9220# a_10676_9339# a_10884_9339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X335 a_853_9334# a_432_9334# a_116_9215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X336 a_1902_n5908# a_1481_n5908# a_1808_n5908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X337 a_10887_n1764# a_11618_n2074# a_11826_n2074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X338 a_11512_5213# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X339 a_30651_4908# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X340 vdd d4 a_18118_5281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X341 a_25888_5493# a_25675_5493# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X342 vdd a_24265_6056# a_24057_6056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X343 a_21994_n5889# a_21667_n8089# a_21989_n7912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X344 a_13854_1304# a_10153_1170# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X345 a_29065_4081# a_29068_3350# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X346 gnd d1 a_33358_n3171# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X347 gnd d1 a_8197_n4329# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X348 a_38157_3776# a_38414_3586# a_38016_4368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X349 vdd d0 a_9135_5013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X350 gnd d0 a_19166_n2987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X351 vout a_19119_n829# a_19416_288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X352 a_37066_n6508# a_36645_n6508# a_36127_n6198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X353 a_35706_5498# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X354 a_16880_4724# a_16813_4132# a_16897_3161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X355 vdd d4 a_3031_5235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X356 a_21042_n1740# a_20621_n1740# a_19886_n1571# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X357 a_34038_n6220# a_34043_n5483# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X358 gnd a_34294_n8442# a_34086_n8442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X359 a_31801_6870# a_31588_6870# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X360 a_2747_n4676# a_3000_n4880# a_2778_n3560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X361 a_15942_n4011# a_15521_n4011# a_15206_n4015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X362 a_2885_1543# a_3872_1109# a_3827_1122# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X363 a_17974_4721# a_18958_5018# a_18909_5208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X364 gnd d0 a_14110_2217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X365 a_21667_n8089# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X366 a_20619_5452# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X367 a_2772_n8160# a_2791_n7086# a_2742_n7070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X368 a_21043_n2294# a_20622_n2294# a_20306_n2203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X369 vdd d1 a_38412_6895# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X370 a_24865_n10698# a_25122_n10714# a_24964_n10698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X371 gnd a_19166_n6850# a_18958_n6850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X372 a_24013_n4375# a_24009_n4563# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X373 vdd d2 a_28241_6379# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X374 a_35392_3497# a_35920_3292# a_36128_3292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X375 a_29062_n7359# a_29068_n6622# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X376 a_33106_1352# a_34090_1649# a_34045_1662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X377 a_5172_n10171# a_9133_n10154# a_7941_n9640# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X378 a_1792_n7584# a_1371_n7584# a_853_n7274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X379 a_17970_4898# a_18227_4708# a_17834_4210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X380 a_32995_n5746# a_33248_n5950# a_32790_n10642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X381 a_30865_n4505# a_30652_n4505# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X382 a_11514_n3701# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X383 a_12805_n3753# a_12824_n2679# a_12775_n2663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X384 vdd a_18225_n9849# a_18017_n9849# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X385 a_31072_n2848# a_31803_n3158# a_32011_n3158# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X386 vdd d0 a_4081_n2392# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X387 a_25675_n6193# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X388 a_5911_n4006# a_6642_n4316# a_6850_n4316# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X389 gnd a_34296_n5687# a_34088_n5687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X390 a_35393_1521# a_35393_1291# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X391 a_10151_1728# a_10680_1618# a_10888_1618# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X392 a_11616_5786# a_11403_5786# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X393 gnd a_14110_4977# a_13902_4977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X394 a_38154_n9814# a_38411_n9830# a_38018_n9115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X395 a_10149_n6826# a_10676_n7279# a_10884_n7279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X396 vdd a_29322_n1860# a_29114_n1860# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X397 a_32993_7446# a_33007_8549# a_32962_8562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X398 a_35922_1640# a_35709_1640# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X399 a_35390_n7305# a_35918_n7301# a_36126_n7301# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X400 vdd a_23185_6338# a_22977_6338# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X401 a_21557_7968# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X402 a_36645_5808# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X403 a_38047_n3775# a_38304_n3791# a_38047_n5975# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X404 a_854_8231# a_433_8231# a_117_8341# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X405 a_20619_n6152# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X406 gnd d6 a_35153_n10719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X407 vdd a_29321_3337# a_29113_3337# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X408 a_16895_n5954# a_16568_n8154# a_16895_n8154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X409 a_30333_n9929# a_30333_n9700# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X410 a_12773_n7075# a_12963_n6499# a_12918_n6295# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X411 a_648_2716# a_435_2716# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X412 a_30652_3805# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X413 a_10149_4808# a_10678_4927# a_10886_4927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X414 a_15519_n8423# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X415 a_10887_n3421# a_11617_n3177# a_11825_n3177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X416 a_24013_2760# a_24009_2937# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X417 a_36787_n2607# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X418 a_35390_n7764# a_35390_n7535# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X419 a_28018_n7994# a_28271_n8198# a_28020_n5782# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X420 a_36643_9117# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X421 a_7940_n4313# a_8197_n4329# a_7799_n4905# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X422 a_25677_n3438# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X423 a_5912_3860# a_5491_3860# a_5175_3970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X424 gnd a_9133_9425# a_8925_9425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X425 a_33106_1352# a_33359_1339# a_32961_2121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X426 a_25359_n9049# a_25886_n9502# a_26094_n9502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X427 a_29070_n2210# a_29066_n2398# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X428 a_12918_5783# a_13171_5770# a_12773_6552# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X429 a_35708_1086# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X430 a_20304_n6386# a_20304_n6156# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X431 a_37076_7435# a_36785_6319# a_37065_6911# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X432 a_5173_n8652# a_5702_n8972# a_5910_n8972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X433 gnd d1 a_38412_n8727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X434 a_10887_3824# a_10466_3824# a_10150_3705# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X435 a_15204_8387# a_15204_8158# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X436 a_30335_n5704# a_30335_n5517# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X437 a_433_n6171# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X438 a_15941_n5114# a_15520_n5114# a_15206_n4661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X439 a_32025_n8094# a_31911_n8094# a_32025_n5894# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X440 a_29067_n8828# a_29320_n9032# a_28128_n8518# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X441 gnd d3 a_3031_n3764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X442 vdd a_28380_9096# a_28172_9096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X443 a_26755_n4808# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X444 gnd a_39353_1136# a_39145_1136# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X445 gnd d1 a_28384_n2104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X446 a_15204_n7970# a_15204_n7783# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X447 a_33105_n4070# a_34089_n4584# a_34040_n4568# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X448 a_15941_7174# a_16671_6930# a_16879_6930# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X449 a_21989_7389# a_21698_6273# a_21979_5762# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X450 a_30335_5205# a_30335_5018# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X451 a_17863_n8018# a_17877_n9338# a_17832_n9134# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X452 a_20832_n6152# a_20619_n6152# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X453 a_15942_n5668# a_15521_n5668# a_15205_n5577# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X454 a_32790_n10642# a_33040_n5950# a_32995_n5746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X455 a_2888_2469# a_3872_2766# a_3827_2779# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X456 a_15734_n2908# a_15521_n2908# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X457 a_10885_7133# a_10464_7133# a_10148_7243# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X458 vdd a_18086_n7132# a_17878_n7132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X459 gnd a_28240_n9314# a_28032_n9314# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X460 a_28129_n5209# a_29113_n5723# a_29068_n5519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X461 a_11545_1885# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X462 a_25676_6047# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X463 a_3825_n7703# a_3821_n7891# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X464 a_24011_n8787# a_24264_n8991# a_23072_n8477# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X465 vdd a_24267_n2373# a_24059_n2373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X466 a_32963_n6868# a_33148_n7583# a_33103_n7379# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X467 a_1793_4678# a_1372_4678# a_855_4922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X468 a_12807_n7977# a_12821_n9297# a_12772_n9281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X469 a_30649_n10020# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X470 a_14710_n10722# a_14967_n10738# a_9776_n10838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X471 a_10149_n6410# a_10678_n6730# a_10886_n6730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X472 a_31071_n6157# a_30650_n6157# a_30335_n5704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X473 a_15207_n2268# a_15207_n2039# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X474 a_21991_2977# a_21700_1861# a_21980_2453# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X475 a_15731_8826# a_15518_8826# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X476 a_21558_n5359# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X477 a_36997_8525# a_36784_8525# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X478 a_28130_n3003# a_29114_n3517# a_29065_n3501# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X479 a_32995_3034# a_33009_4137# a_32964_4150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X480 a_36126_n8404# a_36857_n8714# a_37065_n8714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X481 a_25362_1286# a_25364_1187# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X482 a_22932_6351# a_23117_6849# a_23072_6862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X483 a_31944_n2566# a_31731_n2566# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X484 a_1372_5781# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X485 a_649_1613# a_436_1613# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X486 a_21559_3556# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X487 a_34039_n4014# a_34296_n4030# a_33101_n4258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X488 a_5172_n9525# a_5173_n9068# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X489 a_38020_n4703# a_38273_n4907# a_38051_n3587# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X490 a_39094_n6261# a_39099_n5524# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X491 a_18912_5580# a_19165_5567# a_17970_6001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X492 a_2886_n8496# a_3870_n9010# a_3825_n8806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X493 a_435_1059# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X494 a_36130_1640# a_36860_1396# a_37068_1396# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X495 vdd a_8196_5806# a_7988_5806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X496 a_21979_n6462# a_21558_n6462# a_21040_n6152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X497 a_34043_4971# a_34296_4958# a_33104_4661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X498 a_35389_n9741# a_35918_n10061# a_36126_n10061# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X499 a_36126_6601# a_35705_6601# a_35390_6806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X500 a_30651_n5608# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X501 gnd a_18118_5281# a_17910_5281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X502 a_36784_n9225# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X503 a_7943_n6331# a_8196_n6535# a_7798_n7111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X504 a_37168_527# a_36955_527# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X505 a_31728_8484# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X506 a_5173_n8881# a_5173_n8652# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X507 gnd a_9135_5013# a_8927_5013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X508 a_28016_n5970# a_28273_n5986# a_27815_n10678# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X509 a_10147_8990# a_10675_8785# a_10883_8785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X510 a_11823_n7589# a_11402_n7589# a_10885_n7833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X511 a_35390_7265# a_35390_7036# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X512 a_16879_6930# a_16458_6930# a_15941_7174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X513 a_5175_3741# a_5175_3511# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X514 vdd d0 a_39354_n2419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X515 a_37078_3023# a_36787_1907# a_37067_2499# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X516 vdd d0 a_9133_7768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X517 a_5703_n6766# a_5490_n6766# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X518 a_27246_522# a_28065_5257# a_28016_5447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X519 a_25887_n8399# a_25674_n8399# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X520 gnd d0 a_39351_n5174# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X521 a_27983_n9298# a_28240_n9314# a_28018_n7994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X522 a_6567_8539# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X523 vdd d0 a_29321_n4066# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X524 a_16458_8033# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X525 a_17969_8207# a_18956_7773# a_18907_7963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X526 a_21667_5189# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X527 a_28129_5800# a_29113_6097# a_29068_6110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X528 a_15732_n10080# a_15519_n10080# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X529 a_15731_n9526# a_15518_n9526# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X530 a_118_n5718# a_646_n6171# a_854_n6171# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X531 a_27033_n9812# a_26612_n9812# a_26095_n10056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X532 a_649_n2313# a_436_n2313# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X533 a_26097_n3987# a_25676_n3987# a_25361_n3991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X534 a_31913_2982# a_31700_2982# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X535 a_30336_n3498# a_30864_n3951# a_31072_n3951# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X536 vdd a_4077_7727# a_3869_7727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X537 a_9875_n10838# a_9825_n10854# a_9776_n10838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X538 a_15732_7723# a_15519_7723# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X539 a_857_n2313# a_1587_n2069# a_1795_n2069# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X540 a_32995_n5746# a_33038_n8162# a_32993_n7958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X541 a_36999_n4813# a_36786_n4813# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X542 a_17971_n3215# a_18958_n2987# a_18909_n2971# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X543 a_15733_4414# a_15520_4414# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X544 a_11841_n3701# a_11727_n3701# a_11834_n5736# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X545 a_16460_3621# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X546 a_3824_n8252# a_4077_n8456# a_2882_n8684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X547 a_36999_4113# a_36786_4113# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X548 a_31730_4072# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X549 a_22934_1939# a_23119_2437# a_23074_2450# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X550 vdd a_9133_9425# a_8925_9425# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X551 a_31941_n9184# a_31728_n9184# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X552 vdd a_8057_1986# a_7849_1986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X553 a_13857_n2742# a_14110_n2946# a_12915_n3174# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X554 a_15203_9261# a_15203_9031# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X555 a_12914_5960# a_13171_5770# a_12773_6552# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X556 a_32958_8739# a_33148_7957# a_33099_8147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X557 a_7801_8617# a_8054_8604# a_7832_7501# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X558 a_11834_7413# a_11543_6297# a_11824_5786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X559 a_39096_n1849# a_39097_9424# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X560 a_18914_1168# a_19167_1155# a_17972_1589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X561 a_39096_n9382# a_39349_n9586# a_38154_n9814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X562 gnd a_14110_n6809# a_13902_n6809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X563 vdd a_8198_1394# a_7990_1394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X564 a_5702_7169# a_5489_7169# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X565 a_24010_n7130# a_24006_n7318# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X566 a_10147_n9948# a_10676_n10039# a_10884_n10039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X567 a_16878_n9836# a_16457_n9836# a_15939_n9526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X568 vdd d0 a_39354_1690# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X569 a_39100_n3318# a_39353_n3522# a_38161_n3008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X570 a_24009_n3460# a_24266_n3476# a_23074_n2962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X571 a_15204_n8427# a_15732_n8423# a_15940_n8423# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X572 a_20303_n7718# a_20303_n7489# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X573 vdd a_39353_1136# a_39145_1136# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X574 a_26098_3841# a_25677_3841# a_25361_3722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X575 a_23068_8142# a_24055_7708# a_24006_7898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X576 a_5487_8821# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X577 a_20304_5657# a_20304_5200# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X578 a_21989_5189# a_21880_5189# a_22088_5189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X579 a_10149_4578# a_10677_4373# a_10885_4373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X580 a_15206_3746# a_15206_3516# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X581 a_3826_n5497# a_4079_n5701# a_2887_n5187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X582 a_32011_3561# a_31943_4072# a_32027_3101# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X583 a_1584_7987# a_1371_7987# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X584 vdd d0 a_24266_n4579# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X585 a_15205_n5348# a_15205_n5118# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X586 gnd d0 a_39353_n4625# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X587 gnd d0 a_4078_5521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X588 a_2772_n8160# a_2791_n7086# a_2746_n6882# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X589 gnd d0 a_24263_n7334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X590 a_36130_n2340# a_35709_n2340# a_35393_n2020# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X591 a_38161_2496# a_39145_2793# a_39100_2806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X592 a_30866_1599# a_30653_1599# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X593 a_30334_n7264# a_30862_n7260# a_31070_n7260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X594 a_10463_n7279# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X595 a_2573_n10656# a_2830_n10672# a_2672_n10656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X596 a_35705_n7301# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X597 a_6738_541# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X598 a_6569_4127# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X599 vdd a_9134_n5188# a_8926_n5188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X600 a_34038_8457# a_34041_7726# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X601 a_15522_2762# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X602 a_10883_8785# a_11614_9095# a_11822_9095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X603 a_37066_4705# a_36645_4705# a_36128_4949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X604 a_25887_n10056# a_25674_n10056# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X605 gnd a_23327_n3166# a_23119_n3166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X606 a_17971_3795# a_18958_3361# a_18909_3551# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X607 gnd d0 a_9134_7219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X608 a_20831_n10015# a_20618_n10015# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X609 a_20305_n3493# a_20305_n3306# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X610 vdd a_39352_n2968# a_39144_n2968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X611 a_25359_n8403# a_25359_n7946# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X612 vdd d1 a_3138_n9803# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X613 a_6864_n5949# a_6537_n8149# a_6859_n7972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X614 a_7801_n9129# a_7986_n9844# a_7941_n9640# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X615 a_2884_3749# a_3871_3315# a_3822_3505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X616 a_30863_n7814# a_30650_n7814# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X617 a_15734_3311# a_15521_3311# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X618 a_5172_9485# a_5172_9256# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X619 a_25673_n9502# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X620 a_18913_3374# a_18909_3551# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X621 vdd a_18118_5281# a_17910_5281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X622 a_25675_5493# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X623 a_21981_1350# a_21560_1350# a_21042_1040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X624 a_24005_9001# a_24262_8811# a_23067_9245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X625 a_5489_n8972# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X626 a_2745_n9088# a_2930_n9803# a_2881_n9787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X627 a_13853_n6793# a_14110_n6809# a_12918_n6295# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X628 a_10885_n5073# a_10464_n5073# a_10150_n4620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X629 gnd d2 a_28240_8585# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X630 a_15204_7055# a_15204_6825# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X631 vdd a_9135_5013# a_8927_5013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X632 a_1793_n6481# a_1372_n6481# a_855_n6725# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X633 a_31698_n8094# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X634 a_5703_6066# a_5490_6066# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X635 a_2774_n5948# a_2823_n3764# a_2774_n3748# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X636 a_435_n3416# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X637 a_12916_1548# a_13173_1358# a_12775_2140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X638 gnd d1 a_3142_n2082# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X639 a_7803_4205# a_8056_4192# a_7834_3089# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X640 a_7800_n2699# a_7990_n2123# a_7941_n2107# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X641 a_10678_n2867# a_10465_n2867# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X642 a_15940_9380# a_15519_9380# a_15203_9261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X643 a_10678_6030# a_10465_6030# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X644 a_15207_1769# a_15736_1659# a_15944_1659# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X645 a_16672_5827# a_16459_5827# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X646 vdd d0 a_34293_n9545# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X647 vdd a_38412_6895# a_38204_6895# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X648 a_18909_n4074# a_18914_n3337# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X649 gnd d1 a_38414_n3212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X650 a_23070_3730# a_24057_3296# a_24008_3486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X651 a_24011_n8787# a_24007_n8975# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X652 gnd a_23184_8544# a_22976_8544# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X653 a_31942_6278# a_31729_6278# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X654 a_31070_6560# a_30649_6560# a_30334_6765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X655 a_12035_505# a_11926_505# a_12134_505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X656 a_17969_8207# a_18956_7773# a_18911_7786# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X657 a_16673_2518# a_16460_2518# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X658 a_6864_n8149# a_6567_n9239# a_6847_n9831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X659 a_21040_7109# a_20619_7109# a_20303_6990# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X660 a_1586_3575# a_1373_3575# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X661 gnd a_29320_5543# a_29112_5543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X662 a_6866_n3737# a_6752_n3737# a_6859_n5772# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X663 a_8876_9615# a_8879_8884# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X664 a_10465_n6730# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X665 vdd d0 a_19165_n7953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X666 a_21669_2977# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X667 a_26828_n4297# a_26615_n4297# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X668 a_15205_4849# a_15734_4968# a_15942_4968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X669 vdd a_9136_n4639# a_8928_n4639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X670 gnd a_13169_9079# a_12961_9079# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X671 a_13854_4064# a_14111_3874# a_12919_3577# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X672 a_1370_n9790# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X673 a_34042_n6032# a_34038_n6220# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X674 a_18912_n4989# a_19165_n5193# a_17970_n5421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X675 a_13858_n1639# a_13854_n1827# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X676 a_2103_500# a_1682_500# a_1902_5208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X677 a_32008_9076# a_31587_9076# a_31070_9320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X678 vdd d2 a_18088_n2720# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X679 vdd d0 a_39349_8857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X680 a_23070_n4253# a_23327_n4269# a_22929_n4845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X681 a_11403_5786# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X682 a_25360_5241# a_25888_5493# a_26096_5493# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X683 a_2772_7637# a_3029_7447# a_2778_5248# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X684 gnd d0 a_14109_n7912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X685 a_3822_n6788# a_3825_n6046# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X686 a_6430_n2110# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X687 gnd d0 a_19165_n6296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X688 a_29066_n7171# a_29062_n7359# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X689 a_435_2716# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X690 a_38051_n5787# a_38304_n5991# a_37846_n10683# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X691 a_116_n10130# a_4077_n10113# a_2885_n9599# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X692 a_16570_n3742# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X693 a_18910_1345# a_19167_1155# a_17972_1589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X694 a_2884_n4272# a_3871_n4044# a_3822_n4028# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X695 a_36128_n2889# a_36859_n3199# a_37067_n3199# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X696 a_32009_n7570# a_31588_n7570# a_31070_n7260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X697 a_27050_n8130# a_26753_n9220# a_27033_n9812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X698 a_30861_8766# a_30648_8766# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X699 vdd a_17917_n10718# a_17709_n10718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X700 vdd a_4079_4972# a_3871_4972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X701 a_25677_1081# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X702 a_24007_4589# a_24264_4399# a_23069_4833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X703 a_431_n9480# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X704 a_39097_1880# a_39100_1149# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X705 a_27989_n4698# a_28174_n5413# a_28125_n5397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X706 a_25361_n2888# a_25889_n2884# a_26097_n2884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X707 gnd d2 a_28242_4173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X708 a_29068_n6622# a_29064_n6810# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X709 a_25361_n3118# a_25890_n3438# a_26098_n3438# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X710 vdd d0 a_4078_5521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X711 a_26936_n5930# a_26723_n5930# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X712 a_10675_n9485# a_10462_n9485# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X713 a_12807_7465# a_13060_7452# a_12809_5253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X714 a_21977_n9771# a_21556_n9771# a_21039_n10015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X715 a_26097_6047# a_26827_5803# a_27035_5803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X716 gnd d1 a_23326_n5372# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X717 a_34043_3314# a_34296_3301# a_33101_3735# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X718 a_25887_7699# a_25674_7699# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X719 a_16674_1415# a_16461_1415# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X720 a_32989_7623# a_33008_6343# a_32959_6533# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X721 a_21041_6006# a_20620_6006# a_20304_6116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X722 a_30651_n3951# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X723 gnd a_23186_4132# a_22978_4132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X724 a_31072_2148# a_30651_2148# a_30336_2353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X725 a_17971_3795# a_18958_3361# a_18913_3374# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X726 vdd a_8197_n3226# a_7989_n3226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X727 a_16879_6930# a_16812_6338# a_16890_7454# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X728 a_26094_8802# a_26825_9112# a_27033_9112# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X729 a_18914_n4440# a_19167_n4644# a_17975_n4130# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X730 a_11514_n3701# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X731 a_30336_n4414# a_30336_n4185# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X732 a_39099_5012# a_39352_4999# a_38160_4702# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X733 a_34037_n7323# a_34294_n7339# a_33099_n7567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X734 a_37081_n8135# a_36967_n8135# a_37081_n5935# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X735 a_5912_n4560# a_6642_n4316# a_6850_n4316# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X736 vdd d3 a_23215_7428# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X737 a_2884_3749# a_3871_3315# a_3826_3328# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X738 gnd d2 a_18087_n4926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X739 a_20618_7658# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X740 vdd a_2830_n10672# a_2622_n10672# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X741 a_25364_1187# a_25890_1081# a_26098_1081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X742 a_39095_5189# a_39098_4458# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X743 a_36130_n2340# a_36860_n2096# a_37068_n2096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X744 a_36784_8525# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X745 a_17969_n7627# a_18226_n7643# a_17833_n6928# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X746 a_5909_n7315# a_5488_n7315# a_5173_n7319# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X747 vdd d0 a_14109_n5152# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X748 vdd d2 a_28240_8585# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X749 a_35391_5703# a_35919_5498# a_36127_5498# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X750 gnd d2 a_38271_n9319# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X751 a_436_1613# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X752 a_10463_n10039# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X753 a_647_n5622# a_434_n5622# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X754 vdd a_29323_n2414# a_29115_n2414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X755 a_38019_n6909# a_38204_n7624# a_38159_n7420# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X756 a_15519_n8423# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X757 a_21040_n5049# a_21771_n5359# a_21979_n5359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X758 a_17969_7104# a_18226_6914# a_17833_6416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X759 a_10150_n4620# a_10150_n4433# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X760 a_10151_n2227# a_10680_n2318# a_10888_n2318# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X761 vdd d1 a_28381_7993# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X762 vdd a_33358_n4274# a_33150_n4274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X763 a_2882_8161# a_3139_7971# a_2741_8753# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X764 a_21560_n2050# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X765 a_30863_4354# a_30650_4354# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X766 a_16892_n3565# a_16601_n2626# a_16881_n3218# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X767 gnd d0 a_34297_n4584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X768 vdd a_19166_n4090# a_18958_n4090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X769 a_16460_n4321# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X770 gnd a_29320_n6272# a_29112_n6272# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X771 a_16895_7573# a_16598_8544# a_16879_8033# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X772 a_15207_n2455# a_15207_n2268# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X773 a_25358_n9506# a_25886_n9502# a_26094_n9502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X774 a_855_n3965# a_434_n3965# a_119_n3969# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X775 a_35921_3846# a_35708_3846# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X776 vdd a_23184_8544# a_22976_8544# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X777 gnd d1 a_23327_3540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X778 a_5173_n8881# a_5702_n8972# a_5910_n8972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X779 gnd a_39350_n10140# a_39142_n10140# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X780 a_38020_n4703# a_38205_n5418# a_38156_n5402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X781 a_12920_1371# a_13904_1668# a_13859_1681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X782 a_10677_n8936# a_10464_n8936# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X783 a_20302_9425# a_20302_9196# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X784 vdd a_9133_7768# a_8925_7768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X785 vdd a_29320_5543# a_29112_5543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X786 a_120_n1763# gnd gnd sky130_fd_pr__res_generic_nd w=17 l=81
X787 a_10149_5037# a_10149_4808# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X788 a_39098_n6073# a_39094_n6261# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X789 vdd a_34296_n2927# a_34088_n2927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X790 a_854_7128# a_433_7128# a_117_7009# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X791 a_15204_6825# a_15732_6620# a_15940_6620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X792 a_6864_n5949# a_6750_n5949# a_6958_n5949# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X793 a_1793_n5378# a_1726_n4786# a_1810_n3696# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X794 a_12809_3053# a_13062_3040# a_12805_5430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X795 vdd d1 a_13169_n9808# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X796 a_29062_7939# a_29067_7213# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X797 a_855_n5622# a_1585_n5378# a_1793_n5378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X798 a_25889_3287# a_25676_3287# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X799 a_8881_4472# a_8877_4649# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X800 a_22933_4145# a_23118_4643# a_23069_4833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X801 a_13850_n9548# a_14107_n9564# a_12912_n9792# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X802 a_6642_n4316# a_6429_n4316# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X803 vdd d3 a_13062_n3769# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X804 gnd a_8196_n5432# a_7988_n5432# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X805 a_1805_2996# a_1514_1880# a_1795_1369# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X806 a_31700_2982# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X807 a_34038_n7877# a_34041_n7135# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X808 a_35390_7452# a_35390_7265# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X809 a_5172_9485# a_5701_9375# a_5909_9375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X810 a_38014_8780# a_38204_7998# a_38155_8188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X811 gnd a_28273_n3786# a_28065_n3786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X812 a_31802_4664# a_31589_4664# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X813 gnd a_33216_n7072# a_33008_n7072# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X814 a_23073_n6271# a_24057_n6785# a_24008_n6769# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X815 a_11404_n4280# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X816 a_15520_4414# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X817 a_29067_4453# a_29320_4440# a_28125_4874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X818 a_36127_n8958# a_36857_n8714# a_37065_n8714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X819 a_21994_7508# a_21697_8479# a_21978_7968# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X820 a_36786_4113# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X821 a_2744_n2658# a_2934_n2082# a_2885_n2066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X822 a_24006_9555# a_24009_8824# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X823 a_18912_7237# a_18908_7414# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X824 a_31944_n2566# a_31731_n2566# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X825 a_27045_5230# a_26936_5230# a_27144_5230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X826 a_10884_9339# a_10463_9339# a_10147_9449# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X827 a_13853_5167# a_13856_4436# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X828 vdd d2 a_28242_4173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X829 a_35393_1291# a_35921_1086# a_36129_1086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X830 a_25361_2619# a_25890_2738# a_26098_2738# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X831 vdd d1 a_23325_7952# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X832 a_22931_n9069# a_23116_n9784# a_23071_n9580# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X833 a_17835_n2516# a_18088_n2720# a_17861_n3794# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X834 gnd d0 a_9134_5562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X835 a_37066_n6508# a_36645_n6508# a_36128_n6752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X836 a_29063_n6256# a_29320_n6272# a_28125_n6500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X837 a_17971_2692# a_18228_2502# a_17835_2004# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X838 a_21042_n1740# a_20621_n1740# a_20306_n1744# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X839 a_22960_n5929# a_23009_n3745# a_22964_n3541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X840 a_33102_n2052# a_34089_n1824# a_34044_n1620# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X841 vdd a_39354_1690# a_39146_1690# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X842 a_12803_7642# a_13060_7452# a_12809_5253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X843 a_38047_n3775# a_38066_n2701# a_38017_n2685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X844 a_17832_8622# a_18017_9120# a_17968_9310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X845 a_32989_7623# a_33008_6343# a_32963_6356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X846 a_30334_n7494# a_30334_n7264# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X847 a_17973_n7439# a_18957_n7953# a_18912_n7749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X848 a_21912_n4767# a_21699_n4767# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X849 vdd a_23186_4132# a_22978_4132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X850 a_1371_7987# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X851 a_648_3819# a_435_3819# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X852 a_38154_9291# a_38411_9101# a_38018_8603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X853 gnd a_4078_5521# a_3870_5521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X854 a_15203_n9760# a_15203_n9530# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X855 a_855_6025# a_434_6025# a_118_6135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X856 a_34045_n2174# a_34298_n2378# a_33106_n1864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X857 a_22930_n2639# a_23120_n2063# a_23071_n2047# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X858 a_30653_1599# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X859 a_1374_n2069# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X860 a_17835_n2516# a_18020_n3231# a_17975_n3027# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X861 a_39100_n1661# a_39096_n1849# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X862 a_36125_8807# a_35704_8807# a_35389_9012# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X863 a_12917_n7398# a_13901_n7912# a_13852_n7896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X864 a_29065_n3501# a_29322_n3517# a_28130_n3003# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X865 gnd d2 a_33218_n2660# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X866 gnd a_8057_n2715# a_7849_n2715# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X867 a_20533_n10895# a_20790_n10911# a_19441_n829# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X868 a_12918_n6295# a_13171_n6499# a_12773_n7075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X869 a_17970_n6524# a_18957_n6296# a_18908_n6280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X870 a_5174_n5572# a_5174_n5343# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X871 a_33100_n5361# a_33357_n5377# a_32964_n4662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X872 gnd a_9134_7219# a_8926_7219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X873 a_15731_n9526# a_15518_n9526# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X874 a_27033_n9812# a_26612_n9812# a_26094_n9502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X875 a_35392_2394# a_35393_1937# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X876 a_20303_n7905# a_20303_n7718# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X877 a_3822_3505# a_3827_2779# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X878 a_5173_8153# a_5702_8272# a_5910_8272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X879 a_8883_n4435# a_8879_n4623# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X880 a_12919_3577# a_13172_3564# a_12774_4346# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X881 vdd d0 a_29322_n4620# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X882 a_30336_n3955# a_30864_n3951# a_31072_n3951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X883 a_31803_3561# a_31590_3561# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X884 a_6639_9131# a_6426_9131# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X885 gnd d0 a_29319_n7375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X886 vdd d1 a_33357_n6480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X887 a_10888_1618# a_10467_1618# a_10151_1499# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X888 a_21040_5452# a_20619_5452# a_20304_5200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X889 a_26826_n7606# a_26613_n7606# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X890 vdd d6 a_25122_n10714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X891 a_15521_3311# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X892 a_25676_n2884# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X893 a_31073_n1745# a_30652_n1745# a_30337_n1749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X894 a_15942_4968# a_16672_4724# a_16880_4724# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X895 gnd d0 a_9133_n10154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X896 a_4778_n10717# a_4728_n10733# a_4679_n10717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X897 a_25677_n3438# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X898 a_20306_n2203# a_20306_n1974# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X899 a_28128_8006# a_29112_8303# a_29067_8316# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X900 a_10886_4927# a_10465_4927# a_10149_5037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X901 a_3821_7368# a_4078_7178# a_2886_6881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X902 vdd a_18229_n2128# a_18021_n2128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X903 a_1696_n3696# a_1483_n3696# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X904 vdd d1 a_23327_3540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X905 a_5490_6066# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X906 a_17832_n9134# a_18085_n9338# a_17863_n8018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X907 a_20308_1146# a_20834_1040# a_21042_1040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X908 gnd d0 a_9136_1150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X909 a_645_n10034# a_432_n10034# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X910 a_10885_n5073# a_11616_n5383# a_11824_n5383# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X911 vdd d3 a_8087_n3805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X912 a_26967_n7014# a_26754_n7014# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X913 a_17861_3271# a_17880_1991# a_17831_2181# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X914 a_12805_3230# a_13062_3040# a_12805_5430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X915 a_10465_6030# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X916 a_3824_9397# a_5172_9485# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X917 a_12773_6552# a_12963_5770# a_12914_5960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X918 a_5912_n4560# a_5491_n4560# a_5175_n4240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X919 a_33106_n1864# a_34090_n2378# a_34045_n2174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X920 a_36998_6319# a_36785_6319# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X921 a_5704_n1800# a_5491_n1800# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X922 gnd d1 a_8195_n7638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X923 a_29065_2978# a_29068_2247# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X924 a_22933_4145# a_23118_4643# a_23073_4656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X925 a_16460_2518# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X926 a_1373_3575# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X927 a_36754_n8135# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X928 vdd a_34295_n8996# a_34087_n8996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X929 a_12913_8166# a_13170_7976# a_12772_8758# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X930 a_21040_n5049# a_20619_n5049# a_20305_n4596# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X931 a_5705_n2354# a_5492_n2354# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X932 a_16879_6930# a_16458_6930# a_15940_6620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X933 a_21868_481# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X934 a_36127_4395# a_35706_4395# a_35391_4600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X935 a_29068_n5519# a_29321_n5723# a_28129_n5209# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X936 gnd d2 a_33215_n9278# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X937 vdd d0 a_39353_3896# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X938 a_24985_n1506# a_25890_n1781# a_26098_n1781# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X939 gnd d1 a_33359_1339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X940 a_12914_n5380# a_13901_n5152# a_13856_n4948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X941 a_29063_4630# a_29320_4440# a_28125_4874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X942 a_17829_n7116# a_18019_n6540# a_17970_n6524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X943 a_20833_n2843# a_20620_n2843# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X944 a_29066_9419# a_29319_9406# a_28127_9109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X945 vdd d1 a_18226_8017# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X946 a_10148_6784# a_10676_6579# a_10884_6579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X947 a_21558_n5359# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X948 a_119_n3325# a_119_n3096# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X949 a_11836_n3524# a_11545_n2585# a_11825_n3177# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X950 a_10467_n2318# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X951 a_32010_5767# a_31942_6278# a_32020_7394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X952 gnd d0 a_29321_n6826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X953 a_24013_n3272# a_24009_n3460# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X954 a_18911_1899# a_19168_1709# a_17976_1412# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X955 gnd d0 a_4077_7727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X956 gnd a_4078_n6250# a_3870_n6250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X957 vdd d0 a_9134_5562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X958 vdd a_39353_n3522# a_39145_n3522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X959 a_21913_1861# a_21700_1861# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X960 a_30863_n7814# a_30650_n7814# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X961 a_21042_1040# a_20621_1040# a_20308_1146# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X962 vdd d0 a_4079_n5701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X963 a_26095_9356# a_25674_9356# a_25358_9466# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X964 a_25673_n9502# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X965 a_15942_3311# a_16673_3621# a_16881_3621# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X966 a_29965_345# a_29752_345# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X967 a_5909_n7315# a_6640_n7625# a_6848_n7625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X968 gnd a_13171_n5396# a_12963_n5396# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X969 a_31590_n3158# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X970 a_20620_n6706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X971 vdd d0 a_24264_7159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X972 a_31070_n8363# a_30649_n8363# a_30334_n8367# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X973 a_5489_n8972# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X974 a_17832_8622# a_18017_9120# a_17972_9133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X975 a_39094_8498# a_39351_8308# a_38159_8011# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X976 gnd a_39350_n7380# a_39142_n7380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X977 vdd a_28380_n9825# a_28172_n9825# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X978 a_17970_6001# a_18957_5567# a_18908_5757# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X979 gnd a_28242_4173# a_28034_4173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X980 vdd d0 a_39353_n1865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X981 a_32989_n8146# a_33008_n7072# a_32963_n6868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X982 vdd d2 a_28243_n2696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X983 a_435_n3416# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X984 a_35918_6601# a_35705_6601# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X985 a_5488_n10075# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X986 a_1513_n4786# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X987 a_24011_8275# a_24007_8452# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X988 a_36647_n2096# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X989 a_12776_n9093# a_12961_n9808# a_12916_n9604# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X990 vdd a_4078_5521# a_3870_5521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X991 gnd a_25122_n10714# a_24914_n10714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X992 a_10678_n2867# a_10465_n2867# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X993 a_25360_5241# a_25360_5054# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X994 a_1586_n4275# a_1373_n4275# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X995 a_13859_1681# a_14112_1668# a_12920_1371# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X996 a_15733_5517# a_15520_5517# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X997 a_10883_8785# a_10462_8785# a_10148_8533# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X998 a_12805_n5953# a_12854_n3769# a_12809_n3565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X999 gnd d0 a_9136_2807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1000 gnd d0 a_39350_6651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1001 a_31073_2702# a_30652_2702# a_30336_2812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1002 gnd a_28381_n7619# a_28173_n7619# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1003 a_25674_7699# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1004 a_25361_n4450# a_25361_n4221# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1005 a_16461_1415# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1006 a_15734_2208# a_15521_2208# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1007 a_21980_3556# a_21559_3556# a_21041_3246# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1008 a_33100_4838# a_33357_4648# a_32964_4150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1009 a_5701_n8418# a_5488_n8418# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1010 gnd a_28384_n2104# a_28176_n2104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1011 a_12915_3754# a_13172_3564# a_12774_4346# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1012 gnd d3 a_8085_n8217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1013 a_7802_6411# a_8055_6398# a_7828_7678# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1014 a_25888_n5090# a_25675_n5090# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1015 a_16890_5254# a_16781_5254# a_16989_5254# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1016 a_20304_n5283# a_20304_n5053# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1017 vdd a_23215_7428# a_23007_7428# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1018 vdd d0 a_4080_3869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1019 a_15204_7284# a_15204_7055# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1020 gnd a_4080_2766# a_3872_2766# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1021 a_35920_n6752# a_35707_n6752# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1022 a_1793_5781# a_1372_5781# a_855_6025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1023 a_10149_5224# a_10677_5476# a_10885_5476# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1024 gnd d1 a_28382_n5413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1025 a_10677_8236# a_10464_8236# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1026 a_33103_n7379# a_34087_n7893# a_34038_n7877# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1027 a_854_5471# a_433_5471# a_118_5219# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1028 a_20830_n9461# a_20617_n9461# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1029 a_25889_n5644# a_25676_n5644# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1030 a_26099_1635# a_25678_1635# a_25362_1516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1031 a_7629_n10697# a_7886_n10713# a_4679_n10717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1032 a_5488_6615# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1033 a_120_n2409# a_647_n2862# a_855_n2862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1034 a_10150_2372# a_10678_2167# a_10886_2167# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1035 a_1803_5208# a_1694_5208# a_1902_5208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1036 gnd d1 a_28383_3581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1037 a_5490_n2903# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1038 gnd a_29319_7749# a_29111_7749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1039 vdd a_24265_n5682# a_24057_n5682# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1040 a_645_6574# a_432_6574# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1041 a_16570_n3742# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1042 vdd d0 a_9136_1150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1043 a_35389_9242# a_35918_9361# a_36126_9361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1044 a_39093_n7364# a_39350_n7380# a_38155_n7608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1045 a_10148_n9032# a_10148_n8845# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1046 a_26097_4944# a_25676_4944# a_25360_5054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1047 a_30650_4354# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1048 a_23074_3553# a_24058_3850# a_24013_3863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1049 a_25359_7447# a_25887_7699# a_26095_7699# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1050 a_10884_6579# a_11615_6889# a_11823_6889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1051 a_21042_2697# a_20621_2697# a_20305_2578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1052 a_12773_6552# a_12963_5770# a_12918_5783# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1053 a_37067_2499# a_36646_2499# a_36129_2743# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1054 a_7832_7501# a_7846_8604# a_7797_8794# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1055 a_17972_1589# a_18959_1155# a_18910_1345# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1056 a_24008_3486# a_24013_2760# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1057 vdd d0 a_39350_n8483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1058 gnd a_23327_3540# a_23119_3540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1059 a_25361_3035# a_25361_2848# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1060 a_13855_n2381# a_13858_n1639# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1061 a_34045_n2174# a_34041_n2362# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1062 a_32221_486# a_32112_486# a_32320_486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1063 a_31071_7114# a_31801_6870# a_32009_6870# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1064 vdd a_4080_1109# a_3872_1109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1065 a_21977_n9771# a_21556_n9771# a_21038_n9461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1066 a_32965_n2456# a_33150_n3171# a_33101_n3155# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1067 a_15207_n2268# a_15736_n2359# a_15944_n2359# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1068 vdd a_38414_n4315# a_38206_n4315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1069 a_15735_1105# a_15522_1105# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1070 a_10885_4373# a_10464_4373# a_10150_4121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1071 a_20303_n8362# a_20831_n8358# a_21039_n8358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1072 a_36130_n2340# a_35709_n2340# a_35393_n2249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1073 a_30335_n6807# a_30862_n7260# a_31070_n7260# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1074 a_7941_n9640# a_8194_n9844# a_7801_n9129# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1075 a_15205_n5118# a_15733_n5114# a_15941_n5114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1076 gnd d0 a_4080_1109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1077 a_31801_n8673# a_31588_n8673# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1078 a_25676_3287# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1079 a_30335_n6161# a_30335_n5704# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1080 a_30651_n3951# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1081 a_24006_6795# a_24263_6605# a_23068_7039# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1082 gnd d0 a_9136_n3536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1083 gnd d2 a_28241_6379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1084 a_5173_n7778# a_5173_n7549# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1085 a_14663_485# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1086 a_7828_n8201# a_8085_n8217# a_7834_n5801# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1087 a_33106_1352# a_34090_1649# a_34041_1839# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1088 a_30334_8514# a_30334_8327# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1089 gnd d4 a_13062_n5969# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1090 a_37081_7554# a_36967_7435# a_37081_5354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1091 vdd d0 a_39352_n5728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1092 a_7804_1999# a_8057_1986# a_7830_3266# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1093 a_5701_n10075# a_5488_n10075# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1094 a_5175_2638# a_5175_2408# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1095 a_18911_9443# a_20302_9425# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1096 a_36858_4705# a_36645_4705# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1097 a_3820_n8440# a_3825_n7703# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1098 a_10150_2372# a_10151_1915# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1099 a_20832_n8912# a_20619_n8912# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1100 a_15941_7174# a_15520_7174# a_15204_7055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1101 gnd d0 a_29320_7200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1102 a_853_n8377# a_1584_n8687# a_1792_n8687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1103 a_5489_5512# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1104 a_12776_n9093# a_13029_n9297# a_12807_n7977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1105 gnd a_3141_n4288# a_2933_n4288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1106 a_10153_1170# a_10679_1064# a_10887_1064# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1107 a_35393_1750# a_35922_1640# a_36130_1640# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1108 a_34042_5520# a_34295_5507# a_33100_5941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1109 a_32993_7446# a_33007_8549# a_32958_8739# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1110 a_5909_n7315# a_5488_n7315# a_5174_n6862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1111 gnd a_23185_6338# a_22977_6338# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1112 a_32022_2982# a_31731_1866# a_32012_1355# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1113 vdd a_28242_4173# a_28034_4173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1114 a_27035_n6503# a_26967_n7014# a_27045_n7953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1115 a_1725_n6992# a_1512_n6992# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1116 a_647_n5622# a_434_n5622# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1117 a_1587_1369# a_1374_1369# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1118 vdd a_23325_7952# a_23117_7952# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1119 a_20306_1245# a_20308_1146# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1120 gnd a_9134_5562# a_8926_5562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1121 gnd a_29321_3337# a_29113_3337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1122 a_11823_7992# a_11402_7992# a_10884_7682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1123 a_24005_n9524# a_24262_n9540# a_23067_n9768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1124 a_6850_n3213# a_6429_n3213# a_5912_n3457# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1125 a_647_2162# a_434_2162# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1126 a_28130_n3003# a_28383_n3207# a_27990_n2492# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1127 vdd d1 a_8195_6909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1128 a_6866_3156# a_6569_4127# a_6850_3616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1129 a_13856_n7708# a_13852_n7896# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1130 a_16892_n3565# a_16601_n2626# a_16882_n2115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1131 a_3821_n8994# a_4078_n9010# a_2886_n8496# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1132 a_16460_n4321# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1133 a_3826_n3840# a_3822_n4028# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1134 a_22759_n10637# a_23009_n5945# a_22960_n5929# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1135 vdd d0 a_39350_6651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1136 a_21979_n6462# a_21911_n6973# a_21989_n7912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1137 a_25361_3035# a_25889_3287# a_26097_3287# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1138 a_855_n3965# a_434_n3965# a_119_n3512# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1139 a_12775_2140# a_12965_1358# a_12920_1371# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1140 a_7834_3089# a_7848_4192# a_7799_4382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1141 a_32958_n9262# a_33148_n8686# a_33099_n8670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1142 a_6849_4719# a_6428_4719# a_5911_4963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1143 a_435_3819# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1144 a_10677_n8936# a_10464_n8936# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1145 a_18910_n1868# a_19167_n1884# a_17972_n2112# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1146 a_25677_n1781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1147 a_26095_n7296# a_25674_n7296# a_25360_n6843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1148 vdd a_23326_n6475# a_23118_n6475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1149 gnd a_34296_n4030# a_34088_n4030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1150 a_30862_6560# a_30649_6560# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1151 a_6428_5822# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1152 vdd a_4080_2766# a_3872_2766# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1153 a_12912_n9792# a_13899_n9564# a_13850_n9548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1154 gnd a_19168_n2438# a_18960_n2438# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1155 a_30337_n1749# a_30041_n1547# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1156 a_24008_2383# a_24265_2193# a_23070_2627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1157 a_6642_n4316# a_6429_n4316# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1158 a_3824_9397# a_4077_9384# a_2885_9087# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1159 gnd d2 a_28243_1967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1160 a_117_8341# a_646_8231# a_854_8231# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1161 a_23067_9245# a_24054_8811# a_24005_9001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1162 gnd d1 a_23326_5746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1163 a_20304_4554# a_20305_4097# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1164 vdd d0 a_24264_n7888# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1165 a_8881_n8847# a_8877_n9035# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1166 a_15206_2643# a_15206_2413# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1167 a_12919_3577# a_13903_3874# a_13858_3887# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1168 gnd d0 a_39351_n7934# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1169 vdd d1 a_28383_3581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1170 a_11834_n5736# a_11725_n5913# a_11933_n5913# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1171 a_2884_n4272# a_3141_n4288# a_2743_n4864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1172 a_37083_3142# a_36969_3023# a_37076_5235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1173 a_31590_3561# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1174 a_6426_9131# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1175 a_15942_6071# a_15521_6071# a_15205_6181# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1176 vdd a_18227_n5437# a_18019_n5437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1177 a_27986_n2680# a_28176_n2104# a_28131_n1900# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1178 vdd d0 a_34297_n1824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1179 a_15203_9031# a_15731_8826# a_15939_8826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1180 a_26097_n3987# a_26828_n4297# a_27036_n4297# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1181 a_37078_n3546# a_36969_n3723# a_37076_n5758# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1182 a_32009_n7570# a_31588_n7570# a_31071_n7814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1183 a_117_n8611# a_646_n8931# a_854_n8931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1184 a_29962_n10819# a_34945_n10719# a_32889_n10642# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1185 a_34044_1108# a_34297_1095# a_33102_1529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1186 a_38156_n5402# a_38413_n5418# a_38020_n4703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1187 a_12775_2140# a_13032_1950# a_12805_3230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1188 a_32995_3034# a_33009_4137# a_32960_4327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1189 a_10149_n6410# a_10149_n6180# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1190 a_20306_1475# a_20835_1594# a_21043_1594# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1191 a_34038_7354# a_34041_6623# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1192 a_34042_5520# a_34038_5697# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1193 a_4778_n10717# a_10033_n10854# a_9875_n10838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1194 gnd a_23187_1926# a_22979_1926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1195 a_17972_1589# a_18959_1155# a_18914_1168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1196 vdd a_23327_3540# a_23119_3540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1197 a_14876_485# a_14663_485# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1198 gnd a_9136_1150# a_8928_1150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1199 a_11825_3580# a_11404_3580# a_10886_3270# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1200 a_14830_n1530# a_15735_n1805# a_15943_n1805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1201 a_32025_n8094# a_31728_n9184# a_32008_n9776# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1202 a_25359_n7300# a_25360_n6843# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1203 vdd d1 a_23328_n2063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1204 a_26095_6596# a_26826_6906# a_27034_6906# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1205 a_15206_n4245# a_15206_n4015# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1206 vdd d1 a_38413_n6521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1207 vdd d1 a_8197_2497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1208 vdd d3 a_3029_7447# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1209 a_26936_n5930# a_26723_n5930# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1210 gnd d4 a_8087_n6005# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1211 a_35917_n9507# a_35704_n9507# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1212 vdd d0 a_39352_2239# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1213 a_39092_9047# a_39098_8321# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1214 a_21912_n4767# a_21699_n4767# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1215 a_5175_n3137# a_5704_n3457# a_5912_n3457# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1216 a_18913_2271# a_18909_2448# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1217 a_36785_6319# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1218 gnd d0 a_4077_n10113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1219 a_16812_n7038# a_16599_n7038# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1220 a_26096_4390# a_25675_4390# a_25361_4138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1221 a_18907_n8486# a_19164_n8502# a_17969_n8730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1222 a_12809_5253# a_12852_7452# a_12803_7642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1223 a_5910_8272# a_6640_8028# a_6848_8028# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1224 gnd d1 a_3140_n5391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1225 gnd d0 a_9133_7768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1226 a_27035_5803# a_26614_5803# a_26096_5493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1227 a_21698_6273# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1228 a_435_n1759# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1229 a_23070_n4253# a_24057_n4025# a_24012_n3821# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1230 a_32027_n3682# a_31913_n3682# a_32020_n5717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1231 vdd a_14108_n7358# a_13900_n7358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1232 a_28020_n3582# a_28034_n4902# a_27985_n4886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1233 vdd a_39353_3896# a_39145_3896# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1234 a_34036_n9529# a_34042_n8792# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1235 a_30864_2148# a_30651_2148# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1236 gnd d0 a_24263_9365# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1237 vdd d0 a_34295_8267# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1238 vdd a_18088_n2720# a_17880_n2720# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1239 a_32027_3101# a_31913_2982# a_32020_5194# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1240 a_27033_9112# a_26612_9112# a_26095_9356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1241 vdd a_18226_8017# a_18018_8017# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1242 a_3826_4985# a_4079_4972# a_2887_4675# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1243 a_18909_n2971# a_18915_n2234# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1244 a_117_n7737# a_117_n7508# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1245 gnd d1 a_23328_1334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1246 a_24011_n7684# a_24007_n7872# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1247 a_24013_n4375# a_24266_n4579# a_23074_n4065# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1248 a_30333_n9929# a_30862_n10020# a_31070_n10020# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1249 gnd a_4077_7727# a_3869_7727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1250 a_23071_n2047# a_24058_n1819# a_24009_n1803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1251 a_15204_7471# a_15732_7723# a_15940_7723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1252 vdd a_9134_5562# a_8926_5562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1253 a_21700_1861# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1254 a_26826_n7606# a_26613_n7606# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1255 a_38156_n6505# a_39143_n6277# a_39094_n6261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1256 a_27983_n9298# a_28173_n8722# a_28128_n8518# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1257 vdd a_9134_n7948# a_8926_n7948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1258 gnd d2 a_23186_n4861# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1259 a_15205_4619# a_15733_4414# a_15941_4414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1260 a_10151_n1998# a_10680_n2318# a_10888_n2318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1261 a_31073_n1745# a_30652_n1745# a_30041_n1547# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1262 a_35920_4949# a_35707_4949# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1263 vdd a_24264_7159# a_24056_7159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1264 vdd d0 a_4077_n7353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1265 a_27983_8775# a_28173_7993# a_28128_8006# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1266 a_23068_n7562# a_23325_n7578# a_22932_n6863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1267 a_38159_n7420# a_38412_n7624# a_38019_n6909# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1268 a_34042_n4929# a_34038_n5117# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1269 a_36128_n3992# a_36859_n4302# a_37067_n4302# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1270 a_22934_1939# a_23119_2437# a_23070_2627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1271 a_31074_n2299# a_30653_n2299# a_30337_n2208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1272 a_35705_6601# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1273 a_852_8780# a_1583_9090# a_1791_9090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1274 gnd d0 a_19163_n9605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1275 a_39097_n2403# a_39100_n1661# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1276 a_20618_n8358# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1277 a_2885_n9599# a_3138_n9803# a_2745_n9088# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1278 vdd a_3141_n3185# a_2933_n3185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1279 a_30337_1709# a_30866_1599# a_31074_1599# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1280 a_5173_7279# a_5702_7169# a_5910_7169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1281 gnd a_9134_n6291# a_8926_n6291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1282 a_2888_n4084# a_3872_n4598# a_3827_n4394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1283 a_30333_8971# a_30334_8514# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1284 a_31802_5767# a_31589_5767# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1285 vdd d1 a_23325_n8681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1286 a_6428_n6522# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1287 a_15520_5517# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1288 a_116_n10130# a_116_n9943# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1289 a_7944_n3022# a_8928_n3536# a_8879_n3520# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1290 a_31803_2458# a_31590_2458# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1291 gnd a_9136_2807# a_8928_2807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1292 a_7945_n1919# a_8198_n2123# a_7800_n2699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1293 a_6859_n5772# a_6750_n5949# a_6958_n5949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1294 a_29068_2247# a_29321_2234# a_28126_2668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1295 a_15521_2208# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1296 a_15206_4162# a_15206_3975# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1297 a_25359_n8862# a_25359_n8633# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1298 a_12604_n10661# a_12854_n5969# a_12805_n5953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1299 gnd a_29321_n2963# a_29113_n2963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1300 a_11825_n3177# a_11404_n3177# a_10887_n3421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1301 a_18911_n2422# a_18914_n1680# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1302 a_36787_1907# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1303 gnd d1 a_18227_5811# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1304 a_6850_2513# a_6429_2513# a_5911_2203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1305 a_13850_9025# a_13856_8299# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1306 a_3820_9574# a_4077_9384# a_2885_9087# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1307 a_12805_5430# a_12854_3040# a_12805_3230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1308 vdd d1 a_23326_5746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1309 a_29068_n5519# a_29064_n5707# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1310 a_5175_2638# a_5704_2757# a_5912_2757# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1311 vdd d1 a_3139_7971# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1312 gnd d0 a_9135_3356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1313 a_5705_n2354# a_5492_n2354# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1314 a_15940_n7320# a_15519_n7320# a_15205_n6867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1315 a_35391_n6202# a_35391_n5745# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1316 a_3820_9574# a_3823_8843# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1317 a_20302_n9695# a_20302_n9465# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1318 a_35393_n2020# a_35393_n1790# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1319 a_17861_n5994# a_17910_n3810# a_17865_n3606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1320 a_8883_n1675# a_8879_n1863# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1321 gnd d0 a_24265_4953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1322 a_26754_n7014# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1323 a_10150_2831# a_10679_2721# a_10887_2721# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1324 a_20833_n2843# a_20620_n2843# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1325 a_10464_8236# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1326 a_17833_6416# a_18018_6914# a_17969_7104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1327 a_5909_9375# a_5488_9375# a_5172_9256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1328 gnd a_18087_n4926# a_17879_n4926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1329 a_15733_n5114# a_15520_n5114# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1330 a_25361_n4637# a_25361_n4450# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1331 a_36644_6911# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1332 a_10148_n8386# a_10676_n8382# a_10884_n8382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1333 a_20834_n3397# a_20621_n3397# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1334 gnd d0 a_9136_n1879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1335 gnd a_4079_3315# a_3871_3315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1336 a_23068_n8665# a_24055_n8437# a_24006_n8421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1337 a_432_6574# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1338 vdd a_9136_1150# a_8928_1150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1339 a_18912_n7749# a_19165_n7953# a_17973_n7439# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1340 a_21698_n6973# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1341 a_5175_n3137# a_5175_n2907# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1342 a_5910_n7869# a_6640_n7625# a_6848_n7625# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1343 a_25359_8363# a_25359_8134# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1344 a_20620_n6706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1345 a_31070_n8363# a_30649_n8363# a_30334_n7910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1346 a_30336_n3311# a_30336_n3082# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1347 a_3826_n3840# a_4079_n4044# a_2884_n4272# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1348 a_15204_7471# a_15204_7284# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1349 a_33105_2455# a_33358_2442# a_32965_1944# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1350 a_11839_n5913# a_11512_n8113# a_11834_n7936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1351 a_34044_n1620# a_34297_n1824# a_33102_n2052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1352 a_5174_5947# a_5703_6066# a_5911_6066# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1353 a_22958_n8141# a_23215_n8157# a_22964_n5741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1354 a_18910_4105# a_19167_3915# a_17975_3618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1355 a_12920_1371# a_13173_1358# a_12775_2140# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1356 a_13853_n6793# a_13856_n6051# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1357 a_12809_5253# a_12852_7452# a_12807_7465# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1358 a_34043_n6586# a_34039_n6774# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1359 a_29064_n2947# a_29321_n2963# a_28126_n3191# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1360 a_31804_1355# a_31591_1355# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1361 a_1586_n4275# a_1373_n4275# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1362 gnd d0 a_4081_1663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1363 a_21041_3246# a_20620_3246# a_20305_2994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1364 a_25677_3841# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1365 vdd a_33356_n7583# a_33148_n7583# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1366 a_39092_n9570# a_39098_n8833# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1367 a_15522_1105# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1368 a_15207_1956# a_15207_1769# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1369 vdd a_8195_n8741# a_7987_n8741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1370 vdd a_29321_n6826# a_29113_n6826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1371 a_26969_n2602# a_26756_n2602# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1372 a_15941_5517# a_16672_5827# a_16880_5827# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1373 a_31804_n2055# a_31591_n2055# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1374 gnd d0 a_34295_n7893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1375 vdd d0 a_24263_9365# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1376 gnd a_29318_n9581# a_29110_n9581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1377 a_11512_n5913# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1378 a_15943_2762# a_16673_2518# a_16881_2518# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1379 gnd a_29322_n3517# a_29114_n3517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1380 a_18907_n10143# a_19164_n10159# a_17972_n9645# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1381 a_36756_n3723# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1382 a_24012_3309# a_24008_3486# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1383 a_35917_8807# a_35704_8807# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1384 a_26615_n4297# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1385 vdd d1 a_23328_1334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1386 vdd d1 a_3141_3559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1387 a_20303_6990# a_20303_6760# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1388 a_35920_n6752# a_35707_n6752# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1389 a_23075_1347# a_24059_1644# a_24010_1834# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1390 a_36126_9361# a_36856_9117# a_37064_9117# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1391 a_39098_n4970# a_39094_n5158# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1392 a_20830_n9461# a_20617_n9461# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1393 a_12774_4346# a_12964_3564# a_12915_3754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1394 a_32020_n7917# a_31729_n6978# a_32009_n7570# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1395 a_25889_n5644# a_25676_n5644# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1396 a_2776_7460# a_3029_7447# a_2778_5248# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1397 a_119_n2866# a_647_n2862# a_855_n2862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1398 a_33099_7044# a_33356_6854# a_32963_6356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1399 a_29062_6836# a_29068_6110# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1400 a_6640_n7625# a_6427_n7625# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1401 a_5490_n2903# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1402 a_26096_n6193# a_25675_n6193# a_25360_n6197# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1403 a_1374_1369# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1404 a_16811_8544# a_16598_8544# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1405 a_18911_6683# a_19164_6670# a_17969_7104# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1406 gnd d0 a_9133_n8497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1407 a_34041_9383# a_34037_9560# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1408 a_434_2162# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1409 a_39100_n4421# a_39096_n4609# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1410 vdd a_8195_6909# a_7987_6909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1411 a_30334_8514# a_30861_8766# a_31069_8766# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1412 a_30865_n3402# a_30652_n3402# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1413 a_5491_n3457# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1414 a_1725_6292# a_1512_6292# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1415 a_32960_n4850# a_33217_n4866# a_32995_n3546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1416 a_5911_n4006# a_5490_n4006# a_5175_n3553# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1417 a_36128_2189# a_35707_2189# a_35392_2394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1418 a_11402_n7589# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1419 a_3824_n8252# a_3820_n8440# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1420 a_853_7677# a_432_7677# a_117_7425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1421 a_38156_n5402# a_39143_n5174# a_39098_n4970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1422 a_29064_2424# a_29321_2234# a_28126_2668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1423 a_2747_n4676# a_2932_n5391# a_2883_n5375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1424 a_13855_n2381# a_14112_n2397# a_12920_n1883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1425 a_34041_n8238# a_34294_n8442# a_33099_n8670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1426 a_5912_n4560# a_5491_n4560# a_5175_n4469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1427 a_6781_n7033# a_6568_n7033# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1428 a_28123_9286# a_29110_8852# a_29061_9042# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1429 gnd d1 a_28382_5787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1430 a_11542_8503# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1431 a_11823_n8692# a_11402_n8692# a_10884_n8382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1432 a_12805_5430# a_12854_3040# a_12809_3053# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1433 a_644_8780# a_431_8780# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1434 a_37064_n9817# a_36643_n9817# a_36126_n10061# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1435 vdd d0 a_9135_3356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1436 a_17973_n8542# a_18226_n8746# a_17828_n9322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1437 a_26096_7150# a_25675_7150# a_25359_7260# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1438 a_33100_n5361# a_34087_n5133# a_34042_n4929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1439 gnd d0 a_14109_n6255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1440 a_9987_364# a_19208_288# a_19416_288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1441 a_31801_n8673# a_31588_n8673# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1442 vdd a_33246_n8162# a_33038_n8162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1443 a_25239_461# a_24818_461# a_25140_461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1444 a_12772_8758# a_12962_7976# a_12917_7989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1445 a_39095_6292# a_39352_6102# a_38160_5805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1446 gnd a_28243_1967# a_28035_1967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1447 gnd a_23326_5746# a_23118_5746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1448 a_8880_7781# a_8876_7958# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1449 a_35919_4395# a_35706_4395# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1450 a_10467_n2318# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1451 a_34043_n5483# a_34296_n5687# a_33104_n5173# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1452 vdd d0 a_19167_n3541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1453 a_2882_n7581# a_3869_n7353# a_3824_n7149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1454 vdd a_4079_3315# a_3871_3315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1455 a_33101_n3155# a_34088_n2927# a_34039_n2911# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1456 a_25239_461# a_29965_345# a_19317_288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1457 a_25358_9237# a_25358_9007# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1458 a_36126_7704# a_36857_8014# a_37065_8014# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1459 a_20832_n8912# a_20619_n8912# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1460 gnd d3 a_23215_7428# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1461 a_1372_n5378# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1462 a_10886_2167# a_11617_2477# a_11825_2477# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1463 a_10884_6579# a_10463_6579# a_10149_6327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1464 gnd d0 a_39351_4445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1465 vdd a_13172_n3190# a_12964_n3190# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1466 a_17968_n9833# a_18955_n9605# a_18906_n9589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1467 a_38047_n5975# a_38096_n3791# a_38051_n3587# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1468 a_21880_n5889# a_21667_n5889# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1469 gnd d0 a_14111_n3500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1470 a_33101_2632# a_33358_2442# a_32965_1944# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1471 a_12809_n3565# a_13062_n3769# a_12805_n5953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1472 a_25887_9356# a_25674_9356# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1473 a_16813_4132# a_16600_4132# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1474 vdd d0 a_29320_n7929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1475 a_32962_8562# a_33147_9060# a_33098_9250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1476 a_6850_n3213# a_6429_n3213# a_5911_n2903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1477 gnd a_4079_n2941# a_3871_n2941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1478 a_8883_n3332# a_8879_n3520# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1479 vdd a_8197_2497# a_7989_2497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1480 a_30336_4102# a_30863_4354# a_31071_4354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1481 vdd d1 a_33355_n9789# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1482 vdd d0 a_4081_1663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1483 a_21978_n7565# a_21911_n6973# a_21989_n7912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1484 gnd d0 a_29319_9406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1485 vdd d3 a_33248_n3750# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1486 vdd a_8087_n3805# a_7879_n3805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1487 vdd a_39352_2239# a_39144_2239# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1488 a_5488_7718# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1489 a_28020_5270# a_28063_7469# a_28018_7482# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1490 a_10150_3018# a_10678_3270# a_10886_3270# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1491 a_35391_n5745# a_35919_n6198# a_36127_n6198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1492 a_35392_3956# a_35921_3846# a_36129_3846# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1493 a_855_3265# a_434_3265# a_119_3013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1494 gnd a_39351_7205# a_39143_7205# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1495 a_16879_n8733# a_16811_n9244# a_16895_n8154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1496 a_1794_n3172# a_1373_n3172# a_855_n2862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1497 a_5489_4409# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1498 a_5701_n8418# a_5488_n8418# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1499 gnd d5 a_12861_n10677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1500 gnd d1 a_28384_1375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1501 a_39095_3532# a_39100_2806# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1502 a_20618_9315# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1503 a_11544_4091# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1504 a_12920_1371# a_13904_1668# a_13855_1858# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1505 gnd d8 a_20790_n10911# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1506 gnd a_9133_7768# a_8925_7768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1507 vdd d1 a_28384_n2104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1508 a_646_4368# a_433_4368# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1509 gnd a_13031_n4885# a_12823_n4885# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1510 a_30865_2702# a_30652_2702# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1511 a_10677_n5073# a_10464_n5073# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1512 a_35390_7036# a_35919_7155# a_36127_7155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1513 gnd d1 a_33359_n2068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1514 vdd d2 a_18085_8609# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1515 a_16769_546# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1516 a_30651_2148# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1517 gnd a_24263_9365# a_24055_9365# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1518 a_5909_n10075# a_5488_n10075# a_5172_n9984# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1519 a_10680_1618# a_10467_1618# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1520 vdd a_34295_8267# a_34087_8267# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1521 a_23075_1347# a_24059_1644# a_24014_1657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1522 a_13856_n7708# a_14109_n7912# a_12917_n7398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1523 a_10463_n8382# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1524 a_7941_n2107# a_8928_n1879# a_8879_n1863# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1525 a_5910_n7869# a_5489_n7869# a_5173_n7549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1526 a_12774_4346# a_12964_3564# a_12919_3577# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1527 a_5702_n5109# a_5489_n5109# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1528 a_7828_7678# a_7847_6398# a_7798_6588# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1529 a_119_4116# a_119_3929# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1530 a_16989_5254# a_16568_5254# a_16895_5373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1531 gnd a_23328_1334# a_23120_1334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1532 a_11839_n5913# a_11725_n5913# a_11933_n5913# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1533 vdd a_13170_n8705# a_12962_n8705# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1534 a_20303_n8362# a_20303_n7905# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1535 a_27985_4363# a_28175_3581# a_28126_3771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1536 a_18907_6860# a_19164_6670# a_17969_7104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1537 a_31072_4908# a_31802_4664# a_32010_4664# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1538 a_10885_5476# a_10464_5476# a_10149_5681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1539 a_5703_n5663# a_5490_n5663# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1540 a_27035_5803# a_26967_6314# a_27045_7430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1541 a_37083_n3723# a_36969_n3723# a_37076_n5758# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1542 a_7798_n7111# a_8055_n7127# a_7828_n8201# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1543 gnd d3 a_23217_3016# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1544 a_5704_3860# a_5491_3860# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1545 a_32020_5194# a_31700_2982# a_32027_3101# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1546 vdd d4 a_28273_5257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1547 a_1902_5208# a_1481_5208# a_1808_5327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1548 a_10886_2167# a_10465_2167# a_10151_1915# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1549 a_117_n8840# a_646_n8931# a_854_n8931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1550 a_34040_n9341# a_34036_n9529# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1551 a_17832_n9134# a_18017_n9849# a_17968_n9833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1552 a_19416_288# a_18995_288# a_9987_364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1553 a_25889_4944# a_25676_4944# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1554 a_31073_n1745# a_31804_n2055# a_32012_n2055# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1555 a_15207_n1809# a_15735_n1805# a_15943_n1805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1556 a_17861_5471# a_17910_3081# a_17861_3271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1557 a_3820_n10097# a_3823_n9355# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1558 a_38021_n2497# a_38206_n3212# a_38161_n3008# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1559 a_18913_n2783# a_18909_n2971# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1560 a_28127_n2088# a_29114_n1860# a_29065_n1844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1561 gnd a_4076_n9559# a_3868_n9559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1562 a_20302_n10111# a_24263_n10094# a_23071_n9580# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1563 a_15941_8277# a_15520_8277# a_15204_8387# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1564 a_33104_n6276# a_33357_n6480# a_32959_n7056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1565 gnd a_18086_6403# a_17878_6403# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1566 a_17865_n3606# a_17879_n4926# a_17834_n4722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1567 a_36859_2499# a_36646_2499# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1568 a_19441_n829# a_19332_n829# vout vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1569 a_31590_2458# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1570 a_35917_n9507# a_35704_n9507# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1571 a_10886_n6730# a_10465_n6730# a_10149_n6410# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1572 a_15207_n2039# a_15736_n2359# a_15944_n2359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1573 gnd d0 a_29321_4994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1574 a_15206_2872# a_15735_2762# a_15943_2762# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1575 gnd d0 a_34296_6061# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1576 a_20303_n7905# a_20831_n8358# a_21039_n8358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1577 vdd d0 a_9133_n7394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1578 a_5175_n3366# a_5704_n3457# a_5912_n3457# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1579 a_28016_5447# a_28065_3057# a_28020_3070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1580 gnd a_18227_5811# a_18019_5811# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1581 a_18909_n6834# a_18912_n6092# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1582 a_12774_n4869# a_13031_n4885# a_12809_n3565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1583 a_32009_6870# a_31588_6870# a_31070_6560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1584 a_32009_n7570# a_31942_n6978# a_32020_n7917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1585 a_20305_3681# a_20834_3800# a_21042_3800# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1586 vdd d4 a_18118_n6010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1587 a_10679_n4524# a_10466_n4524# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1588 vdd a_23326_5746# a_23118_5746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1589 gnd a_9135_3356# a_8927_3356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1590 a_11824_5786# a_11403_5786# a_10885_5476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1591 vdd d1 a_28381_n8722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1592 a_13853_3510# a_13858_2784# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1593 a_29064_6287# a_29067_5556# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1594 vdd d1 a_8196_4703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1595 a_24011_7172# a_24007_7349# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1596 a_1584_n7584# a_1371_n7584# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1597 a_13853_5167# a_14110_4977# a_12918_4680# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1598 gnd a_8085_n8217# a_7877_n8217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1599 a_20304_n5053# a_20832_n5049# a_21040_n5049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1600 vdd d2 a_18087_4197# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1601 gnd a_24265_4953# a_24057_4953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1602 vdd d1 a_13171_n5396# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1603 a_34041_1839# a_34298_1649# a_33106_1352# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1604 vdd d0 a_39351_4445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1605 a_17660_n10702# a_17910_n6010# a_17861_n5994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1606 a_7938_n8725# a_8925_n8497# a_8876_n8481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1607 a_38161_2496# a_38414_2483# a_38021_1985# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1608 a_13852_n5136# a_14109_n5152# a_12914_n5380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1609 a_7830_3266# a_7849_1986# a_7800_2176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1610 gnd a_28382_n5413# a_28174_n5413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1611 a_26095_6596# a_25674_6596# a_25360_6344# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1612 a_31072_3251# a_31803_3561# a_32011_3561# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1613 a_32991_n3734# a_33010_n2660# a_32961_n2644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1614 a_32962_8562# a_33147_9060# a_33102_9073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1615 a_18909_2448# a_19166_2258# a_17971_2692# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1616 a_10887_1064# a_10466_1064# a_10151_1269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1617 a_27037_1391# a_26969_1902# a_27047_3018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1618 a_21697_8479# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1619 gnd d2 a_18086_n7132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1620 a_23075_n1859# a_24059_n2373# a_24010_n2357# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1621 vdd a_23016_n10653# a_22808_n10653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1622 a_6429_3616# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1623 a_36129_n4546# a_36859_n4302# a_37067_n4302# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1624 a_8878_n5726# a_9135_n5742# a_7943_n5228# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1625 a_37081_n5935# a_36754_n8135# a_37081_n8135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1626 a_3825_7191# a_4078_7178# a_2886_6881# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1627 a_118_6135# a_647_6025# a_855_6025# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1628 gnd d1 a_3140_5765# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1629 a_22933_n4657# a_23118_n5372# a_23073_n5168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1630 a_21042_3800# a_20621_3800# a_20305_3681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1631 vdd d1 a_28384_1375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1632 a_12914_n6483# a_13901_n6255# a_13852_n6239# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1633 a_6427_6925# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1634 a_28124_n8706# a_29111_n8478# a_29062_n8462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1635 a_1793_n6481# a_1725_n6992# a_1803_n7931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1636 a_6428_n6522# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1637 a_31591_1355# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1638 a_35392_3727# a_35392_3497# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1639 a_11926_505# a_11713_505# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1640 a_5910_5512# a_5489_5512# a_5174_5717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1641 vdd d0 a_9135_n6845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1642 gnd a_18088_1991# a_17880_1991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1643 gnd a_13171_5770# a_12963_5770# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1644 a_12912_n9792# a_13169_n9808# a_12776_n9093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1645 a_28131_1388# a_29115_1685# a_29066_1875# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1646 a_10148_n7929# a_10148_n7742# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1647 vdd a_19165_n6296# a_18957_n6296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1648 a_5911_2203# a_5490_2203# a_5176_1951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1649 a_8882_n3881# a_9135_n4085# a_7940_n4313# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1650 vdd a_24263_9365# a_24055_9365# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1651 a_25359_8550# a_25359_8363# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1652 a_854_n6171# a_433_n6171# a_118_n6175# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1653 a_17975_n3027# a_18959_n3541# a_18914_n3337# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1654 a_24009_n1803# a_24266_n1819# a_23071_n2047# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1655 a_39100_n1661# a_39353_n1865# a_38158_n2093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1656 a_26924_522# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1657 gnd d0 a_4079_n6804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1658 a_35704_8807# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1659 vdd a_23328_1334# a_23120_1334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1660 a_22858_n10637# a_22808_n10653# a_22759_n10637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1661 a_16882_n2115# a_16461_n2115# a_15943_n1805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1662 a_11826_1374# a_11405_1374# a_10887_1064# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1663 a_35390_n8867# a_35919_n8958# a_36127_n8958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1664 gnd d5 a_7886_n10713# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1665 a_27985_4363# a_28175_3581# a_28130_3594# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1666 a_15205_n5577# a_15734_n5668# a_15942_n5668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1667 a_23072_7965# a_23325_7952# a_22927_8734# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1668 a_2883_4852# a_3870_4418# a_3825_4431# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1669 vdd a_38412_n7624# a_38204_n7624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1670 a_15520_n8977# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1671 a_6537_5249# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1672 a_118_n5072# a_119_n4615# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1673 a_12919_n2986# a_13903_n3500# a_13854_n3484# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1674 a_3824_1853# a_3827_1122# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1675 a_2885_9087# a_3869_9384# a_3820_9574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1676 vdd d3 a_23217_3016# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1677 a_12920_n1883# a_13173_n2087# a_12775_n2663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1678 a_20617_8761# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1679 a_39096_n9382# a_39092_n9570# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1680 a_27035_n5400# a_26614_n5400# a_26096_n5090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1681 gnd d1 a_18226_8017# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1682 a_36128_n6752# a_35707_n6752# a_35391_n6661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1683 a_28125_n6500# a_28382_n6516# a_27984_n7092# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1684 a_26097_2184# a_25676_2184# a_25362_1932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1685 a_21981_1350# a_21913_1861# a_21991_2977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1686 a_15939_8826# a_15518_8826# a_15204_8574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1687 a_21698_n6973# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1688 a_29065_1321# a_25364_1187# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1689 a_17861_5471# a_17910_3081# a_17865_3094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1690 gnd a_38413_n5418# a_38205_n5418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1691 a_24008_n2906# a_24014_n2169# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1692 a_39098_n8833# a_39094_n9021# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1693 a_12916_9092# a_13900_9389# a_13855_9402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1694 a_1512_6292# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1695 a_21699_4067# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1696 a_35706_n6198# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1697 a_12805_3230# a_12824_1950# a_12779_1963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1698 a_16598_n9244# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1699 a_29065_2978# a_29322_2788# a_28130_2491# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1700 gnd d0 a_24264_7159# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1701 a_10149_5037# a_10678_4927# a_10886_4927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1702 gnd a_3139_n7597# a_2931_n7597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1703 vdd d0 a_34296_6061# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1704 vdd d1 a_3142_n2082# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1705 a_27034_6906# a_26613_6906# a_26096_7150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1706 vdd d0 a_9136_3910# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1707 vdd d1 a_8196_n5432# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1708 a_35393_n2249# a_35393_n2020# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1709 gnd d1 a_3142_1353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1710 a_29066_6659# a_29062_6836# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1711 a_36128_6052# a_35707_6052# a_35391_5933# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1712 a_431_8780# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1713 a_15205_5265# a_15733_5517# a_15941_5517# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1714 vdd a_9135_3356# a_8927_3356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1715 gnd d0 a_14107_8835# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1716 a_26969_n2602# a_26756_n2602# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1717 a_39101_1703# a_39354_1690# a_38162_1393# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1718 gnd d7 a_10033_n10854# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1719 a_435_n1759# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1720 a_25888_4390# a_25675_4390# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1721 a_11512_n5913# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1722 a_22960_n3729# a_22979_n2655# a_22934_n2451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1723 gnd a_24265_n6785# a_24057_n6785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1724 a_33104_4661# a_33357_4648# a_32964_4150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1725 a_38157_2673# a_38414_2483# a_38021_1985# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1726 a_6537_7449# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1727 a_33103_7970# a_34087_8267# a_34042_8280# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1728 a_1694_7408# a_1481_7408# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1729 a_39097_n8279# a_39350_n8483# a_38155_n8711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1730 a_36756_n3723# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1731 a_35706_4395# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1732 a_38018_8603# a_38203_9101# a_38154_9291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1733 a_29066_n7171# a_29319_n7375# a_28124_n7603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1734 a_11823_n7589# a_11756_n6997# a_11834_n7936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1735 gnd a_34294_n7339# a_34086_n7339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1736 vdd a_23324_n9784# a_23116_n9784# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1737 a_25360_n6427# a_25360_n6197# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1738 gnd a_23215_7428# a_23007_7428# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1739 a_1793_5781# a_1725_6292# a_1803_7408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1740 a_3827_n4394# a_4080_n4598# a_2888_n4084# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1741 vdd a_23217_n3745# a_23009_n3745# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1742 a_16672_n6527# a_16459_n6527# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1743 a_31591_n2055# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1744 a_6850_3616# a_6429_3616# a_5912_3860# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1745 vdd a_38302_n8203# a_38094_n8203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1746 a_5174_5947# a_5174_5717# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1747 gnd a_19166_n5747# a_18958_n5747# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1748 gnd a_38274_n2701# a_38066_n2701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1749 a_37277_527# a_37168_527# a_35171_466# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1750 a_10149_5681# a_10149_5224# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1751 a_28128_n8518# a_28381_n8722# a_27983_n9298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1752 a_6640_n7625# a_6427_n7625# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1753 a_37846_n10683# a_38096_n5991# a_38047_n5975# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1754 gnd d2 a_3000_n4880# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1755 a_9779_364# a_9566_364# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1756 a_2884_n4272# a_3871_n4044# a_3826_n3840# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1757 a_25674_9356# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1758 a_16600_4132# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1759 vdd d1 a_3140_5765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1760 a_7938_n7622# a_8925_n7394# a_8880_n7190# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1761 a_20618_n8358# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1762 a_30865_n3402# a_30652_n3402# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1763 a_38157_n3196# a_39144_n2968# a_39095_n2952# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1764 a_5491_n3457# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1765 a_34045_1662# a_34041_1839# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1766 a_8881_n7744# a_8877_n7932# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1767 a_10150_3705# a_10679_3824# a_10887_3824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1768 vdd d0 a_34295_n5133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1769 a_11839_7532# a_11725_7413# a_11839_5332# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1770 a_5911_n2903# a_6642_n3213# a_6850_n3213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1771 vdd a_13171_5770# a_12963_5770# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1772 a_13851_n8445# a_13856_n7708# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1773 gnd d0 a_29319_n10135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1774 a_28131_1388# a_29115_1685# a_29070_1698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1775 a_11616_4683# a_11403_4683# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1776 vdd d1 a_3139_n8700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1777 gnd d4 a_33248_n5950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1778 gnd a_8087_n6005# a_7879_n6005# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1779 a_11834_n5736# a_11514_n3701# a_11841_n3701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1780 a_21557_6865# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1781 a_36645_4705# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1782 a_34042_4417# a_34038_4594# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1783 a_20619_n5049# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1784 a_37064_n9817# a_36643_n9817# a_36125_n9507# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1785 a_12778_n4681# a_12963_n5396# a_12918_n5192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1786 gnd d0 a_34296_n2927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1787 a_433_4368# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1788 gnd a_9135_n2982# a_8927_n2982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1789 a_30652_2702# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1790 vdd d1 a_38411_n9830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1791 a_31913_n3682# a_31700_n3682# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1792 a_33100_n6464# a_34087_n6236# a_34038_n6220# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1793 a_34040_n1808# a_35016_n1511# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1794 a_26966_n9220# a_26753_n9220# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1795 a_1724_8498# a_1511_8498# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1796 a_15206_n3142# a_15206_n2912# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1797 a_15940_n7320# a_15519_n7320# a_15204_n7324# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1798 a_432_n8377# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1799 a_37078_3023# a_36787_1907# a_37068_1396# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1800 a_11616_n6486# a_11403_n6486# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1801 a_30337_1709# a_30337_1480# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1802 a_2885_9087# a_3869_9384# a_3824_9397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1803 vdd d3 a_38304_n3791# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1804 a_7940_n3210# a_8197_n3226# a_7804_n2511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1805 a_22962_n7953# a_22976_n9273# a_22931_n9069# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1806 a_28124_n7603# a_29111_n7375# a_29066_n7171# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1807 a_5912_2757# a_5491_2757# a_5175_2867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1808 vdd a_3001_n2674# a_2793_n2674# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1809 a_6539_3037# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1810 a_120_1494# a_120_1264# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1811 a_29064_n2947# a_29070_n2210# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1812 gnd d3 a_28271_n8198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1813 vdd d0 a_29318_8852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1814 a_10887_2721# a_10466_2721# a_10150_2602# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1815 a_3827_n4394# a_3823_n4582# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1816 a_433_n5068# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1817 a_25362_1516# a_25362_1286# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1818 a_5491_3860# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1819 a_25678_1635# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1820 gnd a_23217_3016# a_23009_3016# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1821 a_20303_7863# a_20303_7406# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1822 vdd a_28273_5257# a_28065_5257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1823 gnd a_23186_n4861# a_22978_n4861# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1824 a_33105_n2967# a_34089_n3481# a_34040_n3465# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1825 a_20305_n3306# a_20834_n3397# a_21042_n3397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1826 a_1512_n6992# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1827 a_28016_3247# a_28035_1967# a_27990_1980# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1828 gnd d0 a_29320_n9032# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1829 a_7943_n6331# a_8927_n6845# a_8882_n6641# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1830 gnd a_14111_n1843# a_13903_n1843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1831 a_25676_4944# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1832 a_24011_n7684# a_24264_n7888# a_23072_n7374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1833 vdd d1 a_3142_1353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1834 a_32025_5313# a_31698_7394# a_32020_7394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1835 a_647_n3965# a_434_n3965# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1836 a_11841_3120# a_11727_3001# a_11834_5213# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1837 a_10149_n5307# a_10678_n5627# a_10886_n5627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1838 a_31071_n5054# a_30650_n5054# a_30336_n4601# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1839 a_15203_n10176# a_18907_n10143# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1840 gnd a_4080_n3495# a_3872_n3495# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1841 gnd a_34296_6061# a_34088_6061# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1842 a_30335_5018# a_30335_4789# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1843 a_21558_5762# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1844 a_17975_3618# a_18959_3915# a_18914_3928# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1845 a_16878_n9836# a_16811_n9244# a_16895_n8154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1846 gnd d0 a_24264_n8991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1847 a_12775_2140# a_12965_1358# a_12916_1548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1848 a_36646_3602# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1849 a_36126_n7301# a_36857_n7611# a_37065_n7611# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1850 a_32993_n7958# a_33007_n9278# a_32962_n9074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1851 a_35706_n8958# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1852 a_25674_n10056# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1853 gnd a_18227_n6540# a_18019_n6540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1854 a_21559_2453# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1855 a_34039_n2911# a_34296_n2927# a_33101_n3155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1856 a_6783_n2621# a_6570_n2621# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1857 a_16812_6338# a_16599_6338# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1858 a_30335_5892# a_30864_6011# a_31072_6011# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1859 a_18912_4477# a_19165_4464# a_17970_4898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1860 a_2886_n7393# a_3870_n7907# a_3825_n7703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1861 gnd a_9132_n9600# a_8924_n9600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1862 a_15206_3516# a_15734_3311# a_15942_3311# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1863 vdd a_8196_4703# a_7988_4703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1864 a_21979_n5359# a_21558_n5359# a_21040_n5049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1865 a_30335_6308# a_30862_6560# a_31070_6560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1866 a_6426_n9831# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1867 a_1726_4086# a_1513_4086# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1868 a_7943_n5228# a_8196_n5432# a_7803_n4717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1869 a_31803_n4261# a_31590_n4261# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1870 a_25359_n7946# a_25887_n8399# a_26095_n8399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1871 gnd d2 a_38273_n4907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1872 a_32320_486# a_31899_486# a_32119_5194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1873 a_3827_3882# a_3823_4059# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1874 vdd a_2998_n9292# a_2790_n9292# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1875 a_19119_n829# d9 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1876 a_25359_n7759# a_25359_n7530# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1877 vdd a_14111_3874# a_13903_3874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1878 a_38014_8780# a_38271_8590# a_38049_7487# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1879 a_11543_6297# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1880 vdd a_33216_n7072# a_33008_n7072# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1881 a_35920_2189# a_35707_2189# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1882 a_5703_n5663# a_5490_n5663# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1883 vdd d4 a_28273_n5986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1884 a_2744_n2658# a_2934_n2082# a_2889_n1878# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1885 a_35391_n5099# a_35392_n4642# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1886 a_855_n3965# a_1586_n4275# a_1794_n4275# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1887 a_13854_n1827# a_14111_n1843# a_12916_n2071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1888 vdd d0 a_19164_n10159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1889 a_9776_n10838# a_14759_n10738# a_12703_n10661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1890 a_36998_n7019# a_36785_n7019# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1891 a_17969_7104# a_18956_6670# a_18907_6860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1892 a_35062_466# a_34849_466# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1893 a_1727_n2580# a_1514_n2580# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1894 gnd d3 a_18116_7493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1895 gnd a_14108_n8461# a_13900_n8461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1896 a_26097_n2884# a_25676_n2884# a_25361_n2888# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1897 vdd d2 a_28240_n9314# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1898 a_25361_n3534# a_25361_n3347# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1899 a_3823_n3479# a_4080_n3495# a_2888_n2981# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1900 a_27984_6569# a_28174_5787# a_28125_5977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1901 a_18906_9066# a_19163_8876# a_17968_9310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1902 a_13858_2784# a_14111_2771# a_12919_2474# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1903 a_27034_8009# a_26966_8520# a_27050_7549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1904 gnd d3 a_3029_7447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1905 a_36126_n10061# a_35705_n10061# a_35389_n9970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1906 a_39093_9601# a_39096_8870# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1907 gnd a_39351_n9037# a_39143_n9037# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1908 a_28131_n1900# a_29115_n2414# a_29066_n2398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1909 a_5910_n6212# a_5489_n6212# a_5174_n6216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1910 a_3824_n7149# a_4077_n7353# a_2882_n7581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1911 a_21981_n2050# a_21913_n2561# a_21991_n3500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1912 gnd d0 a_39352_2239# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1913 vdd d2 a_23187_1926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1914 a_22930_n2639# a_23120_n2063# a_23075_n1859# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1915 gnd a_13060_7452# a_12852_7452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1916 gnd d0 a_24264_5502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1917 a_10679_n4524# a_10466_n4524# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1918 a_25888_7150# a_25675_7150# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1919 a_12914_4857# a_13171_4667# a_12778_4169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1920 a_16814_1926# a_16601_1926# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1921 a_5701_9375# a_5488_9375# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1922 a_32963_6356# a_33148_6854# a_33099_7044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1923 gnd d0 a_4077_n8456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1924 a_23072_n8477# a_23325_n8681# a_22927_n9257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1925 a_36858_n6508# a_36645_n6508# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1926 a_13853_n5690# a_13856_n4948# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1927 a_34043_n5483# a_34039_n5671# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1928 gnd a_18085_8609# a_17877_8609# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1929 vdd a_23217_3016# a_23009_3016# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1930 a_15204_n7324# a_15732_n7320# a_15940_n7320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1931 gnd d0 a_14110_n2946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1932 a_21669_2977# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1933 gnd d0 a_34295_8267# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1934 a_15205_5078# a_15734_4968# a_15942_4968# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1935 a_8882_6129# a_8878_6306# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1936 a_17861_n3794# a_18118_n3810# a_17861_n5994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1937 a_23068_7039# a_24055_6605# a_24006_6795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1938 a_856_1059# a_435_1059# a_122_1165# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1939 gnd a_18226_8017# a_18018_8017# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1940 a_30333_n9470# a_30334_n9013# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1941 a_117_n9027# a_644_n9480# a_852_n9480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1942 a_1584_6884# a_1371_6884# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1943 vdd d0 a_24266_n3476# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1944 a_10147_9449# a_10147_9220# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1945 a_15940_n10080# a_15519_n10080# a_15203_n9760# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1946 gnd d0 a_39353_n3522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1947 a_31911_7394# a_31698_7394# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1948 a_20619_7109# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1949 a_11545_1885# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1950 a_28124_7080# a_28381_6890# a_27988_6392# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1951 a_24012_2206# a_24008_2383# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1952 a_6568_6333# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1953 a_35391_4830# a_35920_4949# a_36128_4949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1954 a_2741_n9276# a_2931_n8700# a_2886_n8496# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1955 a_30648_n9466# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1956 vdd d2 a_18086_6403# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1957 a_34040_4045# a_34297_3855# a_33105_3558# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1958 gnd a_24264_7159# a_24056_7159# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1959 a_25359_8550# a_25886_8802# a_26094_8802# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1960 vdd a_34296_6061# a_34088_6061# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1961 a_38160_4702# a_38413_4689# a_38020_4191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1962 gnd d3 a_18118_3081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1963 a_6750_7449# a_6537_7449# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1964 a_1724_n9198# a_1511_n9198# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1965 vdd a_9136_3910# a_8928_3910# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1966 a_10884_n7279# a_10463_n7279# a_10148_n7283# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1967 a_31071_5457# a_31802_5767# a_32010_5767# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1968 a_35391_n6661# a_35391_n6432# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1969 gnd a_3142_1353# a_2934_1353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1970 a_31942_n6978# a_31729_n6978# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1971 a_27986_2157# a_28176_1375# a_28127_1565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1972 a_31073_2702# a_31803_2458# a_32011_2458# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1973 a_18908_4654# a_19165_4464# a_17970_4898# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1974 a_18907_n8486# a_18912_n7749# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1975 a_2884_2646# a_3871_2212# a_3822_2402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1976 a_10886_3270# a_10465_3270# a_10150_3475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1977 gnd a_14107_8835# a_13899_8835# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1978 vdd a_13032_n2679# a_12824_n2679# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1979 a_16568_7454# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1980 a_27036_3597# a_26968_4108# a_27052_3137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1981 gnd d3 a_3031_3035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1982 gnd a_19164_n10159# a_18956_n10159# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1983 a_5705_1654# a_5492_1654# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1984 a_25675_4390# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1985 vdd a_38271_n9319# a_38063_n9319# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1986 a_8880_9438# a_8876_9615# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1987 a_35393_n2436# a_35920_n2889# a_36128_n2889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1988 a_13851_9579# a_13854_8848# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1989 a_34038_n8980# a_34295_n8996# a_33103_n8482# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1990 a_3824_n7149# a_3820_n7337# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1991 a_13853_n5690# a_14110_n5706# a_12918_n5192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1992 a_7799_n4905# a_7989_n4329# a_7944_n4125# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1993 gnd d0 a_24266_1090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1994 a_1481_7408# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1995 a_5910_n7869# a_5489_n7869# a_5173_n7778# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1996 a_5703_4963# a_5490_4963# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X1997 a_35393_n2436# a_35393_n2249# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X1998 a_19208_288# a_18995_288# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1999 vdd d0 a_4076_8830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2000 a_15520_n8977# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2001 vdd d0 a_14110_n6809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2002 a_15206_3746# a_15735_3865# a_15943_3865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2003 gnd a_18087_4197# a_17879_4197# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2004 a_15940_n8423# a_16671_n8733# a_16879_n8733# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2005 a_3826_n6600# a_3822_n6788# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2006 a_2672_n10656# a_2622_n10672# a_1902_n5908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2007 a_5910_4409# a_5489_4409# a_5175_4157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2008 gnd d0 a_34297_3855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2009 a_16672_4724# a_16459_4724# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2010 a_36128_n6752# a_35707_n6752# a_35391_n6432# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2011 a_23070_2627# a_24057_2193# a_24008_2383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2012 gnd a_23217_n5945# a_23009_n5945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2013 a_17969_7104# a_18956_6670# a_18911_6683# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2014 gnd a_33356_n8686# a_33148_n8686# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2015 a_1586_2472# a_1373_2472# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2016 gnd a_29320_4440# a_29112_4440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2017 a_31913_2982# a_31700_2982# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2018 a_10465_n5627# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2019 a_26828_n3194# a_26615_n3194# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2020 a_16598_n9244# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2021 a_27985_n4886# a_28175_n4310# a_28130_n4106# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2022 vdd a_9136_n3536# a_8928_n3536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2023 a_5173_n8422# a_5173_n7965# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2024 a_13854_2961# a_14111_2771# a_12919_2474# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2025 vdd d2 a_18088_1991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2026 a_23070_n3150# a_23327_n3166# a_22934_n2451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2027 a_11403_4683# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2028 a_34041_9383# a_35389_9471# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2029 a_30863_n6157# a_30650_n6157# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2030 a_26096_n8953# a_25675_n8953# a_25359_n8862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2031 a_10886_n6730# a_10465_n6730# a_10149_n6639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2032 a_5175_n4010# a_5703_n4006# a_5911_n4006# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2033 a_5178_1206# a_5704_1100# a_5912_1100# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2034 a_33104_5764# a_34088_6061# a_34039_6251# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2035 a_20306_n1744# a_20834_n1740# a_21042_n1740# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2036 a_6752_3037# a_6539_3037# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2037 vdd a_13060_7452# a_12852_7452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2038 a_1791_n9790# a_1370_n9790# a_853_n10034# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2039 gnd d0 a_19165_n5193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2040 a_10147_n9719# a_10147_n9489# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2041 a_15206_n3558# a_15734_n4011# a_15942_n4011# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2042 vdd d1 a_23327_n4269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2043 a_25674_n8399# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2044 a_20306_n1974# a_20835_n2294# a_21043_n2294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2045 a_1511_8498# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2046 vdd a_28384_n2104# a_28176_n2104# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2047 vdd a_38411_9101# a_38203_9101# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2048 gnd d1 a_18228_3605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2049 gnd d0 a_4080_n1838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2050 a_7798_n7111# a_7988_n6535# a_7939_n6519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2051 gnd d0 a_24263_n10094# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2052 gnd a_19165_n9056# a_18957_n9056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2053 gnd d4 a_38304_n5991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2054 a_16890_n5777# a_16570_n3742# a_16897_n3742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2055 a_7800_2176# a_7990_1394# a_7945_1407# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2056 a_34040_8829# a_34293_8816# a_33098_9250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2057 a_12918_4680# a_13902_4977# a_13857_4990# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2058 a_1584_7987# a_1371_7987# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2059 gnd d1 a_3141_3559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2060 a_36127_8258# a_35706_8258# a_35390_8139# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2061 vdd a_29318_8852# a_29110_8852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2062 a_39095_2429# a_39101_1703# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2063 vdd d0 a_4078_4418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2064 a_23069_n6459# a_24056_n6231# a_24011_n6027# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2065 a_17834_4210# a_18019_4708# a_17970_4898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2066 a_5911_3306# a_5490_3306# a_5175_3511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2067 a_16989_n5954# a_17917_n10718# a_14710_n10722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2068 a_28014_n8182# a_28033_n7108# a_27984_n7092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2069 a_26097_4944# a_26827_4700# a_27035_4700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2070 a_31943_4072# a_31730_4072# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2071 a_16672_n6527# a_16459_n6527# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2072 a_25887_6596# a_25674_6596# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2073 a_8879_n9396# a_8875_n9584# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2074 a_29063_7390# a_29066_6659# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2075 a_21041_4903# a_20620_4903# a_20304_5013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2076 a_16879_8033# a_16811_8544# a_16895_7573# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2077 a_17971_2692# a_18958_2258# a_18913_2271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2078 a_20306_1891# a_20306_1704# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2079 a_22088_n5889# a_21667_n5889# a_21989_n5712# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2080 vdd d3 a_18118_3081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2081 vdd a_3142_1353# a_2934_1353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2082 a_25889_n3987# a_25676_n3987# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2083 vdd d0 a_14108_9389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2084 a_18914_n3337# a_19167_n3541# a_17975_n3027# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2085 gnd d0 a_34295_n6236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2086 gnd d2 a_23185_n7067# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2087 a_5912_n3457# a_6642_n3213# a_6850_n3213# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2088 a_27986_2157# a_28176_1375# a_28131_1388# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2089 a_20303_n7259# a_20304_n6802# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2090 a_1792_7987# a_1724_8498# a_1808_7527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2091 a_20622_n2294# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2092 a_2884_2646# a_3871_2212# a_3826_2225# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2093 vdd a_24265_n4025# a_24057_n4025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2094 vdd d3 a_3031_3035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2095 a_20618_6555# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2096 gnd a_28242_n4902# a_28034_n4902# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2097 a_1696_2996# a_1483_2996# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2098 a_24011_n6027# a_24007_n6215# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2099 gnd d0 a_19167_n4644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2100 a_11834_n5736# a_11514_n3701# a_11836_n3524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2101 a_120_n1993# a_120_n1763# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2102 a_2882_n8684# a_3869_n8456# a_3820_n8440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2103 a_35391_4600# a_35919_4395# a_36127_4395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2104 vdd d2 a_33215_8549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2105 a_5909_9375# a_6639_9131# a_6847_9131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2106 a_15519_n7320# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2107 a_12915_n3174# a_13902_n2946# a_13853_n2930# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2108 gnd a_13172_n4293# a_12964_n4293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2109 vdd d1 a_18226_n7643# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2110 a_5174_6176# a_5174_5947# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2111 a_33102_n9585# a_33355_n9789# a_32962_n9074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2112 vdd a_33358_n3171# a_33150_n3171# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2113 gnd a_24266_n1819# a_24058_n1819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2114 a_2882_7058# a_3139_6868# a_2746_6370# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2115 a_1513_4086# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2116 a_432_n8377# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2117 a_35390_n8638# a_35919_n8958# a_36127_n8958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2118 a_10884_n10039# a_10463_n10039# a_10147_n9719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2119 a_15205_n5348# a_15734_n5668# a_15942_n5668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2120 a_10149_n5077# a_10150_n4620# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2121 gnd d0 a_34297_n3481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2122 vdd a_19166_n2987# a_18958_n2987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2123 vdd a_13170_7976# a_12962_7976# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2124 gnd a_29320_n5169# a_29112_n5169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2125 a_32995_n3546# a_33248_n3750# a_32991_n5934# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2126 a_855_n2862# a_434_n2862# a_119_n2866# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2127 a_37076_n5758# a_36967_n5935# a_37175_n5935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2128 a_35921_2743# a_35708_2743# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2129 a_12912_9269# a_13899_8835# a_13854_8848# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2130 a_21981_n2050# a_21560_n2050# a_21042_n1740# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2131 a_5173_n7778# a_5702_n7869# a_5910_n7869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2132 a_18909_n5731# a_18912_n4989# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2133 vdd d0 a_9137_1704# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2134 vdd a_8085_7488# a_7877_7488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2135 a_10677_n7833# a_10464_n7833# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2136 a_853_9334# a_432_9334# a_116_9444# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2137 vdd a_29320_4440# a_29112_4440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2138 a_16881_n4321# a_16460_n4321# a_15943_n4565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2139 a_29064_5184# a_29067_4453# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2140 a_35922_n2340# a_35709_n2340# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2141 a_13853_2407# a_13859_1681# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2142 a_35389_n9511# a_35390_n9054# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2143 a_32022_n3505# a_31731_n2566# a_32011_n3158# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2144 a_25889_2184# a_25676_2184# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2145 gnd a_18086_n7132# a_17878_n7132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2146 a_7834_5289# a_8087_5276# a_7060_541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2147 a_6642_n3213# a_6429_n3213# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2148 a_16881_3621# a_16813_4132# a_16897_3161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2149 gnd a_18116_7493# a_17908_7493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2150 a_33104_5764# a_34088_6061# a_34043_6074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2151 a_22934_n2451# a_23187_n2655# a_22960_n3729# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2152 a_25359_n7946# a_25359_n7759# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2153 a_35707_2189# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2154 a_38019_6397# a_38204_6895# a_38155_7085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2155 a_38019_n6909# a_38272_n7113# a_38045_n8187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2156 vdd a_39351_8308# a_39143_8308# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2157 a_10886_4927# a_10465_4927# a_10149_4808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2158 a_647_n3965# a_434_n3965# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2159 a_35707_n2889# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2160 a_20619_5452# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2161 vdd d0 a_14107_n9564# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2162 a_1794_3575# a_1726_4086# a_1810_3115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2163 a_10149_n5536# a_10678_n5627# a_10886_n5627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2164 a_25890_n4541# a_25677_n4541# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2165 a_23073_n5168# a_24057_n5682# a_24008_n5666# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2166 gnd a_39352_2239# a_39144_2239# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2167 a_28020_5270# a_28063_7469# a_28014_7659# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2168 a_36127_n7855# a_36857_n7611# a_37065_n7611# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2169 a_6851_1410# a_6430_1410# a_5913_1654# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2170 a_32025_n5894# a_31911_n5894# a_32119_n5894# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2171 gnd a_24264_5502# a_24056_5502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2172 a_34043_n3826# a_34296_n4030# a_33101_n4258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2173 a_6783_n2621# a_6570_n2621# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2174 vdd d2 a_33217_4137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2175 a_12918_n6295# a_13902_n6809# a_13857_n6605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2176 a_13857_3333# a_14110_3320# a_12915_3754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2177 a_25675_7150# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2178 vdd d1 a_23325_6849# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2179 a_11825_n4280# a_11404_n4280# a_10886_n3970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2180 a_16601_1926# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2181 a_16458_n8733# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2182 a_855_6025# a_1585_5781# a_1793_5781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2183 a_2774_n3748# a_2793_n2674# a_2748_n2470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2184 a_6426_n9831# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2185 a_37066_n5405# a_36645_n5405# a_36128_n5649# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2186 a_29063_n5153# a_29320_n5169# a_28125_n5397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2187 a_32991_n5934# a_33040_n3750# a_32995_n3546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2188 a_11725_n8113# a_11512_n8113# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2189 a_17975_n4130# a_18228_n4334# a_17830_n4910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2190 gnd a_24263_n8437# a_24055_n8437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2191 a_13851_n10102# a_13854_n9360# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2192 a_30333_n10116# a_34037_n10083# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2193 a_35392_2624# a_35392_2394# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2194 a_10151_1499# a_10680_1618# a_10888_1618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2195 a_857_1613# a_436_1613# a_120_1494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2196 a_20832_8212# a_20619_8212# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2197 a_31803_n4261# a_31590_n4261# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2198 gnd a_34295_8267# a_34087_8267# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2199 a_8880_n7190# a_9133_n7394# a_7938_n7622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2200 a_7942_6922# a_8195_6909# a_7802_6411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2201 a_2745_n9088# a_2998_n9292# a_2776_n7972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2202 vdd d0 a_29320_n6272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2203 a_38016_n4891# a_38206_n4315# a_38157_n4299# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2204 a_36645_5808# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2205 a_25359_7447# a_25359_7260# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2206 a_24007_n5112# a_24264_n5128# a_23069_n5356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2207 a_17865_n5806# a_18118_n6010# a_17660_n10702# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2208 a_1371_6884# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2209 a_21558_4659# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2210 a_648_2716# a_435_2716# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2211 a_1803_7408# a_1512_6292# a_1792_6884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2212 a_855_4922# a_434_4922# a_118_5032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2213 a_853_n10034# a_1583_n9790# a_1791_n9790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2214 a_11823_n8692# a_11755_n9203# a_11839_n8113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2215 a_36129_2743# a_36859_2499# a_37067_2499# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2216 a_20834_n4500# a_20621_n4500# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2217 gnd d4 a_28273_5257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2218 a_856_n4519# a_1586_n4275# a_1794_n4275# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2219 a_853_n10034# a_432_n10034# a_116_n9943# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2220 a_21771_n6462# a_21558_n6462# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2221 a_29067_n6068# a_29063_n6256# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2222 a_17970_n5421# a_18957_n5193# a_18908_n5177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2223 gnd a_18118_3081# a_17910_3081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2224 a_1795_n2069# a_1374_n2069# a_857_n2313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2225 vdd d0 a_29321_6097# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2226 a_10887_3824# a_10466_3824# a_10150_3934# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2227 vdd d0 a_29322_n3517# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2228 a_30336_n2852# a_30864_n2848# a_31072_n2848# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2229 a_12919_2474# a_13172_2461# a_12779_1963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2230 a_11839_5332# a_11512_7413# a_11834_7413# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2231 a_22931_n9069# a_23184_n9273# a_22962_n7953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2232 gnd d1 a_13171_n6499# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2233 a_28016_n3770# a_28273_n3786# a_28016_n5970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2234 vdd d0 a_9132_8871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2235 vdd d1 a_33357_n5377# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2236 a_13856_n6051# a_14109_n6255# a_12914_n6483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2237 a_21989_7389# a_21698_6273# a_21978_6865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2238 a_5910_n6212# a_5489_n6212# a_5174_n5759# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2239 a_5492_1654# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2240 a_39098_n7730# a_39094_n7918# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2241 a_21980_n3153# a_21913_n2561# a_21991_n3500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2242 a_26966_n9220# a_26753_n9220# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2243 a_28016_5447# a_28065_3057# a_28016_3247# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2244 a_26826_8009# a_26613_8009# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2245 a_16457_9136# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2246 a_30334_n9013# a_30334_n8826# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2247 a_28128_6903# a_29112_7200# a_29067_7213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2248 gnd a_24266_1090# a_24058_1090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2249 a_6780_n9239# a_6567_n9239# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2250 a_5176_1535# a_5176_1305# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2251 a_5703_n4006# a_5490_n4006# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2252 a_26829_n2091# a_26616_n2091# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2253 vdd d1 a_23327_2437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2254 a_5490_4963# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2255 a_16895_n8154# a_16781_n8154# a_16895_n5954# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2256 a_4799_n1525# a_5704_n1800# a_5912_n1800# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2257 a_2776_n7972# a_2790_n9292# a_2745_n9088# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2258 vdd a_4076_8830# a_3868_8830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2259 vdd a_19165_n9056# a_18957_n9056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2260 a_26829_1391# a_26616_1391# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2261 gnd d1 a_33356_7957# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2262 a_8882_n6641# a_9135_n6845# a_7943_n6331# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2263 a_15731_8826# a_15518_8826# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2264 a_854_n8931# a_433_n8931# a_117_n8840# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2265 a_34045_1662# a_34298_1649# a_33106_1352# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2266 gnd a_34297_3855# a_34089_3855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2267 a_19441_n829# a_20582_n10911# a_9875_n10838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2268 a_22928_n7051# a_23118_n6475# a_23069_n6459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2269 a_21559_3556# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2270 a_36647_1396# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2271 a_38160_5805# a_39144_6102# a_39095_6292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2272 a_15204_n8886# a_15204_n8657# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2273 a_16982_546# a_16769_546# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2274 a_7830_5466# a_8087_5276# a_7060_541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2275 gnd d0 a_24263_7708# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2276 a_1373_2472# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2277 a_20304_6116# a_20304_5887# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2278 a_31700_2982# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2279 a_12913_7063# a_13170_6873# a_12777_6375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2280 a_31070_n10020# a_30649_n10020# a_30333_n9929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2281 a_10151_1728# a_10151_1499# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2282 a_18913_2271# a_19166_2258# a_17971_2692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2283 a_30648_n9466# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2284 vdd a_39351_n6277# a_39143_n6277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2285 a_15207_1310# a_15735_1105# a_15943_1105# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2286 a_17975_n4130# a_18959_n4644# a_18910_n4628# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2287 vdd d0 a_39353_2793# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2288 a_119_n4428# a_648_n4519# a_856_n4519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2289 a_37168_527# a_36955_527# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2290 a_25360_n5324# a_25360_n5094# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2291 a_8883_1163# a_8879_1340# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2292 a_16670_n9836# a_16457_n9836# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2293 a_6866_n3737# a_6569_n4827# a_6849_n5419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2294 a_852_8780# a_431_8780# a_117_8528# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2295 a_17834_n4722# a_18019_n5437# a_17970_n5421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2296 a_26097_4944# a_25676_4944# a_25360_4825# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2297 a_5174_4844# a_5174_4614# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2298 a_10149_4578# a_10150_4121# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2299 gnd d0 a_29321_n5723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2300 a_32112_486# a_31899_486# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2301 a_11834_5213# a_11514_3001# a_11836_3001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2302 a_13853_3510# a_14110_3320# a_12915_3754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2303 a_35706_n8958# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2304 gnd d0 a_4077_6624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2305 gnd a_4078_n5147# a_3870_n5147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2306 vdd d0 a_9134_4459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2307 a_13856_8299# a_14109_8286# a_12917_7989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2308 a_32010_n6467# a_31589_n6467# a_31072_n6711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2309 a_33106_n1864# a_33359_n2068# a_32961_n2644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2310 a_6567_8539# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2311 a_117_7882# a_117_7425# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2312 a_21979_n5359# a_21558_n5359# a_21041_n5603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2313 a_36754_n5935# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2314 a_10888_n2318# a_10467_n2318# a_10151_n1998# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2315 a_16458_8033# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2316 gnd a_18228_3605# a_18020_3605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2317 a_20620_n5603# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2318 a_5489_n7869# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2319 a_18914_3928# a_18910_4105# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2320 a_17970_4898# a_18957_4464# a_18908_4654# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2321 a_13851_n7342# a_13857_n6605# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2322 a_13855_1858# a_13858_1127# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2323 a_1371_7987# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2324 a_21041_n6706# a_20620_n6706# a_20304_n6615# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2325 a_32011_n3158# a_31590_n3158# a_31072_n2848# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2326 a_33104_n6276# a_34088_n6790# a_34043_n6586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2327 vdd d1 a_28383_n4310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2328 vdd a_4078_4418# a_3870_4418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2329 gnd a_13030_n7091# a_12822_n7091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2330 a_1586_n3172# a_1373_n3172# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2331 a_2883_4852# a_3870_4418# a_3821_4608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2332 a_33098_n9773# a_34085_n9545# a_34036_n9529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2333 a_15733_4414# a_15520_4414# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2334 a_15941_n8977# a_16671_n8733# a_16879_n8733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2335 a_31730_4072# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2336 a_11614_n9795# a_11401_n9795# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2337 a_6958_n5949# a_6537_n5949# a_6859_n5772# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2338 a_1810_n3696# a_1513_n4786# a_1794_n4275# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2339 a_25674_6596# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2340 a_21980_2453# a_21559_2453# a_21041_2143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2341 a_1372_n6481# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2342 vdd d2 a_3001_1945# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2343 a_11822_9095# a_11755_8503# a_11839_7532# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2344 gnd d0 a_24265_3296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2345 vdd a_18118_3081# a_17910_3081# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2346 a_10465_n5627# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2347 vdd a_4079_n6804# a_3871_n6804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2348 a_5702_7169# a_5489_7169# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2349 a_12915_2651# a_13172_2461# a_12779_1963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2350 vdd a_14108_9389# a_13900_9389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2351 a_3822_n4028# a_4079_n4044# a_2884_n4272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2352 a_3826_4985# a_3822_5162# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2353 a_7803_n4717# a_8056_n4921# a_7834_n3601# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2354 a_31698_n5894# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2355 a_3827_n3291# a_3823_n3479# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2356 a_26098_3841# a_25677_3841# a_25361_3951# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2357 vout a_19119_n829# a_19441_n829# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2358 a_5487_8821# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2359 a_27050_5349# a_26723_7430# a_27045_7430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2360 a_10150_4121# a_10677_4373# a_10885_4373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2361 a_1483_2996# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2362 a_10677_7133# a_10464_7133# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2363 a_26096_n8953# a_25675_n8953# a_25359_n8633# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2364 vdd a_39351_n7934# a_39143_n7934# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2365 a_23069_4833# a_24056_4399# a_24007_4589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2366 a_35393_1937# a_35393_1750# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2367 a_10885_5476# a_11616_5786# a_11824_5786# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2368 a_17968_9310# a_18955_8876# a_18910_8889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2369 vdd a_33215_8549# a_33007_8549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2370 a_12919_2474# a_13903_2771# a_13854_2961# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2371 a_1585_4678# a_1372_4678# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2372 gnd a_29319_6646# a_29111_6646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2373 a_7938_n8725# a_8195_n8741# a_7797_n9317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2374 a_30335_n6391# a_30335_n6161# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2375 a_6738_541# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2376 a_1694_n8108# a_1481_n8108# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2377 a_22858_n10637# a_25122_n10714# a_24964_n10698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2378 a_31072_n6711# a_30651_n6711# a_30335_n6620# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2379 a_6569_4127# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2380 a_36858_n6508# a_36645_n6508# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2381 a_34041_7726# a_34037_7903# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2382 a_5911_n2903# a_5490_n2903# a_5175_n2907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2383 a_23074_2450# a_24058_2747# a_24013_2760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2384 a_3825_5534# a_3821_5711# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2385 a_25360_6344# a_25887_6596# a_26095_6596# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2386 a_35392_n4226# a_35392_n3996# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2387 a_12778_4169# a_12963_4667# a_12918_4680# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2388 a_15205_n6867# a_15732_n7320# a_15940_n7320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2389 a_8882_n3881# a_8878_n4069# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2390 a_10150_n3974# a_10678_n3970# a_10886_n3970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2391 a_16890_n5777# a_16570_n3742# a_16892_n3565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2392 a_30650_n6157# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2393 a_33103_7970# a_34087_8267# a_34038_8457# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2394 vdd d0 a_39350_n7380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2395 a_15521_n4011# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2396 gnd a_18225_n9849# a_18017_n9849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2397 gnd d0 a_4081_n2392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2398 a_18907_n10143# a_18910_n9401# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2399 vdd a_9137_1704# a_8929_1704# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2400 a_5175_n4469# a_5175_n4240# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2401 a_8881_8335# a_9134_8322# a_7942_8025# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2402 a_20304_n6802# a_20304_n6615# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2403 a_15522_n4565# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2404 vdd a_38414_n3212# a_38206_n3212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2405 gnd a_29322_n1860# a_29114_n1860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2406 a_35389_n10157# a_35389_n9970# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2407 a_38051_n3587# a_38304_n3791# a_38047_n5975# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2408 a_25676_2184# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2409 a_30651_n2848# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2410 a_12773_n7075# a_12963_n6499# a_12914_n6483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2411 a_4679_n10717# a_7678_n10713# a_6958_n5949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2412 gnd d2 a_33216_6343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2413 a_3827_2779# a_3823_2956# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2414 vdd d0 a_4077_6624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2415 a_13852_8476# a_14109_8286# a_12917_7989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2416 a_15207_1540# a_15736_1659# a_15944_1659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2417 a_853_n7274# a_1584_n7584# a_1792_n7584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2418 a_26096_7150# a_26826_6906# a_27034_6906# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2419 a_31942_6278# a_31729_6278# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2420 a_34042_4417# a_34295_4404# a_33100_4838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2421 a_16568_n8154# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2422 a_35707_6052# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2423 a_16673_2518# a_16460_2518# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2424 a_1586_3575# a_1373_3575# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2425 a_30865_n1745# a_30652_n1745# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2426 a_5491_n1800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2427 a_30336_3456# a_30864_3251# a_31072_3251# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2428 a_21040_7109# a_20619_7109# a_20303_7219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2429 gnd d0 a_14110_6080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2430 a_17970_4898# a_18957_4464# a_18912_4477# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2431 vdd a_33217_4137# a_33009_4137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2432 vdd a_23325_6849# a_23117_6849# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2433 a_27990_n2492# a_28243_n2696# a_28016_n3770# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2434 gnd a_29321_2234# a_29113_2234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2435 a_17863_n8018# a_17877_n9338# a_17828_n9322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2436 a_30337_n1979# a_30337_n1749# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2437 a_1902_5208# a_1895_500# a_2103_500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2438 a_11403_n6486# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2439 a_32790_n10642# a_33040_n5950# a_32991_n5934# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2440 a_3821_n7891# a_4078_n7907# a_2886_n7393# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2441 a_36645_n6508# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2442 a_16460_n3218# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2443 a_25362_1932# a_25889_2184# a_26097_2184# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2444 gnd a_24267_n2373# a_24059_n2373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2445 a_855_n2862# a_434_n2862# a_120_n2409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2446 a_32963_n6868# a_33148_n7583# a_33099_n7567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2447 vdd d0 a_24262_n9540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2448 a_37081_n5935# a_36967_n5935# a_37175_n5935# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2449 a_39099_n3867# a_39352_n4071# a_38157_n4299# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2450 a_33105_3558# a_34089_3855# a_34040_4045# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2451 a_10677_n7833# a_10464_n7833# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2452 a_435_2716# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2453 vdd d0 a_4078_n9010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2454 a_12703_n10661# a_14967_n10738# a_9776_n10838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2455 a_16881_n4321# a_16460_n4321# a_15942_n4011# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2456 a_11825_n3177# a_11758_n2585# a_11836_n3524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2457 vdd a_23326_n5372# a_23118_n5372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2458 a_8883_3923# a_9136_3910# a_7944_3613# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2459 a_16781_n8154# a_16568_n8154# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2460 a_120_n2222# a_120_n1993# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2461 vdd d1 a_28380_9096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2462 gnd a_28273_5257# a_28065_5257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2463 a_24014_n2169# a_24010_n2357# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2464 a_3822_n4028# a_3827_n3291# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2465 a_5053_480# a_4632_480# a_4954_480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2466 a_32022_n3505# a_31731_n2566# a_32012_n2055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2467 vdd d0 a_19167_n1884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2468 a_12772_8758# a_13029_8568# a_12807_7465# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2469 a_16674_n2115# a_16461_n2115# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2470 a_6642_n3213# a_6429_n3213# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2471 a_2886_n8496# a_3870_n9010# a_3821_n8994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2472 a_8882_5026# a_8878_5203# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2473 a_18908_4654# a_18914_3928# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2474 a_35920_4949# a_35707_4949# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2475 gnd d2 a_33218_1931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2476 gnd d1 a_23326_4643# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2477 vdd d1 a_28383_2478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2478 a_12919_2474# a_13903_2771# a_13858_2784# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2479 a_19886_n1571# a_20834_n1740# a_21042_n1740# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2480 vdd a_29319_6646# a_29111_6646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2481 vdd a_9132_8871# a_8924_8871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2482 a_25890_n4541# a_25677_n4541# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2483 gnd d1 a_38412_7998# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2484 a_26096_5493# a_26827_5803# a_27035_5803# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2485 a_26097_n2884# a_26828_n3194# a_27036_n3194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2486 a_5912_1100# a_5491_1100# a_5176_1305# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2487 a_26613_8009# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2488 vdd d1 a_3141_n4288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2489 a_30862_n8363# a_30649_n8363# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2490 a_5174_n5759# a_5702_n6212# a_5910_n6212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2491 gnd d1 a_8197_n3226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2492 a_16880_5827# a_16812_6338# a_16890_7454# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2493 a_16458_n8733# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2494 vdd d1 a_33359_n2068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2495 a_6861_3037# a_6570_1921# a_6850_2513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2496 vdd a_23327_2437# a_23119_2437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2497 a_27987_n9110# a_28240_n9314# a_28018_n7994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2498 a_36130_1640# a_35709_1640# a_35393_1750# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2499 a_37066_n5405# a_36645_n5405# a_36127_n5095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2500 a_36787_1907# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2501 vdd a_34297_n4584# a_34089_n4584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2502 a_13855_9402# a_15203_9490# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2503 a_15734_n6771# a_15521_n6771# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2504 a_35391_n5558# a_35391_n5329# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2505 vdd d1 a_38413_n5418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2506 a_26616_1391# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2507 gnd a_33356_7957# a_33148_7957# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2508 a_8877_8512# a_9134_8322# a_7942_8025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2509 a_20618_7658# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2510 a_18907_n7383# a_18913_n6646# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2511 a_20619_4349# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2512 a_20305_n4180# a_20305_n3950# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2513 gnd d1 a_18225_9120# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2514 a_35919_8258# a_35706_8258# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2515 a_24011_n6027# a_24264_n6231# a_23069_n6459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2516 gnd a_24263_7708# a_24055_7708# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2517 a_18907_n7383# a_19164_n7399# a_17969_n7627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2518 a_35392_2394# a_35920_2189# a_36128_2189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2519 a_21994_5308# a_21667_7389# a_21994_7508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2520 vdd d2 a_33216_6343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2521 a_32995_n5746# a_33038_n8162# a_32989_n8146# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2522 a_16890_5254# a_16570_3042# a_16892_3042# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2523 a_854_8231# a_1584_7987# a_1792_7987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2524 gnd d0 a_9133_6665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2525 a_27035_4700# a_26614_4700# a_26096_4390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2526 a_11822_n9795# a_11755_n9203# a_11839_n8113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2527 a_15203_n9989# a_15732_n10080# a_15940_n10080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2528 a_23070_n3150# a_24057_n2922# a_24012_n2718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2529 a_21771_n6462# a_21558_n6462# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2530 vdd a_39353_2793# a_39145_2793# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2531 a_16895_7573# a_16598_8544# a_16878_9136# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2532 a_856_3819# a_435_3819# a_119_3700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2533 a_25358_n9736# a_25358_n9506# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2534 a_2882_n8684# a_3139_n8700# a_2741_n9276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2535 vdd d0 a_19164_n8502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2536 a_39101_n2215# a_39097_n2403# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2537 a_24011_5515# a_24007_5692# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2538 a_35921_3846# a_35708_3846# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2539 a_39097_9424# a_39350_9411# a_38158_9114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2540 a_36126_n10061# a_35705_n10061# a_35389_n9741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2541 a_26099_n2335# a_26829_n2091# a_27037_n2091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2542 a_31698_7394# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2543 a_2883_n6478# a_3870_n6250# a_3825_n6046# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2544 vdd d0 a_14110_6080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2545 gnd a_3029_n8176# a_2821_n8176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2546 a_2741_8753# a_2931_7971# a_2882_8161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2547 vdd a_18228_n4334# a_18020_n4334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2548 a_1808_7527# a_1511_8498# a_1791_9090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2549 gnd a_4077_6624# a_3869_6624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2550 a_854_7128# a_433_7128# a_117_7238# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2551 vdd a_29321_2234# a_29113_2234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2552 a_11823_7992# a_11402_7992# a_10885_8236# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2553 vdd a_9134_4459# a_8926_4459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2554 a_27988_n6904# a_28173_n7619# a_28128_n7415# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2555 a_11615_n8692# a_11402_n8692# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2556 a_15519_n7320# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2557 a_10465_n3970# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2558 a_26098_1081# a_26829_1391# a_27037_1391# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2559 a_29065_8865# a_29318_8852# a_28123_9286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2560 a_12913_8166# a_13900_7732# a_13851_7922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2561 a_5173_n7319# a_5174_n6862# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2562 gnd d0 a_24266_n4579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2563 gnd a_18229_n2128# a_18021_n2128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2564 a_5172_9256# a_5701_9375# a_5909_9375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2565 a_1902_n5908# a_2830_n10672# a_2672_n10656# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2566 vdd d0 a_29320_8303# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2567 a_12918_4680# a_13171_4667# a_12778_4169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2568 vdd d5 a_17917_n10718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2569 gnd a_9134_n5188# a_8926_n5188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2570 a_31802_4664# a_31589_4664# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2571 vdd d1 a_23325_n7578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2572 a_5173_n7549# a_5702_n7869# a_5910_n7869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2573 gnd d1 a_38412_n7624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2574 a_35921_n1786# a_35708_n1786# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2575 a_23068_8142# a_24055_7708# a_24010_7721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2576 a_38162_n1905# a_38415_n2109# a_38017_n2685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2577 a_15520_4414# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2578 a_854_n8931# a_433_n8931# a_117_n8611# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2579 gnd a_39352_n2968# a_39144_n2968# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2580 a_21994_7508# a_21697_8479# a_21977_9071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2581 a_34038_n5117# a_34044_n4380# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2582 a_21039_n8358# a_20618_n8358# a_20303_n7905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2583 a_35922_n2340# a_35709_n2340# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2584 a_24009_8824# a_24005_9001# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2585 gnd d1 a_3138_n9803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2586 a_18909_n6834# a_19166_n6850# a_17974_n6336# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2587 a_7801_n9129# a_7986_n9844# a_7937_n9828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2588 a_20832_n5049# a_20619_n5049# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2589 a_6849_n6522# a_6428_n6522# a_5911_n6766# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2590 a_28127_9109# a_29111_9406# a_29066_9419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2591 a_32020_7394# a_31911_7394# a_32025_5313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2592 gnd a_24265_3296# a_24057_3296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2593 a_27137_522# a_26924_522# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2594 a_13858_1127# a_14111_1114# a_12916_1548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2595 vdd d1 a_23326_4643# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2596 vdd a_33218_n2660# a_33010_n2660# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2597 vdd d1 a_3139_6868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2598 a_7834_n5801# a_7877_n8217# a_7832_n8013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2599 a_28127_n9621# a_29111_n10135# a_29062_n10119# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2600 a_856_3819# a_1586_3575# a_1794_3575# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2601 a_38160_n6317# a_39144_n6831# a_39099_n6627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2602 gnd d0 a_9135_2253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2603 a_38156_5982# a_38413_5792# a_38015_6574# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2604 a_38154_n9814# a_39141_n9586# a_39092_n9570# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2605 a_13857_n6605# a_14110_n6809# a_12918_n6295# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2606 a_26828_3597# a_26615_3597# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2607 a_7060_541# a_7879_5276# a_7830_5466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2608 a_20833_6006# a_20620_6006# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2609 a_16670_n9836# a_16457_n9836# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2610 a_6866_n3737# a_6569_n4827# a_6850_n4316# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2611 a_10464_7133# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2612 gnd a_23185_n7067# a_22977_n7067# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2613 a_13857_n6605# a_13853_n6793# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2614 a_6864_7568# a_6750_7449# a_6864_5368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2615 a_26096_n8953# a_26826_n8709# a_27034_n8709# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2616 a_10886_n6730# a_11616_n6486# a_11824_n6486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2617 a_15205_n5577# a_15205_n5348# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2618 a_38159_8011# a_39143_8308# a_39094_8498# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2619 a_10147_n10135# a_13851_n10102# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2620 gnd a_14110_n4049# a_13902_n4049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2621 a_1372_4678# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2622 a_10148_n7283# a_10676_n7279# a_10884_n7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2623 a_1810_3115# a_1513_4086# a_1793_4678# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2624 vdd d0 a_34296_n6790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2625 gnd a_4079_2212# a_3871_2212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2626 a_32010_n6467# a_31589_n6467# a_31071_n6157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2627 vdd a_3031_n5964# a_2823_n5964# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2628 a_8878_n4069# a_9135_n4085# a_7940_n4313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2629 vdd a_29319_n8478# a_29111_n8478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2630 a_27987_n9110# a_28172_n9825# a_28123_n9809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2631 gnd d0 a_34293_n9545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2632 a_36754_n5935# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2633 a_646_n6171# a_433_n6171# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2634 a_20620_n5603# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2635 a_31070_n7260# a_30649_n7260# a_30335_n6807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2636 a_28020_n5782# a_28063_n8198# a_28018_n7994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2637 a_12915_3754# a_13902_3320# a_13853_3510# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2638 gnd d0 a_19165_n7953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2639 a_8880_n8293# a_8876_n8481# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2640 vdd d1 a_18225_9120# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2641 a_5174_4844# a_5703_4963# a_5911_4963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2642 gnd a_9136_n4639# a_8928_n4639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2643 a_24011_n4924# a_24007_n5112# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2644 a_21041_n6706# a_20620_n6706# a_20304_n6386# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2645 a_10888_1618# a_10467_1618# a_10151_1728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2646 a_18910_3002# a_19167_2812# a_17975_2515# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2647 a_21040_5452# a_20619_5452# a_20304_5657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2648 a_16892_n3565# a_16783_n3742# a_16890_n5777# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2649 a_12916_n2071# a_13173_n2087# a_12775_n2663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2650 a_23074_n4065# a_23327_n4269# a_22929_n4845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2651 a_17972_n2112# a_18959_n1884# a_18914_n1680# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2652 a_7802_6411# a_7987_6909# a_7938_7099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2653 vdd d0 a_9133_6665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2654 a_6750_n8149# a_6537_n8149# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2655 a_21041_2143# a_20620_2143# a_20306_1891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2656 a_25887_n7296# a_25674_n7296# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2657 vdd a_8195_n7638# a_7987_n7638# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2658 a_15941_4414# a_16672_4724# a_16880_4724# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2659 vdd d3 a_23215_n8157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2660 a_39094_5738# a_39099_5012# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2661 a_20306_n1974# a_20306_n1744# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2662 a_6640_8028# a_6427_8028# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2663 vdd d0 a_29321_n2963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2664 a_39093_9601# a_39350_9411# a_38158_9114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2665 a_38017_2162# a_38274_1972# a_38047_3252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2666 a_32022_2982# a_31913_2982# a_32020_5194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2667 gnd a_33216_6343# a_33008_6343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2668 a_28129_4697# a_29113_4994# a_29068_5007# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2669 a_119_n4615# a_646_n5068# a_854_n5068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2670 a_2747_4164# a_3000_4151# a_2778_3048# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2671 vdd a_33215_n9278# a_33007_n9278# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2672 a_26615_n3194# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2673 a_23072_n8477# a_24056_n8991# a_24011_n8787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2674 a_38049_7487# a_38063_8590# a_38014_8780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2675 a_30337_n2395# a_30864_n2848# a_31072_n2848# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2676 vdd a_4077_6624# a_3869_6624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2677 a_11933_n5913# a_11512_n5913# a_11839_n5913# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2678 a_2743_n4864# a_2933_n4288# a_2888_n4084# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2679 a_5175_n4656# a_5175_n4469# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2680 a_15732_6620# a_15519_6620# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2681 a_5489_n6212# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2682 a_35920_n5649# a_35707_n5649# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2683 a_27036_n4297# a_26615_n4297# a_26098_n4541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2684 a_12779_1963# a_12964_2461# a_12915_2651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2685 a_31911_n5894# a_31698_n5894# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2686 a_16460_2518# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2687 a_12913_8166# a_13900_7732# a_13855_7745# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2688 a_1373_3575# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2689 a_6866_3156# a_6752_3037# a_6859_5249# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2690 a_38161_3599# a_39145_3896# a_39096_4086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2691 a_35389_9012# a_35390_8555# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2692 vdd a_38103_n10699# a_37895_n10699# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2693 a_38051_n3587# a_38065_n4907# a_38020_n4703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2694 a_6780_n9239# a_6567_n9239# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2695 a_31072_n6711# a_30651_n6711# a_30335_n6391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2696 gnd a_14110_n5706# a_13902_n5706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2697 vdd d0 a_4079_4972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2698 a_5911_n2903# a_5490_n2903# a_5176_n2450# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2699 a_39094_n5158# a_39100_n4421# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2700 a_15519_9380# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2701 vdd a_29319_n10135# a_29111_n10135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2702 a_10149_6327# a_10676_6579# a_10884_6579# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2703 a_10676_9339# a_10463_9339# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2704 a_853_6574# a_432_6574# a_118_6322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2705 vdd d0 a_24266_3850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2706 a_26098_2738# a_25677_2738# a_25361_2619# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2707 a_17829_6593# a_18019_5811# a_17974_5824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2708 vdd a_14110_4977# a_13902_4977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2709 a_34041_n7135# a_34294_n7339# a_33099_n7567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2710 a_5912_n3457# a_5491_n3457# a_5175_n3366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2711 a_15519_n10080# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2712 a_35390_8139# a_35390_7909# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2713 gnd d1 a_28382_4684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2714 a_12916_n9604# a_13900_n10118# a_10147_n10135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2715 vdd d2 a_33217_n4866# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2716 vdd a_8056_n4921# a_7848_n4921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2717 a_7942_8025# a_8195_8012# a_7797_8794# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2718 a_26723_n8130# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2719 a_30335_5662# a_30335_5205# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2720 a_11823_n7589# a_11402_n7589# a_10884_n7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2721 a_13854_1304# a_14111_1114# a_12916_1548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2722 gnd d0 a_4078_4418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2723 a_17969_n8730# a_18956_n8502# a_18911_n8298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2724 gnd a_2830_n10672# a_2622_n10672# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2725 a_15522_n4565# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2726 a_21043_n2294# a_21773_n2050# a_21981_n2050# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2727 a_29965_345# a_29752_345# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2728 vdd d0 a_9135_2253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2729 vdd d0 a_14112_n2397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2730 a_17973_n7439# a_18226_n7643# a_17833_n6928# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2731 a_26616_n2091# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2732 gnd a_29320_n7929# a_29112_n7929# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2733 a_118_n6634# a_118_n6405# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2734 a_24012_n6581# a_24008_n6769# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2735 a_15942_n4011# a_16673_n4321# a_16881_n4321# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2736 a_17976_n1924# a_18960_n2438# a_18915_n2234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2737 gnd d0 a_14109_n5152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2738 a_7060_541# a_7879_5276# a_7834_5289# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2739 a_31801_n7570# a_31588_n7570# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2740 gnd a_18229_1399# a_18021_1399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2741 a_23073_4656# a_24057_4953# a_24012_4966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2742 a_36129_3846# a_36859_3602# a_37067_3602# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2743 a_119_n4199# a_648_n4519# a_856_n4519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2744 gnd a_29323_n2414# a_29115_n2414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2745 vdd a_4080_n1838# a_3872_n1838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2746 a_12777_6375# a_12962_6873# a_12917_6886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2747 a_13852_5716# a_13857_4990# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2748 a_39095_5189# a_39352_4999# a_38160_4702# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2749 a_17971_2692# a_18958_2258# a_18909_2448# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2750 gnd a_33218_1931# a_33010_1931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2751 gnd a_23326_4643# a_23118_4643# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2752 gnd d1 a_18226_n8746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2753 gnd a_33358_n4274# a_33150_n4274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2754 a_34043_n3826# a_34039_n4014# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2755 vdd a_4079_2212# a_3871_2212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2756 a_36126_6601# a_36857_6911# a_37065_6911# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2757 gnd a_38412_7998# a_38204_7998# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2758 a_20832_n7809# a_20619_n7809# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2759 a_25889_4944# a_25676_4944# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2760 a_15734_2208# a_15521_2208# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2761 a_21980_3556# a_21559_3556# a_21042_3800# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2762 a_3823_8843# a_4076_8830# a_2881_9264# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2763 vdd d0 a_19165_8327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2764 a_30865_n1745# a_30652_n1745# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2765 a_26098_n4541# a_25677_n4541# a_25361_n4450# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2766 a_11757_n4791# a_11544_n4791# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2767 a_10888_n2318# a_10467_n2318# a_10151_n2227# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2768 a_21978_n8668# a_21910_n9179# a_21994_n8089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2769 a_12915_3754# a_13902_3320# a_13857_3333# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2770 a_4632_480# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2771 a_5489_n7869# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2772 a_29067_n4965# a_29063_n5153# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2773 gnd d2 a_33215_8549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2774 a_1793_n5378# a_1372_n5378# a_855_n5622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2775 a_30866_n2299# a_30653_n2299# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2776 gnd d1 a_13169_n9808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2777 a_35389_n9970# a_35389_n9741# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2778 a_13854_n9360# a_14107_n9564# a_12912_n9792# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2779 a_10677_8236# a_10464_8236# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2780 a_854_5471# a_433_5471# a_118_5676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2781 gnd d3 a_13062_n3769# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2782 a_37081_5354# a_36967_5235# a_37175_5235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2783 a_26099_1635# a_25678_1635# a_25362_1745# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2784 gnd d0 a_34294_9370# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2785 a_5488_6615# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2786 a_10151_1915# a_10678_2167# a_10886_2167# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2787 a_35392_n4642# a_35919_n5095# a_36127_n5095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2788 a_35392_2853# a_35921_2743# a_36129_2743# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2789 a_855_2162# a_434_2162# a_120_1910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2790 a_6958_n5949# a_6537_n5949# a_6864_n5949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2791 gnd a_18225_9120# a_18017_9120# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2792 a_35706_8258# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2793 a_35391_5933# a_35391_5703# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2794 a_20303_n8592# a_20303_n8362# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2795 gnd d0 a_14109_8286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2796 a_5701_n7315# a_5488_n7315# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2797 vdd a_33216_6343# a_33008_6343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2798 a_30334_n7910# a_30334_n7723# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2799 a_2743_4341# a_3000_4151# a_2778_3048# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2800 gnd a_9133_6665# a_8925_6665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2801 a_21040_n8912# a_21770_n8668# a_21978_n8668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2802 a_17828_n9322# a_18018_n8746# a_17973_n8542# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2803 a_26613_n8709# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2804 a_35391_n5745# a_35391_n5558# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2805 a_34039_5148# a_34296_4958# a_33104_4661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2806 a_11839_7532# a_11542_8503# a_11823_7992# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2807 a_38014_8780# a_38204_7998# a_38159_8011# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2808 a_17863_n8018# a_18116_n8222# a_17865_n5806# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2809 a_10463_n7279# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2810 vdd a_13062_n5969# a_12854_n5969# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2811 a_25361_4138# a_25888_4390# a_26096_4390# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2812 vdd a_4077_n8456# a_3869_n8456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2813 a_22931_n9069# a_23116_n9784# a_23067_n9768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2814 a_27036_2494# a_26969_1902# a_27047_3018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2815 a_29067_n6068# a_29320_n6272# a_28125_n6500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2816 a_12779_1963# a_12964_2461# a_12919_2474# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2817 a_30337_n2208# a_30337_n1979# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2818 a_22960_n5929# a_23009_n3745# a_22960_n3729# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2819 a_15204_n7783# a_15204_n7554# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2820 a_6537_n8149# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2821 vdd a_13170_n7602# a_12962_n7602# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2822 a_1682_500# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2823 gnd d0 a_24262_8811# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2824 a_26936_7430# a_26723_7430# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2825 a_11618_n2074# a_11405_n2074# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2826 a_31587_9076# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2827 a_28124_8183# a_29111_7749# a_29066_7762# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2828 a_10885_4373# a_10464_4373# a_10149_4578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2829 a_10884_n8382# a_10463_n8382# a_10148_n7929# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2830 a_20305_3681# a_20305_3451# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2831 vdd a_39349_n9586# a_39141_n9586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2832 a_8882_6129# a_9135_6116# a_7943_5819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2833 a_17973_n7439# a_18957_n7953# a_18908_n7937# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2834 a_117_n7737# a_646_n7828# a_854_n7828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2835 a_6427_6925# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2836 a_15943_3865# a_15522_3865# a_15206_3746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2837 a_30862_n8363# a_30649_n8363# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2838 a_5174_n6216# a_5702_n6212# a_5910_n6212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2839 a_29064_3527# a_29069_2801# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2840 a_119_3929# a_119_3700# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2841 gnd a_4936_n10733# a_4728_n10733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2842 a_5172_n10171# a_8876_n10138# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2843 a_37076_7435# a_36967_7435# a_37081_5354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2844 gnd d2 a_33217_4137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2845 vdd d2 a_8055_n7127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2846 a_10150_n3517# a_10678_n3970# a_10886_n3970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2847 a_116_9444# a_645_9334# a_853_9334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2848 a_35392_n3996# a_35920_n3992# a_36128_n3992# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2849 a_34043_6074# a_34039_6251# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2850 vdd d1 a_28382_4684# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2851 a_7938_8202# a_8195_8012# a_7797_8794# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2852 a_9875_n10838# a_20790_n10911# a_19441_n829# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2853 a_15734_n6771# a_15521_n6771# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2854 a_20303_8322# a_20832_8212# a_21040_8212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2855 a_15941_7174# a_15520_7174# a_15204_7284# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2856 a_33104_n5173# a_33357_n5377# a_32964_n4662# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2857 a_37076_n7958# a_36785_n7019# a_37066_n6508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2858 a_35392_n4226# a_35921_n4546# a_36129_n4546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2859 vdd a_28383_n4310# a_28175_n4310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2860 a_20304_n6802# a_20831_n7255# a_21039_n7255# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2861 a_117_6779# a_118_6322# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2862 a_32022_2982# a_31731_1866# a_32011_2458# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2863 a_34043_2211# a_34296_2198# a_33101_2632# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2864 a_30337_1250# a_30865_1045# a_31073_1045# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2865 a_30651_n2848# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2866 a_1587_1369# a_1374_1369# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2867 gnd d1 a_33357_n6480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2868 a_20305_2578# a_20834_2697# a_21042_2697# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2869 a_7942_8025# a_8926_8322# a_8877_8512# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2870 gnd d0 a_14111_3874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2871 gnd d6 a_25122_n10714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2872 a_39099_n3867# a_39095_n4055# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2873 a_10679_n3421# a_10466_n3421# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2874 vdd a_23326_4643# a_23118_4643# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2875 a_6866_3156# a_6569_4127# a_6849_4719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2876 a_4954_480# a_6738_541# a_7060_541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2877 gnd a_9135_2253# a_8927_2253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2878 a_11824_4683# a_11403_4683# a_10885_4373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2879 vdd d1 a_28381_n7619# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2880 a_33102_n9585# a_34086_n10099# a_30333_n10116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2881 a_38051_3075# a_38065_4178# a_38020_4191# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2882 a_23070_n4253# a_24057_n4025# a_24008_n4009# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2883 a_32958_8739# a_33148_7957# a_33103_7970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2884 vdd d2 a_13031_n4885# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2885 a_26615_3597# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2886 a_20620_6006# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2887 a_1370_n9790# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2888 a_6850_n4316# a_6782_n4827# a_6866_n3737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2889 gnd d3 a_8087_n3805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2890 a_31588_7973# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2891 vdd a_39351_n9037# a_39143_n9037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2892 vdd a_4077_n10113# a_3869_n10113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2893 a_25888_n6193# a_25675_n6193# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2894 a_1795_1369# a_1727_1880# a_1805_2996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2895 a_27034_6906# a_26613_6906# a_26095_6596# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2896 a_28126_3771# a_29113_3337# a_29068_3350# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2897 a_23071_n9580# a_24055_n10094# a_24006_n10078# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2898 a_33106_n1864# a_34090_n2378# a_34041_n2362# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2899 a_6428_5822# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2900 a_10148_7887# a_10148_7430# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2901 vdd a_13060_n8181# a_12852_n8181# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2902 a_31071_n6157# a_31802_n6467# a_32010_n6467# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2903 vdd a_24264_n6231# a_24056_n6231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2904 a_6429_2513# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2905 a_36129_n3443# a_36859_n3199# a_37067_n3199# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2906 a_36645_n6508# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2907 vdd d0 a_34294_9370# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2908 a_16460_n3218# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2909 a_117_8112# a_646_8231# a_854_8231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2910 a_34040_1285# a_30339_1151# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2911 a_34044_3868# a_34040_4045# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2912 vdd a_18225_9120# a_18017_9120# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2913 a_37078_3023# a_36969_3023# a_37076_5235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2914 a_116_n9484# a_117_n9027# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2915 a_12920_n1883# a_13904_n2397# a_13859_n2193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2916 gnd d1 a_3140_4662# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2917 gnd d1 a_23327_2437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2918 a_36126_9361# a_35705_9361# a_35389_9242# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2919 vdd d0 a_14109_8286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2920 a_12914_n5380# a_13901_n5152# a_13852_n5136# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2921 a_6428_n5419# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2922 a_15204_8574# a_15731_8826# a_15939_8826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2923 vdd a_9133_6665# a_8925_6665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2924 a_8884_1717# a_8880_1894# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2925 a_20304_n6386# a_20833_n6706# a_21041_n6706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2926 vdd d0 a_9135_n5742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2927 a_31073_n3402# a_31803_n3158# a_32011_n3158# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2928 a_30333_9430# a_30333_9201# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2929 a_36856_n9817# a_36643_n9817# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2930 a_26097_3287# a_26828_3597# a_27036_3597# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2931 a_30335_n5288# a_30335_n5058# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2932 a_10151_n2227# a_10151_n1998# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2933 a_36126_n8404# a_35705_n8404# a_35390_n8408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2934 a_27987_8598# a_28172_9096# a_28127_9109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2935 a_34041_6623# a_34037_6800# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2936 a_6849_n6522# a_6428_n6522# a_5910_n6212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2937 a_3825_4431# a_3821_4608# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2938 a_35392_n3123# a_35392_n2893# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2939 a_7944_3613# a_8928_3910# a_8879_4100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2940 gnd d0 a_4079_n5701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2941 a_10676_7682# a_10463_7682# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2942 a_27050_7549# a_26753_8520# a_27034_8009# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2943 gnd d1 a_28380_n9825# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2944 gnd d0 a_9135_n4085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2945 a_30336_3915# a_30336_3686# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2946 a_31801_6870# a_31588_6870# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2947 a_27990_1980# a_28175_2478# a_28130_2491# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2948 a_21697_n9179# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2949 a_15520_n7874# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2950 a_8878_6306# a_9135_6116# a_7943_5819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2951 gnd d0 a_39353_n1865# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2952 vdd d0 a_24266_n1819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2953 a_20304_n5699# a_20304_n5512# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2954 a_3825_8294# a_3821_8471# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2955 a_22759_n10637# a_23016_n10653# a_22858_n10637# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2956 a_8884_n2229# a_8880_n2417# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2957 a_5174_5260# a_5174_5073# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2958 a_12776_n9093# a_12961_n9808# a_12912_n9792# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2959 gnd d1 a_18226_6914# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2960 a_5909_7718# a_6640_8028# a_6848_8028# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2961 a_15941_n8977# a_15520_n8977# a_15204_n8886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2962 a_27035_5803# a_26614_5803# a_26097_6047# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2963 a_12805_n5953# a_12854_n3769# a_12805_n3753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2964 a_21698_6273# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2965 a_28128_n8518# a_29112_n9032# a_29067_n8828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2966 gnd d1 a_13173_n2087# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2967 gnd d0 a_9134_4459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2968 vdd d2 a_13029_8568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2969 a_35706_n5095# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2970 gnd d0 a_14108_7732# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2971 vdd a_19163_n9605# a_18955_n9605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2972 a_10463_9339# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2973 a_21880_7389# a_21667_7389# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2974 a_13858_n3296# a_13854_n3484# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2975 a_35922_1640# a_35709_1640# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2976 vdd a_24266_3850# a_24058_3850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2977 vdd a_34295_n6236# a_34087_n6236# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2978 a_5176_n2450# a_5703_n2903# a_5911_n2903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2979 a_21557_n8668# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2980 a_852_n9480# a_431_n9480# a_116_n9484# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2981 a_16895_n8154# a_16598_n9244# a_16878_n9836# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2982 vdd d0 a_9136_2807# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2983 a_7942_8025# a_8926_8322# a_8881_8335# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2984 a_16897_n3742# a_16783_n3742# a_16890_n5777# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2985 gnd a_4078_4418# a_3870_4418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2986 a_15206_4162# a_15733_4414# a_15941_4414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2987 a_20835_1594# a_20622_1594# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2988 vdd a_9135_2253# a_8927_2253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2989 a_10149_5911# a_10149_5681# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X2990 a_8884_n2229# a_9137_n2433# a_7945_n1919# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2991 a_35390_7909# a_35918_7704# a_36126_7704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2992 a_6958_n5949# a_7886_n10713# a_4679_n10717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2993 a_11401_n9795# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2994 a_8879_8884# a_9132_8871# a_7937_9305# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2995 vdd a_38271_8590# a_38063_8590# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2996 a_30650_n8917# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2997 a_12918_n5192# a_13171_n5396# a_12778_n4681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X2998 a_7798_6588# a_8055_6398# a_7828_7678# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2999 a_12914_5960# a_13901_5526# a_13852_5716# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3000 gnd a_24265_n5682# a_24057_n5682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3001 a_24012_n2718# a_24265_n2922# a_23070_n3150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3002 a_39097_n7176# a_39350_n7380# a_38155_n7608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3003 a_28123_n9809# a_28380_n9825# a_27987_n9110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3004 a_5173_7050# a_5702_7169# a_5910_7169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3005 a_10678_3270# a_10465_3270# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3006 a_34041_n8238# a_34037_n8426# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3007 a_11933_n5913# a_11512_n5913# a_11834_n5736# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3008 a_31803_2458# a_31590_2458# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3009 a_23069_5936# a_24056_5502# a_24011_5515# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3010 a_5489_n6212# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3011 gnd d0 a_4080_2766# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3012 a_25676_4944# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3013 a_21040_4349# a_20619_4349# a_20305_4097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3014 a_15521_2208# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3015 a_21772_n3153# a_21559_n3153# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3016 gnd d0 a_39350_n8483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3017 a_7828_n8201# a_7847_n7127# a_7802_n6923# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3018 a_10465_n3970# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3019 a_5175_3054# a_5175_2867# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3020 vdd a_19165_8327# a_18957_8327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3021 a_18914_n1680# a_18910_n1868# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3022 a_16672_n5424# a_16459_n5424# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3023 a_35707_n3992# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3024 gnd a_38411_n9830# a_38203_n9830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3025 a_3822_n2925# a_3828_n2188# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3026 a_6850_2513# a_6429_2513# a_5912_2757# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3027 vdd a_9136_n1879# a_8928_n1879# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3028 gnd d0 a_24267_1644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3029 a_28128_n7415# a_28381_n7619# a_27988_n6904# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3030 gnd a_14111_2771# a_13903_2771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3031 a_29065_n9377# a_29061_n9565# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3032 a_2884_n3169# a_3871_n2941# a_3826_n2737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3033 gnd a_33215_8549# a_33007_8549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3034 gnd a_38414_n4315# a_38206_n4315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3035 a_27037_1391# a_26616_1391# a_26099_1635# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3036 a_15734_6071# a_15521_6071# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3037 a_13856_5539# a_13852_5716# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3038 a_35708_n4546# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3039 vdd d1 a_3140_4662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3040 a_20618_n7255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3041 a_32012_n2055# a_31591_n2055# a_31074_n2299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3042 a_857_1613# a_1587_1369# a_1795_1369# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3043 a_10150_2602# a_10679_2721# a_10887_2721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3044 a_10464_8236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3045 a_23074_2450# a_24058_2747# a_24009_2937# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3046 a_5909_9375# a_5488_9375# a_5172_9485# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3047 gnd a_34294_9370# a_34086_9370# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3048 vdd a_13171_4667# a_12963_4667# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3049 a_12778_4169# a_12963_4667# a_12914_4857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3050 vdd d1 a_3139_n7597# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3051 a_21039_n8358# a_20618_n8358# a_20303_n8362# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3052 a_5173_n9068# a_5700_n9521# a_5908_n9521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3053 a_5912_n3457# a_5491_n3457# a_5175_n3137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3054 a_12809_n3565# a_12823_n4885# a_12778_n4681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3055 a_28014_n8182# a_28033_n7108# a_27988_n6904# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3056 vdd d0 a_4080_1109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3057 vdd a_34295_n7893# a_34087_n7893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3058 a_33100_n5361# a_34087_n5133# a_34038_n5117# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3059 a_15943_n4565# a_16673_n4321# a_16881_n4321# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3060 a_8881_n8847# a_9134_n9051# a_7942_n8537# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3061 a_13858_2784# a_13854_2961# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3062 a_7800_n2699# a_8057_n2715# a_7830_n3789# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3063 gnd d0 a_19166_6121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3064 a_432_n7274# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3065 a_11616_n5383# a_11403_n5383# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3066 a_6569_n4827# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3067 vdd a_28381_6890# a_28173_6890# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3068 a_39099_n6627# a_39352_n6831# a_38160_n6317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3069 a_12916_1548# a_13903_1114# a_13854_1304# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3070 a_5174_n6446# a_5174_n6216# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3071 a_24009_n9336# a_24262_n9540# a_23067_n9768# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3072 vdd d2 a_23185_n7067# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3073 a_26095_n8399# a_26826_n8709# a_27034_n8709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3074 a_24014_1657# a_24010_1834# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3075 a_3825_n8806# a_4078_n9010# a_2886_n8496# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3076 vdd a_4081_n2392# a_3873_n2392# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3077 a_34038_5697# a_34295_5507# a_33100_5941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3078 a_25677_3841# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3079 a_31589_n6467# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3080 a_21041_3246# a_20620_3246# a_20305_3451# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3081 gnd a_24262_8811# a_24054_8811# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3082 a_26723_7430# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3083 a_18907_7963# a_18912_7237# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3084 a_23071_1524# a_24058_1090# a_24013_1103# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3085 a_25359_8363# a_25888_8253# a_26096_8253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3086 a_6864_5368# a_6537_7449# a_6859_7449# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3087 a_15942_2208# a_16673_2518# a_16881_2518# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3088 vdd d0 a_14108_7732# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3089 a_26098_n4541# a_25677_n4541# a_25361_n4221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3090 a_18914_n1680# a_19167_n1884# a_17972_n2112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3091 a_26825_9112# a_26612_9112# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3092 a_31070_n7260# a_30649_n7260# a_30334_n7264# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3093 a_36128_6052# a_36858_5808# a_37066_5808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3094 a_7944_3613# a_8197_3600# a_7799_4382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3095 vdd a_35153_n10719# a_34945_n10719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3096 vdd a_9133_n8497# a_8925_n8497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3097 a_39094_7395# a_39351_7205# a_38159_6908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3098 a_24011_4412# a_24007_4589# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3099 gnd a_23326_n6475# a_23118_n6475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3100 gnd a_33217_4137# a_33009_4137# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3101 a_7943_n5228# a_8927_n5742# a_8882_n5538# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3102 a_36967_n8135# a_36754_n8135# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3103 a_2748_1958# a_3001_1945# a_2774_3225# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3104 a_30337_n2395# a_30337_n2208# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3105 a_38045_7664# a_38064_6384# a_38015_6574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3106 gnd d1 a_33355_9060# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3107 a_36125_8807# a_36856_9117# a_37064_9117# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3108 a_1803_n7931# a_1512_n6992# a_1792_n7584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3109 a_647_n2862# a_434_n2862# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3110 a_15206_n4661# a_15206_n4474# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3111 a_34044_2765# a_34297_2752# a_33105_2455# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3112 a_22088_5189# a_22081_481# a_22289_481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3113 a_16814_1926# a_16601_1926# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3114 gnd d1 a_13170_7976# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3115 gnd d0 a_24264_n7888# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3116 a_17975_2515# a_18959_2812# a_18914_2825# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3117 a_2888_n4084# a_3141_n4288# a_2743_n4864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3118 a_12914_5960# a_13901_5526# a_13856_5539# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3119 a_7940_n4313# a_8927_n4085# a_8878_n4069# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3120 a_1374_1369# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3121 a_21039_9315# a_21769_9071# a_21977_9071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3122 vdd d3 a_28271_7469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3123 a_119_n3969# a_119_n3512# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3124 a_5701_n7315# a_5488_n7315# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3125 gnd a_18227_n5437# a_18019_n5437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3126 a_29068_3350# a_29064_3527# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3127 vdd d3 a_3029_n8176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3128 a_39097_n8279# a_39093_n8467# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3129 a_28125_5977# a_29112_5543# a_29063_5733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3130 a_434_n6725# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3131 a_7797_n9317# a_8054_n9333# a_7832_n8013# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3132 vdd d0 a_4080_2766# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3133 a_853_7677# a_432_7677# a_117_7882# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3134 a_12776_8581# a_13029_8568# a_12807_7465# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3135 a_25360_n6843# a_25887_n7296# a_26095_n7296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3136 a_35920_n5649# a_35707_n5649# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3137 a_24009_n1803# a_24985_n1506# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3138 a_11825_2477# a_11758_1885# a_11836_3001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3139 a_38015_n7097# a_38272_n7113# a_38045_n8187# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3140 a_12775_n2663# a_12965_n2087# a_12916_n2071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3141 a_854_4368# a_433_4368# a_119_4116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3142 a_35391_5059# a_35920_4949# a_36128_4949# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3143 vdd d0 a_24267_1644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3144 a_6847_n9831# a_6426_n9831# a_5909_n10075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3145 a_5176_n2034# a_5176_n1804# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3146 vdd a_14111_2771# a_13903_2771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3147 gnd d1 a_28383_2478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3148 a_3821_n6234# a_4078_n6250# a_2883_n6478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3149 a_28126_n4294# a_29113_n4066# a_29064_n4050# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3150 a_1795_n2069# a_1727_n2580# a_1805_n3519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3151 a_7802_n6923# a_8055_n7127# a_7828_n8201# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3152 a_27045_n7953# a_26936_n8130# a_27050_n5930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3153 a_855_n2862# a_1586_n3172# a_1794_n3172# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3154 a_18911_n8298# a_19164_n8502# a_17969_n8730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3155 a_25239_461# a_24818_461# a_22289_481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3156 vdd a_34294_9370# a_34086_9370# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3157 a_10884_n10039# a_11614_n9795# a_11822_n9795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3158 a_39096_1326# a_35395_1192# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3159 a_15206_2872# a_15206_2643# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3160 a_32008_n9776# a_31941_n9184# a_32025_n8094# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3161 a_13857_n5502# a_13853_n5690# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3162 gnd a_14108_n7358# a_13900_n7358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3163 gnd a_23327_2437# a_23119_2437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3164 vdd d0 a_14111_n1843# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3165 a_30074_345# a_29965_345# a_19317_288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3166 vdd d0 a_34294_n10099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3167 a_38047_3252# a_38066_1972# a_38017_2162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3168 a_27989_4186# a_28174_4684# a_28125_4874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3169 a_32959_6533# a_33149_5751# a_33100_5941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3170 a_10884_6579# a_10463_6579# a_10148_6784# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3171 vdd a_18116_n8222# a_17908_n8222# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3172 a_35392_n4455# a_35921_n4546# a_36129_n4546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3173 a_18914_n3337# a_18910_n3525# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3174 a_11405_n2074# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3175 a_32009_7973# a_31941_8484# a_32025_7513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3176 a_36129_n1786# a_35708_n1786# a_35016_n1511# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3177 a_15203_9031# a_15204_8574# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3178 a_5703_4963# a_5490_4963# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3179 a_30333_n9700# a_30333_n9470# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3180 a_21981_1350# a_21560_1350# a_21043_1594# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3181 a_20303_n7259# a_20831_n7255# a_21039_n7255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3182 vdd a_30219_n10835# a_30011_n10835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3183 a_7797_8794# a_7987_8012# a_7938_8202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3184 vdd d0 a_19166_6121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3185 a_31801_n7570# a_31588_n7570# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3186 a_12916_1548# a_13903_1114# a_13858_1127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3187 vdd d3 a_28273_3057# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3188 a_30333_n10116# a_30333_n9929# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3189 a_6430_n2110# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3190 gnd a_9134_n7948# a_8926_n7948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3191 a_35390_n7535# a_35390_n7305# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3192 a_10679_n3421# a_10466_n3421# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3193 a_34044_1108# a_34040_1285# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3194 a_10463_7682# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3195 a_8880_n7190# a_8876_n7378# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3196 a_8884_1717# a_9137_1704# a_7945_1407# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3197 a_28127_1565# a_29114_1131# a_29065_1321# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3198 a_23072_n7374# a_23325_n7578# a_22932_n6863# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3199 gnd d0 a_4077_n7353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3200 a_15940_9380# a_15519_9380# a_15203_9490# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3201 a_11834_n7936# a_11543_n6997# a_11824_n6486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3202 a_25360_n6427# a_25889_n6747# a_26097_n6747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3203 a_10678_6030# a_10465_6030# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3204 a_18910_3002# a_18913_2271# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3205 a_855_3265# a_434_3265# a_119_3470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3206 a_35392_3727# a_35921_3846# a_36129_3846# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3207 a_15204_8158# a_15204_7928# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3208 a_20832_n7809# a_20619_n7809# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3209 gnd d0 a_34295_7164# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3210 gnd a_3141_n3185# a_2933_n3185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3211 a_27045_5230# a_26725_3018# a_27047_3018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3212 a_5489_4409# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3213 a_8882_n6641# a_8878_n6829# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3214 a_2888_n4084# a_3872_n4598# a_3823_n4582# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3215 gnd a_18226_6914# a_18018_6914# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3216 a_39094_4635# a_39100_3909# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3217 gnd d1 a_23325_n8681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3218 a_24865_n10698# a_27864_n10694# a_27144_n5930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3219 a_6849_n5419# a_6782_n4827# a_6866_n3737# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3220 gnd a_3139_7971# a_2931_7971# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3221 vdd a_14109_n9015# a_13901_n9015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3222 a_22289_481# a_21868_481# a_22088_5189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3223 a_2881_9264# a_3868_8830# a_3819_9020# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3224 gnd a_9134_4459# a_8926_4459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3225 a_29062_9596# a_29065_8865# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3226 a_11823_6889# a_11402_6889# a_10884_6579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3227 a_38045_7664# a_38064_6384# a_38019_6397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3228 a_1792_n8687# a_1724_n9198# a_1808_n8108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3229 vdd d3 a_18118_n3810# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3230 a_16769_546# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3231 a_30337_1250# a_30339_1151# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3232 a_2746_n6882# a_2931_n7597# a_2886_n7393# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3233 vdd d1 a_33355_9060# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3234 a_5487_n9521# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3235 a_31072_n6711# a_31802_n6467# a_32010_n6467# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3236 gnd a_14108_7732# a_13900_7732# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3237 a_32020_n5717# a_31700_n3682# a_32022_n3505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3238 a_5175_n3553# a_5175_n3366# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3239 a_34040_2942# a_34297_2752# a_33105_2455# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3240 a_1584_n8687# a_1371_n8687# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3241 a_33102_9073# a_34086_9370# a_34037_9560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3242 a_11825_n4280# a_11757_n4791# a_11841_n3701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3243 vdd a_9136_2807# a_8928_2807# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3244 a_31071_4354# a_31802_4664# a_32010_4664# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3245 a_10148_7430# a_10676_7682# a_10884_7682# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3246 a_16600_n4832# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3247 a_12134_505# a_14876_485# a_9888_364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3248 a_31069_8766# a_30648_8766# a_30334_8514# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3249 a_17861_n5994# a_17910_n3810# a_17861_n3794# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3250 a_646_n8931# a_433_n8931# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3251 a_20622_1594# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3252 a_28125_5977# a_29112_5543# a_29067_5556# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3253 a_31070_n10020# a_30649_n10020# a_30333_n9700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3254 a_20304_n6615# a_20833_n6706# a_21041_n6706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3255 a_36856_n9817# a_36643_n9817# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3256 a_11404_n3177# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3257 a_10886_2167# a_10465_2167# a_10150_2372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3258 a_36126_n8404# a_35705_n8404# a_35390_n7951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3259 a_21039_n8358# a_21770_n8668# a_21978_n8668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3260 a_29065_n1844# a_30041_n1547# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3261 a_26613_n8709# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3262 a_21667_7389# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3263 a_6428_4719# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3264 gnd d0 a_29323_1685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3265 a_15944_1659# a_15523_1659# a_15207_1540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3266 a_7804_n2511# a_7989_n3226# a_7944_n3022# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3267 a_10465_3270# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3268 a_117_7238# a_646_7128# a_854_7128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3269 a_21041_4903# a_20620_4903# a_20304_4784# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3270 a_38014_n9303# a_38204_n8727# a_38155_n8711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3271 a_2884_n3169# a_3141_n3185# a_2748_n2470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3272 a_31590_2458# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3273 gnd d2 a_13030_6362# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3274 a_15520_n7874# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3275 a_15942_4968# a_15521_4968# a_15205_5078# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3276 a_30335_4559# a_30336_4102# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3277 vdd d0 a_14110_n5706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3278 a_20304_6116# a_20833_6006# a_21041_6006# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3279 a_15206_2643# a_15735_2762# a_15943_2762# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3280 a_28020_n5782# a_28273_n5986# a_27815_n10678# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3281 a_22962_n7953# a_23215_n8157# a_22964_n5741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3282 a_28130_2491# a_29114_2788# a_29065_2978# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3283 a_118_n5531# a_118_n5302# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3284 a_117_n7508# a_646_n7828# a_854_n7828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3285 gnd a_24267_1644# a_24059_1644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3286 a_36128_n5649# a_35707_n5649# a_35391_n5329# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3287 a_29068_n2759# a_29321_n2963# a_28126_n3191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3288 a_15941_n8977# a_15520_n8977# a_15204_n8657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3289 a_33102_n2052# a_33359_n2068# a_32961_n2644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3290 gnd a_33356_n7583# a_33148_n7583# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3291 a_32119_n5894# a_31698_n5894# a_32025_n5894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3292 a_11544_n4791# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3293 a_7943_5819# a_8927_6116# a_8878_6306# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3294 gnd d0 a_4079_3315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3295 a_37065_8014# a_36644_8014# a_36126_7704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3296 a_15521_6071# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3297 gnd a_8195_n8741# a_7987_n8741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3298 a_27990_n2492# a_28175_n3207# a_28130_n3003# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3299 a_11825_2477# a_11404_2477# a_10886_2167# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3300 a_27989_4186# a_28174_4684# a_28129_4697# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3301 a_23071_9068# a_23324_9055# a_22931_8557# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3302 a_32959_6533# a_33149_5751# a_33104_5764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3303 gnd a_14110_3320# a_13902_3320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3304 a_3826_3328# a_3822_3505# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3305 a_15203_n10176# a_19164_n10159# a_17972_n9645# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3306 a_2778_n5760# a_2821_n8176# a_2776_n7972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3307 a_30863_n5054# a_30650_n5054# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3308 a_10886_n5627# a_10465_n5627# a_10149_n5536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3309 a_5175_n2907# a_5703_n2903# a_5911_n2903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3310 a_7797_8794# a_7987_8012# a_7942_8025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3311 vdd a_13030_n7091# a_12822_n7091# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3312 a_16895_n8154# a_16598_n9244# a_16879_n8733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3313 a_21770_7968# a_21557_7968# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3314 a_20620_n3946# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3315 a_34041_7726# a_34294_7713# a_33099_8147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3316 a_21697_8479# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3317 a_39094_5738# a_39351_5548# a_38156_5982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3318 vdd d1 a_23327_n3166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3319 a_25674_n7296# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3320 a_13851_n10102# a_14108_n10118# a_12916_n9604# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3321 a_28127_1565# a_29114_1131# a_29069_1144# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3322 a_6429_3616# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3323 a_856_n4519# a_435_n4519# a_119_n4199# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3324 gnd a_19166_6121# a_18958_6121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3325 a_39093_n10124# a_39350_n10140# a_38158_n9626# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3326 a_30650_n8917# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3327 gnd d1 a_18228_2502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3328 a_7803_n4717# a_7988_n5432# a_7939_n5416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3329 a_18911_n2422# a_19168_n2438# a_17976_n1924# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3330 vdd d0 a_34295_7164# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3331 a_118_5906# a_647_6025# a_855_6025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3332 a_1514_n2580# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3333 a_1803_n7931# a_1694_n8108# a_1808_n5908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3334 gnd d2 a_2999_n7086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3335 a_20303_n7489# a_20303_n7259# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3336 a_11926_505# a_11713_505# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3337 a_1584_6884# a_1371_6884# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3338 gnd d1 a_3141_2456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3339 a_36127_7155# a_35706_7155# a_35390_7036# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3340 a_24013_n3272# a_24266_n3476# a_23074_n2962# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3341 a_38162_n1905# a_39146_n2419# a_39101_n2215# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3342 gnd d2 a_13032_1950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3343 a_15205_6368# a_15732_6620# a_15940_6620# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3344 gnd d1 a_38411_9101# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3345 a_38156_n5402# a_39143_n5174# a_39094_n5158# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3346 a_13859_n2193# a_14112_n2397# a_12920_n1883# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3347 a_5911_2203# a_5490_2203# a_5175_2408# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3348 a_24010_9378# a_25358_9466# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3349 a_9888_364# a_14663_485# a_12134_505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3350 a_39100_2806# a_39353_2793# a_38161_2496# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3351 a_25362_n2431# a_25362_n2244# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3352 a_16672_n5424# a_16459_n5424# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3353 vdd a_14108_7732# a_13900_7732# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3354 a_26612_9112# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3355 a_29064_n6810# a_29321_n6826# a_28129_n6312# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3356 a_28126_n4294# a_29113_n4066# a_29068_n3862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3357 a_12916_n2071# a_13903_n1843# a_13858_n1639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3358 a_7797_8794# a_8054_8604# a_7832_7501# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3359 a_1805_2996# a_1514_1880# a_1794_2472# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3360 a_33099_n8670# a_33356_n8686# a_32958_n9262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3361 a_33102_9073# a_34086_9370# a_34041_9383# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3362 a_10149_6140# a_10149_5911# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3363 a_35708_n4546# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3364 a_35920_n3992# a_35707_n3992# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3365 a_11826_1374# a_11405_1374# a_10888_1618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3366 a_10677_5476# a_10464_5476# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3367 vdd d0 a_34298_n2378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3368 vdd a_9137_n2433# a_8929_n2433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3369 a_27045_7430# a_26754_6314# a_27035_5803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3370 a_20618_n7255# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3371 a_25889_n2884# a_25676_n2884# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3372 a_6537_5249# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3373 gnd d0 a_34295_n5133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3374 gnd a_33355_9060# a_33147_9060# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3375 gnd a_33246_n8162# a_33038_n8162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3376 a_2888_n2981# a_3872_n3495# a_3827_n3291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3377 a_1694_5208# a_1481_5208# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3378 a_20617_8761# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3379 a_6428_n5419# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3380 a_1374_n2069# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3381 vdd d1 a_28382_5787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3382 a_16601_1926# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3383 a_20305_2578# a_20305_2348# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3384 vdd a_24265_n2922# a_24057_n2922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3385 a_5172_9256# a_5172_9026# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3386 a_35918_9361# a_35705_9361# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3387 a_5172_n9525# a_5700_n9521# a_5908_n9521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3388 a_13854_n4587# a_13857_n3845# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3389 gnd d0 a_19167_n3541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3390 a_34044_n4380# a_34040_n4568# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3391 a_2882_n7581# a_3869_n7353# a_3820_n7337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3392 vdd d0 a_29323_1685# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3393 a_15939_8826# a_15518_8826# a_15203_9031# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3394 a_25676_n6747# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3395 a_21043_n2294# a_20622_n2294# a_20306_n1974# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3396 a_119_2826# a_119_2597# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3397 a_27036_3597# a_26615_3597# a_26098_3841# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3398 a_15733_8277# a_15520_8277# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3399 a_10147_n10135# a_10147_n9948# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3400 a_21699_4067# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3401 a_21980_n4256# a_21559_n4256# a_21042_n4500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3402 gnd a_13172_n3190# a_12964_n3190# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3403 a_39096_4086# a_39099_3355# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3404 a_34043_4971# a_34039_5148# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3405 a_38047_n5975# a_38096_n3791# a_38047_n3775# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3406 vdd d2 a_13030_6362# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3407 a_432_n7274# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3408 a_6569_n4827# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3409 a_855_4922# a_434_4922# a_118_4803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3410 a_35390_n7535# a_35919_n7855# a_36127_n7855# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3411 a_14710_n10722# a_17709_n10718# a_17660_n10702# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3412 a_10884_n8382# a_11615_n8692# a_11823_n8692# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3413 vdd a_13170_6873# a_12962_6873# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3414 a_30649_9320# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3415 a_26966_8520# a_26753_8520# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3416 vdd a_24267_1644# a_24059_1644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3417 a_11839_5332# a_11725_5213# a_11933_5213# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3418 a_1511_n9198# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3419 a_36128_6052# a_35707_6052# a_35391_6162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3420 gnd d1 a_33355_n9789# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3421 vdd d2 a_18085_n9338# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3422 a_24011_8275# a_24264_8262# a_23072_7965# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3423 a_31589_n6467# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3424 a_38161_n4111# a_39145_n4625# a_39096_n4609# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3425 a_23074_n4065# a_24058_n4579# a_24013_n4375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3426 a_7943_5819# a_8927_6116# a_8882_6129# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3427 vdd d0 a_4079_3315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3428 gnd d3 a_33248_n3750# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3429 gnd a_8087_n3805# a_7879_n3805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3430 a_23068_n7562# a_24055_n7334# a_24006_n7318# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3431 a_38015_6574# a_38205_5792# a_38156_5982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3432 gnd a_28383_3581# a_28175_3581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3433 a_8879_8884# a_8875_9061# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3434 gnd a_39349_8857# a_39141_8857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3435 a_20305_n2847# a_20306_n2390# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3436 a_23067_9245# a_23324_9055# a_22931_8557# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3437 gnd d0 a_19165_8327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3438 vdd a_14110_3320# a_13902_3320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3439 a_11614_9095# a_11401_9095# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3440 a_1694_7408# a_1481_7408# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3441 a_7799_4382# a_8056_4192# a_7834_3089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3442 a_10150_3934# a_10150_3705# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3443 a_12913_n8689# a_13900_n8461# a_13855_n8257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3444 a_21557_n8668# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3445 a_10679_1064# a_10466_1064# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3446 vdd d2 a_28243_1967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3447 a_8877_n6275# a_9134_n6291# a_7939_n6519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3448 a_34037_7903# a_34294_7713# a_33099_8147# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3449 vdd d5 a_23016_n10653# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3450 a_3825_n6046# a_3821_n6234# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3451 a_31074_n2299# a_30653_n2299# a_30337_n1979# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3452 a_647_n2862# a_434_n2862# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3453 a_23070_3730# a_24057_3296# a_24012_3309# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3454 vdd a_39352_n6831# a_39144_n6831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3455 a_37000_n2607# a_36787_n2607# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3456 a_5490_4963# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3457 vdd a_33248_n5950# a_33040_n5950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3458 a_39095_n4055# a_39352_n4071# a_38157_n4299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3459 a_25677_2738# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3460 a_31069_n9466# a_31800_n9776# a_32008_n9776# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3461 a_10148_6784# a_10149_6327# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3462 a_35391_6349# a_35391_6162# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3463 vdd a_29321_n5723# a_29113_n5723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3464 vdd a_19166_6121# a_18958_6121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3465 a_32995_5234# a_33038_7433# a_32989_7623# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3466 gnd a_13170_n8705# a_12962_n8705# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3467 a_36643_n9817# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3468 a_9779_364# a_9566_364# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3469 gnd d2 a_38272_n7113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3470 a_7943_5819# a_8196_5806# a_7798_6588# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3471 a_1726_n4786# a_1513_n4786# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3472 vdd a_28273_3057# a_28065_3057# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3473 a_12918_n5192# a_13902_n5706# a_13857_n5502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3474 a_39100_1149# a_39096_1326# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3475 a_26725_n3718# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3476 a_5702_5512# a_5489_5512# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3477 a_434_n6725# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3478 a_7937_9305# a_8924_8871# a_8875_9061# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3479 vdd d1 a_3141_2456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3480 a_11834_7413# a_11725_7413# a_11839_5332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3481 a_7828_7678# a_7847_6398# a_7802_6411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3482 a_17975_n3027# a_18228_n3231# a_17835_n2516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3483 a_13854_4064# a_13857_3333# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3484 a_10677_n6176# a_10464_n6176# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3485 gnd d2 a_2998_8563# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3486 a_10465_6030# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3487 a_30336_3915# a_30865_3805# a_31073_3805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3488 gnd a_34295_7164# a_34087_7164# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3489 a_32119_5194# a_31698_5194# a_32020_5194# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3490 a_16879_n8733# a_16458_n8733# a_15941_n8977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3491 a_21557_6865# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3492 vdd d0 a_29320_n5169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3493 a_38021_n2497# a_38206_n3212# a_38157_n3196# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3494 a_36645_4705# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3495 a_6847_n9831# a_6426_n9831# a_5908_n9521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3496 gnd d1 a_18228_n4334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3497 a_19416_288# a_19332_n829# vout gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3498 a_24013_3863# a_24266_3850# a_23074_3553# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3499 a_26096_n5090# a_25675_n5090# a_25360_n5094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3500 gnd d0 a_9133_n7394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3501 a_28124_8183# a_29111_7749# a_29062_7939# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3502 a_38017_2162# a_38207_1380# a_38158_1570# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3503 a_5489_8272# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3504 a_118_5676# a_646_5471# a_854_5471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3505 vdd a_33355_9060# a_33147_9060# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3506 a_12778_n4681# a_13031_n4885# a_12809_n3565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3507 gnd d4 a_33248_5221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3508 vdd d0 a_24264_n5128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3509 gnd d4 a_18118_n6010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3510 vdd a_2999_6357# a_2791_6357# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3511 gnd d0 a_19167_3915# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3512 a_5173_n7965# a_5173_n7778# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3513 a_30336_n4185# a_30336_n3955# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3514 a_1696_2996# a_1483_2996# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3515 a_3825_7191# a_3821_7368# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3516 a_34040_n4568# a_34297_n4584# a_33105_n4070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3517 a_12604_n10661# a_12861_n10677# a_12703_n10661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3518 a_25888_n8953# a_25675_n8953# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3519 a_39098_4458# a_39094_4635# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3520 a_10887_2721# a_10466_2721# a_10150_2831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3521 a_21042_1040# a_20621_1040# a_20306_1245# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3522 a_25678_1635# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3523 a_34039_3491# a_34296_3301# a_33101_3735# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3524 a_12913_n8689# a_13170_n8705# a_12772_n9281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3525 vdd a_24264_n8991# a_24056_n8991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3526 a_25360_6157# a_25889_6047# a_26097_6047# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3527 a_13856_n4948# a_14109_n5152# a_12914_n5380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3528 a_5176_n2263# a_5176_n2034# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3529 a_1481_n8108# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3530 a_29061_n9565# a_29318_n9581# a_28123_n9809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3531 vdd d3 a_28273_n3786# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3532 gnd a_29323_1685# a_29115_1685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3533 a_7945_1407# a_8198_1394# a_7800_2176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3534 gnd a_23016_n10653# a_22808_n10653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3535 a_5704_1100# a_5491_1100# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3536 a_24007_8452# a_24264_8262# a_23072_7965# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3537 a_38051_3075# a_38065_4178# a_38016_4368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3538 a_11836_3001# a_11727_3001# a_11834_5213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3539 a_25360_n6656# a_25889_n6747# a_26097_n6747# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3540 vdd a_38273_n4907# a_38065_n4907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3541 gnd d1 a_33356_6854# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3542 a_8882_n5538# a_9135_n5742# a_7943_n5228# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3543 a_26097_n3987# a_25676_n3987# a_25361_n3534# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3544 vdd d2 a_2999_n7086# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3545 a_24818_461# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3546 vdd a_28383_3581# a_28175_3581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3547 a_10149_4808# a_10149_4578# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3548 a_116_n9943# a_116_n9714# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3549 a_22933_n4657# a_23118_n5372# a_23069_n5356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3550 a_21559_2453# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3551 gnd d0 a_24263_6605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3552 a_32020_n7917# a_31729_n6978# a_32010_n6467# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3553 gnd d0 a_9135_n6845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3554 a_30336_n4185# a_30865_n4505# a_31073_n4505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3555 a_12916_n9604# a_13169_n9808# a_12776_n9093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3556 a_15206_3059# a_15734_3311# a_15942_3311# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3557 a_5173_8569# a_5173_8382# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3558 a_39097_7767# a_39350_7754# a_38155_8188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3559 a_15204_n8657# a_15733_n8977# a_15941_n8977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3560 a_28126_3771# a_29113_3337# a_29064_3527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3561 a_31941_n9184# a_31728_n9184# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3562 a_34041_n7135# a_34037_n7323# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3563 a_7799_4382# a_7989_3600# a_7940_3790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3564 a_5487_n9521# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3565 a_17975_n3027# a_18959_n3541# a_18910_n3525# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3566 a_29066_1875# a_29069_1144# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3567 vdd d1 a_8194_n9844# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3568 a_16890_n5777# a_16781_n5954# a_16989_n5954# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3569 a_32995_5234# a_33038_7433# a_32993_7446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3570 a_38158_n2093# a_38415_n2109# a_38017_n2685# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3571 a_33099_n8670# a_34086_n8442# a_34041_n8238# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3572 a_16600_n4832# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3573 a_10150_n3974# a_10150_n3517# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3574 a_38049_n7999# a_38063_n9319# a_38014_n9303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3575 a_13853_2407# a_14110_2217# a_12915_2651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3576 a_35706_n7855# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3577 a_646_n8931# a_433_n8931# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3578 a_26827_n5400# a_26614_n5400# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3579 a_15736_n2359# a_15523_n2359# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3580 a_13856_7196# a_14109_7183# a_12917_6886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3581 a_13856_4436# a_13852_4613# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3582 a_32010_n5364# a_31589_n5364# a_31072_n5608# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3583 a_18910_n4628# a_18913_n3886# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3584 a_31911_5194# a_31698_5194# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3585 a_21977_9071# a_21556_9071# a_21038_8761# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3586 gnd a_18228_2502# a_18020_2502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3587 vdd d2 a_2998_8563# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3588 vdd a_34295_7164# a_34087_7164# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3589 gnd a_8054_n9333# a_7846_n9333# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3590 a_5172_n10171# a_5172_n9984# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3591 a_12912_9269# a_13169_9079# a_12776_8581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3592 a_35390_n8408# a_35390_n7951# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3593 a_1371_6884# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3594 a_31070_6560# a_31801_6870# a_32009_6870# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3595 a_21041_n5603# a_20620_n5603# a_20304_n5512# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3596 a_33104_n5173# a_34088_n5687# a_34043_n5483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3597 vdd d1 a_28383_n3207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3598 vdd a_23185_n7067# a_22977_n7067# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3599 gnd a_13032_1950# a_12824_1950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3600 a_27990_1980# a_28175_2478# a_28126_2668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3601 a_6750_5249# a_6537_5249# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3602 a_11836_3001# a_11545_1885# a_11826_1374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3603 a_15941_n7874# a_16671_n7630# a_16879_n7630# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3604 a_38017_2162# a_38207_1380# a_38162_1393# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3605 a_25360_n6843# a_25360_n6656# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3606 vdd a_14110_n4049# a_13902_n4049# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3607 a_5704_2757# a_5491_2757# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3608 vdd d4 a_33248_5221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3609 a_1372_n5378# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3610 a_16568_5254# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3611 a_25361_4138# a_25361_3951# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3612 gnd d0 a_24265_2193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3613 a_10464_5476# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3614 a_5174_n5343# a_5174_n5113# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3615 vdd a_4079_n5701# a_3871_n5701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3616 a_31899_486# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3617 a_39099_3355# a_39352_3342# a_38157_3776# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3618 a_31587_n9776# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3619 a_3822_n2925# a_4079_n2941# a_2884_n3169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3620 a_32020_n7917# a_31911_n8094# a_32025_n5894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3621 a_1793_n6481# a_1372_n6481# a_854_n6171# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3622 a_22960_n3729# a_22979_n2655# a_22930_n2639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3623 gnd d2 a_13029_8568# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3624 a_1481_5208# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3625 a_32320_486# a_35062_466# a_30074_345# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3626 vdd a_18226_n8746# a_18018_n8746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3627 a_18907_6860# a_18913_6134# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3628 a_21994_7508# a_21880_7389# a_21994_5308# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3629 a_35393_1521# a_35922_1640# a_36130_1640# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3630 a_856_1059# a_435_1059# a_120_1264# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3631 a_26096_n7850# a_25675_n7850# a_25359_n7530# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3632 a_10886_n5627# a_10465_n5627# a_10149_n5307# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3633 a_18995_288# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3634 a_16989_5254# a_16982_546# a_14985_485# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3635 gnd d0 a_34296_4958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3636 gnd d0 a_4079_n4044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3637 a_35705_9361# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3638 a_13852_n8999# a_13855_n8257# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3639 a_34042_n8792# a_34038_n8980# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3640 vdd a_29323_1685# a_29115_1685# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3641 a_10885_4373# a_11616_4683# a_11824_4683# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3642 gnd d2 a_8056_n4921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3643 a_20620_n3946# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3644 a_38155_n8711# a_38412_n8727# a_38014_n9303# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3645 gnd a_23324_n9784# a_23116_n9784# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3646 a_10149_n5723# a_10677_n6176# a_10885_n6176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3647 gnd d7 a_30219_n10835# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3648 a_35391_n6202# a_35919_n6198# a_36127_n6198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3649 a_15520_n6217# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3650 a_15520_8277# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3651 a_29067_8316# a_29320_8303# a_28128_8006# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3652 vdd a_12861_n10677# a_12653_n10677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3653 a_7938_n7622# a_8195_n7638# a_7802_n6923# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3654 gnd a_23217_n3745# a_23009_n3745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3655 gnd a_38302_n8203# a_38094_n8203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3656 a_20621_n4500# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3657 a_36858_n5405# a_36645_n5405# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3658 a_10888_n2318# a_11618_n2074# a_11826_n2074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3659 gnd a_14109_5526# a_13901_5526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3660 a_25887_n10056# a_25674_n10056# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3661 a_15203_n10176# a_15203_n9989# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3662 a_15206_n3558# a_15206_n3371# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3663 a_7945_1407# a_8929_1704# a_8880_1894# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3664 a_26753_8520# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3665 a_6750_7449# a_6537_7449# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3666 a_7938_n7622# a_8925_n7394# a_8876_n7378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3667 a_30650_n5054# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3668 a_33103_6867# a_34087_7164# a_34038_7354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3669 a_15521_n2908# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3670 a_31072_6011# a_30651_6011# a_30335_5892# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3671 a_31072_2148# a_31803_2458# a_32011_2458# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3672 a_16568_7454# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3673 gnd a_39350_9411# a_39142_9411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3674 a_29068_2247# a_29064_2424# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3675 a_39093_7944# a_39350_7754# a_38155_8188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3676 a_39097_n7176# a_39093_n7364# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3677 a_5705_1654# a_5492_1654# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3678 gnd d1 a_3139_n8700# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3679 a_15522_n3462# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3680 a_26938_3018# a_26725_3018# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3681 a_11839_n8113# a_11542_n9203# a_11822_n9795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3682 a_15942_n4011# a_15521_n4011# a_15206_n3558# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3683 gnd a_19165_8327# a_18957_8327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3684 a_22964_5229# a_23217_5216# a_22190_481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3685 a_11401_9095# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3686 gnd d1 a_18227_4708# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3687 a_1481_7408# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3688 gnd a_34295_n8996# a_34087_n8996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3689 a_6849_n6522# a_6781_n7033# a_6859_n7972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3690 a_15943_n4565# a_15522_n4565# a_15206_n4474# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3691 a_16812_n7038# a_16599_n7038# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3692 a_15735_n1805# a_15522_n1805# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3693 a_31944_1866# a_31731_1866# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3694 a_10466_1064# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3695 a_28130_n4106# a_29114_n4620# a_29069_n4416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3696 vdd a_28243_1967# a_28035_1967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3697 a_17861_3271# a_17880_1991# a_17835_2004# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3698 a_1583_9090# a_1370_9090# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3699 a_24010_7721# a_24006_7898# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3700 a_3819_n9543# a_4076_n9559# a_2881_n9787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3701 a_37067_n4302# a_36999_n4813# a_37083_n3723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3702 gnd d3 a_38304_n3791# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3703 a_28124_n7603# a_29111_n7375# a_29062_n7359# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3704 a_22962_n7953# a_22976_n9273# a_22927_n9257# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3705 gnd d2 a_13031_4156# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3706 a_32959_n7056# a_33149_n6480# a_33104_n6276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3707 a_119_n3096# a_119_n2866# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3708 a_13852_7373# a_14109_7183# a_12917_6886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3709 gnd a_3001_n2674# a_2793_n2674# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3710 a_5910_4409# a_5489_4409# a_5174_4614# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3711 gnd a_24265_n4025# a_24057_n4025# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3712 a_6861_3037# a_6570_1921# a_6851_1410# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3713 gnd a_13171_4667# a_12963_4667# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3714 a_15204_n8427# a_15204_n7970# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3715 a_32889_n10642# a_32839_n10658# a_32119_n5894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3716 vdd a_19165_n5193# a_18957_n5193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3717 a_10884_7682# a_10463_7682# a_10148_7887# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3718 a_10675_n9485# a_10462_n9485# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3719 a_1586_2472# a_1373_2472# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3720 a_20303_8509# a_20303_8322# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3721 a_854_n5068# a_433_n5068# a_118_n5072# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3722 a_25676_n6747# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3723 a_10151_1269# a_10153_1170# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3724 a_11825_3580# a_11404_3580# a_10887_3824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3725 a_29069_3904# a_29322_3891# a_28130_3594# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3726 a_21980_n4256# a_21559_n4256# a_21041_n3946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3727 a_7832_7501# a_8085_7488# a_7834_5289# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3728 a_16895_n5954# a_16568_n8154# a_16890_n7977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3729 vdd a_3140_n6494# a_2932_n6494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3730 a_21880_n8089# a_21667_n8089# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3731 a_5912_n1800# a_5491_n1800# a_5176_n1804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3732 a_29062_9596# a_29319_9406# a_28127_9109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3733 a_35390_n7764# a_35919_n7855# a_36127_n7855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3734 a_11403_n5383# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3735 a_23072_6862# a_23325_6849# a_22932_6351# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3736 vdd a_38304_n5991# a_38096_n5991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3737 a_36127_n5095# a_35706_n5095# a_35392_n4642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3738 gnd a_2998_8563# a_2790_8563# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3739 gnd d4 a_38304_5262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3740 gnd a_14111_1114# a_13903_1114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3741 a_7943_n6331# a_8927_n6845# a_8878_n6829# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3742 a_30652_n4505# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3743 a_21773_n2050# a_21560_n2050# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3744 gnd d2 a_28243_n2696# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3745 a_10149_n5536# a_10149_n5307# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3746 a_6752_3037# a_6539_3037# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3747 a_36128_n5649# a_35707_n5649# a_35391_n5558# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3748 a_28125_n5397# a_28382_n5413# a_27989_n4698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3749 a_11824_n6486# a_11403_n6486# a_10886_n6730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3750 a_25361_n4221# a_25361_n3991# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3751 vdd d0 a_4078_n7907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3752 a_16881_n3218# a_16460_n3218# a_15942_n2908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3753 a_16568_n5954# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3754 a_39095_3532# a_39352_3342# a_38157_3776# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3755 gnd a_33248_5221# a_33040_5221# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3756 gnd d0 a_39352_n4071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3757 a_32993_n7958# a_33007_n9278# a_32958_n9262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3758 gnd a_19167_3915# a_18959_3915# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3759 a_12134_505# a_11713_505# a_12035_505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3760 vdd a_14967_n10738# a_14759_n10738# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3761 a_1483_2996# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3762 a_29069_3904# a_29065_4081# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3763 a_36857_8014# a_36644_8014# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3764 a_20832_n6152# a_20619_n6152# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3765 a_2886_n7393# a_3870_n7907# a_3821_n7891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3766 a_2744_n2658# a_3001_n2674# a_2774_n3748# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3767 a_21043_1594# a_20622_1594# a_20306_1704# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3768 a_36127_8258# a_35706_8258# a_35390_8368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3769 a_15732_n8423# a_15519_n8423# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3770 a_28129_n6312# a_29113_n6826# a_29064_n6810# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3771 a_13852_n6239# a_13857_n5502# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3772 a_37000_n2607# a_36787_n2607# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3773 a_25890_n3438# a_25677_n3438# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3774 gnd d1 a_38412_6895# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3775 vdd a_19167_n4644# a_18959_n4644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3776 a_26094_8802# a_25673_8802# a_25359_8550# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3777 gnd a_28382_5787# a_28174_5787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3778 gnd a_2998_n9292# a_2790_n9292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3779 a_31070_n10020# a_31800_n9776# a_32008_n9776# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3780 a_36643_n9817# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3781 a_856_n4519# a_435_n4519# a_119_n4428# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3782 vdd a_14109_5526# a_13901_5526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3783 a_15206_n4015# a_15206_n3558# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3784 a_39096_n4609# a_39353_n4625# a_38161_n4111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3785 gnd d3 a_28271_7469# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3786 a_38158_n2093# a_39145_n1865# a_39100_n1661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3787 a_33103_6867# a_34087_7164# a_34042_7177# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3788 a_16458_n7630# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3789 a_24006_n7318# a_24263_n7334# a_23068_n7562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3790 a_28016_n3770# a_28035_n2696# a_27990_n2492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3791 a_37064_9117# a_36997_8525# a_37081_7554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3792 a_13858_n1639# a_14111_n1843# a_12916_n2071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3793 a_5491_1100# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3794 gnd d0 a_19164_n10159# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3795 vdd a_34297_n3481# a_34089_n3481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3796 a_7834_3089# a_8087_3076# a_7830_5466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3797 a_6848_8028# a_6427_8028# a_5909_7718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3798 a_27052_3137# a_26755_4108# a_27036_3597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3799 a_5911_6066# a_6641_5822# a_6849_5822# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3800 a_9776_n10838# a_14759_n10738# a_14710_n10722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3801 vdd a_39350_9411# a_39142_9411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3802 a_20302_n9924# a_20831_n10015# a_21039_n10015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3803 gnd a_33356_6854# a_33148_6854# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3804 a_8877_7409# a_9134_7219# a_7942_6922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3805 a_20302_n10111# a_20302_n9924# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3806 a_20618_6555# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3807 gnd a_3000_4151# a_2792_4151# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3808 a_16879_n8733# a_16458_n8733# a_15940_n8423# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3809 a_39101_n2215# a_39354_n2419# a_38162_n1905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3810 gnd d2 a_28240_n9314# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3811 a_3827_n3291# a_4080_n3495# a_2888_n2981# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3812 a_22960_5406# a_23217_5216# a_22190_481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3813 a_11757_4091# a_11544_4091# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3814 a_35919_7155# a_35706_7155# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3815 a_31698_n8094# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3816 a_24011_n4924# a_24264_n5128# a_23069_n5356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3817 a_18909_6311# a_18912_5580# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3818 a_5908_8821# a_6639_9131# a_6847_9131# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3819 gnd a_24263_6605# a_24055_6605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3820 vdd d0 a_39350_n10140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3821 a_854_7128# a_1584_6884# a_1792_6884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3822 a_5701_7718# a_5488_7718# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3823 gnd d0 a_24264_n6231# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3824 a_7832_7501# a_7846_8604# a_7801_8617# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3825 vdd d2 a_13031_4156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3826 a_21771_n5359# a_21558_n5359# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3827 a_7834_n3601# a_7848_n4921# a_7799_n4905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3828 a_17976_1412# a_18960_1709# a_18911_1899# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3829 a_20831_9315# a_20618_9315# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3830 a_10464_n6176# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3831 a_856_2716# a_435_2716# a_119_2597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3832 vdd d0 a_19164_n7399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3833 a_2882_n7581# a_3139_n7597# a_2746_n6882# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3834 a_15519_7723# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3835 a_35706_n6198# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3836 a_35921_2743# a_35708_2743# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3837 a_27984_6569# a_28174_5787# a_28129_5800# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3838 a_26967_6314# a_26754_6314# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3839 a_25888_n8953# a_25675_n8953# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3840 gnd a_23328_n2063# a_23120_n2063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3841 a_2883_n5375# a_3870_n5147# a_3825_n4943# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3842 a_118_n6175# a_646_n6171# a_854_n6171# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3843 vdd a_18228_n3231# a_18020_n3231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3844 a_24012_6069# a_24265_6056# a_23073_5759# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3845 a_5174_5073# a_5703_4963# a_5911_4963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3846 a_7797_n9317# a_7987_n8741# a_7942_n8537# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3847 a_38016_4368# a_38206_3586# a_38157_3776# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3848 a_17865_n3606# a_18118_n3810# a_17861_n5994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3849 a_117_7882# a_645_7677# a_853_7677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3850 gnd a_28384_1375# a_28176_1375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3851 a_18908_n9040# a_18911_n8298# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3852 a_30864_n6711# a_30651_n6711# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3853 a_5490_n6766# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3854 a_6752_n3737# a_6539_n3737# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3855 vdd d4 a_38304_5262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3856 vdd a_14111_1114# a_13903_1114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3857 vdd a_2998_8563# a_2790_8563# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3858 a_24008_n6769# a_24265_n6785# a_23073_n6271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3859 a_3826_2225# a_3822_2402# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3860 gnd d3 a_28273_3057# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3861 vdd a_18085_8609# a_17877_8609# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3862 a_38155_n8711# a_39142_n8483# a_39097_n8279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3863 a_10886_n3970# a_10465_n3970# a_10150_n3517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3864 a_2741_n9276# a_2931_n8700# a_2882_n8684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3865 gnd d0 a_34296_3301# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3866 vdd d0 a_29320_7200# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3867 a_37066_4705# a_36999_4113# a_37083_3142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3868 a_436_n2313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3869 a_5913_1654# a_6643_1410# a_6851_1410# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3870 a_854_n7828# a_433_n7828# a_117_n7508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3871 a_11933_5213# a_11512_5213# a_11834_5213# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3872 a_10679_n1764# a_10466_n1764# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3873 a_6568_n7033# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3874 a_5491_2757# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3875 vdd a_33248_5221# a_33040_5221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3876 a_39098_n8833# a_39351_n9037# a_38159_n8523# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3877 a_30334_7868# a_30334_7411# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3878 a_32011_n4261# a_31943_n4772# a_32027_n3682# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3879 a_38017_n2685# a_38274_n2701# a_38047_n3775# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3880 a_18909_n5731# a_19166_n5747# a_17974_n5233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3881 a_21991_n3500# a_21700_n2561# a_21980_n3153# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3882 a_24005_n9524# a_24011_n8787# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3883 vdd d0 a_34294_n8442# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3884 a_36786_n4813# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3885 a_30336_n4414# a_30865_n4505# a_31073_n4505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3886 gnd d1 a_38415_n2109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3887 gnd a_13032_n2679# a_12824_n2679# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3888 gnd a_24265_2193# a_24057_2193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3889 gnd d0 a_39352_6102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3890 a_5172_n9755# a_5172_n9525# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3891 a_15204_n8886# a_15733_n8977# a_15941_n8977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3892 a_38160_n5214# a_39144_n5728# a_39099_n5524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3893 a_856_2716# a_1586_2472# a_1794_2472# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3894 a_5703_3306# a_5490_3306# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3895 a_38156_4879# a_38413_4689# a_38020_4191# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3896 a_20832_8212# a_20619_8212# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3897 a_857_1613# a_436_1613# a_120_1723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3898 vdd d0 a_19166_n6850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3899 a_7834_3089# a_7848_4192# a_7803_4205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3900 a_1696_n3696# a_1483_n3696# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3901 a_26828_2494# a_26615_2494# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3902 a_16895_n5954# a_16781_n5954# a_16989_n5954# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3903 a_1371_n8687# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3904 a_18913_n3886# a_19166_n4090# a_17971_n4318# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3905 gnd a_34296_4958# a_34088_4958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3906 a_21558_4659# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3907 a_10886_n5627# a_11616_n5383# a_11824_n5383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3908 a_5175_n2907# a_5176_n2450# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3909 a_7830_n5989# a_8087_n6005# a_7629_n10697# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3910 a_36646_2499# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3911 a_38159_6908# a_39143_7205# a_39094_7395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3912 a_2772_n8160# a_3029_n8176# a_2778_n5760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3913 gnd d0 a_14110_n6809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3914 a_35706_n7855# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3915 vdd d0 a_34296_n5687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3916 a_21991_n3500# a_21882_n3677# a_21989_n5712# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3917 a_2672_n10656# a_2622_n10672# a_2573_n10656# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3918 a_32010_n5364# a_31589_n5364# a_31071_n5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3919 a_8878_n2966# a_9135_n2982# a_7940_n3210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3920 a_30335_4789# a_30864_4908# a_31072_4908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3921 a_26725_n3718# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3922 a_7830_3266# a_8087_3076# a_7830_5466# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3923 a_15206_2413# a_15734_2208# a_15942_2208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3924 a_119_3470# a_647_3265# a_855_3265# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3925 a_7798_6588# a_7988_5806# a_7939_5996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3926 a_36129_n1786# a_36860_n2096# a_37068_n2096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3927 a_117_8341# a_117_8112# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3928 vdd a_3000_4151# a_2792_4151# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3929 a_31803_n3158# a_31590_n3158# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3930 vdd d0 a_9135_n4085# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3931 a_27985_n4886# a_28175_n4310# a_28126_n4294# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3932 a_11839_5332# a_11512_7413# a_11839_7532# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3933 vdd a_18087_4197# a_17879_4197# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3934 a_25362_n1785# a_25890_n1781# a_26098_n1781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3935 a_16459_5827# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3936 a_21041_n5603# a_20620_n5603# a_20304_n5283# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3937 a_28130_3594# a_29114_3891# a_29069_3904# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3938 a_22930_2116# a_23120_1334# a_23071_1524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3939 a_15205_6368# a_15205_6181# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3940 a_13855_9402# a_14108_9389# a_12916_9092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3941 a_853_7677# a_1584_7987# a_1792_7987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3942 a_34040_1285# a_34297_1095# a_33102_1529# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3943 a_5492_1654# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3944 vdd a_18085_n9338# a_17877_n9338# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3945 a_25362_n2015# a_25891_n2335# a_26099_n2335# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3946 a_11836_n3524# a_11545_n2585# a_11826_n2074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3947 a_26725_3018# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3948 a_27052_n3718# a_26755_n4808# a_27036_n4297# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3949 a_39096_2983# a_39099_2252# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3950 a_10676_n8382# a_10463_n8382# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3951 a_26826_8009# a_26613_8009# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3952 a_16457_9136# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3953 gnd a_18227_4708# a_18019_4708# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3954 a_36127_7155# a_36857_6911# a_37065_6911# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3955 a_22929_n4845# a_23186_n4861# a_22964_n3541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3956 vdd d1 a_13173_n2087# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3957 a_29062_7939# a_29319_7749# a_28124_8183# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3958 a_38014_n9303# a_38271_n9319# a_38049_n7999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3959 gnd d1 a_23327_n4269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3960 a_24007_n5112# a_24013_n4375# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3961 vdd a_14111_n4603# a_13903_n4603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3962 a_31731_1866# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3963 a_23072_n7374# a_24056_n7888# a_24011_n7684# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3964 a_38159_n7420# a_39143_n7934# a_39094_n7918# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3965 a_31587_n9776# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3966 a_1370_9090# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3967 a_24008_6246# a_24265_6056# a_23073_5759# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3968 a_36128_n3992# a_35707_n3992# a_35392_n3996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3969 a_38016_4368# a_38206_3586# a_38161_3599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3970 a_5702_n8972# a_5489_n8972# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3971 a_34038_n6220# a_34295_n6236# a_33100_n6464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3972 a_644_n9480# a_431_n9480# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3973 a_22081_481# a_21868_481# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3974 a_19332_n829# a_19119_n829# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3975 vdd a_28384_1375# a_28176_1375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3976 a_5910_n5109# a_5489_n5109# a_5174_n5113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3977 a_27036_n3194# a_26615_n3194# a_26098_n3438# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3978 a_16982_546# a_16769_546# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3979 a_21039_7658# a_21770_7968# a_21978_7968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3980 a_31911_n8094# a_31698_n8094# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3981 a_12913_7063# a_13900_6629# a_13855_6642# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3982 a_1373_2472# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3983 a_28128_8006# a_28381_7993# a_27983_8775# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3984 a_20304_5887# a_20304_5657# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3985 a_17970_n6524# a_18227_n6540# a_17829_n7116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3986 a_20618_n10015# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3987 a_18908_n6280# a_18913_n5543# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X3988 a_15520_n6217# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3989 gnd d0 a_24264_4399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3990 a_5910_8272# a_5489_8272# a_5173_8153# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3991 a_15209_1211# a_15735_1105# a_15943_1105# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3992 a_39098_5561# a_39351_5548# a_38156_5982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3993 a_8875_n9584# a_9132_n9600# a_7937_n9828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3994 a_31072_n5608# a_30651_n5608# a_30335_n5288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3995 a_36858_n5405# a_36645_n5405# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3996 a_38015_n7097# a_38205_n6521# a_38160_n6317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3997 a_21041_n3946# a_21772_n4256# a_21980_n4256# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3998 gnd a_38304_5262# a_38096_5262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X3999 a_36128_3292# a_35707_3292# a_35392_3040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4000 a_34042_8280# a_34038_8457# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4001 vdd d0 a_24266_2747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4002 a_35391_5246# a_35391_5059# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4003 a_17834_4210# a_18019_4708# a_17974_4721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4004 a_11834_5213# a_11514_3001# a_11841_3120# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4005 a_25359_n8403# a_25887_n8399# a_26095_n8399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4006 a_27144_5230# a_26723_5230# a_27045_5230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4007 a_25359_n8633# a_25359_n8403# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4008 a_432_n10034# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4009 a_17969_n7627# a_18956_n7399# a_18911_n7195# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4010 a_15522_n3462# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4011 a_116_8985# a_117_8528# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4012 vdd a_8196_n6535# a_7988_n6535# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4013 a_11839_n8113# a_11542_n9203# a_11823_n8692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4014 a_22928_6528# a_23185_6338# a_22958_7618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4015 a_1791_9090# a_1370_9090# a_852_8780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4016 a_25358_9007# a_25359_8550# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4017 a_119_n3096# a_648_n3416# a_856_n3416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4018 a_3823_8843# a_3819_9020# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4019 a_1694_n5908# a_1481_n5908# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4020 a_25362_n1785# a_24985_n1506# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4021 gnd d0 a_19163_8876# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4022 a_15943_n4565# a_15522_n4565# a_15206_n4245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4023 a_15735_n1805# a_15522_n1805# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4024 gnd d1 a_18226_n7643# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4025 a_35918_n10061# a_35705_n10061# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4026 gnd a_33358_n3171# a_33150_n3171# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4027 a_27037_n2091# a_26616_n2091# a_26098_n1781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4028 a_31071_8217# a_30650_8217# a_30334_8098# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4029 a_13851_n8445# a_14108_n8461# a_12913_n8689# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4030 gnd a_8197_n4329# a_7989_n4329# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4031 a_15944_1659# a_16674_1415# a_16882_1415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4032 a_37846_n10683# a_38103_n10699# a_34896_n10703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4033 a_37066_n5405# a_36999_n4813# a_37083_n3723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4034 gnd a_19166_n2987# a_18958_n2987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4035 a_5704_3860# a_5491_3860# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4036 a_15736_n2359# a_15523_n2359# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4037 a_8880_9438# a_9133_9425# a_7941_9128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4038 gnd a_38412_6895# a_38204_6895# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4039 a_21980_2453# a_21559_2453# a_21042_2697# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4040 a_37078_n3546# a_36787_n2607# a_37067_n3199# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4041 a_12915_2651# a_13902_2217# a_13857_2230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4042 a_11823_7992# a_11755_8503# a_11839_7532# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4043 a_25359_8134# a_25359_7904# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4044 a_10679_3824# a_10466_3824# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4045 a_34038_n7877# a_34295_n7893# a_33103_n7379# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4046 a_30336_n3082# a_30336_n2852# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4047 a_15204_8387# a_15733_8277# a_15941_8277# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4048 a_8877_n9035# a_9134_n9051# a_7942_n8537# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4049 a_4679_n10717# a_4936_n10733# a_4778_n10717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4050 a_34039_n4014# a_34044_n3277# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4051 vdd d1 a_8198_n2123# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4052 a_39100_1149# a_39353_1136# a_38158_1570# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4053 a_22930_2116# a_23120_1334# a_23075_1347# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4054 a_22927_n9257# a_23117_n8681# a_23072_n8477# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4055 a_10677_7133# a_10464_7133# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4056 a_13856_n6051# a_13852_n6239# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4057 a_30652_n4505# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4058 a_15940_n7320# a_16671_n7630# a_16879_n7630# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4059 a_16881_3621# a_16460_3621# a_15942_3311# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4060 a_32009_6870# a_31588_6870# a_31071_7114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4061 a_29063_n5153# a_29069_n4416# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4062 a_35706_7155# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4063 a_1585_4678# a_1372_4678# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4064 a_854_n8931# a_1584_n8687# a_1792_n8687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4065 a_17974_n6336# a_18958_n6850# a_18913_n6646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4066 gnd d0 a_14109_7183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4067 a_8878_2443# a_8884_1717# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4068 gnd d0 a_14107_n9564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4069 a_16568_n5954# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4070 a_29068_6110# a_29321_6097# a_28129_5800# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4071 a_116_n9484# a_644_n9480# a_852_n9480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4072 a_25358_n9965# a_25887_n10056# a_26095_n10056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4073 a_11617_n4280# a_11404_n4280# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4074 a_31588_7973# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4075 a_12918_n6295# a_13902_n6809# a_13853_n6793# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4076 a_21669_n3677# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4077 a_39101_1703# a_39097_1880# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4078 vdd d1 a_13169_9079# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4079 a_26754_6314# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4080 a_29067_n4965# a_29320_n5169# a_28125_n5397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4081 a_32991_n5934# a_33040_n3750# a_32991_n3734# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4082 a_2774_n3748# a_2793_n2674# a_2744_n2658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4083 a_26096_n7850# a_25675_n7850# a_25359_n7759# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4084 a_37068_1396# a_36647_1396# a_36129_1086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4085 a_15732_n8423# a_15519_n8423# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4086 a_33104_4661# a_34088_4958# a_34039_5148# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4087 a_27034_n8709# a_26613_n8709# a_26095_n8399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4088 a_17865_5294# a_18118_5281# a_17091_546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4089 a_117_7009# a_117_6779# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4090 gnd d3 a_18116_n8222# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4091 a_10884_n7279# a_10463_n7279# a_10149_n6826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4092 a_5173_7466# a_5173_7279# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4093 a_8882_5026# a_9135_5013# a_7943_4716# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4094 gnd a_38412_n8727# a_38204_n8727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4095 gnd d0 a_29320_n6272# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4096 a_35920_3292# a_35707_3292# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4097 a_39097_7767# a_39093_7944# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4098 a_7940_n4313# a_8927_n4085# a_8882_n3881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4099 a_26827_n6503# a_26614_n6503# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4100 a_25677_n1781# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4101 vdd a_38304_5262# a_38096_5262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4102 a_2778_5248# a_3031_5235# a_2004_500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4103 a_37081_n8135# a_36784_n9225# a_37064_n9817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4104 a_30862_n7260# a_30649_n7260# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4105 a_15943_2762# a_15522_2762# a_15206_2643# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4106 a_11825_3580# a_11757_4091# a_11841_3120# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4107 vdd a_13029_n9297# a_12821_n9297# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4108 gnd a_28273_3057# a_28065_3057# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4109 a_10151_n2414# a_10678_n2867# a_10886_n2867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4110 a_25678_n2335# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4111 a_5174_5717# a_5702_5512# a_5910_5512# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4112 a_21042_3800# a_20621_3800# a_20305_3910# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4113 a_35392_n2893# a_35920_n2889# a_36128_n2889# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4114 gnd a_34296_3301# a_34088_3301# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4115 a_15521_n2908# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4116 a_32964_n4662# a_33217_n4866# a_32995_n3546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4117 a_15734_n5668# a_15521_n5668# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4118 a_10150_n2871# a_10151_n2414# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4119 a_12775_n2663# a_12965_n2087# a_12920_n1883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4120 a_35392_n3123# a_35921_n3443# a_36129_n3443# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4121 vdd a_28383_n3207# a_28175_n3207# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4122 a_35707_6052# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4123 a_30336_2999# a_30864_3251# a_31072_3251# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4124 a_30864_6011# a_30651_6011# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4125 a_3820_7917# a_4077_7727# a_2882_8161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4126 a_22960_n5929# a_23217_n5945# a_22759_n10637# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4127 gnd d1 a_33357_n5377# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4128 a_26098_n4541# a_26828_n4297# a_27036_n4297# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4129 gnd a_39352_6102# a_39144_6102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4130 a_27050_n5930# a_26723_n8130# a_27050_n8130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4131 a_31731_n2566# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4132 a_5490_3306# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4133 a_21771_5762# a_21558_5762# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4134 a_26615_2494# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4135 a_8876_9615# a_9133_9425# a_7941_9128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4136 a_17830_n4910# a_18020_n4334# a_17971_n4318# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4137 a_7800_2176# a_8057_1986# a_7830_3266# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4138 gnd a_2999_6357# a_2791_6357# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4139 a_32025_n8094# a_31728_n9184# a_32009_n8673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4140 a_29069_n4416# a_29322_n4620# a_28130_n4106# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4141 a_25360_n5740# a_25360_n5553# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4142 a_11756_6297# a_11543_6297# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4143 a_2776_n7972# a_2790_n9292# a_2741_n9276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4144 a_24012_6069# a_24008_6246# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4145 a_39095_n4055# a_39100_n3318# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4146 a_21559_n4256# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4147 a_3820_6814# a_3826_6088# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4148 a_118_n6175# a_118_n5718# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4149 a_1791_n9790# a_1370_n9790# a_852_n9480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4150 a_19441_n829# a_20582_n10911# a_20533_n10895# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4151 a_39096_1326# a_39353_1136# a_38158_1570# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4152 vdd a_39354_n2419# a_39146_n2419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4153 a_6752_n3737# a_6539_n3737# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4154 a_22088_5189# a_21667_5189# a_21994_5308# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4155 a_30864_n6711# a_30651_n6711# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4156 a_5490_n6766# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4157 a_25674_n8399# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4158 a_31071_n5054# a_31802_n5364# a_32010_n5364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4159 vdd d0 a_4080_n4598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4160 a_5910_n6212# a_6641_n6522# a_6849_n6522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4161 a_13855_7745# a_13851_7922# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4162 a_36645_n5405# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4163 a_37277_527# a_38096_5262# a_38047_5452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4164 a_7834_5289# a_7877_7488# a_7828_7678# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4165 gnd a_39351_n6277# a_39143_n6277# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4166 vdd a_28381_n8722# a_28173_n8722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4167 a_10148_n9032# a_10675_n9485# a_10883_n9485# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4168 a_34042_n7689# a_34038_n7877# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4169 vdd d0 a_14109_7183# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4170 a_2745_8576# a_2930_9074# a_2881_9264# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4171 a_436_n2313# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4172 a_31698_5194# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4173 a_16881_n3218# a_16460_n3218# a_15943_n3462# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4174 a_11822_9095# a_11401_9095# a_10884_9339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4175 a_20304_n5283# a_20833_n5603# a_21041_n5603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4176 a_10679_n1764# a_10466_n1764# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4177 a_26097_2184# a_26828_2494# a_27036_2494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4178 vdd d0 a_24263_7708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4179 a_26613_8009# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4180 a_36126_n7301# a_35705_n7301# a_35390_n7305# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4181 a_32010_n5364# a_31943_n4772# a_32027_n3682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4182 a_21991_n3500# a_21700_n2561# a_21981_n2050# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4183 a_36860_1396# a_36647_1396# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4184 a_36786_n4813# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4185 a_6849_n5419# a_6428_n5419# a_5910_n5109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4186 a_24010_9378# a_24006_9555# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4187 gnd d0 a_34295_5507# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4188 vdd d0 a_29319_9406# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4189 a_37065_6911# a_36998_6319# a_37076_7435# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4190 a_21773_1350# a_21560_1350# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4191 a_17861_5471# a_18118_5281# a_17091_546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4192 a_23067_9245# a_24054_8811# a_24009_8824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4193 a_5912_3860# a_6642_3616# a_6850_3616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4194 gnd d0 a_19168_1709# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4195 vdd a_39351_7205# a_39143_7205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4196 a_8878_5203# a_9135_5013# a_7943_4716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4197 a_20619_4349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4198 a_25890_n3438# a_25677_n3438# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4199 gnd a_3001_1945# a_2793_1945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4200 a_35919_8258# a_35706_8258# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4201 a_27985_n4886# a_28242_n4902# a_28020_n3582# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4202 vdd d1 a_18229_n2128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4203 a_2774_5425# a_3031_5235# a_2004_500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4204 a_33104_n6276# a_34088_n6790# a_34039_n6774# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4205 gnd d1 a_28383_n4310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4206 a_16890_5254# a_16570_3042# a_16897_3161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4207 a_5909_6615# a_6640_6925# a_6848_6925# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4208 a_15941_n7874# a_15520_n7874# a_15204_n7783# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4209 a_8878_n2966# a_8884_n2229# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4210 gnd a_24264_4399# a_24056_4399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4211 a_21996_n3677# a_21882_n3677# a_21989_n5712# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4212 a_15732_9380# a_15519_9380# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4213 a_25886_8802# a_25673_8802# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4214 gnd d0 a_39351_8308# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4215 a_28128_n7415# a_29112_n7929# a_29067_n7725# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4216 a_13857_2230# a_14110_2217# a_12915_2651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4217 vdd a_23187_1926# a_22979_1926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4218 a_16458_n7630# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4219 a_10463_n10039# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4220 a_855_4922# a_1585_4678# a_1793_4678# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4221 a_12915_n4277# a_13172_n4293# a_12774_n4869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4222 gnd a_39353_n4625# a_39145_n4625# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4223 vdd a_24266_n4579# a_24058_n4579# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4224 a_38155_7085# a_38412_6895# a_38019_6397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4225 a_32020_5194# a_31911_5194# a_32119_5194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4226 a_856_3819# a_435_3819# a_119_3929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4227 a_32962_n9074# a_33147_n9789# a_33102_n9585# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4228 a_22931_8557# a_23184_8544# a_22962_7441# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4229 a_3823_n9355# a_3819_n9543# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4230 gnd a_24263_n7334# a_24055_n7334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4231 a_39094_n6261# a_39351_n6277# a_38156_n6505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4232 a_27984_6569# a_28241_6379# a_28014_7659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4233 a_20832_7109# a_20619_7109# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4234 a_10148_n8616# a_10677_n8936# a_10885_n8936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4235 gnd a_4079_n6804# a_3871_n6804# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4236 a_15204_n7324# a_15205_n6867# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4237 vdd a_24266_2747# a_24058_2747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4238 a_26968_4108# a_26755_4108# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4239 a_7830_5466# a_7879_3076# a_7830_3266# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4240 a_6781_6333# a_6568_6333# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4241 a_35392_n4642# a_35392_n4455# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4242 a_25674_n10056# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4243 a_12916_9092# a_13169_9079# a_12776_8581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4244 a_36860_n2096# a_36647_n2096# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4245 a_20303_7406# a_20303_7219# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4246 a_7942_6922# a_8926_7219# a_8881_7232# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4247 a_31943_n4772# a_31730_n4772# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4248 a_6864_5368# a_6750_5249# a_6958_5249# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4249 a_10150_3018# a_10150_2831# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4250 a_26096_5493# a_25675_5493# a_25360_5698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4251 a_25362_n2244# a_25891_n2335# a_26099_n2335# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4252 vdd a_3138_n9803# a_2930_n9803# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4253 a_35390_6806# a_35918_6601# a_36126_6601# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4254 a_21978_n8668# a_21557_n8668# a_21039_n8358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4255 a_20834_n3397# a_20621_n3397# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4256 a_32961_n2644# a_33151_n2068# a_33102_n2052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4257 a_15205_n6680# a_15205_n6451# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4258 gnd d0 a_19164_9430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4259 a_29067_5556# a_29063_5733# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4260 a_119_3470# a_119_3013# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4261 vdd a_3031_n3764# a_2823_n3764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4262 a_30650_n7814# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4263 a_21771_n5359# a_21558_n5359# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4264 a_30335_n5704# a_30863_n6157# a_31071_n6157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4265 a_10680_n2318# a_10467_n2318# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4266 a_12914_4857# a_13901_4423# a_13852_4613# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4267 a_7942_n8537# a_8195_n8741# a_7797_n9317# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4268 a_7941_n9640# a_8925_n10154# a_5172_n10171# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4269 gnd a_19163_8876# a_18955_8876# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4270 a_17865_n5806# a_17908_n8222# a_17859_n8206# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4271 a_25031_461# a_24818_461# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4272 a_21989_5189# a_21669_2977# a_21996_3096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4273 gnd d0 a_9137_n2433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4274 vdd a_18086_6403# a_17878_6403# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4275 a_11822_n9795# a_11401_n9795# a_10884_n10039# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4276 vdd a_7886_n10713# a_7678_n10713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4277 gnd d0 a_34297_1095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4278 vdd d0 a_29321_4994# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4279 a_3822_5162# a_4079_4972# a_2887_4675# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4280 a_25361_n3118# a_25361_n2888# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4281 gnd d1 a_13171_n5396# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4282 a_23069_4833# a_24056_4399# a_24011_4412# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4283 a_5491_3860# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4284 gnd d2 a_38271_8590# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4285 a_5702_n8972# a_5489_n8972# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4286 a_12777_n6887# a_13030_n7091# a_12803_n8165# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4287 gnd d0 a_24265_n2922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4288 gnd a_3142_n2082# a_2934_n2082# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4289 gnd d0 a_39350_n7380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4290 a_10465_n2867# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4291 a_35707_n2889# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4292 a_6750_n5949# a_6537_n5949# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4293 a_2886_7984# a_3870_8281# a_3821_8471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4294 a_10466_3824# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4295 a_27137_522# a_26924_522# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4296 a_37277_527# a_38096_5262# a_38051_5275# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4297 a_29069_2801# a_29065_2978# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4298 vdd a_34293_n9545# a_34085_n9545# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4299 gnd a_38414_n3212# a_38206_n3212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4300 a_855_3265# a_1586_3575# a_1794_3575# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4301 a_648_n4519# a_435_n4519# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4302 a_35708_n3443# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4303 gnd d0 a_39353_3896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4304 a_10886_n3970# a_10465_n3970# a_10150_n3974# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4305 a_2745_8576# a_2930_9074# a_2885_9087# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4306 a_33101_3735# a_34088_3301# a_34039_3491# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4307 a_21042_n4500# a_21772_n4256# a_21980_n4256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4308 a_15940_7723# a_15519_7723# a_15204_7471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4309 a_20833_6006# a_20620_6006# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4310 a_24006_n8421# a_24263_n8437# a_23068_n8665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4311 a_116_n9714# a_645_n10034# a_853_n10034# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4312 a_22933_4145# a_23186_4132# a_22964_3029# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4313 vdd a_19165_n7953# a_18957_n7953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4314 a_10464_7133# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4315 a_26615_n4297# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4316 a_21994_n5889# a_21667_n8089# a_21994_n8089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4317 a_4679_n10717# a_7678_n10713# a_7629_n10697# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4318 a_6859_7449# a_6750_7449# a_6864_5368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4319 a_11756_n6997# a_11543_n6997# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4320 a_854_n7828# a_433_n7828# a_117_n7737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4321 a_36998_n7019# a_36785_n7019# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4322 a_1372_4678# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4323 a_21039_n7255# a_20618_n7255# a_20303_n7259# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4324 a_39094_n7918# a_39351_n7934# a_38159_n7420# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4325 a_15206_n2912# a_15207_n2455# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4326 a_38160_4702# a_39144_4999# a_39095_5189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4327 vdd d1 a_18227_5811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4328 a_26098_1081# a_25677_1081# a_25362_1286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4329 gnd a_19165_n6296# a_18957_n6296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4330 a_30335_6121# a_30335_5892# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4331 a_15943_n3462# a_16673_n3218# a_16881_n3218# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4332 a_26096_n6193# a_25675_n6193# a_25360_n5740# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4333 vdd a_39351_n5174# a_39143_n5174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4334 a_120_1264# a_648_1059# a_856_1059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4335 a_36127_5498# a_35706_5498# a_35391_5246# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4336 a_119_n3325# a_648_n3416# a_856_n3416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4337 a_34043_3314# a_34039_3491# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4338 a_39099_n5524# a_39352_n5728# a_38160_n5214# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4339 gnd d4 a_13062_5240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4340 vdd d0 a_24265_4953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4341 a_17833_6416# a_18018_6914# a_17973_6927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4342 gnd d0 a_9134_n9051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4343 a_26095_n7296# a_26826_n7606# a_27034_n7606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4344 vdd a_18088_1991# a_17880_1991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4345 vdd d2 a_8057_n2715# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4346 a_7941_9128# a_8194_9115# a_7801_8617# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4347 a_3825_n7703# a_4078_n7907# a_2886_n7393# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4348 a_8875_n9584# a_8881_n8847# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4349 a_18909_5208# a_18912_4477# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4350 a_31589_n5364# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4351 a_21041_2143# a_20620_2143# a_20305_2348# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4352 gnd d0 a_39352_n6831# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4353 a_25359_7260# a_25888_7150# a_26096_7150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4354 a_117_n8381# a_117_n7924# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4355 gnd d0 a_24262_n9540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4356 a_26723_n5930# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4357 a_28129_n6312# a_28382_n6516# a_27984_n7092# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4358 a_6640_8028# a_6427_8028# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4359 a_22927_8734# a_23184_8544# a_22962_7441# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4360 a_10462_n9485# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4361 a_37078_n3546# a_36787_n2607# a_37068_n2096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4362 a_16458_6930# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4363 vdd d0 a_14108_6629# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4364 a_26098_n3438# a_25677_n3438# a_25361_n3118# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4365 gnd d0 a_4078_n9010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4366 a_1805_n3519# a_1696_n3696# a_1803_n5731# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4367 a_36128_4949# a_36858_4705# a_37066_4705# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4368 a_8876_7958# a_9133_7768# a_7938_8202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4369 gnd a_23326_n5372# a_23118_n5372# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4370 a_30074_345# a_34849_466# a_35171_466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4371 a_7830_5466# a_7879_3076# a_7834_3089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4372 a_30336_3456# a_30336_2999# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4373 a_27034_n7606# a_26967_n7014# a_27045_n7953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4374 gnd d0 a_19167_n1884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4375 a_14985_485# a_16769_546# a_17091_546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4376 a_646_8231# a_433_8231# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4377 a_15942_3311# a_15521_3311# a_15206_3059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4378 a_5176_n1804# a_5704_n1800# a_5912_n1800# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4379 a_1727_1880# a_1514_1880# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4380 a_30651_6011# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4381 a_27052_n3718# a_26755_n4808# a_27035_n5400# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4382 a_6861_3037# a_6752_3037# a_6859_5249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4383 vdd d0 a_19164_9430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4384 gnd d1 a_13170_6873# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4385 a_18908_n7937# a_18911_n7195# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4386 a_35918_n8404# a_35705_n8404# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4387 a_24006_n10078# a_24263_n10094# a_23071_n9580# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4388 a_12914_4857# a_13901_4423# a_13856_4436# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4389 a_5176_n2034# a_5705_n2354# a_5913_n2354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4390 a_30649_7663# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4391 a_5911_6066# a_5490_6066# a_5174_5947# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4392 a_28125_4874# a_29112_4440# a_29063_4630# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4393 a_434_n5622# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4394 gnd d1 a_3141_n4288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4395 a_10676_9339# a_10463_9339# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4396 a_853_6574# a_432_6574# a_117_6779# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4397 a_36129_1086# a_35708_1086# a_35395_1192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4398 a_21669_n3677# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4399 a_26098_2738# a_25677_2738# a_25361_2848# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4400 a_16880_5827# a_16459_5827# a_15941_5517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4401 gnd a_34297_n4584# a_34089_n4584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4402 a_34896_n10703# a_35153_n10719# a_29962_n10819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4403 vdd d1 a_38412_7998# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4404 a_2886_7984# a_3870_8281# a_3825_8294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4405 a_30334_6765# a_30335_6308# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4406 a_39097_1880# a_39354_1690# a_38162_1393# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4407 vdd d2 a_8054_n9333# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4408 a_13859_n2193# a_13855_n2381# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4409 a_3821_n5131# a_4078_n5147# a_2883_n5375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4410 a_10464_n8936# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4411 vdd d2 a_38272_n7113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4412 a_21978_7968# a_21557_7968# a_21040_8212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4413 a_26827_n6503# a_26614_n6503# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4414 a_31072_n5608# a_30651_n5608# a_30335_n5517# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4415 vdd d0 a_29319_7749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4416 a_36128_3292# a_36859_3602# a_37067_3602# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4417 a_22929_4322# a_23186_4132# a_22964_3029# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4418 a_37081_n8135# a_36784_n9225# a_37065_n8714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4419 a_18911_n7195# a_19164_n7399# a_17969_n7627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4420 a_38018_8603# a_38203_9101# a_38158_9114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4421 vdd a_39351_5548# a_39143_5548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4422 vdd d2 a_18087_n4926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4423 a_3825_5534# a_4078_5521# a_2883_5955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4424 vdd d0 a_4078_n6250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4425 gnd d2 a_8055_n7127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4426 a_38160_n6317# a_38413_n6521# a_38015_n7097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4427 a_10150_n2871# a_10678_n2867# a_10886_n2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4428 a_25678_n2335# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4429 a_25890_n1781# a_25677_n1781# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4430 vdd a_13062_n3769# a_12854_n3769# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4431 gnd d0 a_19164_n8502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4432 a_2886_n8496# a_3139_n8700# a_2741_n9276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4433 a_28123_9286# a_29110_8852# a_29065_8865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4434 a_35392_n3352# a_35921_n3443# a_36129_n3443# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4435 vdd a_24263_7708# a_24055_7708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4436 a_8881_7232# a_9134_7219# a_7942_6922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4437 a_10150_2602# a_10150_2372# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4438 a_2883_n6478# a_3870_n6250# a_3821_n6234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4439 a_7945_n1919# a_8929_n2433# a_8880_n2417# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4440 a_26936_5230# a_26723_5230# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4441 vdd d0 a_19166_5018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4442 a_15942_4968# a_15521_4968# a_15205_4849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4443 a_11824_5786# a_11756_6297# a_11834_7413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4444 a_117_7238# a_117_7009# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4445 a_12778_n4681# a_12963_n5396# a_12914_n5380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4446 a_20832_5452# a_20619_5452# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4447 vdd d4 a_13062_5240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4448 a_1694_n5908# a_1481_n5908# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4449 a_25360_n5094# a_25888_n5090# a_26096_n5090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4450 a_11826_n2074# a_11405_n2074# a_10888_n2318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4451 a_5173_7923# a_5701_7718# a_5909_7718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4452 a_39094_8498# a_39097_7767# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4453 a_31731_n2566# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4454 gnd a_34295_5507# a_34087_5507# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4455 a_20306_1475# a_20306_1245# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4456 a_3823_n1822# a_4799_n1525# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4457 a_22958_7618# a_22977_6338# a_22932_6351# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4458 a_7937_9305# a_8194_9115# a_7801_8617# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4459 a_32025_7513# a_31728_8484# a_32009_7973# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4460 a_21560_1350# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4461 a_29066_n8274# a_29062_n8462# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4462 gnd a_19168_1709# a_18960_1709# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4463 a_37076_5235# a_36967_5235# a_37175_5235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4464 a_20302_9425# a_20831_9315# a_21039_9315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4465 a_15205_5265# a_15205_5078# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4466 a_25360_n5324# a_25889_n5644# a_26097_n5644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4467 a_27987_8598# a_28240_8585# a_28018_7482# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4468 vdd d2 a_38273_4178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4469 a_20533_n10895# a_30011_n10835# a_29962_n10819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4470 a_10678_4927# a_10465_4927# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4471 a_35392_2624# a_35921_2743# a_36129_2743# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4472 a_855_2162# a_434_2162# a_119_2367# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4473 a_35706_8258# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4474 vdd d1 a_33356_7957# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4475 a_30863_8217# a_30650_8217# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4476 a_16882_1415# a_16461_1415# a_15943_1105# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4477 a_20834_n1740# a_20621_n1740# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4478 gnd d1 a_23325_n7578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4479 a_30336_2353# a_30864_2148# a_31072_2148# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4480 vdd a_14109_n7912# a_13901_n7912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4481 a_21559_n4256# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4482 a_15734_n4011# a_15521_n4011# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4483 a_7941_9128# a_8925_9425# a_8876_9615# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4484 gnd d0 a_14110_4977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4485 a_25673_8802# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4486 a_13857_2230# a_13853_2407# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4487 a_20835_n2294# a_20622_n2294# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4488 a_21770_7968# a_21557_7968# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4489 a_18913_n6646# a_19166_n6850# a_17974_n6336# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4490 a_11839_7532# a_11542_8503# a_11822_9095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4491 a_31072_n5608# a_31802_n5364# a_32010_n5364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4492 vdd d0 a_29321_3337# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4493 a_31589_5767# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4494 a_5911_n6766# a_6641_n6522# a_6849_n6522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4495 a_10148_8346# a_10148_8117# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4496 a_36645_n5405# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4497 vdd d5 a_38103_n10699# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4498 gnd a_33218_n2660# a_33010_n2660# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4499 a_1584_n7584# a_1371_n7584# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4500 a_29962_n10819# a_30219_n10835# a_20533_n10895# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4501 a_24013_1103# a_24009_1280# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4502 a_26755_4108# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4503 a_35390_n9054# a_35390_n8867# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4504 a_17968_n9833# a_18225_n9849# a_17832_n9134# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4505 a_5908_n9521# a_5487_n9521# a_5172_n9525# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4506 a_31587_9076# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4507 a_20304_4784# a_20304_4554# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4508 a_28125_4874# a_29112_4440# a_29067_4453# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4509 a_20304_n5512# a_20833_n5603# a_21041_n5603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4510 vdd a_29322_n4620# a_29114_n4620# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4511 a_38018_n9115# a_38203_n9830# a_38158_n9626# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4512 a_29065_n1844# a_29322_n1860# a_28127_n2088# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4513 a_35921_1086# a_35708_1086# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4514 a_36126_n7301# a_35705_n7301# a_35391_n6848# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4515 a_21039_n7255# a_21770_n7565# a_21978_n7565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4516 gnd a_19164_9430# a_18956_9430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4517 a_15943_3865# a_15522_3865# a_15206_3975# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4518 a_7942_n8537# a_8926_n9051# a_8877_n9035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4519 vdd a_33357_n6480# a_33149_n6480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4520 a_26613_n7606# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4521 a_16897_n3742# a_16600_n4832# a_16880_n5424# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4522 a_7830_n3789# a_7849_n2715# a_7804_n2511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4523 gnd d0 a_34296_n6790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4524 gnd a_3031_n5964# a_2823_n5964# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4525 a_11826_1374# a_11758_1885# a_11836_3001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4526 a_116_9215# a_645_9334# a_853_9334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4527 gnd a_29319_n8478# a_29111_n8478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4528 a_34042_7177# a_34038_7354# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4529 a_11825_n3177# a_11404_n3177# a_10886_n2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4530 a_20834_1040# a_20621_1040# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4531 a_5175_3511# a_5703_3306# a_5911_3306# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4532 gnd a_34297_1095# a_34089_1095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4533 a_20303_8093# a_20832_8212# a_21040_8212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4534 a_27034_n8709# a_26613_n8709# a_26096_n8953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4535 a_28020_n5782# a_28063_n8198# a_28014_n8182# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4536 a_25359_n7530# a_25359_n7300# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4537 a_1483_n3696# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4538 a_13852_8476# a_13855_7745# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4539 a_38159_8011# a_39143_8308# a_39098_8321# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4540 a_27989_4186# a_28242_4173# a_28020_3070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4541 a_26096_4390# a_26827_4700# a_27035_4700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4542 a_26094_n9502# a_25673_n9502# a_25358_n9506# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4543 a_1792_n7584# a_1725_n6992# a_1803_n7931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4544 a_30339_1151# a_30865_1045# a_31073_1045# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4545 a_26754_n7014# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4546 a_20831_n8358# a_20618_n8358# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4547 vdd d1 a_3141_n3185# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4548 a_17972_n2112# a_18959_n1884# a_18910_n1868# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4549 a_3821_5711# a_4078_5521# a_2883_5955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4550 a_15941_n7874# a_15520_n7874# a_15204_n7554# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4551 a_30862_n7260# a_30649_n7260# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4552 a_15733_n5114# a_15520_n5114# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4553 a_5175_n4656# a_5702_n5109# a_5910_n5109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4554 a_120_n1763# a_648_n1759# a_856_n1759# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4555 a_4954_480# a_6738_541# a_6958_5249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4556 a_32025_n5894# a_31698_n8094# a_32020_n7917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4557 a_7943_4716# a_8927_5013# a_8878_5203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4558 a_28128_n8518# a_29112_n9032# a_29063_n9016# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4559 a_6641_n6522# a_6428_n6522# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4560 gnd d4 a_28273_n5986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4561 gnd d0 a_4079_2212# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4562 a_10675_8785# a_10462_8785# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4563 a_5491_n1800# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4564 gnd a_39353_3896# a_39145_3896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4565 gnd d3 a_23215_n8157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4566 gnd a_8195_n7638# a_7987_n7638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4567 a_21772_3556# a_21559_3556# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4568 a_2004_500# a_2823_5235# a_2774_5425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4569 a_20620_6006# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4570 a_15734_n5668# a_15521_n5668# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4571 a_11841_3120# a_11544_4091# a_11824_4683# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4572 a_32964_4150# a_33149_4648# a_33104_4661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4573 gnd d0 a_29321_n2963# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4574 a_17829_n7116# a_18086_n7132# a_17859_n8206# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4575 a_5492_n2354# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4576 a_10148_n8845# a_10677_n8936# a_10885_n8936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4577 a_23072_n8477# a_24056_n8991# a_24007_n8975# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4578 gnd a_33215_n9278# a_33007_n9278# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4579 a_24010_n2357# a_24267_n2373# a_23075_n1859# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4580 a_39096_8870# a_39092_9047# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4581 a_2743_n4864# a_2933_n4288# a_2884_n4272# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4582 a_20620_n2843# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4583 gnd d1 a_3138_9074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4584 a_31943_n4772# a_31730_n4772# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4585 vdd d2 a_23187_n2655# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4586 a_22958_7618# a_23215_7428# a_22964_5229# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4587 a_31941_8484# a_31728_8484# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4588 vdd a_18227_5811# a_18019_5811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4589 a_13857_n3845# a_14110_n4049# a_12915_n4277# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4590 a_34041_6623# a_34294_6610# a_33099_7044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4591 a_120_1723# a_649_1613# a_857_1613# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4592 a_35390_8555# a_35390_8368# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4593 a_1585_5781# a_1372_5781# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4594 a_34039_n2911# a_34045_n2174# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4595 a_2774_n5948# a_3031_n5964# a_2573_n10656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4596 a_15205_5722# a_15205_5265# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4597 a_37065_n8714# a_36644_n8714# a_36127_n8958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4598 a_6429_2513# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4599 a_2882_8161# a_3869_7727# a_3824_7740# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4600 vdd d3 a_18116_7493# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4601 a_27983_8775# a_28240_8585# a_28018_7482# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4602 a_30650_n7814# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4603 a_21041_n3946# a_20620_n3946# a_20305_n3950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4604 a_31074_1599# a_31804_1355# a_32012_1355# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4605 gnd a_38103_n10699# a_37895_n10699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4606 a_33101_n4258# a_34088_n4030# a_34043_n3826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4607 a_7832_n8013# a_7846_n9333# a_7801_n9129# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4608 a_38051_n3587# a_38065_n4907# a_38016_n4891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4609 a_13856_n4948# a_13852_n5136# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4610 a_29066_7762# a_29319_7749# a_28124_8183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4611 a_24008_n5666# a_24011_n4924# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4612 gnd a_13062_5240# a_12854_5240# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4613 a_118_4803# a_647_4922# a_855_4922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4614 vdd a_24265_4953# a_24057_4953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4615 vdd d0 a_14108_n10118# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4616 a_36126_9361# a_35705_9361# a_35389_9471# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4617 a_6780_8539# a_6567_8539# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4618 a_21911_n6973# a_21698_n6973# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4619 a_16671_8033# a_16458_8033# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4620 vdd a_39353_n1865# a_39145_n1865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4621 a_7941_9128# a_8925_9425# a_8880_9438# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4622 a_21880_5189# a_21667_5189# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4623 a_7830_3266# a_7849_1986# a_7804_1999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4624 a_2746_6370# a_2931_6868# a_2882_7058# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4625 vdd a_28243_n2696# a_28035_n2696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4626 vdd d0 a_4079_n4044# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4627 a_26095_7699# a_25674_7699# a_25359_7904# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4628 vdd d0 a_19168_n2438# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4629 a_20834_2697# a_20621_2697# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4630 a_16598_8544# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4631 a_11823_6889# a_11402_6889# a_10885_7133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4632 a_27815_n10678# a_28065_n5986# a_28020_n5782# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4633 a_13858_n4399# a_13854_n4587# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4634 a_10147_9220# a_10147_8990# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4635 a_1805_n3519# a_1514_n2580# a_1794_n3172# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4636 a_35389_9012# a_35917_8807# a_36125_8807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4637 a_11615_n7589# a_11402_n7589# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4638 a_7828_n8201# a_7847_n7127# a_7798_n7111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4639 a_10465_n2867# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4640 vdd d0 a_24264_5502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4641 a_1373_n4275# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4642 a_23074_3553# a_23327_3540# a_22929_4322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4643 vdd a_14108_6629# a_13900_6629# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4644 a_12913_7063# a_13900_6629# a_13851_6819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4645 gnd d0 a_24266_n3476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4646 a_17969_n8730# a_18956_n8502# a_18907_n8486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4647 a_18915_n2234# a_18911_n2422# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4648 gnd d0 a_14112_n2397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4649 a_35708_n3443# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4650 a_10677_4373# a_10464_4373# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4651 a_17976_n1924# a_18960_n2438# a_18911_n2422# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4652 a_28018_n7994# a_28032_n9314# a_27987_n9110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4653 a_32011_3561# a_31590_3561# a_31072_3251# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4654 a_6847_9131# a_6426_9131# a_5908_8821# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4655 vdd d0 a_29321_n6826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4656 a_35390_n9054# a_35917_n9507# a_36125_n9507# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4657 a_433_8231# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4658 a_23068_7039# a_24055_6605# a_24010_6618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4659 gnd a_4080_n1838# a_3872_n1838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4660 a_35391_n6432# a_35391_n6202# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4661 a_3824_9397# a_3820_9574# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4662 vdd d1 a_33356_n8686# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4663 a_8881_n6087# a_8877_n6275# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4664 gnd d6 a_4936_n10733# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4665 a_26825_n9812# a_26612_n9812# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4666 a_1514_1880# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4667 a_15519_n10080# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4668 a_25675_n5090# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4669 a_39097_6664# a_39093_6841# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4670 a_38158_n9626# a_39142_n10140# a_35389_n10157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4671 vdd a_19164_9430# a_18956_9430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4672 a_37081_5354# a_36754_7435# a_37076_7435# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4673 a_21039_n7255# a_20618_n7255# a_20304_n6802# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4674 a_31072_n3951# a_30651_n3951# a_30336_n3955# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4675 gnd d0 a_24266_2747# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4676 a_34037_7903# a_34042_7177# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4677 vdd d0 a_34298_1649# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4678 a_20303_n9008# a_20303_n8821# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4679 a_25676_n5644# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4680 a_6849_n5419# a_6428_n5419# a_5911_n5663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4681 a_1795_n2069# a_1374_n2069# a_856_n1759# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4682 vdd d2 a_23184_n9273# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4683 vdd a_18229_1399# a_18021_1399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4684 a_27036_2494# a_26615_2494# a_26098_2738# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4685 a_13854_8848# a_13850_9025# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4686 a_15733_7174# a_15520_7174# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4687 a_5700_8821# a_5487_8821# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4688 a_21980_n3153# a_21559_n3153# a_21042_n3397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4689 a_33100_5941# a_34087_5507# a_34038_5697# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4690 a_8877_5752# a_8882_5026# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4691 a_22932_6351# a_23185_6338# a_22958_7618# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4692 a_34042_n8792# a_34295_n8996# a_33103_n8482# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4693 a_13857_n5502# a_14110_n5706# a_12918_n5192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4694 a_10463_9339# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4695 a_27985_4363# a_28242_4173# a_28020_3070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4696 gnd a_39350_7754# a_39142_7754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4697 a_23068_8142# a_23325_7952# a_22927_8734# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4698 a_8881_5575# a_9134_5562# a_7939_5996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4699 a_11615_7992# a_11402_7992# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4700 vdd a_38412_7998# a_38204_7998# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4701 a_6782_4127# a_6569_4127# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4702 a_26096_n7850# a_26826_n7606# a_27034_n7606# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4703 a_31589_n5364# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4704 a_38161_n3008# a_39145_n3522# a_39096_n3506# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4705 a_23074_n2962# a_24058_n3476# a_24013_n3272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4706 a_7943_4716# a_8927_5013# a_8882_5026# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4707 a_10148_7014# a_10148_6784# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4708 vdd d0 a_4079_2212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4709 a_35390_7452# a_35918_7704# a_36126_7704# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4710 a_3827_3882# a_4080_3869# a_2888_3572# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4711 vdd a_29319_n7375# a_29111_n7375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4712 a_26097_3287# a_25676_3287# a_25361_3492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4713 a_116_8985# a_644_8780# a_852_8780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4714 a_2004_500# a_2823_5235# a_2778_5248# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4715 a_1808_n8108# a_1511_n9198# a_1791_n9790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4716 a_20305_4097# a_20305_3910# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4717 a_646_n5068# a_433_n5068# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4718 vdd d0 a_24266_1090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4719 gnd d0 a_19165_7224# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4720 a_29067_n7725# a_29320_n7929# a_28128_n7415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4721 vdd a_14110_2217# a_13902_2217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4722 gnd d0 a_4078_8281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4723 a_17830_4387# a_18020_3605# a_17971_3795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4724 a_31913_n3682# a_31700_n3682# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4725 a_12913_n7586# a_13900_n7358# a_13855_n7154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4726 a_12915_2651# a_13902_2217# a_13853_2407# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4727 a_3823_n1822# a_4080_n1838# a_2885_n2066# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4728 gnd a_9136_n3536# a_8928_n3536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4729 a_24012_4966# a_24008_5143# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4730 a_21557_n7565# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4731 vdd d1 a_3138_9074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4732 a_22962_7441# a_22976_8544# a_22927_8734# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4733 a_11841_n3701# a_11544_n4791# a_11824_n5383# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4734 a_39095_n2952# a_39101_n2215# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4735 a_35707_3292# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4736 a_8877_n5172# a_9134_n5188# a_7939_n5416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4737 a_17861_n3794# a_17880_n2720# a_17835_n2516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4738 a_34037_6800# a_34294_6610# a_33099_7044# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4739 a_21040_4349# a_20619_4349# a_20304_4554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4740 gnd a_13062_n5969# a_12854_n5969# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4741 a_23074_n2962# a_23327_n3166# a_22934_n2451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4742 a_23070_2627# a_24057_2193# a_24012_2206# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4743 a_8875_9061# a_8881_8335# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4744 vdd a_39352_n5728# a_39144_n5728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4745 a_25358_9466# a_25887_9356# a_26095_9356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4746 gnd d2 a_38272_6384# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4747 a_30862_n10020# a_30649_n10020# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4748 a_39095_n2952# a_39352_n2968# a_38157_n3196# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4749 a_20618_n10015# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4750 vdd a_19166_5018# a_18958_5018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4751 a_26723_5230# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4752 a_35918_n8404# a_35705_n8404# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4753 a_21978_n8668# a_21557_n8668# a_21040_n8912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4754 a_5908_n9521# a_6639_n9831# a_6847_n9831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4755 vdd d0 a_14107_8835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4756 gnd a_13170_n7602# a_12962_n7602# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4757 a_5172_n9755# a_5701_n10075# a_5909_n10075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4758 vdd d0 a_9134_n6291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4759 a_37076_5235# a_36756_3023# a_37078_3023# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4760 a_7943_4716# a_8196_4703# a_7803_4205# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4761 a_10884_n10039# a_10463_n10039# a_10147_n9948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4762 a_5176_n2263# a_5705_n2354# a_5913_n2354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4763 a_6958_5249# a_6537_5249# a_6859_5249# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4764 a_10680_n2318# a_10467_n2318# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4765 a_13855_6642# a_13851_6819# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4766 a_2887_5778# a_3871_6075# a_3822_6265# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4767 a_15734_6071# a_15521_6071# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4768 a_10467_1618# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4769 a_25888_5493# a_25675_5493# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4770 vdd a_13062_5240# a_12854_5240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4771 vdd d0 a_39352_n4071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4772 a_119_n4428# a_119_n4199# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4773 a_856_1059# a_1587_1369# a_1795_1369# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4774 a_434_n5622# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4775 a_1512_n6992# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4776 a_33102_1529# a_34089_1095# a_34040_1285# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4777 a_15941_5517# a_15520_5517# a_15205_5265# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4778 gnd d0 a_29320_5543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4779 vdd a_38273_4178# a_38065_4178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4780 a_10677_n5073# a_10464_n5073# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4781 a_2748_n2470# a_2933_n3185# a_2888_n2981# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4782 a_22934_1939# a_23187_1926# a_22960_3206# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4783 a_10465_4927# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4784 a_1585_n6481# a_1372_n6481# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4785 a_5489_n5109# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4786 a_21882_2977# a_21669_2977# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4787 vdd a_33356_7957# a_33148_7957# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4788 a_30336_2812# a_30865_2702# a_31073_2702# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4789 a_30650_8217# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4790 a_23070_3730# a_23327_3540# a_22929_4322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4791 a_8883_1163# a_9136_1150# a_7941_1584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4792 gnd d1 a_13169_9079# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4793 a_11617_3580# a_11404_3580# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4794 a_6750_n5949# a_6537_n5949# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4795 gnd d1 a_18228_n3231# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4796 gnd a_28383_n4310# a_28175_n4310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4797 vdd d1 a_18228_3605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4798 a_35392_3040# a_35920_3292# a_36128_3292# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4799 a_28124_7080# a_29111_6646# a_29062_6836# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4800 a_10464_n8936# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4801 a_648_n4519# a_435_n4519# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4802 a_25360_6344# a_25360_6157# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4803 a_35171_466# a_36955_527# a_37277_527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4804 a_5173_6820# a_5174_6363# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4805 gnd d0 a_19167_2812# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4806 a_852_8780# a_431_8780# a_116_8985# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4807 gnd a_29320_8303# a_29112_8303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4808 a_34040_n3465# a_34297_n3481# a_33105_n2967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4809 a_26827_5803# a_26614_5803# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4810 a_16458_6930# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4811 a_8879_n4623# a_9136_n4639# a_7944_n4125# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4812 a_25890_1081# a_25677_1081# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4813 gnd d2 a_13031_n4885# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4814 a_18906_9066# a_18912_8340# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4815 a_22964_3029# a_22978_4132# a_22929_4322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4816 a_27037_n2091# a_26969_n2602# a_27047_n3541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4817 a_39096_4086# a_39353_3896# a_38161_3599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4818 a_34040_2942# a_34043_2211# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4819 a_25359_8134# a_25888_8253# a_26096_8253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4820 a_18906_n9589# a_18912_n8852# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4821 a_31074_n2299# a_31804_n2055# a_32012_n2055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4822 a_6864_5368# a_6537_7449# a_6864_7568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4823 a_22929_n4845# a_23119_n4269# a_23074_n4065# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4824 a_34039_2388# a_34296_2198# a_33101_2632# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4825 a_12913_n7586# a_13170_n7602# a_12777_n6887# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4826 vdd a_24264_n7888# a_24056_n7888# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4827 gnd d2 a_38274_1972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4828 a_26825_9112# a_26612_9112# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4829 a_17969_8207# a_18226_8017# a_17828_8799# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4830 gnd d1 a_33357_5751# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4831 a_36127_5498# a_36858_5808# a_37066_5808# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4832 a_15942_n2908# a_16673_n3218# a_16881_n3218# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4833 vdd a_34297_n1824# a_34089_n1824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4834 vdd a_39350_7754# a_39142_7754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4835 a_3824_7740# a_4077_7727# a_2882_8161# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4836 vdd d1 a_13170_n8705# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4837 a_8877_5752# a_9134_5562# a_7939_5996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4838 a_20621_1040# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4839 a_37067_n3199# a_36646_n3199# a_36129_n3443# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4840 gnd a_13060_n8181# a_12852_n8181# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4841 a_21041_6006# a_21771_5762# a_21979_5762# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4842 a_35392_n3539# a_35392_n3352# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4843 a_1808_n5908# a_1481_n8108# a_1808_n8108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4844 a_24007_7349# a_24264_7159# a_23072_6862# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4845 a_35919_5498# a_35706_5498# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4846 vdd d0 a_29318_n9581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4847 a_25360_n5553# a_25889_n5644# a_26097_n5644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4848 a_26097_n2884# a_25676_n2884# a_25362_n2431# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4849 a_647_6025# a_434_6025# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4850 vdd a_23328_n2063# a_23120_n2063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4851 gnd d0 a_29322_1131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4852 a_15943_1105# a_15522_1105# a_15209_1211# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4853 a_10148_n8386# a_10148_n7929# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4854 vdd a_28383_2478# a_28175_2478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4855 vdd a_38413_n6521# a_38205_n6521# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4856 a_21989_n5712# a_21880_n5889# a_22088_n5889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4857 a_12920_n1883# a_13904_n2397# a_13855_n2381# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4858 a_21038_8761# a_21769_9071# a_21977_9071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4859 vdd d0 a_19165_7224# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4860 a_30334_n9013# a_30861_n9466# a_31069_n9466# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4861 a_26723_n5930# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4862 a_7801_8617# a_7986_9115# a_7937_9305# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4863 vdd d0 a_4078_8281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4864 a_29067_4453# a_29063_4630# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4865 a_31074_1599# a_30653_1599# a_30337_1480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4866 a_119_2367# a_120_1910# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4867 a_35704_n9507# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4868 a_26098_n3438# a_25677_n3438# a_25361_n3347# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4869 gnd d0 a_9135_n5742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4870 a_30336_n3082# a_30865_n3402# a_31073_n3402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4871 a_20831_7658# a_20618_7658# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4872 a_21769_n9771# a_21556_n9771# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4873 a_10462_8785# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4874 a_12703_n10661# a_12653_n10677# a_11933_n5913# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4875 a_8883_2820# a_9136_2807# a_7944_2510# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4876 a_39097_6664# a_39350_6651# a_38155_7085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4877 a_22962_7441# a_22976_8544# a_22931_8557# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4878 a_15204_n7554# a_15733_n7874# a_15941_n7874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4879 a_28126_2668# a_29113_2234# a_29064_2424# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4880 a_7938_8202# a_8925_7768# a_8880_7781# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4881 a_27050_5349# a_26723_7430# a_27050_7549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4882 vdd d2 a_38272_6384# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4883 a_854_4368# a_433_4368# a_118_4573# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4884 a_11543_n6997# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4885 a_33099_n7567# a_34086_n7339# a_34041_n7135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4886 a_5908_n9521# a_5487_n9521# a_5173_n9068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4887 gnd a_3138_9074# a_2930_9074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4888 a_2887_5778# a_3871_6075# a_3826_6088# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4889 a_37081_n5935# a_36754_n8135# a_37076_n7958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4890 a_646_n7828# a_433_n7828# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4891 vdd d1 a_8197_n4329# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4892 a_1372_5781# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4893 a_39094_n9021# a_39351_n9037# a_38159_n8523# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4894 a_22088_n5889# a_23016_n10653# a_22858_n10637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4895 a_37068_n2096# a_36647_n2096# a_36129_n1786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4896 a_21040_n7809# a_21770_n7565# a_21978_n7565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4897 a_17833_n6928# a_18018_n7643# a_17973_n7439# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4898 vdd d1 a_38415_n2109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4899 vdd a_18116_7493# a_17908_7493# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4900 a_26613_n7606# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4901 vdd d0 a_29320_5543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4902 a_36129_1086# a_36860_1396# a_37068_1396# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4903 a_10150_3475# a_10150_3018# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4904 a_12803_n8165# a_13060_n8181# a_12809_n5765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4905 a_16897_n3742# a_16600_n4832# a_16881_n4321# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4906 a_13854_n9360# a_13850_n9548# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4907 a_29066_n2398# a_29323_n2414# a_28131_n1900# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4908 a_3826_3328# a_4079_3315# a_2884_3749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4909 vdd a_4077_n7353# a_3869_n7353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4910 a_8879_1340# a_9136_1150# a_7941_1584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4911 a_854_n6171# a_433_n6171# a_118_n5718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4912 a_31070_9320# a_30649_9320# a_30333_9201# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4913 a_33101_n4258# a_33358_n4274# a_32960_n4850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4914 a_21043_1594# a_21773_1350# a_21981_1350# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4915 a_24005_9001# a_24011_8275# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4916 a_16814_n2626# a_16601_n2626# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4917 a_10148_8533# a_10675_8785# a_10883_8785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4918 a_18909_n4074# a_19166_n4090# a_17971_n4318# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4919 a_30335_n5517# a_30335_n5288# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4920 gnd a_19163_n9605# a_18955_n9605# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4921 a_20621_2697# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4922 a_28124_7080# a_29111_6646# a_29066_6659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4923 a_13856_n8811# a_13852_n8999# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4924 a_26094_n9502# a_25673_n9502# a_25359_n9049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4925 vdd a_23325_n8681# a_23117_n8681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4926 a_30334_n8597# a_30863_n8917# a_31071_n8917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4927 a_34043_n2723# a_34039_n2911# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4928 vdd a_24264_5502# a_24056_5502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4929 vdd a_14110_n2946# a_13902_n2946# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4930 a_3822_5162# a_3825_4431# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4931 a_34043_2211# a_34039_2388# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4932 gnd d0 a_29322_2788# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4933 a_18913_n6646# a_18909_n6834# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4934 a_15203_9490# a_15732_9380# a_15940_9380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4935 a_6641_n6522# a_6428_n6522# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4936 a_20833_3246# a_20620_3246# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4937 a_10464_4373# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4938 a_21977_n9771# a_21910_n9179# a_21994_n8089# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4939 a_21667_5189# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4940 a_2772_7637# a_2791_6357# a_2746_6370# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4941 a_22964_3029# a_22978_4132# a_22933_4145# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4942 a_1793_n5378# a_1372_n5378# a_854_n5068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4943 a_7939_n6519# a_8926_n6291# a_8881_n6087# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4944 a_30866_n2299# a_30653_n2299# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4945 a_5492_n2354# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4946 a_20303_7219# a_20832_7109# a_21040_7109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4947 vdd d6 a_35153_n10719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4948 a_27988_6392# a_28241_6379# a_28014_7659# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4949 a_27045_5230# a_26725_3018# a_27052_3137# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4950 vdd d0 a_34296_n4030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4951 a_117_n7278# a_118_n6821# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4952 a_10886_n3970# a_11617_n4280# a_11825_n4280# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4953 vdd d1 a_33357_5751# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4954 a_6848_6925# a_6781_6333# a_6859_7449# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4955 a_25361_3951# a_25361_3722# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4956 a_32008_n9776# a_31587_n9776# a_31070_n10020# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4957 gnd a_24266_2747# a_24058_2747# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4958 a_28020_n3582# a_28273_n3786# a_28016_n5970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4959 a_20620_n2843# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4960 vdd a_34298_1649# a_34090_1649# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4961 a_10150_n4620# a_10677_n5073# a_10885_n5073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4962 a_7942_6922# a_8926_7219# a_8877_7409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4963 a_15520_n5114# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4964 a_15520_7174# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4965 a_29067_7213# a_29320_7200# a_28128_6903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4966 gnd d1 a_8196_n6535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4967 a_35392_n3996# a_35392_n3539# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4968 a_37064_9117# a_36643_9117# a_36125_8807# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4969 a_32963_n6868# a_33216_n7072# a_32989_n8146# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4970 a_30336_2353# a_30337_1896# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4971 a_37065_n8714# a_36644_n8714# a_36126_n8404# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4972 a_20621_n3397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4973 a_2004_500# a_1895_500# a_2103_500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4974 gnd a_9136_n1879# a_8928_n1879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4975 a_21041_n3946# a_20620_n3946# a_20305_n3493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4976 a_11834_7413# a_11543_6297# a_11823_6889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4977 a_32963_6356# a_33148_6854# a_33103_6867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4978 vdd d1 a_38412_n8727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4979 gnd a_14109_4423# a_13901_4423# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4980 a_2884_n3169# a_3871_n2941# a_3822_n2925# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4981 vdd d0 a_29322_1131# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4982 a_25359_6801# a_25360_6344# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4983 a_15941_n6217# a_15520_n6217# a_15205_n6221# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4984 a_5909_7718# a_5488_7718# a_5173_7466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4985 a_11402_7992# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4986 a_7801_8617# a_7986_9115# a_7941_9128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4987 a_28125_n6500# a_29112_n6272# a_29067_n6068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4988 a_21042_n4500# a_20621_n4500# a_20305_n4409# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4989 a_31069_8766# a_30648_8766# a_30333_8971# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4990 a_21911_n6973# a_21698_n6973# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4991 a_20834_n1740# a_20621_n1740# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4992 a_5174_n6862# a_5174_n6675# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X4993 a_21039_9315# a_20618_9315# a_20302_9196# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4994 a_16811_n9244# a_16598_n9244# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4995 a_39093_6841# a_39350_6651# a_38155_7085# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4996 a_119_3929# a_648_3819# a_856_3819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4997 a_25888_n5090# a_25675_n5090# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X4998 gnd d1 a_3139_n7597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4999 a_28126_2668# a_29113_2234# a_29068_2247# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5000 a_6428_4719# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5001 a_5053_480# a_4632_480# a_2103_500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5002 a_1373_n4275# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5003 a_15942_n2908# a_15521_n2908# a_15207_n2455# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5004 vdd a_24266_1090# a_24058_1090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5005 gnd a_19165_7224# a_18957_7224# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5006 a_15944_1659# a_15523_1659# a_15207_1769# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5007 a_12809_n3565# a_12823_n4885# a_12774_n4869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5008 gnd a_4078_8281# a_3870_8281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5009 a_26756_n2602# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5010 a_20306_n2203# a_20835_n2294# a_21043_n2294# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5011 a_31591_n2055# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5012 gnd a_34295_n7893# a_34087_n7893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5013 a_117_7009# a_646_7128# a_854_7128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5014 a_15943_n3462# a_15522_n3462# a_15206_n3371# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5015 vdd a_18087_n4926# a_17879_n4926# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5016 vdd a_3138_9074# a_2930_9074# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5017 gnd a_28241_n7108# a_28033_n7108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5018 a_28130_n3003# a_29114_n3517# a_29069_n3313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5019 a_7804_n2511# a_8057_n2715# a_7830_n3789# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5020 a_35389_n9511# a_35917_n9507# a_36125_n9507# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5021 a_20304_5887# a_20833_6006# a_21041_6006# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5022 a_32964_n4662# a_33149_n5377# a_33104_n5173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5023 gnd a_38272_6384# a_38064_6384# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5024 a_38160_5805# a_39144_6102# a_39099_6115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5025 a_12772_n9281# a_12962_n8705# a_12917_n8501# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5026 a_26825_n9812# a_26612_n9812# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5027 a_3828_1676# a_3824_1853# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5028 a_27990_1980# a_28243_1967# a_28016_3247# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5029 a_23073_5759# a_23326_5746# a_22928_6528# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5030 vdd a_14107_8835# a_13899_8835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5031 a_10150_n4204# a_10679_n4524# a_10887_n4524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5032 a_31072_n3951# a_30651_n3951# a_30336_n3498# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5033 gnd a_4081_n2392# a_3873_n2392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5034 vdd d0 a_4076_n9559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5035 a_15521_6071# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5036 a_38158_n9626# a_38411_n9830# a_38018_n9115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5037 a_37065_8014# a_36644_8014# a_36127_8258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5038 a_25675_5493# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5039 a_3822_3505# a_4079_3315# a_2884_3749# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5040 a_7939_n6519# a_8196_n6535# a_7798_n7111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5041 a_25676_n5644# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5042 a_11825_2477# a_11404_2477# a_10887_2721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5043 a_117_n8840# a_117_n8611# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5044 a_10676_6579# a_10463_6579# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5045 a_24006_n7318# a_24012_n6581# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5046 a_21667_n5889# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5047 a_32010_5767# a_31589_5767# a_31071_5457# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5048 a_4845_480# a_4632_480# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5049 vdd a_3140_n5391# a_2932_n5391# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5050 gnd a_9133_n8497# a_8925_n8497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5051 a_11836_3001# a_11545_1885# a_11825_2477# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5052 vdd d1 a_28381_6890# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5053 a_25889_n3987# a_25676_n3987# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5054 a_7943_n5228# a_8927_n5742# a_8878_n5726# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5055 a_30652_n3402# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5056 a_17972_n2112# a_18229_n2128# a_17831_n2704# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5057 a_11404_3580# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5058 a_7944_n4125# a_8197_n4329# a_7799_n4905# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5059 a_20831_n8358# a_20618_n8358# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5060 a_11824_n5383# a_11403_n5383# a_10886_n5627# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5061 vdd d0 a_34297_3855# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5062 gnd a_648_n1759# a_856_n1759# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5063 a_27035_4700# a_26614_4700# a_26097_4944# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5064 vdd a_18228_3605# a_18020_3605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5065 a_39094_7395# a_39097_6664# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5066 a_39095_2429# a_39352_2239# a_38157_2673# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5067 a_119_n4615# a_119_n4428# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5068 a_5704_n4560# a_5491_n4560# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5069 a_36129_3846# a_35708_3846# a_35392_3727# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5070 gnd d1 a_38413_5792# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5071 gnd a_19167_2812# a_18959_2812# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5072 gnd d0 a_14108_6629# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5073 a_20305_n3306# a_20305_n3077# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5074 a_8880_7781# a_9133_7768# a_7938_8202# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5075 a_16989_n5954# a_16568_n5954# a_16895_n5954# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5076 a_20832_n5049# a_20619_n5049# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5077 a_26614_5803# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5078 a_36127_7155# a_35706_7155# a_35390_7265# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5079 a_21557_n7565# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5080 vdd d0 a_19165_5567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5081 a_28129_n5209# a_29113_n5723# a_29064_n5707# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5082 a_26098_n1781# a_25677_n1781# a_25362_n1785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5083 a_24010_9378# a_24263_9365# a_23071_9068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5084 a_3824_n2376# a_4081_n2392# a_2889_n1878# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5085 a_16599_6338# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5086 vdd a_19167_n3541# a_18959_n3541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5087 gnd a_38274_1972# a_38066_1972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5088 a_18909_3551# a_18914_2825# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5089 a_26612_9112# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5090 gnd a_28382_4684# a_28174_4684# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5091 gnd a_33357_5751# a_33149_5751# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5092 vdd d2 a_3001_n2674# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5093 a_5909_n10075# a_6639_n9831# a_6847_n9831# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5094 a_11758_n2585# a_11545_n2585# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5095 a_1895_500# a_1682_500# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5096 a_23075_1347# a_23328_1334# a_22930_2116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5097 vdd d0 a_24265_3296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5098 a_856_n3416# a_435_n3416# a_119_n3325# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5099 vdd a_14109_4423# a_13901_4423# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5100 a_10148_7243# a_10148_7014# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5101 a_3825_n6046# a_4078_n6250# a_2883_n6478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5102 a_39096_n3506# a_39353_n3522# a_38161_n3008# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5103 a_10677_5476# a_10464_5476# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5104 a_25677_1081# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5105 gnd d3 a_33246_7433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5106 a_27045_7430# a_26754_6314# a_27034_6906# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5107 a_5053_480# a_9779_364# a_9987_364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5108 a_10678_2167# a_10465_2167# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5109 a_1694_5208# a_1481_5208# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5110 a_35390_n7951# a_35390_n7764# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5111 a_35706_5498# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5112 a_32012_1355# a_31591_1355# a_31073_1045# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5113 a_34036_9006# a_34293_8816# a_33098_9250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5114 a_434_6025# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5115 vdd d0 a_39353_n4625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5116 gnd a_29322_1131# a_29114_1131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5117 a_5175_n4240# a_5175_n4010# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5118 a_35918_9361# a_35705_9361# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5119 vdd a_33355_n9789# a_33147_n9789# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5120 a_16879_n7630# a_16458_n7630# a_15940_n7320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5121 vdd d0 a_24263_n7334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5122 a_21697_n9179# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5123 vdd a_19165_7224# a_18957_7224# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5124 gnd d0 a_14111_n1843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5125 vdd a_4078_8281# a_3870_8281# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5126 a_15203_n9989# a_15203_n9760# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5127 a_15204_8574# a_15204_8387# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5128 vdd a_33248_n3750# a_33040_n3750# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5129 vdd a_28072_n10694# a_27864_n10694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5130 a_15733_8277# a_15520_8277# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5131 a_25887_7699# a_25674_7699# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5132 a_17833_6416# a_18086_6403# a_17859_7683# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5133 a_8878_n5726# a_8881_n4984# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5134 a_117_n7924# a_645_n8377# a_853_n8377# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5135 a_5701_6615# a_5488_6615# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5136 gnd d0 a_39354_n2419# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5137 gnd a_28381_7993# a_28173_7993# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5138 gnd d0 a_24264_n5128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5139 a_13854_n1827# a_14830_n1530# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5140 a_17974_5824# a_18227_5811# a_17829_6593# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5141 gnd d0 a_29319_7749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5142 a_6851_n2110# a_6430_n2110# a_5913_n2354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5143 a_13852_7373# a_13855_6642# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5144 vdd a_38272_6384# a_38064_6384# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5145 a_30649_n8363# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5146 a_28131_n1900# a_28384_n2104# a_27986_n2680# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5147 gnd d1 a_38415_1380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5148 a_10464_n5073# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5149 a_15519_6620# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5150 a_11834_5213# a_11725_5213# a_11933_5213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5151 a_30335_5018# a_30864_4908# a_31072_4908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5152 a_15207_1310# a_15209_1211# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5153 gnd a_39351_5548# a_39143_5548# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5154 a_23069_5936# a_23326_5746# a_22928_6528# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5155 a_8882_3369# a_9135_3356# a_7940_3790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5156 a_11616_5786# a_11403_5786# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5157 a_25888_n7850# a_25675_n7850# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5158 a_118_n5072# a_646_n5068# a_854_n5068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5159 a_27036_n3194# a_26969_n2602# a_27047_n3541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5160 a_24012_4966# a_24265_4953# a_23073_4656# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5161 a_10885_n6176# a_10464_n6176# a_10149_n6180# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5162 a_852_n9480# a_431_n9480# a_117_n9027# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5163 a_35391_5246# a_35919_5498# a_36127_5498# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5164 vdd a_23187_n2655# a_22979_n2655# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5165 a_7802_n6923# a_7987_n7638# a_7942_n7434# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5166 a_38021_1985# a_38206_2483# a_38157_2673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5167 a_5488_9375# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5168 gnd d0 a_34293_8816# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5169 a_36967_7435# a_36754_7435# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5170 a_117_6779# a_645_6574# a_853_6574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5171 a_24865_n10698# a_27864_n10694# a_27815_n10678# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5172 a_20303_8093# a_20303_7863# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5173 a_5490_n5663# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5174 gnd a_14109_n9015# a_13901_n9015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5175 gnd d0 a_19166_5018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5176 a_17831_2181# a_18021_1399# a_17972_1589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5177 a_24008_n5666# a_24265_n5682# a_23073_n5168# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5178 a_20304_5657# a_20832_5452# a_21040_5452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5179 a_35016_n1511# a_35921_n1786# a_36129_n1786# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5180 a_10679_1064# a_10466_1064# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5181 a_38155_n7608# a_39142_n7380# a_39097_n7176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5182 a_16881_n4321# a_16813_n4832# a_16897_n3742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5183 gnd d3 a_18118_n3810# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5184 gnd d3 a_33248_3021# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5185 a_2746_n6882# a_2931_n7597# a_2882_n7581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5186 a_3824_n2376# a_3827_n1634# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5187 a_27047_3018# a_26756_1902# a_27036_2494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5188 a_853_9334# a_1583_9090# a_1791_9090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5189 a_32991_3211# a_33010_1931# a_32961_2121# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5190 a_5911_n6766# a_5490_n6766# a_5174_n6675# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5191 a_2776_7460# a_2790_8563# a_2741_8753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5192 a_22958_7618# a_22977_6338# a_22928_6528# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5193 a_35708_1086# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5194 a_34038_4594# a_34295_4404# a_33100_4838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5195 a_25677_2738# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5196 vdd d0 a_24265_n6785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5197 a_7939_5996# a_8926_5562# a_8877_5752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5198 gnd d2 a_38273_4178# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5199 a_30334_8327# a_30863_8217# a_31071_8217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5200 a_30333_n9470# a_30861_n9466# a_31069_n9466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5201 a_15205_4619# a_15206_4162# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5202 a_20834_3800# a_20621_3800# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5203 a_35704_n9507# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5204 gnd a_29322_2788# a_29114_2788# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5205 vdd d0 a_34294_n7339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5206 vdd a_9133_n7394# a_8925_n7394# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5207 a_7944_2510# a_8197_2497# a_7804_1999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5208 a_2888_3572# a_3872_3869# a_3823_4059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5209 a_30336_n3311# a_30865_n3402# a_31073_n3402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5210 a_21769_n9771# a_21556_n9771# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5211 a_25889_3287# a_25676_3287# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5212 a_5702_5512# a_5489_5512# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5213 a_38157_n4299# a_38414_n4315# a_38016_n4891# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5214 a_17835_2004# a_18088_1991# a_17861_3271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5215 a_20620_3246# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5216 a_21040_8212# a_21770_7968# a_21978_7968# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5217 a_15204_n7783# a_15733_n7874# a_15941_n7874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5218 a_6859_n7972# a_6568_n7033# a_6848_n7625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5219 vdd a_18118_n6010# a_17910_n6010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5220 gnd d0 a_39351_n9037# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5221 a_5703_2203# a_5490_2203# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5222 a_24006_9555# a_24263_9365# a_23071_9068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5223 a_10466_n4524# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5224 vdd d2 a_38274_n2701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5225 vdd d0 a_19166_n5747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5226 a_2881_n9787# a_3868_n9559# a_3823_n9355# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5227 a_30336_3686# a_30865_3805# a_31073_3805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5228 gnd d0 a_29321_3337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5229 vdd a_28382_4684# a_28174_4684# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5230 a_1371_n7584# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5231 vdd a_33357_5751# a_33149_5751# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5232 a_2884_3749# a_3141_3559# a_2743_4341# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5233 a_23071_1524# a_23328_1334# a_22930_2116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5234 a_11618_1374# a_11405_1374# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5235 a_2888_n2981# a_3141_n3185# a_2748_n2470# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5236 a_20304_5200# a_20304_5013# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5237 a_22927_8734# a_23117_7952# a_23068_8142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5238 vdd d3 a_33246_7433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5239 a_27033_n9812# a_26966_n9220# a_27050_n8130# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5240 a_16897_3161# a_16600_4132# a_16881_3621# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5241 a_5489_8272# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5242 a_118_5219# a_646_5471# a_854_5471# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5243 a_1792_n8687# a_1371_n8687# a_854_n8931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5244 a_10150_n4433# a_10150_n4204# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5245 gnd d0 a_19166_n4090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5246 a_35395_1192# a_35921_1086# a_36129_1086# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5247 vdd a_23184_n9273# a_22976_n9273# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5248 a_36969_3023# a_36756_3023# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5249 a_119_2367# a_647_2162# a_855_2162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5250 a_7803_4205# a_7988_4703# a_7939_4893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5251 vdd a_29322_1131# a_29114_1131# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5252 a_27045_n7953# a_26754_n7014# a_27034_n7606# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5253 a_35391_n5329# a_35391_n5099# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5254 gnd a_29321_6097# a_29113_6097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5255 vdd a_14109_n6255# a_13901_n6255# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5256 a_35919_n5095# a_35706_n5095# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5257 a_8881_n4984# a_8877_n5172# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5258 vdd d0 a_9135_n2982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5259 a_23067_n9768# a_24054_n9540# a_24009_n9336# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5260 a_20305_n3493# a_20833_n3946# a_21041_n3946# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5261 a_31728_8484# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5262 a_27990_n2492# a_28175_n3207# a_28126_n3191# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5263 a_6641_5822# a_6428_5822# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5264 a_16459_4724# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5265 a_16814_n2626# a_16601_n2626# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5266 a_28130_2491# a_29114_2788# a_29069_2801# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5267 a_34037_6800# a_34043_6074# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5268 a_2778_3048# a_2792_4151# a_2743_4341# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5269 a_21039_n10015# a_20618_n10015# a_20302_n9924# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5270 a_22960_3206# a_22979_1926# a_22930_2116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5271 gnd d4 a_8087_5276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5272 a_25360_5928# a_25889_6047# a_26097_6047# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5273 a_853_6574# a_1584_6884# a_1792_6884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5274 a_21989_n7912# a_21698_n6973# a_21978_n7565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5275 a_30334_n8826# a_30863_n8917# a_31071_n8917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5276 a_7941_1584# a_8928_1150# a_8879_1340# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5277 a_26826_6906# a_26613_6906# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5278 a_39097_9424# a_39093_9601# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5279 a_29752_345# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5280 gnd d1 a_33358_3545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5281 a_8877_4649# a_8883_3923# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5282 vdd a_9135_n6845# a_8927_n6845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5283 vdd d1 a_38415_1380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5284 a_23069_n6459# a_23326_n6475# a_22928_n7051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5285 vdd a_14111_n3500# a_13903_n3500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5286 a_8878_3546# a_9135_3356# a_7940_3790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5287 a_38162_1393# a_39146_1690# a_39097_1880# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5288 a_21996_3096# a_21699_4067# a_21980_3556# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5289 a_35389_n10157# a_39350_n10140# a_38158_n9626# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5290 a_21042_3800# a_21772_3556# a_21980_3556# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5291 gnd a_3031_5235# a_2823_5235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5292 vdd d2 a_38271_n9319# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5293 a_18915_n2234# a_19168_n2438# a_17976_n1924# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5294 a_24818_461# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5295 a_32964_4150# a_33149_4648# a_33100_4838# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5296 a_38021_1985# a_38206_2483# a_38161_2496# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5297 vdd a_33359_1339# a_33151_1339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5298 a_32008_n9776# a_31587_n9776# a_31069_n9466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5299 gnd d2 a_18088_n2720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5300 a_20305_2994# a_20305_2807# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5301 a_28128_6903# a_28381_6890# a_27988_6392# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5302 a_17970_n5421# a_18227_n5437# a_17834_n4722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5303 a_22962_7441# a_23215_7428# a_22964_5229# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5304 gnd d1 a_8195_6909# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5305 a_32961_n2644# a_33151_n2068# a_33106_n1864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5306 vdd d3 a_33248_3021# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5307 a_6537_n8149# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5308 a_37076_n5758# a_36756_n3723# a_37083_n3723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5309 a_34040_n3465# a_34043_n2723# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5310 a_10463_6579# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5311 a_39098_4458# a_39351_4445# a_38156_4879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5312 a_2776_7460# a_2790_8563# a_2745_8576# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5313 a_15206_n4015# a_15734_n4011# a_15942_n4011# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5314 a_12916_n2071# a_13903_n1843# a_13854_n1827# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5315 a_38020_n4703# a_38205_n5418# a_38160_n5214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5316 a_2882_8161# a_3869_7727# a_3820_7917# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5317 a_35390_7909# a_35390_7452# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5318 a_21041_n2843# a_21772_n3153# a_21980_n3153# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5319 a_7939_5996# a_8926_5562# a_8881_5575# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5320 vdd d1 a_18227_n6540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5321 gnd a_17917_n10718# a_17709_n10718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5322 a_21039_n10015# a_20618_n10015# a_20302_n9695# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5323 a_15941_n6217# a_15520_n6217# a_15205_n5764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5324 a_21911_6273# a_21698_6273# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5325 a_15206_n4245# a_15735_n4565# a_15943_n4565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5326 a_21979_5762# a_21558_5762# a_21040_5452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5327 gnd d0 a_34298_n2378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5328 a_6847_9131# a_6780_8539# a_6864_7568# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5329 vdd d0 a_9132_n9600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5330 a_15941_8277# a_16671_8033# a_16879_8033# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5331 a_2888_n2981# a_3872_n3495# a_3823_n3479# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5332 a_6643_1410# a_6430_1410# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5333 a_21994_5308# a_21880_5189# a_22088_5189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5334 vdd a_3142_n2082# a_2934_n2082# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5335 vdd a_34297_3855# a_34089_3855# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5336 gnd d0 a_19164_7773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5337 gnd a_3139_6868# a_2931_6868# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5338 a_12773_n7075# a_13030_n7091# a_12803_n8165# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5339 a_16811_n9244# a_16598_n9244# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5340 vdd a_8196_n5432# a_7988_n5432# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5341 a_21977_9071# a_21556_9071# a_21039_9315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5342 a_117_n9027# a_117_n8840# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5343 a_37066_n6508# a_36998_n7019# a_37076_n7958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5344 a_3821_n5131# a_3827_n4394# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5345 a_30866_1599# a_30653_1599# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5346 gnd a_38413_5792# a_38205_5792# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5347 a_1794_n3172# a_1727_n2580# a_1805_n3519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5348 gnd a_14108_6629# a_13900_6629# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5349 a_34036_n9529# a_34293_n9545# a_33098_n9773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5350 a_26756_n2602# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5351 a_21868_481# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5352 a_35391_5059# a_35391_4830# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5353 a_7944_2510# a_8928_2807# a_8879_2997# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5354 a_13855_9402# a_13851_9579# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5355 a_15943_n3462# a_15522_n3462# a_15206_n3142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5356 a_10884_9339# a_11614_9095# a_11822_9095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5357 a_30336_4102# a_30336_3915# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5358 gnd d3 a_38302_7474# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5359 a_31071_7114# a_30650_7114# a_30334_6995# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5360 vdd a_19165_5567# a_18957_5567# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5361 a_13851_n7342# a_14108_n7358# a_12913_n7586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5362 a_26936_7430# a_26723_7430# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5363 a_6750_5249# a_6537_5249# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5364 a_646_n7828# a_433_n7828# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5365 a_5704_2757# a_5491_2757# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5366 a_17831_n2704# a_18088_n2720# a_17861_n3794# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5367 a_21994_n8089# a_21880_n8089# a_21994_n5889# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5368 a_35708_n1786# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5369 vdd d0 a_14108_n8461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5370 vdd a_24265_3296# a_24057_3296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5371 a_16568_5254# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5372 a_10150_n4433# a_10679_n4524# a_10887_n4524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5373 a_3819_9020# a_3825_8294# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5374 gnd d2 a_18085_n9338# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5375 a_23074_n4065# a_24058_n4579# a_24009_n4563# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5376 a_36128_n6752# a_36858_n6508# a_37066_n6508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5377 a_10679_2721# a_10466_2721# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5378 a_10464_5476# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5379 gnd d0 a_34298_1649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5380 gnd a_33246_7433# a_33038_7433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5381 a_15204_7284# a_15733_7174# a_15941_7174# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5382 a_8877_n7932# a_9134_n7948# a_7942_n7434# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5383 a_5172_9026# a_5700_8821# a_5908_8821# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5384 a_22964_3029# a_23217_3016# a_22960_5406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5385 a_28016_5447# a_28273_5257# a_27246_522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5386 a_37000_1907# a_36787_1907# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5387 a_10465_2167# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5388 a_1481_5208# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5389 a_35171_466# a_35062_466# a_30074_345# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5390 a_2778_3048# a_2792_4151# a_2747_4164# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5391 a_22932_n6863# a_23117_n7578# a_23072_n7374# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5392 vdd d4 a_8087_5276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5393 a_38019_n6909# a_38204_n7624# a_38155_n7608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5394 a_12913_n8689# a_13900_n8461# a_13851_n8445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5395 a_37067_n4302# a_36646_n4302# a_36129_n4546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5396 a_6427_n8728# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5397 a_17091_546# a_16982_546# a_14985_485# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5398 a_7941_1584# a_8928_1150# a_8883_1163# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5399 a_5173_n8652# a_5173_n8422# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5400 vdd d0 a_9134_n9051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5401 a_30652_n3402# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5402 a_35705_9361# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5403 a_30862_9320# a_30649_9320# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5404 vdd a_34295_n5133# a_34087_n5133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5405 vdd d1 a_33358_3545# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5406 a_10883_8785# a_10462_8785# a_10147_8990# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5407 a_6849_4719# a_6782_4127# a_6866_3156# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5408 a_8881_n6087# a_9134_n6291# a_7939_n6519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5409 gnd d5 a_23016_n10653# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5410 a_15520_8277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5411 a_25674_7699# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5412 a_854_n7828# a_1584_n7584# a_1792_n7584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5413 a_17974_n5233# a_18958_n5747# a_18913_n5543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5414 a_21913_n2561# a_21700_n2561# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5415 gnd d0 a_19166_3361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5416 a_10148_7430# a_10148_7243# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5417 gnd a_33248_n5950# a_33040_n5950# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5418 a_29068_5007# a_29321_4994# a_28129_4697# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5419 vdd a_3031_5235# a_2823_5235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5420 a_11617_n3177# a_11404_n3177# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5421 a_31588_6870# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5422 gnd a_34296_n2927# a_34088_n2927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5423 gnd a_38415_1380# a_38207_1380# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5424 a_31700_n3682# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5425 a_1791_n9790# a_1724_n9198# a_1808_n8108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5426 gnd a_14110_2217# a_13902_2217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5427 a_26753_n9220# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5428 a_16989_n5954# a_16568_n5954# a_16890_n5777# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5429 a_31072_6011# a_30651_6011# a_30335_6121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5430 a_10148_n7283# a_10149_n6826# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5431 a_11403_5786# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5432 a_25360_5698# a_25888_5493# a_26096_5493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5433 a_11403_n6486# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5434 a_30336_n4601# a_30336_n4414# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5435 a_17971_n4318# a_18958_n4090# a_18909_n4074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5436 vdd a_38304_n3791# a_38096_n3791# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5437 a_15732_n7320# a_15519_n7320# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5438 gnd d3 a_38304_3062# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5439 vdd a_28241_6379# a_28033_6379# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5440 a_39096_n3506# a_39099_n2764# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5441 a_7629_n10697# a_7879_n6005# a_7834_n5801# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5442 a_4778_n10717# a_4728_n10733# a_2672_n10656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5443 a_26938_3018# a_26725_3018# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5444 a_39094_4635# a_39351_4445# a_38156_4879# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5445 gnd a_34293_8816# a_34085_8816# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5446 a_36754_7435# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5447 a_6859_7449# a_6568_6333# a_6849_5822# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5448 gnd d0 a_29320_n5169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5449 a_17834_n4722# a_18087_n4926# a_17865_n3606# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5450 a_7940_n3210# a_8927_n2982# a_8882_n2778# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5451 a_34039_6251# a_34042_5520# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5452 a_856_n3416# a_435_n3416# a_119_n3096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5453 gnd a_19166_5018# a_18958_5018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5454 gnd a_4079_6075# a_3871_6075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5455 a_38049_7487# a_38063_8590# a_38018_8603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5456 a_29067_7213# a_29063_7390# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5457 a_25890_3841# a_25677_3841# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5458 a_36856_9117# a_36643_9117# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5459 a_31944_1866# a_31731_1866# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5460 a_10466_1064# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5461 a_35709_1640# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5462 gnd a_33248_3021# a_33040_3021# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5463 a_8879_4100# a_8882_3369# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5464 a_21042_2697# a_20621_2697# a_20305_2807# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5465 vdd d0 a_19164_7773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5466 a_24008_n4009# a_24013_n3272# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5467 a_21991_2977# a_21882_2977# a_21989_5189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5468 gnd a_38273_4178# a_38065_4178# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5469 a_11725_n8113# a_11512_n8113# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5470 a_34044_n4380# a_34297_n4584# a_33105_n4070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5471 a_21040_n6152# a_20619_n6152# a_20304_n6156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5472 a_33102_n2052# a_34089_n1824# a_34040_n1808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5473 a_22964_n5741# a_23007_n8157# a_22962_n7953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5474 a_11933_n5913# a_12861_n10677# a_12703_n10661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5475 a_26968_n4808# a_26755_n4808# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5476 a_2887_5778# a_3140_5765# a_2742_6547# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5477 a_15942_n2908# a_15521_n2908# a_15206_n2912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5478 a_20621_3800# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5479 a_434_n3965# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5480 a_29064_n5707# a_29321_n5723# a_28129_n5209# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5481 gnd d2 a_33217_n4866# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5482 a_118_n6405# a_118_n6175# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5483 a_22964_n3541# a_22978_n4861# a_22933_n4657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5484 a_28126_n3191# a_29113_n2963# a_29068_n2759# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5485 a_12917_n8501# a_13170_n8705# a_12772_n9281# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5486 a_26098_n3438# a_26828_n3194# a_27036_n3194# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5487 gnd a_24264_n8991# a_24056_n8991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5488 a_25676_3287# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5489 a_27050_7549# a_26753_8520# a_27033_9112# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5490 a_33099_n7567# a_33356_n7583# a_32963_n6868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5491 vdd d3 a_38302_7474# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5492 a_117_n8381# a_645_n8377# a_853_n8377# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5493 a_35920_n2889# a_35707_n2889# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5494 a_118_5676# a_118_5219# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5495 a_29066_7762# a_29062_7939# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5496 a_14663_485# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5497 a_5490_2203# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5498 a_6570_n2621# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5499 a_29065_n9377# a_29318_n9581# a_28123_n9809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5500 a_5910_7169# a_6640_6925# a_6848_6925# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5501 vdd d4 a_23217_n5945# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5502 a_30649_n8363# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5503 a_17835_n2516# a_18020_n3231# a_17971_n3215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5504 a_29069_n3313# a_29322_n3517# a_28130_n3003# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5505 a_25362_1286# a_25890_1081# a_26098_1081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5506 a_11405_1374# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5507 a_16671_n8733# a_16458_n8733# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5508 a_31590_n4261# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5509 gnd a_38273_n4907# a_38065_n4907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5510 a_18907_9620# a_18910_8889# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5511 vdd a_33246_7433# a_33038_7433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5512 a_21559_n3153# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5513 a_17832_8622# a_18085_8609# a_17863_7506# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5514 a_18913_n5543# a_18909_n5731# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5515 gnd d0 a_29322_n4620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5516 a_22960_3206# a_23217_3016# a_22960_5406# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5517 a_10148_n8845# a_10148_n8616# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5518 a_36756_3023# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5519 a_7937_n9828# a_8924_n9600# a_8879_n9396# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5520 a_30864_n5608# a_30651_n5608# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5521 a_5490_n5663# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5522 a_12134_505# a_11713_505# a_11933_5213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5523 a_17973_8030# a_18226_8017# a_17828_8799# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5524 a_36857_8014# a_36644_8014# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5525 vdd a_28273_n5986# a_28065_n5986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5526 gnd d1 a_38414_3586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5527 a_35389_n9741# a_35389_n9511# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5528 a_10884_n7279# a_11615_n7589# a_11823_n7589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5529 a_15518_8826# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5530 a_27988_6392# a_28173_6890# a_28128_6903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5531 a_16880_n5424# a_16813_n4832# a_16897_n3742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5532 vdd a_28381_n7619# a_28173_n7619# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5533 vdd a_20790_n10911# a_20582_n10911# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5534 a_36785_n7019# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5535 a_25361_2848# a_25361_2619# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5536 a_36128_4949# a_35707_4949# a_35391_5059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5537 a_5911_n6766# a_5490_n6766# a_5174_n6446# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5538 a_32995_n3546# a_33009_n4866# a_32964_n4662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5539 a_5703_n4006# a_5490_n4006# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5540 vdd d0 a_19166_3361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5541 gnd d1 a_8194_n9844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5542 a_1514_n2580# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5543 a_33105_3558# a_34089_3855# a_34044_3868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5544 a_24011_7172# a_24264_7159# a_23072_6862# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5545 a_26094_8802# a_25673_8802# a_25358_9007# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5546 a_21989_5189# a_21669_2977# a_21991_2977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5547 a_35392_n2893# a_35393_n2436# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5548 a_38020_4191# a_38205_4689# a_38156_4879# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5549 a_26613_6906# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5550 vdd d3 a_8085_n8217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5551 gnd a_28383_2478# a_28175_2478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5552 a_33099_n8670# a_34086_n8442# a_34037_n8426# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5553 a_5704_n4560# a_5491_n4560# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5554 gnd a_33358_3545# a_33150_3545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5555 vdd a_38415_1380# a_38207_1380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5556 a_8879_4100# a_9136_3910# a_7944_3613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5557 a_31729_n6978# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5558 a_2889_1366# a_3142_1353# a_2744_2135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5559 a_2778_5248# a_2821_7447# a_2776_7460# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5560 a_11615_n8692# a_11402_n8692# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5561 a_20303_7863# a_20831_7658# a_21039_7658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5562 a_25361_n3534# a_25889_n3987# a_26097_n3987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5563 a_28123_n9809# a_29110_n9581# a_29065_n9377# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5564 a_37065_8014# a_36997_8525# a_37081_7554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5565 a_13854_8848# a_14107_8835# a_12912_9269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5566 a_30334_8327# a_30334_8098# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5567 a_10678_3270# a_10465_3270# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5568 a_27052_3137# a_26755_4108# a_27035_4700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5569 a_17828_n9322# a_18018_n8746# a_17969_n8730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5570 vdd a_3000_n4880# a_2792_n4880# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5571 a_6848_8028# a_6427_8028# a_5910_8272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5572 a_21667_n8089# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5573 vdd d3 a_38304_3062# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5574 a_5910_5512# a_6641_5822# a_6849_5822# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5575 gnd d0 a_34295_4404# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5576 a_5174_n5759# a_5174_n5572# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5577 a_10466_n4524# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5578 vdd d2 a_33218_1931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5579 a_32989_n8146# a_33246_n8162# a_32995_n5746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5580 a_5912_2757# a_6642_2513# a_6850_2513# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5581 a_7938_8202# a_8925_7768# a_8876_7958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5582 gnd a_4077_n8456# a_3869_n8456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5583 a_35919_7155# a_35706_7155# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5584 a_33104_n5173# a_34088_n5687# a_34039_n5671# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5585 gnd d1 a_28383_n3207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5586 vdd a_4079_6075# a_3871_6075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5587 a_25358_n10152# a_29062_n10119# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5588 a_5701_7718# a_5488_7718# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5589 gnd a_8195_6909# a_7987_6909# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5590 vdd a_33248_3021# a_33040_3021# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5591 a_17834_4210# a_18087_4197# a_17865_3094# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5592 gnd a_39349_n9586# a_39141_n9586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5593 gnd d0 a_39351_7205# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5594 a_7942_n8537# a_8926_n9051# a_8881_n8847# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5595 a_29064_n4050# a_29069_n3313# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5596 a_5702_4409# a_5489_4409# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5597 vdd d2 a_28242_n4902# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5598 a_12915_n3174# a_13172_n3190# a_12779_n2475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5599 vdd d0 a_14112_1668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5600 a_5175_4157# a_5175_3970# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5601 a_30333_n10116# a_34294_n10099# a_33102_n9585# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5602 gnd a_39353_n3522# a_39145_n3522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5603 vdd a_24266_n3476# a_24058_n3476# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5604 a_20306_n2390# a_20306_n2203# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5605 a_20831_9315# a_20618_9315# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5606 a_856_2716# a_435_2716# a_119_2826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5607 a_15519_7723# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5608 a_26967_6314# a_26754_6314# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5609 a_25358_n9736# a_25887_n10056# a_26095_n10056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5610 a_10148_n7513# a_10677_n7833# a_10885_n7833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5611 a_20305_n3950# a_20833_n3946# a_21041_n3946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5612 gnd a_4079_n5701# a_3871_n5701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5613 a_2883_5955# a_3140_5765# a_2742_6547# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5614 a_16879_n7630# a_16458_n7630# a_15941_n7874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5615 vdd d1 a_13172_n4293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5616 a_3826_n2737# a_4079_n2941# a_2884_n3169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5617 gnd a_28380_n9825# a_28172_n9825# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5618 a_6430_1410# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5619 a_15205_n5764# a_15733_n6217# a_15941_n6217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5620 gnd a_19164_7773# a_18956_7773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5621 vdd d0 a_39351_n6277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5622 a_16890_7454# a_16599_6338# a_16880_5827# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5623 a_1511_n9198# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5624 a_21989_n7912# a_21698_n6973# a_21979_n6462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5625 a_7830_n3789# a_8087_n3805# a_7830_n5989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5626 a_117_7425# a_645_7677# a_853_7677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5627 vdd a_28271_n8198# a_28063_n8198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5628 vdd d0 a_29322_3891# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5629 a_36127_n6198# a_35706_n6198# a_35391_n6202# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5630 a_30653_1599# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5631 a_5489_7169# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5632 a_1586_n3172# a_1373_n3172# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5633 a_118_4573# a_646_4368# a_854_4368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5634 a_17859_7683# a_17878_6403# a_17829_6593# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5635 a_30336_n4601# a_30863_n5054# a_31071_n5054# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5636 a_24009_4040# a_24012_3309# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5637 gnd a_12861_n10677# a_12653_n10677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5638 a_7942_n7434# a_8195_n7638# a_7802_n6923# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5639 a_20305_3451# a_20833_3246# a_21041_3246# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5640 gnd a_38302_7474# a_38094_7474# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5641 a_37067_3602# a_36999_4113# a_37083_3142# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5642 a_25888_n7850# a_25675_n7850# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5643 a_26723_7430# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5644 a_2772_7637# a_2791_6357# a_2742_6547# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5645 a_11933_5213# a_11512_5213# a_11839_5332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5646 a_5491_2757# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5647 a_2741_8753# a_2931_7971# a_2886_7984# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5648 a_5702_n7869# a_5489_n7869# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5649 vdd d6 a_14967_n10738# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5650 a_7940_3790# a_8927_3356# a_8878_3546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5651 a_119_n3512# a_119_n3325# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5652 a_33098_9250# a_34085_8816# a_34036_9006# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5653 vdd a_33047_n10658# a_32839_n10658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5654 a_10151_n1768# a_9855_n1566# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5655 a_13853_n4033# a_14110_n4049# a_12915_n4277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5656 vdd d1 a_38414_3586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5657 a_854_n6171# a_1585_n6481# a_1793_n6481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5658 a_29061_9042# a_29318_8852# a_28123_9286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5659 a_10466_2721# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5660 a_36997_n9225# a_36784_n9225# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5661 a_11545_n2585# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5662 gnd a_34298_1649# a_34090_1649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5663 a_11834_n7936# a_11725_n8113# a_11839_n5913# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5664 gnd d2 a_13030_n7091# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5665 a_37076_n5758# a_36756_n3723# a_37078_n3546# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5666 a_5703_3306# a_5490_3306# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5667 a_855_2162# a_1586_2472# a_1794_2472# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5668 a_10886_n2867# a_10465_n2867# a_10150_n2871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5669 a_15940_6620# a_15519_6620# a_15205_6368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5670 a_20833_4903# a_20620_4903# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5671 a_27050_n8130# a_26936_n8130# a_27050_n5930# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5672 a_26615_n3194# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5673 a_30337_1480# a_30866_1599# a_31074_1599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5674 a_15206_n4474# a_15735_n4565# a_15943_n4565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5675 a_26969_1902# a_26756_1902# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5676 a_18909_2448# a_18915_1722# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5677 vdd a_33358_3545# a_33150_3545# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5678 a_2885_1543# a_3142_1353# a_2744_2135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5679 a_3823_n9355# a_4076_n9559# a_2881_n9787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5680 a_856_n1759# a_435_n1759# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5681 a_28127_9109# a_28380_9096# a_27987_8598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5682 a_20302_9196# a_20302_8966# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5683 gnd a_28240_8585# a_28032_8585# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5684 vdd d0 a_24263_n8437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5685 a_32959_n7056# a_33149_n6480# a_33100_n6464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5686 a_30650_n6157# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5687 gnd a_19166_3361# a_18958_3361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5688 a_27036_n4297# a_26615_n4297# a_26097_n3987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5689 vdd d1 a_18227_4708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5690 a_10678_n6730# a_10465_n6730# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5691 a_31911_n5894# a_31698_n5894# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5692 a_15207_1956# a_15734_2208# a_15942_2208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5693 a_32889_n10642# a_32839_n10658# a_32790_n10642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5694 a_119_3013# a_647_3265# a_855_3265# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5695 a_26936_n8130# a_26723_n8130# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5696 gnd a_19165_n5193# a_18957_n5193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5697 vdd d0 a_39351_n7934# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5698 vdd a_23327_n4269# a_23119_n4269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5699 a_116_9444# a_116_9215# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5700 a_7804_1999# a_7989_2497# a_7940_2687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5701 a_36127_4395# a_35706_4395# a_35392_4143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5702 a_21910_8479# a_21697_8479# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5703 a_21978_7968# a_21557_7968# a_21039_7658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5704 a_16459_5827# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5705 gnd a_3140_n6494# a_2932_n6494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5706 a_13859_1681# a_13855_1858# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5707 gnd a_38304_3062# a_38096_3062# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5708 a_31729_6278# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5709 a_6642_3616# a_6429_3616# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5710 a_7832_n8013# a_8085_n8217# a_7834_n5801# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5711 gnd a_38304_n5991# a_38096_n5991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5712 a_26725_3018# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5713 a_27034_n8709# a_26966_n9220# a_27050_n8130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5714 a_2774_3225# a_2793_1945# a_2744_2135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5715 gnd d0 a_39352_n5728# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5716 a_2743_4341# a_2933_3559# a_2888_3572# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5717 a_28129_n5209# a_28382_n5413# a_27989_n4698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5718 a_6640_6925# a_6427_6925# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5719 a_26098_n1781# a_26829_n2091# a_27037_n2091# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5720 gnd d0 a_4078_n7907# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5721 a_22289_481# a_25031_461# a_25239_461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5722 vdd a_39349_8857# a_39141_8857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5723 a_7828_7678# a_8085_7488# a_7834_5289# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5724 a_10149_6140# a_10678_6030# a_10886_6030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5725 a_31731_1866# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5726 gnd d1 a_13171_5770# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5727 vdd a_19164_7773# a_18956_7773# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5728 gnd d1 a_8198_n2123# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5729 a_10883_n9485# a_10462_n9485# a_10147_n9489# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5730 a_37067_n4302# a_36646_n4302# a_36128_n3992# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5731 gnd a_14967_n10738# a_14759_n10738# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5732 a_25676_n3987# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5733 a_17863_7506# a_18116_7493# a_17865_5294# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5734 gnd a_34295_n6236# a_34087_n6236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5735 a_2748_n2470# a_3001_n2674# a_2774_n3748# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5736 a_35918_n7301# a_35705_n7301# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5737 a_21913_n2561# a_21700_n2561# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5738 a_5910_8272# a_5489_8272# a_5173_8382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5739 a_10678_4927# a_10465_4927# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5740 a_20830_8761# a_20617_8761# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5741 a_27050_7549# a_26936_7430# a_27050_5349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5742 vdd a_38302_7474# a_38094_7474# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5743 gnd a_19167_n4644# a_18959_n4644# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5744 a_30649_6560# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5745 a_18908_n6280# a_19165_n6296# a_17970_n6524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5746 a_6951_541# a_6738_541# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5747 a_20304_n5053# a_20305_n4596# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5748 a_39099_2252# a_39352_2239# a_38157_2673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5749 vdd d5 a_2830_n10672# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5750 vdd d0 a_24263_n10094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5751 a_8879_n1863# a_9855_n1566# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5752 a_6859_n7972# a_6750_n8149# a_6864_n5949# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5753 a_2883_n6478# a_3140_n6494# a_2742_n7070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5754 a_16781_n8154# a_16568_n8154# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5755 a_23071_n2047# a_24058_n1819# a_24013_n1615# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5756 a_24011_5515# a_24264_5502# a_23069_5936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5757 a_38158_n2093# a_39145_n1865# a_39096_n1849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5758 a_7940_3790# a_8927_3356# a_8882_3369# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5759 vdd a_18226_n7643# a_18018_n7643# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5760 a_16880_4724# a_16459_4724# a_15941_4414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5761 a_21912_4067# a_21699_4067# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5762 a_16674_n2115# a_16461_n2115# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5763 a_5912_n1800# a_6643_n2110# a_6851_n2110# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5764 a_1793_5781# a_1372_5781# a_854_5471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5765 gnd a_34297_n3481# a_34089_n3481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5766 a_2886_6881# a_3870_7178# a_3825_7191# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5767 a_36127_n8958# a_35706_n8958# a_35390_n8638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5768 vdd a_28382_5787# a_28174_5787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5769 gnd d0 a_19165_5567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5770 a_38155_n7608# a_38412_n7624# a_38019_n6909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5771 a_15205_n6221# a_15205_n5764# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5772 a_10464_n7833# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5773 a_27984_n7092# a_28174_n6516# a_28129_n6312# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5774 a_26827_n5400# a_26614_n5400# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5775 a_12774_n4869# a_12964_n4293# a_12919_n4089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5776 gnd d0 a_34297_n1824# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5777 gnd a_38414_3586# a_38206_3586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5778 a_1725_6292# a_1512_6292# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5779 gnd d0 a_39350_n10140# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5780 vdd d0 a_4078_n5147# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5781 a_29962_n10819# a_34945_n10719# a_34896_n10703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5782 a_31071_8217# a_30650_8217# a_30334_8327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5783 a_25359_7904# a_25887_7699# a_26095_7699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5784 a_38160_n5214# a_38413_n5418# a_38020_n4703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5785 a_15943_1105# a_16674_1415# a_16882_1415# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5786 a_37067_2499# a_36646_2499# a_36128_2189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5787 a_10885_n8936# a_10464_n8936# a_10148_n8845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5788 vdd a_28240_8585# a_28032_8585# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5789 vdd a_19166_3361# a_18958_3361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5790 gnd d0 a_19164_n7399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5791 a_2886_n7393# a_3139_n7597# a_2746_n6882# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5792 a_32119_5194# a_32112_486# a_32320_486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5793 a_15207_1769# a_15207_1540# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5794 gnd d1 a_38413_n6521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5795 a_5174_n6446# a_5703_n6766# a_5911_n6766# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5796 a_6864_7568# a_6567_8539# a_6848_8028# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5797 a_10150_n3330# a_10150_n3101# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5798 a_2883_n5375# a_3870_n5147# a_3821_n5131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5799 a_17865_3094# a_18118_3081# a_17861_5471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5800 a_16879_8033# a_16458_8033# a_15940_7723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5801 a_434_n3965# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5802 a_10679_3824# a_10466_3824# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5803 vdd a_14107_n9564# a_13899_n9564# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5804 a_11725_7413# a_11512_7413# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5805 a_15204_8158# a_15733_8277# a_15941_8277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5806 a_19317_288# a_19208_288# a_19416_288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5807 a_7797_n9317# a_7987_n8741# a_7938_n8725# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5808 a_10465_3270# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5809 a_17976_1412# a_18960_1709# a_18915_1722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5810 a_35708_3846# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5811 a_15204_7928# a_15204_7471# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5812 a_5173_6820# a_5701_6615# a_5909_6615# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5813 a_24006_n10078# a_24009_n9336# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5814 vdd a_38304_3062# a_38096_3062# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5815 gnd a_34295_4404# a_34087_4404# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5816 a_2778_3048# a_3031_3035# a_2774_5425# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5817 a_38051_5275# a_38094_7474# a_38045_7664# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5818 a_6570_n2621# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5819 vdd a_33218_1931# a_33010_1931# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5820 a_24012_n6581# a_24265_n6785# a_23073_n6271# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5821 a_16881_3621# a_16460_3621# a_15943_3865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5822 a_38155_n8711# a_39142_n8483# a_39093_n8467# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5823 a_24013_1103# a_24266_1090# a_23071_1524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5824 a_35706_7155# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5825 a_11512_n8113# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5826 a_12803_n8165# a_12822_n7091# a_12773_n7075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5827 a_30863_7114# a_30650_7114# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5828 a_16671_n8733# a_16458_n8733# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5829 a_31590_n4261# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5830 a_3819_9020# a_4076_8830# a_2881_9264# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5831 a_23067_n9768# a_23324_n9784# a_22931_n9069# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5832 gnd a_18088_n2720# a_17880_n2720# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5833 vdd d1 a_13171_5770# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5834 gnd d2 a_8054_8604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5835 a_1808_n8108# a_1694_n8108# a_1808_n5908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5836 gnd d0 a_19167_1155# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5837 a_18911_1899# a_18914_1168# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5838 a_36127_n6198# a_36858_n6508# a_37066_n6508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5839 a_22960_n3729# a_23217_n3745# a_22960_n5929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5840 vdd a_14112_1668# a_13904_1668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5841 a_21770_6865# a_21557_6865# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5842 a_34040_n1808# a_34297_n1824# a_33102_n2052# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5843 a_38045_n8187# a_38302_n8203# a_38051_n5787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5844 a_15207_n1809# a_14830_n1530# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5845 a_15205_5078# a_15205_4849# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5846 a_18913_n5543# a_19166_n5747# a_17974_n5233# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5847 a_38021_n2497# a_38274_n2701# a_38047_n3775# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5848 gnd d1 a_8195_8012# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5849 a_27983_n9298# a_28173_n8722# a_28124_n8706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5850 gnd d0 a_34294_n8442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5851 a_2887_n6290# a_3871_n6804# a_3826_n6600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5852 a_31589_4664# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5853 a_5911_n5663# a_6641_n5419# a_6849_n5419# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5854 a_26754_6314# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5855 a_6427_n8728# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5856 a_20621_n4500# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5857 a_5908_8821# a_5487_8821# a_5173_8569# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5858 a_29063_8493# a_29066_7762# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5859 a_25361_3492# a_25889_3287# a_26097_3287# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5860 gnd d0 a_19166_n6850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5861 a_35705_n10061# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5862 a_118_5032# a_647_4922# a_855_4922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5863 vdd a_29322_n3517# a_29114_n3517# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5864 vdd a_29322_3891# a_29114_3891# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5865 a_7940_3790# a_8197_3600# a_7799_4382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5866 gnd a_29319_n10135# a_29111_n10135# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5867 a_7834_n5801# a_8087_n6005# a_7629_n10697# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5868 vdd d1 a_18225_n9849# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5869 a_11727_n3701# a_11514_n3701# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5870 a_15943_2762# a_15522_2762# a_15206_2872# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5871 a_25888_n6193# a_25675_n6193# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5872 vdd a_33357_n5377# a_33149_n5377# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5873 a_38154_9291# a_39141_8857# a_39092_9047# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5874 a_35390_6806# a_35391_6349# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5875 a_11727_3001# a_11514_3001# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5876 gnd a_4080_3869# a_3872_3869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5877 gnd d3 a_3029_n8176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5878 gnd d0 a_34296_n5687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5879 a_25891_1635# a_25678_1635# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5880 a_5174_5260# a_5702_5512# a_5910_5512# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5881 a_8882_n2778# a_9135_n2982# a_7940_n3210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5882 a_26753_n9220# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5883 vdd d0 a_29322_n1860# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5884 a_8876_7958# a_8881_7232# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5885 a_5175_2408# a_5703_2203# a_5911_2203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5886 a_15732_n7320# a_15519_n7320# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5887 a_17975_3618# a_18228_3605# a_17830_4387# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5888 a_27034_n7606# a_26613_n7606# a_26096_n7850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5889 a_38047_5452# a_38096_3062# a_38047_3252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5890 a_39093_n10124# a_39096_n9382# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5891 a_5490_n4006# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5892 a_26616_n2091# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5893 a_11713_505# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5894 a_30041_n1547# a_30865_n1745# a_31073_n1745# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5895 a_30864_6011# a_30651_6011# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5896 vdd d0 a_24262_8811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5897 a_117_n7924# a_117_n7737# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5898 gnd d1 a_18229_n2128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5899 vdd a_38414_3586# a_38206_3586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5900 a_2888_3572# a_3141_3559# a_2743_4341# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5901 a_3821_4608# a_4078_4418# a_2883_4852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5902 a_32027_n3682# a_31730_n4772# a_32010_n5364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5903 a_1803_n5731# a_1483_n3696# a_1810_n3696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5904 gnd a_18085_n9338# a_17877_n9338# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5905 vdd d1 a_13173_1358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5906 gnd d2 a_8056_4192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5907 a_5490_3306# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5908 a_20306_1704# a_20835_1594# a_21043_1594# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5909 a_21771_5762# a_21558_5762# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5910 a_30336_2999# a_30336_2812# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5911 a_22933_n4657# a_23186_n4861# a_22964_n3541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5912 a_14876_485# a_14663_485# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5913 a_21772_2453# a_21559_2453# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5914 a_20620_4903# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5915 a_5911_4963# a_6641_4719# a_6849_4719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5916 gnd a_14111_n4603# a_13903_n4603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5917 a_646_n6171# a_433_n6171# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5918 a_26756_1902# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5919 a_10148_n7742# a_10677_n7833# a_10885_n7833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5920 a_5912_n1800# a_5491_n1800# a_4799_n1525# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5921 a_17861_3271# a_18118_3081# a_17861_5471# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5922 a_23072_n7374# a_24056_n7888# a_24007_n7872# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5923 vdd a_29320_n9032# a_29112_n9032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5924 a_26968_n4808# a_26755_n4808# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5925 a_13851_9579# a_14108_9389# a_12916_9092# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5926 a_15205_n6221# a_15733_n6217# a_15941_n6217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5927 vdd d0 a_34296_4958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5928 vdd a_18227_4708# a_18019_4708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5929 a_5913_n2354# a_5492_n2354# a_5176_n2263# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5930 a_19332_n829# a_19119_n829# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5931 a_2774_3225# a_3031_3035# a_2774_5425# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5932 a_25359_n9049# a_25359_n8862# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5933 a_38051_5275# a_38094_7474# a_38049_7487# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5934 vdd d0 a_14111_3874# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5935 a_21989_n5712# a_21669_n3677# a_21996_n3677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5936 vdd d0 a_24267_n2373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5937 a_15943_n1805# a_16674_n2115# a_16882_n2115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5938 a_2742_6547# a_2932_5765# a_2883_5955# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5939 a_2778_n3560# a_2792_n4880# a_2747_n4676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5940 a_31070_7663# a_30649_7663# a_30334_7411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5941 a_37065_n7611# a_36644_n7611# a_36127_n7855# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5942 a_11824_5786# a_11403_5786# a_10886_6030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5943 a_17974_n6336# a_18227_n6540# a_17829_n7116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5944 a_21041_n2843# a_20620_n2843# a_20305_n2847# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5945 a_32958_8739# a_33215_8549# a_32993_7446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5946 a_33101_n3155# a_34088_n2927# a_34043_n2723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5947 a_30649_9320# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5948 a_26966_8520# a_26753_8520# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5949 gnd d0 a_14110_n4049# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5950 a_29066_6659# a_29319_6646# a_28124_7080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5951 a_5173_n7549# a_5173_n7319# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5952 a_15205_6181# a_15734_6071# a_15942_6071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5953 a_8879_n9396# a_9132_n9600# a_7937_n9828# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5954 vdd d4 a_3031_n5964# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5955 vdd d0 a_29319_n8478# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5956 vdd d0 a_19167_1155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5957 a_26095_n8399# a_25674_n8399# a_25359_n8403# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5958 vdd d0 a_4079_n2941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5959 a_26095_6596# a_25674_6596# a_25359_6801# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5960 vdd d1 a_8195_8012# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5961 vdd d0 a_24264_4399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5962 a_1373_n3172# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5963 a_13852_n5136# a_13858_n4399# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5964 gnd a_33359_1339# a_33151_1339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5965 a_29065_8865# a_29061_9042# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5966 a_30864_n5608# a_30651_n5608# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5967 a_8880_1894# a_9137_1704# a_7945_1407# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5968 vref a_116_9444# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5969 a_17863_7506# a_17877_8609# a_17828_8799# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5970 a_5701_n10075# a_5488_n10075# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5971 a_32959_n7056# a_33216_n7072# a_32989_n8146# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5972 a_36997_n9225# a_36784_n9225# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5973 a_11401_n9795# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5974 a_17969_n7627# a_18956_n7399# a_18907_n7383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5975 a_37066_5808# a_36998_6319# a_37076_7435# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5976 a_13854_n4587# a_14111_n4603# a_12919_n4089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5977 a_30336_n3498# a_30336_n3311# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5978 a_10886_n2867# a_10465_n2867# a_10151_n2414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5979 gnd d0 a_34296_2198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5980 a_5911_3306# a_6642_3616# a_6850_3616# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5981 a_1794_n4275# a_1373_n4275# a_856_n4519# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5982 a_5172_9026# a_5173_8569# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5983 gnd d3 a_13060_7452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5984 a_21978_6865# a_21911_6273# a_21989_7389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5985 a_13855_n8257# a_14108_n8461# a_12913_n8689# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5986 a_34039_5148# a_34042_4417# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5987 a_37175_n5935# a_38103_n10699# a_34896_n10703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5988 a_9987_364# a_9566_364# a_9888_364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5989 a_10465_4927# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5990 a_25886_8802# a_25673_8802# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5991 a_21882_2977# a_21669_2977# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5992 a_9566_364# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5993 a_854_4368# a_1585_4678# a_1793_4678# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5994 gnd d0 a_39352_4999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X5995 a_5702_n6212# a_5489_n6212# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5996 a_8879_2997# a_8882_2266# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5997 a_3822_n5685# a_3825_n4943# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X5998 a_7944_3613# a_8928_3910# a_8883_3923# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5999 a_38047_5452# a_38096_3062# a_38051_3075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6000 a_5173_8153# a_5173_7923# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6001 a_33100_4838# a_34087_4404# a_34038_4594# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6002 a_2744_2135# a_2934_1353# a_2885_1543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6003 a_31072_3251# a_30651_3251# a_30336_2999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6004 a_20832_7109# a_20619_7109# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6005 a_21039_7658# a_20618_7658# a_20303_7406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6006 a_34042_n7689# a_34295_n7893# a_33103_n7379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6007 a_120_1723# a_120_1494# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6008 a_32960_4327# a_33217_4137# a_32995_3034# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6009 a_1481_n8108# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6010 gnd a_39350_6651# a_39142_6651# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6011 a_23068_7039# a_23325_6849# a_22932_6351# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6012 a_6781_6333# a_6568_6333# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6013 a_26968_4108# a_26755_4108# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6014 vdd a_28241_n7108# a_28033_n7108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6015 a_22927_n9257# a_23117_n8681# a_23068_n8665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6016 a_6859_5249# a_6750_5249# a_6958_5249# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6017 gnd a_19165_5567# a_18957_5567# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6018 a_118_n5302# a_118_n5072# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6019 gnd d0 a_14110_n5706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6020 vdd d1 a_18226_6914# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6021 a_35391_6349# a_35918_6601# a_36126_6601# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6022 vdd a_13171_n6499# a_12963_n6499# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6023 a_26097_2184# a_25676_2184# a_25361_2389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6024 vdd d0 a_29319_n10135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6025 a_118_4573# a_119_4116# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6026 a_17974_n6336# a_18958_n6850# a_18909_n6834# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6027 a_25031_461# a_24818_461# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6028 a_24006_7898# a_24011_7172# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6029 a_1512_6292# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6030 a_17865_3094# a_17879_4197# a_17830_4387# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6031 a_15732_n10080# a_15519_n10080# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6032 a_17835_2004# a_18020_2502# a_17971_2692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6033 a_16781_7454# a_16568_7454# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6034 a_37068_1396# a_37000_1907# a_37078_3023# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6035 a_28020_5270# a_28273_5257# a_27246_522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6036 gnd d0 a_29320_n7929# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6037 gnd d3 a_13062_3040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6038 a_2778_n5760# a_2821_n8176# a_2772_n8160# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6039 a_2742_6547# a_2932_5765# a_2887_5778# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6040 a_30333_9430# a_30862_9320# a_31070_9320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6041 a_10148_n7742# a_10148_n7513# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6042 a_10676_n7279# a_10463_n7279# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6043 a_29064_6287# a_29321_6097# a_28129_5800# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6044 a_10466_3824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6045 a_21978_n7565# a_21557_n7565# a_21040_n7809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6046 a_11512_7413# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6047 a_35918_n7301# a_35705_n7301# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6048 vdd d0 a_9134_n5188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6049 vdd a_8085_n8217# a_7877_n8217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6050 a_20304_n5699# a_20832_n6152# a_21040_n6152# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6051 a_10148_8346# a_10677_8236# a_10885_8236# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6052 a_29062_6836# a_29319_6646# a_28124_7080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6053 a_8875_9061# a_9132_8871# a_7937_9305# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6054 a_2887_4675# a_3871_4972# a_3822_5162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6055 gnd d1 a_23327_n3166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6056 a_12775_n2663# a_13032_n2679# a_12805_n3753# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6057 a_30652_n1745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6058 vdd d0 a_39352_n2968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6059 a_5704_1100# a_5491_1100# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6060 a_116_n10130# a_3820_n10097# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6061 a_15940_7723# a_15519_7723# a_15204_7928# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6062 a_21040_n8912# a_20619_n8912# a_20303_n8821# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6063 a_36128_n2889# a_35707_n2889# a_35392_n2893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6064 a_33103_n8482# a_34087_n8996# a_34042_n8792# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6065 vdd d1 a_28382_n6516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6066 a_645_9334# a_432_9334# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6067 a_15941_4414# a_15520_4414# a_15206_4162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6068 gnd d0 a_29320_4440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6069 gnd a_13029_n9297# a_12821_n9297# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6070 a_5702_n7869# a_5489_n7869# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6071 a_10150_n3517# a_10150_n3330# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6072 a_30650_7114# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6073 a_25886_n9502# a_25673_n9502# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6074 a_6783_1921# a_6570_1921# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6075 a_23070_2627# a_23327_2437# a_22934_1939# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6076 a_2742_6547# a_2999_6357# a_2772_7637# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6077 a_1803_n7931# a_1512_n6992# a_1793_n6481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6078 a_33103_7970# a_33356_7957# a_32958_8739# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6079 gnd a_28241_6379# a_28033_6379# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6080 gnd a_19167_1155# a_18959_1155# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6081 gnd a_8054_8604# a_7846_8604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6082 vdd a_24262_n9540# a_24054_n9540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6083 gnd a_28383_n3207# a_28175_n3207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6084 a_5910_7169# a_5489_7169# a_5173_7050# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6085 a_30334_7224# a_30334_6995# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6086 a_30335_5892# a_30335_5662# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6087 vdd d1 a_18228_2502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6088 a_30648_8766# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6089 a_10464_n7833# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6090 a_648_n3416# a_435_n3416# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6091 a_122_1165# a_648_1059# a_856_1059# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6092 vdd a_4078_n9010# a_3870_n9010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6093 vdd d3 a_13060_7452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6094 gnd a_8195_8012# a_7987_8012# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6095 a_22964_n5741# a_23217_n5945# a_22759_n10637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6096 a_25361_3951# a_25890_3841# a_26098_3841# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6097 a_24010_7721# a_24263_7708# a_23068_8142# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6098 gnd a_29320_7200# a_29112_7200# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6099 a_33103_n8482# a_33356_n8686# a_32958_n9262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6100 a_36128_2189# a_35707_2189# a_35393_1937# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6101 a_17859_n8206# a_17878_n7132# a_17833_n6928# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6102 a_16783_3042# a_16570_3042# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6103 a_10885_n8936# a_10464_n8936# a_10148_n8616# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6104 vdd a_19167_n1884# a_18959_n1884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6105 a_1792_7987# a_1371_7987# a_853_7677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6106 a_26827_4700# a_26614_4700# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6107 a_16461_n2115# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6108 gnd a_29321_n4066# a_29113_n4066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6109 vdd d1 a_38411_9101# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6110 a_10676_n10039# a_10463_n10039# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6111 a_8879_n3520# a_9136_n3536# a_7944_n3022# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6112 a_25359_n7300# a_25887_n7296# a_26095_n7296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6113 a_856_n1759# a_435_n1759# a_120_n1763# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6114 a_39096_2983# a_39353_2793# a_38161_2496# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6115 a_13857_n3845# a_13853_n4033# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6116 a_24009_n4563# a_24012_n3821# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6117 a_22934_n2451# a_23119_n3166# a_23074_n2962# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6118 a_5174_n6675# a_5703_n6766# a_5911_n6766# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6119 a_12915_n4277# a_13902_n4049# a_13853_n4033# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6120 a_38158_9114# a_39142_9411# a_39093_9601# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6121 a_3826_6088# a_3822_6265# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6122 a_10678_n6730# a_10465_n6730# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6123 a_2744_2135# a_2934_1353# a_2889_1366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6124 vdd d0 a_9136_n4639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6125 a_36127_4395# a_36858_4705# a_37066_4705# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6126 a_2573_n10656# a_2823_n5964# a_2778_n5760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6127 a_39099_3355# a_39095_3532# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6128 a_36857_n8714# a_36644_n8714# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6129 a_1583_n9790# a_1370_n9790# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6130 a_11514_3001# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6131 a_1724_8498# a_1511_8498# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6132 vdd a_39350_6651# a_39142_6651# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6133 a_30074_345# a_34849_466# a_32320_486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6134 a_3824_6637# a_4077_6624# a_2882_7058# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6135 vdd d1 a_13170_n7602# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6136 a_11615_7992# a_11402_7992# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6137 a_8877_4649# a_9134_4459# a_7939_4893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6138 gnd d1 a_13172_3564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6139 a_15204_n9073# a_15731_n9526# a_15939_n9526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6140 vdd d0 a_39349_n9586# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6141 a_14985_485# a_16769_546# a_16989_5254# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6142 a_28127_n2088# a_28384_n2104# a_27986_n2680# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6143 a_6643_n2110# a_6430_n2110# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6144 gnd d0 a_4080_n4598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6145 a_646_8231# a_433_8231# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6146 a_36644_8014# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6147 gnd a_8197_n3226# a_7989_n3226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6148 a_15942_3311# a_15521_3311# a_15206_3516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6149 a_35919_4395# a_35706_4395# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6150 gnd d1 a_28381_n8722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6151 a_30651_6011# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6152 a_18912_n8852# a_19165_n9056# a_17973_n8542# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6153 vdd a_24262_8811# a_24054_8811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6154 a_15521_n6771# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6155 a_16783_n3742# a_16570_n3742# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6156 vdd a_38413_n5418# a_38205_n5418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6157 vdd d0 a_4078_7178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6158 a_644_n9480# a_431_n9480# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6159 a_5911_6066# a_5490_6066# a_5174_6176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6160 vdd a_13173_1358# a_12965_1358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6161 a_24009_2937# a_24012_2206# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6162 a_30649_7663# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6163 gnd a_8056_4192# a_7848_4192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6164 a_20831_6555# a_20618_6555# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6165 a_10150_3705# a_10150_3475# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6166 a_7834_5289# a_7877_7488# a_7832_7501# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6167 vdd d3 a_13062_3040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6168 a_2744_2135# a_3001_1945# a_2774_3225# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6169 a_10886_6030# a_10465_6030# a_10149_5911# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6170 a_16880_5827# a_16459_5827# a_15942_6071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6171 a_32025_5313# a_31698_7394# a_32025_7513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6172 a_24012_3309# a_24265_3296# a_23070_3730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6173 a_16890_n7977# a_16599_n7038# a_16879_n7630# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6174 a_16881_2518# a_16460_2518# a_15942_2208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6175 a_1794_3575# a_1373_3575# a_855_3265# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6176 vdd a_19164_n8502# a_18956_n8502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6177 a_38015_6574# a_38205_5792# a_38160_5805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6178 vdd a_34296_4958# a_34088_4958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6179 a_30864_n3951# a_30651_n3951# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6180 a_34038_4594# a_34044_3868# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6181 vdd d1 a_13170_7976# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6182 a_853_n8377# a_432_n8377# a_117_n8381# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6183 a_17865_5294# a_17908_7493# a_17859_7683# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6184 a_24008_n4009# a_24265_n4025# a_23070_n4253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6185 vdd d1 a_8197_n3226# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6186 a_11544_4091# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6187 a_3822_2402# a_3828_1676# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6188 a_27989_n4698# a_28242_n4902# a_28020_n3582# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6189 a_11727_n3701# a_11514_n3701# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6190 vdd d0 a_29320_4440# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6191 vdd a_3029_7447# a_2821_7447# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6192 vdd d0 a_34295_5507# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6193 a_32221_486# a_33040_5221# a_32991_5411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6194 a_11402_n8692# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6195 a_26753_8520# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6196 a_2778_5248# a_2821_7447# a_2772_7637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6197 a_1726_4086# a_1513_4086# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6198 a_12918_n5192# a_13902_n5706# a_13853_n5690# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6199 a_3826_2225# a_4079_2212# a_2884_2646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6200 vdd d0 a_39351_n9037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6201 vdd a_9133_n10154# a_8925_n10154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6202 a_13857_3333# a_13853_3510# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6203 a_12919_n4089# a_13172_n4293# a_12774_n4869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6204 vdd d0 a_19168_1709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6205 gnd a_24266_n4579# a_24058_n4579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6206 a_854_n5068# a_433_n5068# a_119_n4615# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6207 a_32962_n9074# a_33147_n9789# a_33098_n9773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6208 a_33101_n3155# a_33358_n3171# a_32965_n2456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6209 a_24013_n1615# a_24266_n1819# a_23071_n2047# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6210 a_27034_n7606# a_26613_n7606# a_26095_n7296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6211 a_39098_n6073# a_39351_n6277# a_38156_n6505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6212 gnd d1 a_8197_3600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6213 vdd d3 a_13060_n8181# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6214 a_28124_n8706# a_28381_n8722# a_27983_n9298# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6215 a_36127_n8958# a_35706_n8958# a_35390_n8867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6216 vdd a_19167_1155# a_18959_1155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6217 a_10676_n10039# a_10463_n10039# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6218 a_18909_n2971# a_19166_n2987# a_17971_n3215# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6219 vdd d0 a_29323_n2414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6220 a_30337_n1749# a_30865_n1745# a_31073_n1745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6221 a_34849_466# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6222 a_11824_n5383# a_11757_n4791# a_11841_n3701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6223 a_7939_5996# a_8196_5806# a_7798_6588# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6224 vdd a_23325_n7578# a_23117_n7578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6225 a_30334_n7494# a_30863_n7814# a_31071_n7814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6226 a_35920_2189# a_35707_2189# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6227 vdd a_8195_8012# a_7987_8012# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6228 vdd a_24264_4399# a_24056_4399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6229 gnd a_38412_n7624# a_38204_n7624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6230 a_37175_n5935# a_36754_n5935# a_37081_n5935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6231 vdd d1 a_33358_n4274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6232 a_21773_n2050# a_21560_n2050# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6233 vdd d0 a_39351_8308# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6234 a_20832_5452# a_20619_5452# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6235 a_32027_n3682# a_31730_n4772# a_32011_n4261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6236 vdd d0 a_19166_n4090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6237 a_30337_n1979# a_30866_n2299# a_31074_n2299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6238 a_16673_n4321# a_16460_n4321# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6239 a_5173_7466# a_5701_7718# a_5909_7718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6240 gnd d0 a_34297_2752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6241 gnd a_3138_n9803# a_2930_n9803# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6242 a_6641_n5419# a_6428_n5419# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6243 a_20833_2143# a_20620_2143# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6244 a_24964_n10698# a_24914_n10714# a_22858_n10637# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6245 a_29065_n4604# a_29068_n3862# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6246 a_5174_4614# a_5702_4409# a_5910_4409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6247 a_2885_n2066# a_3872_n1838# a_3827_n1634# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6248 a_19416_288# a_18995_288# a_19317_288# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6249 gnd a_34296_2198# a_34088_2198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6250 a_25359_7031# a_25359_6801# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6251 gnd a_3031_n3764# a_2823_n3764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6252 a_20302_9196# a_20831_9315# a_21039_9315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6253 gnd d0 a_14112_1668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6254 a_7941_n9640# a_8925_n10154# a_8876_n10138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6255 a_17833_n6928# a_18086_n7132# a_17859_n8206# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6256 a_7939_n5416# a_8926_n5188# a_8881_n4984# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6257 a_20619_n6152# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6258 a_38158_9114# a_39142_9411# a_39097_9424# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6259 a_30863_8217# a_30650_8217# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6260 a_5175_3511# a_5175_3054# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6261 a_16882_1415# a_16461_1415# a_15944_1659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6262 a_38047_3252# a_38066_1972# a_38021_1985# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6263 a_32963_6356# a_33216_6343# a_32989_7623# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6264 vdd d0 a_34296_n2927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6265 a_36859_2499# a_36646_2499# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6266 gnd a_7886_n10713# a_7678_n10713# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6267 a_35707_4949# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6268 vdd d1 a_33357_4648# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6269 a_10886_n2867# a_11617_n3177# a_11825_n3177# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6270 a_30337_1896# a_30864_2148# a_31072_2148# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6271 a_38045_n8187# a_38064_n7113# a_38015_n7097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6272 a_19317_288# a_29752_345# a_30074_345# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6273 a_25673_8802# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6274 a_3820_6814# a_4077_6624# a_2882_7058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6275 a_18908_5757# a_18913_5031# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6276 vdd d1 a_13172_3564# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6277 a_5913_n2354# a_5492_n2354# a_5176_n2034# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6278 gnd d2 a_8055_6398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6279 a_21910_n9179# a_21697_n9179# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6280 gnd d1 a_8196_n5432# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6281 gnd a_39352_4999# a_39144_4999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6282 a_21989_n5712# a_21669_n3677# a_21991_n3500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6283 a_31589_5767# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6284 a_37065_n7611# a_36644_n7611# a_36126_n7301# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6285 a_21771_4659# a_21558_4659# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6286 vdd a_34296_n6790# a_34088_n6790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6287 a_32119_n5894# a_31698_n5894# a_32020_n5717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6288 gnd d3 a_28273_n3786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6289 a_21041_n2843# a_20620_n2843# a_20306_n2390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6290 a_13857_6093# a_14110_6080# a_12918_5783# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6291 a_33101_n4258# a_34088_n4030# a_34039_n4014# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6292 gnd a_34293_n9545# a_34085_n9545# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6293 a_26755_4108# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6294 a_433_n6171# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6295 a_15941_n5114# a_15520_n5114# a_15205_n5118# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6296 a_5909_6615# a_5488_6615# a_5174_6363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6297 gnd d2 a_33216_n7072# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6298 a_11617_n4280# a_11404_n4280# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6299 a_2774_5425# a_2823_3035# a_2774_3225# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6300 a_28125_n5397# a_29112_n5169# a_29067_n4965# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6301 a_21042_n3397# a_20621_n3397# a_20305_n3306# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6302 a_24010_n8233# a_24263_n8437# a_23068_n8665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6303 a_116_n9714# a_116_n9484# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6304 gnd a_19165_n7953# a_18957_n7953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6305 vdd a_18226_6914# a_18018_6914# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6306 vdd a_3139_7971# a_2931_7971# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6307 a_119_2826# a_648_2716# a_856_2716# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6308 a_8876_n10138# a_8879_n9396# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6309 a_7941_1584# a_8198_1394# a_7800_2176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6310 gnd a_4079_n4044# a_3871_n4044# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6311 a_2881_9264# a_3868_8830# a_3823_8843# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6312 a_23069_n5356# a_24056_n5128# a_24011_n4924# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6313 a_21770_n8668# a_21557_n8668# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6314 vdd d0 a_4080_n3495# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6315 a_25674_n7296# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6316 a_29069_1144# a_29065_1321# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6317 vdd a_23215_n8157# a_23007_n8157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6318 a_5910_n5109# a_6641_n5419# a_6849_n5419# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6319 a_2774_n3748# a_3031_n3764# a_2774_n5948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6320 a_24012_n2718# a_24008_n2906# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6321 a_120_1910# a_120_1723# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6322 a_5175_3054# a_5703_3306# a_5911_3306# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6323 a_31071_n6157# a_30650_n6157# a_30335_n6161# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6324 a_25361_n3347# a_25361_n3118# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6325 gnd a_39351_n5174# a_39143_n5174# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6326 a_1794_n4275# a_1373_n4275# a_855_n3965# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6327 a_16670_9136# a_16457_9136# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6328 a_7944_n4125# a_8928_n4639# a_8883_n4435# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6329 a_20304_4784# a_20833_4903# a_21041_4903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6330 a_17976_1412# a_18229_1399# a_17831_2181# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6331 gnd a_13062_3040# a_12854_3040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6332 a_15206_3516# a_15206_3059# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6333 a_37067_3602# a_36646_3602# a_36128_3292# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6334 a_32012_n2055# a_31591_n2055# a_31073_n1745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6335 vdd a_29321_n4066# a_29113_n4066# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6336 a_38160_4702# a_39144_4999# a_39099_5012# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6337 a_12777_n6887# a_12962_n7602# a_12917_n7398# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6338 a_15205_n5118# a_15206_n4661# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6339 a_32965_1944# a_33218_1931# a_32991_3211# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6340 vdd d0 a_24263_6605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6341 a_15518_n9526# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6342 a_1587_n2069# a_1374_n2069# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6343 a_2745_8576# a_2998_8563# a_2776_7460# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6344 a_23073_4656# a_23326_4643# a_22933_4145# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6345 gnd d2 a_8057_n2715# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6346 a_10150_n3101# a_10679_n3421# a_10887_n3421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6347 a_31072_n2848# a_30651_n2848# a_30337_n2395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6348 a_32221_486# a_33040_5221# a_32995_5234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6349 a_28016_n5970# a_28065_n3786# a_28020_n3582# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6350 a_37065_6911# a_36644_6911# a_36127_7155# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6351 a_7939_n5416# a_8196_n5432# a_7803_n4717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6352 a_3822_2402# a_4079_2212# a_2884_2646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6353 a_38159_8011# a_38412_7998# a_38014_8780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6354 a_7799_4382# a_7989_3600# a_7944_3613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6355 a_5491_1100# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6356 gnd d2 a_8057_1986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6357 a_5702_n6212# a_5489_n6212# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6358 a_21772_3556# a_21559_3556# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6359 a_36859_n3199# a_36646_n3199# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6360 a_32010_4664# a_31589_4664# a_31071_4354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6361 a_35920_n3992# a_35707_n3992# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6362 a_432_9334# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6363 gnd d1 a_38411_n9830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6364 a_25361_n3991# a_25361_n3534# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6365 a_19208_288# a_18995_288# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6366 a_21977_9071# a_21910_8479# a_21994_7508# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6367 a_25889_n2884# a_25676_n2884# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6368 a_31728_n9184# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6369 a_6570_1921# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6370 a_25360_n5740# a_25888_n6193# a_26096_n6193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6371 a_35921_n4546# a_35708_n4546# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6372 a_18908_n9040# a_19165_n9056# a_17973_n8542# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6373 vdd d0 a_34297_2752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6374 a_20831_n7255# a_20618_n7255# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6375 a_120_1494# a_649_1613# a_857_1613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6376 a_37175_5235# a_36754_5235# a_37076_5235# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6377 a_24008_2383# a_24014_1657# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6378 vdd a_18228_2502# a_18020_2502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6379 vdd a_3141_3559# a_2933_3559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6380 a_15204_6825# a_15205_6368# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6381 vdd a_33217_n4866# a_33009_n4866# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6382 a_36129_2743# a_35708_2743# a_35392_2624# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6383 a_2743_4341# a_2933_3559# a_2884_3749# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6384 a_31073_1045# a_31804_1355# a_32012_1355# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6385 a_17972_9133# a_18225_9120# a_17832_8622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6386 a_31071_5457# a_30650_5457# a_30335_5205# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6387 a_39094_n5158# a_39351_n5174# a_38156_n5402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6388 vdd a_14112_n2397# a_13904_n2397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6389 a_32959_6533# a_33216_6343# a_32989_7623# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6390 a_16570_3042# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6391 a_6780_8539# a_6567_8539# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6392 a_8880_6678# a_9133_6665# a_7938_7099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6393 a_26614_4700# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6394 a_16671_8033# a_16458_8033# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6395 a_10885_n8936# a_11615_n8692# a_11823_n8692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6396 a_36125_n9507# a_36856_n9817# a_37064_n9817# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6397 a_16598_8544# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6398 a_33104_4661# a_34088_4958# a_34043_4971# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6399 a_13855_n8257# a_13851_n8445# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6400 a_36967_n8135# a_36754_n8135# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6401 a_24007_n8975# a_24010_n8233# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6402 gnd a_18226_n8746# a_18018_n8746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6403 a_35390_8555# a_35917_8807# a_36125_8807# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6404 a_11755_8503# a_11542_8503# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6405 vdd d0 a_34295_n8996# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6406 a_34038_n5117# a_34295_n5133# a_33100_n5361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6407 a_6782_n4827# a_6569_n4827# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6408 a_26096_4390# a_25675_4390# a_25360_4595# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6409 a_27047_3018# a_26756_1902# a_27037_1391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6410 a_30334_7411# a_30334_7224# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6411 a_6849_5822# a_6428_5822# a_5910_5512# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6412 a_27052_n3718# a_26938_n3718# a_27045_n5753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6413 a_21978_n7565# a_21557_n7565# a_21039_n7255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6414 vdd d0 a_24265_2193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6415 a_18912_n6092# a_18908_n6280# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6416 a_27144_5230# a_27137_522# a_25140_461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6417 a_13853_6270# a_14110_6080# a_12918_5783# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6418 gnd d0 a_4077_9384# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6419 a_1511_8498# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6420 a_3820_n7337# a_3826_n6600# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6421 a_12809_n5765# a_12852_n8181# a_12807_n7977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6422 a_20302_8966# a_20830_8761# a_21038_8761# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6423 a_3825_n4943# a_4078_n5147# a_2883_n5375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6424 a_2774_5425# a_2823_3035# a_2778_3048# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6425 a_11402_7992# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6426 a_10677_4373# a_10464_4373# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6427 gnd a_13172_3564# a_12964_3564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6428 a_31802_n6467# a_31589_n6467# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6429 a_34044_n1620# a_34040_n1808# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6430 a_30652_n1745# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6431 a_32011_3561# a_31590_3561# a_31073_3805# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6432 a_6847_9131# a_6426_9131# a_5909_9375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6433 a_30862_7663# a_30649_7663# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6434 a_34043_n2723# a_34296_n2927# a_33101_n3155# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6435 a_433_8231# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6436 a_5912_1100# a_6643_1410# a_6851_1410# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6437 a_35706_4395# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6438 a_21040_n8912# a_20619_n8912# a_20303_n8592# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6439 a_15735_3865# a_15522_3865# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6440 gnd d0 a_4078_n6250# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6441 a_30653_n2299# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6442 a_17971_n4318# a_18958_n4090# a_18913_n3886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6443 vdd d0 a_39353_n3522# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6444 a_25361_3492# a_25361_3035# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6445 a_1792_6884# a_1725_6292# a_1803_7408# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6446 a_21979_4659# a_21912_4067# a_21996_3096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6447 a_37081_5354# a_36754_7435# a_37081_7554# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6448 a_25886_n9502# a_25673_n9502# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6449 vdd d2 a_13032_1950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6450 a_29068_n2759# a_29064_n2947# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6451 a_34036_9006# a_34042_8280# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6452 a_29063_8493# a_29320_8303# a_28128_8006# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6453 a_20833_n6706# a_20620_n6706# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6454 gnd a_13062_n3769# a_12854_n3769# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6455 a_31803_n3158# a_31590_n3158# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6456 vdd a_4078_7178# a_3870_7178# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6457 a_2886_6881# a_3870_7178# a_3821_7368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6458 a_15733_7174# a_15520_7174# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6459 a_25887_6596# a_25674_6596# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6460 a_5700_8821# a_5487_8821# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6461 a_118_n6821# a_645_n7274# a_853_n7274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6462 a_8876_6855# a_8882_6129# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6463 a_1726_n4786# a_1513_n4786# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6464 a_648_n3416# a_435_n3416# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6465 gnd a_28381_6890# a_28173_6890# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6466 a_7945_1407# a_8929_1704# a_8884_1717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6467 vdd a_13062_3040# a_12854_3040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6468 a_33101_2632# a_34088_2198# a_34039_2388# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6469 gnd d0 a_29319_6646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6470 a_31073_1045# a_30652_1045# a_30339_1151# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6471 gnd d0 a_34294_7713# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6472 a_35389_9471# a_35389_9242# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6473 a_856_n3416# a_1586_n3172# a_1794_n3172# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6474 gnd a_39351_4445# a_39143_4445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6475 a_23069_4833# a_23326_4643# a_22933_4145# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6476 a_6782_4127# a_6569_4127# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6477 a_3822_n6788# a_4079_n6804# a_2887_n6290# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6478 a_2741_8753# a_2998_8563# a_2776_7460# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6479 a_8882_2266# a_9135_2253# a_7940_2687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6480 a_11616_4683# a_11403_4683# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6481 a_21980_n4256# a_21912_n4767# a_21996_n3677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6482 a_10885_n5073# a_10464_n5073# a_10149_n5077# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6483 a_35392_4143# a_35919_4395# a_36127_4395# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6484 a_36857_n8714# a_36644_n8714# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6485 a_11405_n2074# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6486 vdd a_34295_5507# a_34087_5507# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6487 gnd a_14109_n7912# a_13901_n7912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6488 gnd a_29319_9406# a_29111_9406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6489 a_5910_n5109# a_5489_n5109# a_5175_n4656# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6490 a_1513_4086# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6491 vdd a_19168_1709# a_18960_1709# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6492 a_26826_6906# a_26613_6906# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6493 a_15203_n9530# a_15731_n9526# a_15939_n9526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6494 a_27815_n10678# a_28072_n10694# a_24865_n10698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6495 a_30864_3251# a_30651_3251# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6496 gnd a_8197_3600# a_7989_3600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6497 a_5911_n5663# a_5490_n5663# a_5174_n5572# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6498 a_10149_n5307# a_10149_n5077# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6499 vdd a_8055_n7127# a_7847_n7127# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6500 a_5703_n2903# a_5490_n2903# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6501 a_25358_9237# a_25887_9356# a_26095_9356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6502 gnd d5 a_38103_n10699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6503 a_3827_1122# a_3823_1299# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6504 vdd d0 a_24265_n5682# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6505 a_15521_n6771# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6506 a_16783_n3742# a_16570_n3742# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6507 a_17968_9310# a_18225_9120# a_17832_8622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6508 a_30334_7224# a_30863_7114# a_31071_7114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6509 a_37076_5235# a_36756_3023# a_37083_3142# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6510 a_17972_n9645# a_18225_n9849# a_17832_n9134# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6511 a_6958_5249# a_6537_5249# a_6864_5368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6512 a_10467_1618# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6513 gnd a_34297_2752# a_34089_2752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6514 a_8876_6855# a_9133_6665# a_7938_7099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6515 a_118_n6405# a_647_n6725# a_855_n6725# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6516 a_25889_2184# a_25676_2184# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6517 a_38157_n3196# a_38414_n3212# a_38021_n2497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6518 a_29069_n1656# a_29322_n1860# a_28127_n2088# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6519 a_20620_2143# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6520 a_35920_6052# a_35707_6052# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6521 a_29063_n9016# a_29066_n8274# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6522 a_21040_7109# a_21770_6865# a_21978_6865# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6523 gnd a_33357_n6480# a_33149_n6480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6524 a_15941_5517# a_15520_5517# a_15205_5722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6525 gnd a_14112_1668# a_13904_1668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6526 a_6539_n3737# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6527 a_7830_n3789# a_7849_n2715# a_7800_n2699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6528 a_10466_n3421# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6529 a_30336_2583# a_30865_2702# a_31073_2702# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6530 a_646_7128# a_433_7128# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6531 gnd d0 a_29321_2234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6532 a_15942_2208# a_15521_2208# a_15207_1956# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6533 a_30650_8217# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6534 vdd d1 a_38414_n4315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6535 vdd a_33357_4648# a_33149_4648# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6536 a_24007_n6215# a_24012_n5478# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6537 vdd d0 a_4077_9384# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6538 a_30864_n3951# a_30651_n3951# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6539 a_10887_n4524# a_10466_n4524# a_10150_n4433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6540 vdd a_13172_3564# a_12964_3564# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6541 a_853_n8377# a_432_n8377# a_117_n7924# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6542 gnd a_8055_6398# a_7847_6398# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6543 a_7798_n7111# a_7988_n6535# a_7943_n6331# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6544 a_1792_n7584# a_1371_n7584# a_854_n7828# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6545 a_35171_466# a_36955_527# a_37175_5235# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6546 a_25675_n6193# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6547 gnd d1 a_3141_n3185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6548 a_854_5471# a_1585_5781# a_1793_5781# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6549 a_7937_9305# a_8924_8871# a_8879_8884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6550 a_10885_8236# a_10464_8236# a_10148_8117# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6551 a_2885_n9599# a_3869_n10113# a_3820_n10097# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6552 a_5175_3970# a_5704_3860# a_5912_3860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6553 a_25362_1745# a_25891_1635# a_26099_1635# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6554 a_26827_5803# a_26614_5803# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6555 gnd a_29321_4994# a_29113_4994# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6556 vdd a_14109_n5152# a_13901_n5152# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6557 vdd d0 a_14109_n9015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6558 gnd a_38271_n9319# a_38063_n9319# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6559 a_28016_n3770# a_28035_n2696# a_27986_n2680# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6560 a_17660_n10702# a_17917_n10718# a_14710_n10722# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6561 a_8877_8512# a_8880_7781# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6562 a_20306_n2390# a_20833_n2843# a_21041_n2843# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6563 a_32320_486# a_31899_486# a_32221_486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6564 a_27144_5230# a_26723_5230# a_27050_5349# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6565 a_7799_n4905# a_7989_n4329# a_7940_n4313# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6566 a_5700_n9521# a_5487_n9521# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6567 a_11543_6297# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6568 a_18912_5580# a_18908_5757# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6569 a_25360_4825# a_25889_4944# a_26097_4944# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6570 a_24014_n2169# a_24267_n2373# a_23075_n1859# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6571 a_30334_n7723# a_30863_n7814# a_31071_n7814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6572 a_24009_4040# a_24266_3850# a_23074_3553# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6573 a_37175_n5935# a_36754_n5935# a_37076_n5758# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6574 a_38157_n4299# a_39144_n4071# a_39095_n4055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6575 gnd d1 a_33358_2442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6576 vdd d0 a_29319_6646# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6577 vdd a_9135_n5742# a_8927_n5742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6578 a_8877_n5172# a_8883_n4435# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6579 gnd d2 a_23187_n2655# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6580 a_36128_2189# a_36859_2499# a_37067_2499# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6581 a_8880_9438# a_10147_9449# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6582 vdd d0 a_34294_7713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6583 a_37076_n7958# a_36967_n8135# a_37081_n5935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6584 a_16673_n4321# a_16460_n4321# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6585 vdd a_39351_4445# a_39143_4445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6586 a_3825_4431# a_4078_4418# a_2883_4852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6587 a_21040_5452# a_21771_5762# a_21979_5762# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6588 vdd d0 a_19167_3915# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6589 a_23069_n5356# a_23326_n5372# a_22933_n4657# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6590 a_8878_2443# a_9135_2253# a_7940_2687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6591 gnd d1 a_13173_1358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6592 a_2778_n5760# a_3031_n5964# a_2573_n10656# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6593 a_36126_7704# a_35705_7704# a_35390_7452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6594 a_21042_2697# a_21772_2453# a_21980_2453# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6595 a_647_6025# a_434_6025# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6596 gnd d1 a_8196_5806# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6597 a_15943_1105# a_15522_1105# a_15207_1310# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6598 vdd a_13169_n9808# a_12961_n9808# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6599 gnd d0 a_34296_n4030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6600 gnd a_9135_n4085# a_8927_n4085# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6601 a_2889_n1878# a_3873_n2392# a_3828_n2188# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6602 vdd d1 a_23326_n6475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6603 a_15203_n9530# a_15204_n9073# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6604 a_37000_1907# a_36787_1907# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6605 vdd a_24263_6605# a_24055_6605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6606 a_6429_n4316# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6607 a_18914_2825# a_18910_3002# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6608 a_35391_n6848# a_35391_n6661# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6609 a_20305_n4180# a_20834_n4500# a_21042_n4500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6610 vdd a_24266_n1819# a_24058_n1819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6611 gnd a_39353_n1865# a_39145_n1865# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6612 a_20831_7658# a_20618_7658# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6613 a_24006_6795# a_24012_6069# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6614 a_5173_n8422# a_5701_n8418# a_5909_n8418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6615 gnd d0 a_19168_n2438# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6616 a_20832_4349# a_20619_4349# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6617 gnd a_8057_1986# a_7849_1986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6618 a_27052_3137# a_26938_3018# a_27045_5230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6619 gnd a_3140_5765# a_2932_5765# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6620 a_18908_8517# a_19165_8327# a_17973_8030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6621 a_15206_n2912# a_15734_n2908# a_15942_n2908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6622 a_29066_9419# a_29062_9596# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6623 gnd a_13173_n2087# a_12965_n2087# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6624 a_30337_1480# a_30337_1250# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6625 a_2882_7058# a_3869_6624# a_3820_6814# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6626 a_8879_n4623# a_8882_n3881# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6627 a_7939_4893# a_8926_4459# a_8881_4472# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6628 vdd d1 a_18227_n5437# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6629 a_8878_6306# a_8881_5575# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6630 a_32962_8562# a_33215_8549# a_32993_7446# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6631 a_26829_1391# a_26616_1391# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6632 vdd d1 a_33356_6854# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6633 a_35391_n6432# a_35920_n6752# a_36128_n6752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6634 vdd a_28382_n6516# a_28174_n6516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6635 a_15206_n3142# a_15735_n3462# a_15943_n3462# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6636 a_28018_n7994# a_28032_n9314# a_27983_n9298# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6637 a_32011_2458# a_31944_1866# a_32022_2982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6638 a_25359_7260# a_25359_7031# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6639 a_20303_n9008# a_20830_n9461# a_21038_n9461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6640 a_1795_1369# a_1374_1369# a_856_1059# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6641 vdd a_34297_2752# a_34089_2752# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6642 a_10885_8236# a_11615_7992# a_11823_7992# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6643 gnd d0 a_19164_6670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6644 a_38158_n9626# a_39142_n10140# a_39093_n10124# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6645 a_31911_7394# a_31698_7394# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6646 a_35392_4143# a_35392_3956# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6647 a_23069_n6459# a_24056_n6231# a_24007_n6215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6648 vdd d2 a_13030_n7091# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6649 a_29063_n6256# a_29068_n5519# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6650 a_21699_n4767# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6651 vdd d0 a_29321_2234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6652 gnd d2 a_23184_n9273# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6653 vdd d0 a_34296_3301# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6654 a_27050_n5930# a_26723_n8130# a_27045_n7953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6655 gnd d1 a_8198_1394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6656 a_25359_7904# a_25359_7447# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6657 a_32112_486# a_31899_486# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6658 a_30335_4789# a_30335_4559# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6659 a_15518_n9526# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6660 a_648_n1759# a_435_n1759# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6661 vdd d0 a_14108_n7358# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6662 vdd a_24265_2193# a_24057_2193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6663 a_10150_n3330# a_10679_n3421# a_10887_n3421# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6664 vdd d0 a_39352_6102# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6665 a_2776_n7972# a_3029_n8176# a_2778_n5760# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6666 gnd a_4077_9384# a_3869_9384# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6667 a_30334_n8826# a_30334_n8597# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6668 a_17971_n4318# a_18228_n4334# a_17830_n4910# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6669 a_31070_n8363# a_31801_n8673# a_32009_n8673# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6670 a_21996_3096# a_21882_2977# a_21989_5189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6671 a_20833_3246# a_20620_3246# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6672 a_24009_8824# a_24262_8811# a_23067_9245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6673 a_33100_5941# a_34087_5507# a_34042_5520# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6674 a_10464_4373# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6675 a_36644_n8714# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6676 gnd a_29319_n7375# a_29111_n7375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6677 a_26096_8253# a_25675_8253# a_25359_8134# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6678 a_117_8112# a_117_7882# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6679 a_20303_6990# a_20832_7109# a_21040_7109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6680 a_15522_3865# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6681 a_37066_5808# a_36645_5808# a_36127_5498# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6682 a_5172_n9984# a_5701_n10075# a_5909_n10075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6683 a_12913_n7586# a_13900_n7358# a_13851_n7342# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6684 a_24009_n3460# a_24012_n2718# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6685 a_16880_n6527# a_16459_n6527# a_15942_n6771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6686 a_38159_6908# a_39143_7205# a_39098_7218# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6687 a_6849_5822# a_6781_6333# a_6859_7449# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6688 vdd d0 a_9134_n7948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6689 a_17976_n1924# a_18229_n2128# a_17831_n2704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6690 a_3827_n1634# a_4080_n1838# a_2885_n2066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6691 a_25360_5054# a_25360_4825# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6692 a_20303_n8592# a_20832_n8912# a_21040_n8912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6693 a_39100_n3318# a_39096_n3506# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6694 vdd a_13032_1950# a_12824_1950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6695 a_32964_4150# a_33217_4137# a_32995_3034# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6696 vdd d1 a_33358_2442# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6697 a_35921_n4546# a_35708_n4546# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6698 a_39099_2252# a_39095_2429# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6699 a_8881_n4984# a_9134_n5188# a_7939_n5416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6700 a_20831_n7255# a_20618_n7255# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6701 a_15520_7174# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6702 a_25674_6596# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6703 a_38017_n2685# a_38207_n2109# a_38158_n2093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6704 a_37064_9117# a_36643_9117# a_36126_9361# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6705 a_10887_3824# a_11617_3580# a_11825_3580# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6706 a_6848_n8728# a_6427_n8728# a_5909_n8418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6707 a_7798_6588# a_7988_5806# a_7943_5819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6708 a_39099_n2764# a_39352_n2968# a_38157_n3196# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6709 a_33105_2455# a_34089_2752# a_34040_2942# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6710 a_6641_n5419# a_6428_n5419# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6711 a_15205_n6867# a_15205_n6680# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6712 gnd d0 a_9134_n6291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6713 gnd a_34294_7713# a_34086_7713# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6714 a_39099_6115# a_39095_6292# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6715 a_8879_1340# a_5178_1206# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6716 a_5909_7718# a_5488_7718# a_5173_7923# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6717 a_24007_8452# a_24010_7721# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6718 a_16895_7573# a_16781_7454# a_16895_5373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6719 a_13858_3887# a_14111_3874# a_12919_3577# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6720 a_32961_n2644# a_33218_n2660# a_32991_n3734# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6721 a_11403_4683# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6722 a_25360_4595# a_25888_4390# a_26096_4390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6723 a_11403_n5383# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6724 a_21039_9315# a_20618_9315# a_20302_9425# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6725 a_36126_n10061# a_36856_n9817# a_37064_n9817# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6726 a_119_3700# a_648_3819# a_856_3819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6727 a_2748_n2470# a_2933_n3185# a_2884_n3169# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6728 a_1808_7527# a_1694_7408# a_1808_5327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6729 a_34042_n6032# a_34295_n6236# a_33100_n6464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6730 a_6782_n4827# a_6569_n4827# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6731 vdd a_3140_5765# a_2932_5765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6732 a_12917_n8501# a_13901_n9015# a_13856_n8811# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6733 a_22932_n6863# a_23185_n7067# a_22958_n8141# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6734 a_8880_6678# a_8876_6855# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6735 a_36128_4949# a_35707_4949# a_35391_4830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6736 a_11824_n6486# a_11403_n6486# a_10885_n6176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6737 a_2103_500# a_4845_480# a_5053_480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6738 a_2882_7058# a_3869_6624# a_3824_6637# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6739 gnd a_4079_4972# a_3871_4972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6740 gnd a_29321_n6826# a_29113_n6826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6741 a_118_5906# a_118_5676# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6742 a_646_5471# a_433_5471# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6743 a_26967_n7014# a_26754_n7014# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6744 a_31802_n6467# a_31589_n6467# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6745 a_26613_6906# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6746 a_29062_n8462# a_29319_n8478# a_28124_n8706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6747 a_5174_6363# a_5174_6176# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6748 a_30651_3251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6749 vdd d0 a_19164_6670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6750 a_12918_5783# a_13902_6080# a_13853_6270# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6751 a_36754_n8135# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6752 a_28124_8183# a_28381_7993# a_27983_8775# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6753 a_34044_n3277# a_34297_n3481# a_33105_n2967# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6754 a_18911_9443# a_18907_9620# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6755 a_6851_1410# a_6783_1921# a_6861_3037# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6756 a_8883_n4435# a_9136_n4639# a_7944_n4125# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6757 a_2887_4675# a_3140_4662# a_2747_4164# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6758 a_20833_n6706# a_20620_n6706# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6759 a_23074_2450# a_23327_2437# a_22934_1939# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6760 a_2746_6370# a_2999_6357# a_2772_7637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6761 a_434_n2862# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6762 a_21770_n8668# a_21557_n8668# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6763 a_22929_n4845# a_23119_n4269# a_23070_n4253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6764 a_12917_n7398# a_13170_n7602# a_12777_n6887# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6765 gnd a_24264_n7888# a_24056_n7888# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6766 a_25676_2184# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6767 a_10676_6579# a_10463_6579# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6768 a_32010_5767# a_31589_5767# a_31072_6011# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6769 a_117_n7278# a_645_n7274# a_853_n7274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6770 a_21773_1350# a_21560_1350# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6771 a_32011_2458# a_31590_2458# a_31072_2148# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6772 a_39100_3909# a_39096_4086# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6773 a_24008_6246# a_24011_5515# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6774 vdd d0 a_29321_n5723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6775 a_433_7128# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6776 a_30649_n7260# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6777 gnd d1 a_13170_n8705# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6778 a_34041_n2362# a_34044_n1620# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6779 vdd d1 a_33356_n7583# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6780 a_5488_n8418# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6781 a_16897_3161# a_16783_3042# a_16890_5254# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6782 a_1791_9090# a_1724_8498# a_1808_7527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6783 vdd d1 a_8195_n8741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6784 a_32958_n9262# a_33215_n9278# a_32993_n7958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6785 a_35393_1750# a_35393_1521# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6786 a_13857_6093# a_13853_6270# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6787 vdd a_4077_9384# a_3869_9384# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6788 a_21979_n5359# a_21912_n4767# a_21996_n3677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6789 a_31072_n2848# a_30651_n2848# a_30336_n2852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6790 a_6861_n3560# a_6570_n2621# a_6850_n3213# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6791 gnd d0 a_29318_n9581# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6792 a_11725_n5913# a_11512_n5913# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6793 a_36859_3602# a_36646_3602# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6794 a_15732_9380# a_15519_9380# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6795 a_16880_n6527# a_16812_n7038# a_16890_n7977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6796 gnd d0 a_29322_n3517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6797 a_36129_3846# a_35708_3846# a_35392_3956# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6798 vdd d0 a_14110_4977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6799 a_36969_n3723# a_36756_n3723# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6800 a_29065_n3501# a_29068_n2759# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6801 a_35707_n6752# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6802 a_26828_n4297# a_26615_n4297# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6803 gnd a_28380_9096# a_28172_9096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6804 a_20617_n9461# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6805 a_32011_n4261# a_31590_n4261# a_31073_n4505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6806 a_17973_6927# a_18226_6914# a_17833_6416# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6807 a_2886_7984# a_3139_7971# a_2741_8753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6808 a_35391_4600# a_35392_4143# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6809 a_36857_6911# a_36644_6911# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6810 a_3821_5711# a_3826_4985# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6811 a_20305_n3077# a_20305_n2847# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6812 gnd d1 a_38414_2483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6813 a_26614_5803# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6814 a_12703_n10661# a_12653_n10677# a_12604_n10661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6815 a_5175_2408# a_5176_1951# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6816 a_8881_4472# a_9134_4459# a_7939_4893# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6817 a_11615_6889# a_11402_6889# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6818 gnd d1 a_18229_1399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6819 a_5911_n5663# a_5490_n5663# a_5174_n5343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6820 a_5703_n2903# a_5490_n2903# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6821 vdd d0 a_19166_2258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6822 a_13855_7745# a_14108_7732# a_12913_8166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6823 a_32027_3101# a_31730_4072# a_32011_3561# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6824 a_12803_n8165# a_12822_n7091# a_12777_n6887# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6825 a_33105_2455# a_34089_2752# a_34044_2765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6826 a_16599_6338# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6827 a_20304_n6615# a_20304_n6386# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6828 a_29062_n10119# a_29319_n10135# a_28127_n9621# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6829 vdd a_34294_n10099# a_34086_n10099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6830 a_33099_n7567# a_34086_n7339# a_34037_n7323# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6831 a_5704_n3457# a_5491_n3457# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6832 gnd a_33358_2442# a_33150_2442# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6833 vdd a_39350_n8483# a_39142_n8483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6834 gnd a_34294_n10099# a_34086_n10099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6835 vdd a_34294_7713# a_34086_7713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6836 a_7799_n4905# a_8056_n4921# a_7834_n3601# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6837 a_8879_2997# a_9136_2807# a_7944_2510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6838 a_11615_n7589# a_11402_n7589# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6839 a_1805_n3519# a_1514_n2580# a_1795_n2069# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6840 gnd d0 a_4078_7178# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6841 a_20303_6760# a_20831_6555# a_21039_6555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6842 a_36967_5235# a_36754_5235# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6843 a_118_n6634# a_647_n6725# a_855_n6725# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6844 a_25362_n2431# a_25889_n2884# a_26097_n2884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6845 a_9888_364# a_9779_364# a_9987_364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6846 vdd a_19167_3915# a_18959_3915# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6847 gnd a_13173_1358# a_12965_1358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6848 a_10150_4121# a_10150_3934# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6849 a_38051_n5787# a_38094_n8203# a_38049_n7999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6850 a_10678_2167# a_10465_2167# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6851 a_17833_n6928# a_18018_n7643# a_17969_n7627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6852 a_32012_1355# a_31591_1355# a_31074_1599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6853 a_6848_6925# a_6427_6925# a_5910_7169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6854 a_30863_5457# a_30650_5457# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6855 a_434_6025# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6856 gnd a_8196_5806# a_7988_5806# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6857 a_12807_n7977# a_13060_n8181# a_12809_n5765# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6858 a_6539_n3737# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6859 a_10466_n3421# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6860 vdd a_4080_n4598# a_3872_n4598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6861 a_35707_2189# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6862 a_29070_n2210# a_29323_n2414# a_28131_n1900# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6863 a_31588_n8673# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6864 a_15736_1659# a_15523_1659# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6865 a_7938_7099# a_8925_6665# a_8876_6855# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6866 gnd a_4077_n7353# a_3869_n7353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6867 a_13858_3887# a_13854_4064# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6868 gnd d3 a_8085_7488# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6869 a_1793_4678# a_1726_4086# a_1810_3115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6870 a_33105_n4070# a_33358_n4274# a_32960_n4850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6871 a_27047_n3541# a_26938_n3718# a_27045_n5753# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6872 a_20833_4903# a_20620_4903# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6873 a_10887_n4524# a_10466_n4524# a_10150_n4204# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6874 vdd d3 a_33246_n8162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6875 a_25140_461# a_26924_522# a_27246_522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6876 a_5488_n10075# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6877 a_5701_6615# a_5488_6615# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6878 a_15734_4968# a_15521_4968# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6879 a_25888_4390# a_25675_4390# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6880 a_26969_1902# a_26756_1902# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6881 gnd a_23325_n8681# a_23117_n8681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6882 a_7942_n7434# a_8926_n7948# a_8881_n7744# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6883 gnd d1 a_23325_7952# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6884 a_20619_n8912# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6885 a_12918_5783# a_13902_6080# a_13857_6093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6886 a_24014_1657# a_24267_1644# a_23075_1347# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6887 a_21994_n8089# a_21697_n9179# a_21977_n9771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6888 a_21038_8761# a_20617_8761# a_20303_8509# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6889 a_8877_n9035# a_8880_n8293# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6890 a_36646_n3199# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6891 a_15206_2413# a_15207_1956# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6892 a_30333_n9700# a_30862_n10020# a_31070_n10020# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6893 gnd a_3029_7447# a_2821_7447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6894 a_36859_n4302# a_36646_n4302# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6895 vdd a_18118_n3810# a_17910_n3810# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6896 a_1585_n5378# a_1372_n5378# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6897 a_26616_1391# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6898 vdd a_33356_6854# a_33148_6854# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6899 a_20305_n2847# a_20833_n2843# a_21041_n2843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6900 a_2883_4852# a_3140_4662# a_2747_4164# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6901 vdd d1 a_13172_n3190# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6902 a_11617_2477# a_11404_2477# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6903 a_15206_n4661# a_15733_n5114# a_15941_n5114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6904 gnd a_19164_6670# a_18956_6670# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6905 a_7939_n6519# a_8926_n6291# a_8877_n6275# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6906 a_1371_n8687# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6907 a_22931_8557# a_23116_9055# a_23067_9245# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6908 a_5700_n9521# a_5487_n9521# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6909 a_5488_9375# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6910 a_36967_7435# a_36754_7435# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6911 a_1803_7408# a_1512_6292# a_1793_5781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6912 a_5175_3970# a_5175_3741# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6913 a_10149_n6180# a_10149_n5723# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6914 a_118_6322# a_645_6574# a_853_6574# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6915 a_10151_n1998# a_10151_n1768# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6916 a_35393_1937# a_35920_2189# a_36128_2189# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6917 vdd d0 a_29322_2788# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6918 a_36127_n5095# a_35706_n5095# a_35391_n5099# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6919 a_433_n8931# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6920 a_20304_5200# a_20832_5452# a_21040_5452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6921 a_20304_6303# a_20304_6116# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6922 a_25361_n2888# a_25362_n2431# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6923 vdd a_34296_3301# a_34088_3301# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6924 a_31800_9076# a_31587_9076# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6925 a_10151_1915# a_10151_1728# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6926 a_33099_8147# a_34086_7713# a_34037_7903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6927 a_1808_n8108# a_1511_n9198# a_1792_n8687# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6928 a_38156_5982# a_39143_5548# a_39098_5561# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6929 a_20305_2348# a_20833_2143# a_21041_2143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6930 a_6640_6925# a_6427_6925# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6931 a_30865_1045# a_30652_1045# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6932 a_32960_n4850# a_33150_n4274# a_33105_n4070# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6933 a_31698_7394# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6934 a_18913_6134# a_19166_6121# a_17974_5824# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6935 gnd a_8198_1394# a_7990_1394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6936 a_36955_527# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6937 a_25359_7031# a_25888_7150# a_26096_7150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6938 gnd d0 a_39354_1690# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6939 a_16882_1415# a_16814_1926# a_16892_3042# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6940 a_30334_8098# a_30863_8217# a_31071_8217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6941 a_12805_n5953# a_13062_n5969# a_12604_n10661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6942 a_3820_n8440# a_4077_n8456# a_2882_n8684# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6943 a_2746_6370# a_2931_6868# a_2886_6881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6944 a_33102_n9585# a_34086_n10099# a_34037_n10083# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6945 a_28125_n6500# a_29112_n6272# a_29063_n6256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6946 a_1794_n4275# a_1726_n4786# a_1810_n3696# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6947 a_7940_2687# a_8927_2253# a_8878_2443# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6948 a_6429_n4316# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6949 a_17865_n3606# a_17879_n4926# a_17830_n4910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6950 gnd d3 a_8087_3076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6951 gnd d1 a_33357_4648# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6952 a_31071_n8917# a_30650_n8917# a_30334_n8826# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6953 vdd a_39352_6102# a_39144_6102# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6954 a_13853_n2930# a_14110_n2946# a_12915_n3174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6955 vdd d1 a_38414_2483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6956 a_36647_n2096# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6957 a_20620_3246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6958 gnd a_39351_n7934# a_39143_n7934# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6959 a_26095_n10056# a_25674_n10056# a_25358_n9965# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6960 a_10676_n8382# a_10463_n8382# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6961 a_39092_n9570# a_39349_n9586# a_38154_n9814# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6962 a_5703_2203# a_5490_2203# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6963 a_10149_n6180# a_10677_n6176# a_10885_n6176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6964 a_38161_2496# a_39145_2793# a_39096_2983# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6965 a_15203_9490# a_15203_9261# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6966 a_21041_4903# a_21771_4659# a_21979_4659# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6967 a_13851_7922# a_14108_7732# a_12913_8166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6968 vdd d0 a_14110_n4049# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6969 a_13855_n7154# a_13851_n7342# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6970 a_24007_n7872# a_24010_n7130# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6971 a_29070_1698# a_29066_1875# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6972 a_1727_1880# a_1514_1880# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6973 gnd a_3031_3035# a_2823_3035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6974 a_35391_n6661# a_35920_n6752# a_36128_n6752# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6975 a_15206_n3371# a_15735_n3462# a_15943_n3462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6976 a_36128_n3992# a_35707_n3992# a_35392_n3539# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6977 a_11618_1374# a_11405_1374# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6978 vdd a_33358_2442# a_33150_2442# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6979 a_20302_n9465# a_20830_n9461# a_21038_n9461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6980 a_18912_n4989# a_18908_n5177# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6981 a_16897_3161# a_16600_4132# a_16880_4724# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6982 a_33102_9073# a_33355_9060# a_32962_8562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6983 a_15206_3975# a_15206_3746# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X6984 a_31800_n9776# a_31587_n9776# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6985 a_32964_n4662# a_33149_n5377# a_33100_n5361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6986 a_30650_n5054# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6987 a_36647_1396# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6988 a_12772_n9281# a_12962_n8705# a_12913_n8689# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6989 a_27036_n3194# a_26615_n3194# a_26097_n2884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6990 a_36129_n4546# a_35708_n4546# a_35392_n4455# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6991 a_28126_n4294# a_28383_n4310# a_27985_n4886# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6992 a_36969_3023# a_36756_3023# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6993 a_120_1910# a_647_2162# a_855_2162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6994 a_12917_7989# a_13170_7976# a_12772_8758# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6995 a_31801_7973# a_31588_7973# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6996 gnd d0 a_4076_n9559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6997 a_21699_n4767# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6998 vdd a_23327_n3166# a_23119_n3166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X6999 a_28014_7659# a_28271_7469# a_28020_5270# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7000 a_6537_n5949# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7001 a_18914_n4440# a_18910_n4628# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7002 a_7938_7099# a_8925_6665# a_8880_6678# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7003 a_24007_5692# a_24012_4966# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7004 a_25359_n8633# a_25888_n8953# a_26096_n8953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7005 vdd a_10033_n10854# a_9825_n10854# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7006 vdd d5 a_28072_n10694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7007 a_16599_n7038# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7008 a_5176_1764# a_5705_1654# a_5913_1654# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7009 a_6641_5822# a_6428_5822# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7010 a_25361_2389# a_25362_1932# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7011 a_26828_3597# a_26615_3597# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7012 a_21978_6865# a_21557_6865# a_21039_6555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7013 a_16459_4724# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7014 a_32790_n10642# a_33047_n10658# a_32889_n10642# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7015 gnd a_3140_n5391# a_2932_n5391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7016 a_6642_2513# a_6429_2513# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7017 a_15940_9380# a_16670_9136# a_16878_9136# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7018 a_6848_n7625# a_6781_n7033# a_6859_n7972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7019 a_35390_n8638# a_35390_n8408# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7020 a_29752_345# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7021 a_24010_1834# a_24267_1644# a_23075_1347# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7022 a_3823_4059# a_4080_3869# a_2888_3572# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7023 a_18910_4105# a_18913_3374# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7024 a_31071_n8917# a_31801_n8673# a_32009_n8673# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7025 a_23072_7965# a_24056_8262# a_24007_8452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7026 a_433_5471# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7027 a_3820_n10097# a_4077_n10113# a_2885_n9599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7028 a_36644_n8714# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7029 a_35393_n1790# a_35016_n1511# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7030 a_21996_3096# a_21699_4067# a_21979_4659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7031 a_21041_3246# a_21772_3556# a_21980_3556# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7032 a_28130_3594# a_28383_3581# a_27985_4363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7033 vdd a_19164_6670# a_18956_6670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7034 a_39096_8870# a_39349_8857# a_38154_9291# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7035 a_22931_8557# a_23116_9055# a_23071_9068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7036 a_24007_n6215# a_24264_n6231# a_23069_n6459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7037 a_5912_3860# a_5491_3860# a_5175_3741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7038 a_27988_n6904# a_28241_n7108# a_28014_n8182# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7039 a_37067_n3199# a_36646_n3199# a_36128_n2889# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7040 vdd a_34298_n2378# a_34090_n2378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7041 a_16880_n6527# a_16459_n6527# a_15941_n6217# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7042 a_25676_n2884# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7043 a_20303_n8821# a_20832_n8912# a_21040_n8912# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7044 gnd a_34295_n5133# a_34087_n5133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7045 a_26936_5230# a_26723_5230# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7046 a_33099_8147# a_34086_7713# a_34041_7726# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7047 a_21994_n5889# a_21880_n5889# a_22088_n5889# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7048 a_3828_n2188# a_4081_n2392# a_2889_n1878# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7049 a_10463_6579# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7050 gnd a_19167_n3541# a_18959_n3541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7051 gnd d2 a_3001_n2674# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7052 a_21560_1350# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7053 gnd a_3141_3559# a_2933_3559# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7054 a_18909_6311# a_19166_6121# a_17974_5824# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7055 a_2883_n5375# a_3140_n5391# a_2747_n4676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7056 a_21911_6273# a_21698_6273# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7057 a_28016_3247# a_28273_3057# a_28016_5447# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7058 a_21979_5762# a_21558_5762# a_21041_6006# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7059 a_34039_n6774# a_34042_n6032# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7060 a_7940_2687# a_8927_2253# a_8882_2266# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7061 a_6848_8028# a_6780_8539# a_6864_7568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7062 a_35918_7704# a_35705_7704# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7063 a_3827_1122# a_4080_1109# a_2885_1543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7064 vdd d3 a_8087_3076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7065 a_15940_7723# a_16671_8033# a_16879_8033# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7066 a_26096_n5090# a_26827_n5400# a_27035_n5400# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7067 vdd d0 a_19165_n6296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7068 a_17831_n2704# a_18021_n2128# a_17976_n1924# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7069 a_20305_3910# a_20305_3681# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7070 gnd d0 a_19165_4464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7071 vdd d1 a_3140_n6494# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7072 a_10886_6030# a_11616_5786# a_11824_5786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7073 a_5173_n7965# a_5701_n8418# a_5909_n8418# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7074 gnd a_33355_n9789# a_33147_n9789# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7075 a_31073_3805# a_30652_3805# a_30336_3686# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7076 a_29063_n7913# a_29066_n7171# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7077 a_12779_n2475# a_12964_n3190# a_12919_n2986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7078 a_15207_n2455# a_15734_n2908# a_15942_n2908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7079 gnd a_33248_n3750# a_33040_n3750# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7080 gnd a_28072_n10694# a_27864_n10694# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7081 a_15733_n8977# a_15520_n8977# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7082 gnd a_38414_2483# a_38206_2483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7083 vdd d1 a_38412_n7624# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7084 vdd d0 a_34297_1095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7085 vdd a_3031_3035# a_2823_3035# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7086 a_23074_3553# a_24058_3850# a_24009_4040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7087 a_20303_6760# a_20304_6303# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7088 a_31071_7114# a_30650_7114# a_30334_7224# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7089 a_25359_6801# a_25887_6596# a_26095_6596# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7090 a_17973_8030# a_18957_8327# a_18912_8340# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7091 a_30334_7868# a_30862_7663# a_31070_7663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7092 a_11402_6889# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7093 a_10885_n7833# a_10464_n7833# a_10148_n7742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7094 a_16781_n5954# a_16568_n5954# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7095 a_5174_n5113# a_5702_n5109# a_5910_n5109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7096 vdd d2 a_38271_8590# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7097 a_33098_9250# a_33355_9060# a_32962_8562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7098 vdd a_19166_2258# a_18958_2258# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7099 a_18906_n9589# a_19163_n9605# a_17968_n9833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7100 a_7938_7099# a_8195_6909# a_7802_6411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7101 gnd d1 a_38413_n5418# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7102 a_5174_n5343# a_5703_n5663# a_5911_n5663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7103 a_7830_n5989# a_7879_n3805# a_7834_n3601# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7104 a_32012_n2055# a_31944_n2566# a_32022_n3505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7105 a_35919_n6198# a_35706_n6198# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7106 a_34037_9560# a_34040_8829# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7107 a_434_n2862# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7108 a_15204_n8657# a_15204_n8427# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7109 a_10679_2721# a_10466_2721# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7110 gnd a_4078_7178# a_3870_7178# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7111 a_5173_8569# a_5700_8821# a_5908_8821# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7112 a_15204_7055# a_15733_7174# a_15941_7174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7113 a_36754_5235# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7114 a_1810_3115# a_1696_2996# a_1803_5208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7115 a_645_7677# a_432_7677# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7116 a_20834_1040# a_20621_1040# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7117 a_33101_3735# a_34088_3301# a_34043_3314# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7118 gnd a_23187_n2655# a_22979_n2655# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7119 a_7802_n6923# a_7987_n7638# a_7938_n7622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7120 a_120_n2409# a_120_n2222# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7121 a_10465_2167# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7122 a_10151_1499# a_10151_1269# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7123 a_35708_2743# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7124 a_8877_7409# a_8880_6678# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7125 a_26097_6047# a_25676_6047# a_25360_5928# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7126 gnd a_38272_n7113# a_38064_n7113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7127 a_30650_5457# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7128 a_1513_n4786# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7129 vdd d0 a_19163_8876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7130 gnd d0 a_14111_2771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7131 gnd d1 a_28381_7993# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7132 a_12917_7989# a_13901_8286# a_13852_8476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7133 a_24012_n5478# a_24265_n5682# a_23073_n5168# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7134 a_29070_1698# a_29323_1685# a_28131_1388# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7135 a_15523_1659# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7136 a_118_6135# a_118_5906# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7137 a_18912_4477# a_18908_4654# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7138 a_23070_n3150# a_24057_n2922# a_24008_n2906# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7139 a_38155_n7608# a_39142_n7380# a_39093_n7364# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7140 a_6850_3616# a_6782_4127# a_6866_3156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7141 a_27987_n9110# a_28172_n9825# a_28127_n9621# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7142 a_10464_n6176# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7143 a_648_n1759# a_435_n1759# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7144 a_6861_n3560# a_6570_n2621# a_6851_n2110# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7145 a_20620_4903# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7146 a_16671_n7630# a_16458_n7630# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7147 a_23072_7965# a_24056_8262# a_24011_8275# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7148 a_12777_6375# a_13030_6362# a_12803_7642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7149 a_11725_n5913# a_11512_n5913# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7150 a_10887_n4524# a_11617_n4280# a_11825_n4280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7151 a_12915_n4277# a_13902_n4049# a_13857_n3845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7152 vdd d1 a_13171_4667# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7153 gnd d0 a_24265_n6785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7154 a_15521_4968# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7155 a_25675_4390# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7156 a_6958_5249# a_6951_541# a_4954_480# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7157 a_26756_1902# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7158 a_36127_n5095# a_36858_n5405# a_37066_n5405# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7159 a_10888_1618# a_11618_1374# a_11826_1374# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7160 a_28126_3771# a_28383_3581# a_27985_4363# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7161 gnd a_23325_7952# a_23117_7952# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7162 a_11839_n5913# a_11512_n8113# a_11839_n8113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7163 a_35707_n6752# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7164 gnd a_18228_n4334# a_18020_n4334# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7165 a_36969_n3723# a_36756_n3723# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7166 a_17831_2181# a_18021_1399# a_17976_1412# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7167 a_20617_n9461# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7168 a_32011_n4261# a_31590_n4261# a_31072_n3951# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7169 a_8879_n1863# a_9136_n1879# a_7941_n2107# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7170 a_27988_n6904# a_28173_n7619# a_28124_n7603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7171 gnd d0 a_34294_n7339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7172 gnd a_9133_n7394# a_8925_n7394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7173 a_2887_n5187# a_3871_n5701# a_3826_n5497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7174 vdd d1 a_23324_n9784# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7175 a_31911_n8094# a_31698_n8094# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7176 a_6427_n7625# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7177 a_38161_n4111# a_38414_n4315# a_38016_n4891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7178 a_25888_8253# a_25675_8253# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7179 a_13858_1127# a_13854_1304# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7180 vdd a_24264_n5128# a_24056_n5128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7181 a_38155_8188# a_39142_7754# a_39093_7944# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7182 gnd a_18118_n6010# a_17910_n6010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7183 vdd d3 a_23217_n3745# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7184 a_7944_n3022# a_8197_n3226# a_7804_n2511# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7185 a_25361_2389# a_25889_2184# a_26097_2184# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7186 vdd d2 a_23185_6338# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7187 a_31804_n2055# a_31591_n2055# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7188 a_11404_2477# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7189 vdd d3 a_38302_n8203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7190 gnd d2 a_38274_n2701# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7191 gnd d0 a_19166_n5747# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7192 a_36858_5808# a_36645_5808# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7193 a_2881_n9787# a_3868_n9559# a_3819_n9543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7194 a_6848_n8728# a_6427_n8728# a_5910_n8972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7195 a_36754_7435# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7196 a_6859_7449# a_6568_6333# a_6848_6925# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7197 a_25675_n8953# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7198 a_21042_n4500# a_20621_n4500# a_20305_n4180# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7199 gnd d5 a_17917_n10718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7200 vdd a_29322_2788# a_29114_2788# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7201 a_7940_2687# a_8197_2497# a_7804_1999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7202 a_39095_n6815# a_39098_n6073# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7203 a_5704_n3457# a_5491_n3457# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7204 a_25890_3841# a_25677_3841# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7205 a_36856_9117# a_36643_9117# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7206 a_20619_8212# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7207 gnd d1 a_38413_4689# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7208 a_6568_n7033# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7209 a_8879_n3520# a_8882_n2778# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7210 a_8878_5203# a_8881_4472# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7211 a_856_n1759# a_1587_n2069# a_1795_n2069# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7212 a_647_3265# a_434_3265# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7213 a_35391_6162# a_35920_6052# a_36128_6052# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7214 gnd a_23184_n9273# a_22976_n9273# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7215 vdd a_28273_n3786# a_28065_n3786# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7216 a_30652_1045# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7217 a_21769_9071# a_21556_9071# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7218 a_32020_7394# a_31729_6278# a_32010_5767# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7219 vdd d0 a_19165_4464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7220 a_17975_2515# a_18228_2502# a_17835_2004# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7221 a_16895_5373# a_16568_7454# a_16890_7454# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7222 a_12919_3577# a_13903_3874# a_13854_4064# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7223 a_7834_n5801# a_7877_n8217# a_7828_n8201# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7224 a_31588_n8673# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7225 a_17972_n9645# a_18956_n10159# a_15203_n10176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7226 gnd a_14109_n6255# a_13901_n6255# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7227 gnd a_39354_1690# a_39146_1690# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7228 a_38160_n6317# a_39144_n6831# a_39095_n6815# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7229 a_10147_n9489# a_10675_n9485# a_10883_n9485# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7230 gnd d0 a_9135_n2982# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7231 a_23067_n9768# a_24054_n9540# a_24005_n9524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7232 gnd a_33357_4648# a_33149_4648# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7233 vdd a_38414_2483# a_38206_2483# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7234 a_645_n8377# a_432_n8377# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7235 a_2888_2469# a_3141_2456# a_2748_1958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7236 a_34038_8457# a_34295_8267# a_33103_7970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7237 a_1808_5327# a_1481_7408# a_1803_7408# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7238 a_5911_n4006# a_5490_n4006# a_5175_n4010# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7239 a_27037_n2091# a_26616_n2091# a_26099_n2335# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7240 a_12779_1963# a_13032_1950# a_12805_3230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7241 a_38158_9114# a_38411_9101# a_38018_8603# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7242 a_11758_1885# a_11545_1885# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7243 a_5490_2203# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7244 a_20619_n8912# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7245 vdd a_29321_6097# a_29113_6097# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7246 gnd a_9135_n6845# a_8927_n6845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7247 a_6781_n7033# a_6568_n7033# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7248 a_8876_n8481# a_9133_n8497# a_7938_n8725# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7249 a_25358_n10152# a_29319_n10135# a_28127_n9621# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7250 a_21667_n5889# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7251 a_36859_n4302# a_36646_n4302# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7252 gnd a_14111_n3500# a_13903_n3500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7253 a_1514_1880# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7254 a_23073_n6271# a_23326_n6475# a_22928_n7051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7255 a_646_n5068# a_433_n5068# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7256 a_11405_1374# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7257 a_20305_n3950# a_20305_n3493# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7258 vdd a_29320_n7929# a_29112_n7929# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7259 vdd a_8194_n9844# a_7986_n9844# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7260 a_38157_3776# a_39144_3342# a_39095_3532# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7261 a_18910_n9401# a_18906_n9589# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7262 a_30334_n7723# a_30334_n7494# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7263 a_1725_n6992# a_1512_n6992# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7264 a_21994_5308# a_21667_7389# a_21989_7389# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7265 a_36756_3023# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7266 vdd d0 a_14111_2771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7267 a_2747_4164# a_2932_4662# a_2883_4852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7268 a_12917_7989# a_13901_8286# a_13856_8299# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7269 a_433_n8931# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7270 a_17970_n6524# a_18957_n6296# a_18912_n6092# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7271 a_26614_n5400# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7272 a_31070_6560# a_30649_6560# a_30335_6308# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7273 a_15523_n2359# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7274 a_29066_1875# a_29323_1685# a_28131_1388# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7275 a_15518_8826# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7276 a_11824_4683# a_11403_4683# a_10886_4927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7277 a_18912_n8852# a_18908_n9040# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7278 a_17974_n5233# a_18227_n5437# a_17834_n4722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7279 a_30649_n7260# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7280 a_6864_n5949# a_6537_n8149# a_6864_n8149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7281 a_2742_n7070# a_2932_n6494# a_2887_n6290# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7282 a_26615_3597# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7283 a_28128_8006# a_29112_8303# a_29063_8493# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7284 a_5488_n8418# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7285 a_26096_8253# a_26826_8009# a_27034_8009# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7286 a_120_n1993# a_649_n2313# a_857_n2313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7287 a_34896_n10703# a_37895_n10699# a_37175_n5935# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7288 a_12773_6552# a_13030_6362# a_12803_7642# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7289 a_2103_500# a_1682_500# a_2004_500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7290 gnd d1 a_18227_n6540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7291 a_13856_5539# a_14109_5526# a_12914_5960# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7292 a_35919_n8958# a_35706_n8958# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7293 gnd a_33359_n2068# a_33151_n2068# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7294 a_1808_7527# a_1511_8498# a_1792_7987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7295 a_26095_n7296# a_25674_n7296# a_25359_n7300# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7296 a_117_8528# a_644_8780# a_852_8780# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7297 a_37067_2499# a_37000_1907# a_37078_3023# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7298 a_38045_n8187# a_38064_n7113# a_38019_n6909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7299 a_15205_n5764# a_15205_n5577# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7300 gnd d0 a_9132_n9600# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7301 a_6639_n9831# a_6426_n9831# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7302 a_26099_1635# a_26829_1391# a_27037_1391# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7303 a_31071_n8917# a_30650_n8917# a_30334_n8597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7304 a_29062_n10119# a_29065_n9377# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7305 a_5489_n5109# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7306 a_20303_7406# a_20831_7658# a_21039_7658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7307 a_39099_5012# a_39095_5189# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7308 a_24007_7349# a_24010_6618# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7309 a_30334_8098# a_30334_7868# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7310 a_38155_8188# a_39142_7754# a_39097_7767# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7311 a_20304_4554# a_20832_4349# a_21040_4349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7312 a_10148_8117# a_10148_7887# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7313 vdd d2 a_2998_n9292# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7314 a_34039_n6774# a_34296_n6790# a_33104_n6276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7315 a_13854_n3484# a_14111_n3500# a_12919_n2986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7316 a_1794_n3172# a_1373_n3172# a_856_n3416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7317 a_5911_2203# a_6642_2513# a_6850_2513# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7318 a_18912_8340# a_19165_8327# a_17973_8030# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7319 a_34040_n9341# a_34293_n9545# a_33098_n9773# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7320 a_22190_481# a_23009_5216# a_22960_5406# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7321 vdd d2 a_33216_n7072# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7322 a_11822_n9795# a_11401_n9795# a_10883_n9485# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7323 a_7939_4893# a_8926_4459# a_8877_4649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7324 a_29061_9042# a_29067_8316# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7325 a_26723_5230# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7326 a_12807_7465# a_12821_8568# a_12776_8581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7327 a_13855_n7154# a_14108_n7358# a_12913_n7586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7328 vdd d0 a_14111_n4603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7329 a_5173_n9068# a_5173_n8881# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7330 a_27986_2157# a_28243_1967# a_28016_3247# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7331 a_15941_n6217# a_16672_n6527# a_16880_n6527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7332 a_31800_n9776# a_31587_n9776# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7333 a_118_4803# a_118_4573# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7334 a_17859_n8206# a_18116_n8222# a_17865_n5806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7335 a_36129_n4546# a_35708_n4546# a_35392_n4226# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7336 vdd a_4079_n4044# a_3871_n4044# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7337 a_32025_7513# a_31911_7394# a_32025_5313# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7338 a_5702_4409# a_5489_4409# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7339 a_6783_1921# a_6570_1921# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7340 gnd a_8056_n4921# a_7848_n4921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7341 a_39098_5561# a_39094_5738# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7342 gnd d0 a_14108_n8461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7343 gnd d1 a_3139_7971# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7344 a_7944_2510# a_8928_2807# a_8883_2820# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7345 a_10676_7682# a_10463_7682# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7346 a_3828_1676# a_4081_1663# a_2889_1366# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7347 a_21039_6555# a_20618_6555# a_20304_6303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7348 a_25359_n8862# a_25888_n8953# a_26096_n8953# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7349 a_8881_n7744# a_9134_n7948# a_7942_n7434# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7350 a_35705_7704# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7351 a_20831_n10015# a_20618_n10015# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7352 a_28130_3594# a_29114_3891# a_29065_4081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7353 a_11617_3580# a_11404_3580# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7354 a_2884_2646# a_3141_2456# a_2748_1958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7355 a_22932_n6863# a_23117_n7578# a_23068_n7562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7356 a_27050_n5930# a_26936_n5930# a_27144_n5930# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7357 vdd a_3001_1945# a_2793_1945# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7358 a_16890_7454# a_16599_6338# a_16879_6930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7359 gnd a_19165_4464# a_18957_4464# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7360 a_26097_n6747# a_25676_n6747# a_25360_n6656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7361 a_11756_n6997# a_11543_n6997# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7362 a_22932_6351# a_23117_6849# a_23068_7039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7363 a_1808_n5908# a_1481_n8108# a_1803_n7931# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7364 vdd a_4936_n10733# a_4728_n10733# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7365 a_30335_n6391# a_30864_n6711# a_31072_n6711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7366 a_5489_7169# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7367 a_1810_3115# a_1513_4086# a_1794_3575# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7368 vdd a_13171_n5396# a_12963_n5396# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7369 a_119_4116# a_646_4368# a_854_4368# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7370 a_32022_n3505# a_31913_n3682# a_32020_n5717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7371 a_39100_2806# a_39096_2983# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7372 a_24008_5143# a_24011_4412# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7373 a_13852_n8999# a_14109_n9015# a_12917_n8501# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7374 a_17974_n5233# a_18958_n5747# a_18909_n5731# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7375 vdd a_34297_1095# a_34089_1095# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7376 a_20305_2994# a_20833_3246# a_21041_3246# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7377 a_38157_3776# a_39144_3342# a_39099_3355# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7378 a_13857_4990# a_13853_5167# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7379 a_6641_4719# a_6428_4719# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7380 a_21880_7389# a_21667_7389# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7381 a_9855_n1566# a_10679_n1764# a_10887_n1764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7382 a_32995_5234# a_33248_5221# a_32221_486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7383 a_18914_3928# a_19167_3915# a_17975_3618# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7384 a_15522_n1805# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7385 a_2747_4164# a_2932_4662# a_2887_4675# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7386 gnd a_38304_n3791# a_38096_n3791# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7387 a_20835_1594# a_20622_1594# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7388 a_7629_n10697# a_7879_n6005# a_7830_n5989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7389 a_10466_2721# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7390 a_39094_n9021# a_39097_n8279# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7391 a_3821_4608# a_3827_3882# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7392 a_432_7677# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7393 a_10148_7243# a_10677_7133# a_10885_7133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7394 a_20621_1040# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7395 a_10462_n9485# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7396 a_118_n6821# a_118_n6634# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7397 a_7940_n3210# a_8927_n2982# a_8878_n2966# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7398 a_1810_n3696# a_1696_n3696# a_1803_n5731# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7399 a_28129_5800# a_28382_5787# a_27984_6569# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7400 vdd a_19163_8876# a_18955_8876# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7401 a_13852_5716# a_14109_5526# a_12914_5960# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7402 a_20304_n5512# a_20304_n5283# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7403 vdd d2 a_13032_n2679# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7404 a_37081_7554# a_36784_8525# a_37065_8014# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7405 a_17974_5824# a_18958_6121# a_18909_6311# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7406 gnd d2 a_23184_8544# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7407 a_116_n9943# a_645_n10034# a_853_n10034# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7408 a_21560_n2050# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7409 gnd d0 a_14110_3320# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7410 gnd a_28243_n2696# a_28035_n2696# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7411 a_16892_3042# a_16601_1926# a_16881_2518# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7412 a_33103_6867# a_33356_6854# a_32963_6356# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7413 a_27815_n10678# a_28065_n5986# a_28016_n5970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7414 a_27045_n5753# a_26725_n3718# a_27047_n3541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7415 a_6851_n2110# a_6783_n2621# a_6861_n3560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7416 a_22964_n5741# a_23007_n8157# a_22958_n8141# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7417 a_30649_n10020# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7418 vdd a_4078_n7907# a_3870_n7907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7419 a_22190_481# a_23009_5216# a_22964_5229# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7420 a_27050_5349# a_26936_5230# a_27144_5230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7421 a_22964_n3541# a_22978_n4861# a_22929_n4845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7422 a_28126_n3191# a_29113_n2963# a_29064_n2947# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7423 a_15733_n8977# a_15520_n8977# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7424 a_21910_8479# a_21697_8479# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7425 a_24010_6618# a_24263_6605# a_23068_7039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7426 a_25675_8253# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7427 a_118_6322# a_118_6135# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7428 gnd d0 a_4079_6075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7429 a_33103_n7379# a_33356_n7583# a_32963_n6868# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7430 a_31729_6278# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7431 a_25360_n6197# a_25360_n5740# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7432 a_31072_n3951# a_31803_n4261# a_32011_n4261# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7433 gnd a_39352_n4071# a_39144_n4071# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7434 a_6642_3616# a_6429_3616# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7435 a_25362_n2015# a_25362_n1785# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7436 a_21979_4659# a_21558_4659# a_21040_4349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7437 a_10885_n7833# a_10464_n7833# a_10148_n7513# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7438 a_1792_6884# a_1371_6884# a_853_6574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7439 a_16781_n5954# a_16568_n5954# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7440 a_36646_n4302# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7441 gnd d4 a_23217_n5945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7442 gnd a_14110_6080# a_13902_6080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7443 a_5174_5717# a_5174_5260# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7444 a_10148_n7929# a_10676_n8382# a_10884_n8382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7445 gnd d1 a_33356_n8686# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7446 a_5174_n5572# a_5703_n5663# a_5911_n5663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7447 a_10678_n5627# a_10465_n5627# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7448 a_32011_n3158# a_31944_n2566# a_32022_n3505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7449 a_16882_n2115# a_16461_n2115# a_15944_n2359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7450 vdd d1 a_28380_n9825# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7451 a_21882_n3677# a_21669_n3677# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7452 vdd d0 a_9136_n3536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7453 a_25140_461# a_25031_461# a_25239_461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7454 a_3824_1853# a_4081_1663# a_2889_1366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7455 a_36857_n7611# a_36644_n7611# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7456 gnd a_38413_4689# a_38205_4689# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7457 a_34041_1839# a_34044_1108# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7458 a_8877_n7932# a_8880_n7190# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7459 a_6537_n5949# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7460 a_23073_5759# a_24057_6056# a_24008_6246# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7461 a_434_3265# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7462 a_36860_n2096# a_36647_n2096# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7463 a_31070_9320# a_30649_9320# a_30333_9430# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7464 gnd d1 a_13172_2461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7465 a_12772_8758# a_12962_7976# a_12913_8166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7466 a_21042_1040# a_21773_1350# a_21981_1350# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7467 a_34037_n8426# a_34042_n7689# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7468 a_7937_n9828# a_8924_n9600# a_8875_n9584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7469 a_13853_n4033# a_13858_n3296# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7470 a_28131_1388# a_28384_1375# a_27986_2157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7471 a_21556_9071# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7472 vdd a_19165_4464# a_18957_4464# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7473 a_25890_n1781# a_25677_n1781# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7474 gnd d1 a_28381_n7619# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7475 a_5913_1654# a_5492_1654# a_5176_1535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7476 a_25887_n8399# a_25674_n8399# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7477 a_5175_2867# a_5175_2638# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7478 a_18910_n1868# a_19886_n1571# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7479 a_17828_8799# a_18085_8609# a_17863_7506# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7480 vdd d2 a_13029_n9297# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7481 gnd a_20790_n10911# a_20582_n10911# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7482 a_16878_9136# a_16457_9136# a_15939_8826# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7483 a_25891_n2335# a_25678_n2335# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7484 a_37083_3142# a_36786_4113# a_37067_3602# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7485 a_20830_8761# a_20617_8761# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7486 a_29061_n9565# a_29067_n8828# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7487 a_23074_n2962# a_24058_n3476# a_24009_n3460# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7488 a_15203_9261# a_15732_9380# a_15940_9380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7489 gnd d2 a_23186_4132# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7490 a_5911_4963# a_5490_4963# a_5174_5073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7491 a_36128_n5649# a_36858_n5405# a_37066_n5405# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7492 a_6951_541# a_6738_541# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7493 a_35707_4949# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7494 gnd d0 a_19165_n9056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7495 a_11725_5213# a_11512_5213# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7496 a_2888_3572# a_3872_3869# a_3827_3882# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7497 a_15942_n6771# a_15521_n6771# a_15205_n6680# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7498 a_32991_5411# a_33248_5221# a_32221_486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7499 a_12919_n4089# a_13903_n4603# a_13858_n4399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7500 a_28129_n6312# a_29113_n6826# a_29068_n6622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7501 a_120_1264# a_122_1165# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7502 vdd d5 a_33047_n10658# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7503 a_16459_n6527# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7504 a_28123_n9809# a_29110_n9581# a_29061_n9565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7505 a_16880_4724# a_16459_4724# a_15942_4968# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7506 a_21912_4067# a_21699_4067# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7507 a_32958_n9262# a_33148_n8686# a_33103_n8482# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7508 a_6427_n7625# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7509 a_24012_2206# a_24265_2193# a_23070_2627# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7510 gnd a_3000_n4880# a_2792_n4880# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7511 gnd a_24264_n6231# a_24056_n6231# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7512 a_3823_n4582# a_3826_n3840# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7513 a_20306_1245# a_20834_1040# a_21042_1040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7514 a_8880_n2417# a_9137_n2433# a_7945_n1919# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7515 vdd a_19164_n7399# a_18956_n7399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7516 a_22190_481# a_22081_481# a_22289_481# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7517 a_1794_2472# a_1373_2472# a_855_2162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7518 a_38020_4191# a_38205_4689# a_38160_4702# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7519 a_32993_n7958# a_33246_n8162# a_32995_n5746# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7520 a_2746_n6882# a_2999_n7086# a_2772_n8160# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7521 vdd d1 a_13170_6873# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7522 a_853_n7274# a_432_n7274# a_117_n7278# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7523 gnd d0 a_19166_2258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7524 a_25675_n8953# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7525 a_24008_n2906# a_24265_n2922# a_23070_n3150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7526 a_17830_4387# a_18020_3605# a_17975_3618# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7527 a_1808_n5908# a_1694_n5908# a_1902_n5908# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7528 vdd a_3139_n8700# a_2931_n8700# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7529 a_119_n4199# a_119_n3969# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7530 gnd d1 a_8194_9115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7531 gnd a_14108_n10118# a_13900_n10118# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7532 a_35389_n9970# a_35918_n10061# a_36126_n10061# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7533 a_20835_n2294# a_20622_n2294# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7534 a_34043_6074# a_34296_6061# a_33104_5764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7535 a_29069_n4416# a_29065_n4604# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7536 vdd d0 a_24265_n4025# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7537 a_6859_5249# a_6539_3037# a_6861_3037# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7538 a_30651_n6711# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7539 a_21772_n4256# a_21559_n4256# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7540 gnd d0 a_39349_8857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7541 gnd d2 a_28242_n4902# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7542 a_12919_n2986# a_13172_n3190# a_12779_n2475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7543 a_17974_5824# a_18958_6121# a_18913_6134# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7544 a_31072_4908# a_30651_4908# a_30335_5018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7545 vdd d2 a_23184_8544# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7546 a_30335_5662# a_30863_5457# a_31071_5457# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7547 vdd d0 a_14110_3320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7548 vdd a_38411_n9830# a_38203_n9830# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7549 a_28124_n7603# a_28381_n7619# a_27988_n6904# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7550 a_36127_n7855# a_35706_n7855# a_35390_n7764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7551 a_11823_n8692# a_11402_n8692# a_10885_n8936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7552 a_6864_7568# a_6567_8539# a_6847_9131# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7553 a_2885_1543# a_3872_1109# a_3823_1299# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7554 a_16879_8033# a_16458_8033# a_15941_8277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7555 a_7939_4893# a_8196_4703# a_7803_4205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7556 gnd d1 a_13172_n4293# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7557 a_11725_7413# a_11512_7413# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7558 a_17830_4387# a_18087_4197# a_17865_3094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7559 vdd d1 a_33358_n3171# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7560 gnd d0 a_24266_n1819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7561 a_20304_5013# a_20833_4903# a_21041_4903# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7562 a_645_n8377# a_432_n8377# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7563 gnd d0 a_39351_n6277# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7564 vdd d0 a_4079_6075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7565 a_10466_n1764# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7566 a_24007_4589# a_24013_3863# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7567 vdd d0 a_19166_n2987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7568 a_25890_2738# a_25677_2738# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7569 a_35708_3846# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7570 a_5174_6363# a_5701_6615# a_5909_6615# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7571 gnd a_28271_n8198# a_28063_n8198# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7572 a_7834_n3601# a_8087_n3805# a_7830_n5989# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7573 a_30865_3805# a_30652_3805# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7574 a_10149_n6639# a_10149_n6410# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7575 a_33102_1529# a_34089_1095# a_34044_1108# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7576 a_1792_7987# a_1371_7987# a_854_8231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7577 a_35390_8368# a_35919_8258# a_36127_8258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7578 vdd a_34294_n8442# a_34086_n8442# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7579 vdd a_14110_6080# a_13902_6080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7580 a_2743_n4864# a_3000_n4880# a_2778_n3560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7581 gnd a_38415_n2109# a_38207_n2109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7582 a_3823_4059# a_3826_3328# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7583 a_17974_4721# a_18227_4708# a_17834_4210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7584 a_37065_6911# a_36644_6911# a_36126_6601# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7585 a_15206_n4474# a_15206_n4245# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7586 a_30863_7114# a_30650_7114# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7587 vdd a_19166_n6850# a_18958_n6850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7588 a_21040_n5049# a_20619_n5049# a_20304_n5053# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7589 gnd a_29320_n9032# a_29112_n9032# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7590 a_1483_n3696# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7591 a_855_n6725# a_434_n6725# a_118_n6634# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7592 a_23073_5759# a_24057_6056# a_24012_6069# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7593 a_12778_4169# a_13031_4156# a_12809_3053# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7594 a_39093_n8467# a_39098_n7730# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7595 a_8876_n10138# a_9133_n10154# a_7941_n9640# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7596 a_29066_9419# a_30333_9430# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7597 a_7802_6411# a_7987_6909# a_7942_6922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7598 a_39095_n6815# a_39352_n6831# a_38160_n6317# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7599 vdd d1 a_13172_2461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7600 gnd d6 a_14967_n10738# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7601 a_10151_n2414# a_10151_n2227# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7602 a_6570_1921# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7603 a_20305_2807# a_20834_2697# a_21042_2697# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7604 a_21770_6865# a_21557_6865# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7605 a_32991_n5934# a_33248_n5950# a_32790_n10642# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7606 a_38157_n4299# a_39144_n4071# a_39099_n3867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7607 a_12805_n3753# a_12824_n2679# a_12779_n2475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7608 a_4845_480# a_4632_480# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7609 vdd a_29320_8303# a_29112_8303# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7610 a_28127_1565# a_28384_1375# a_27986_2157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7611 a_31589_4664# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7612 gnd a_33047_n10658# a_32839_n10658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7613 a_10463_7682# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7614 vdd a_34296_n5687# a_34088_n5687# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7615 a_5908_8821# a_5487_8821# a_5172_9026# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7616 a_27983_8775# a_28173_7993# a_28124_8183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7617 a_1803_5208# a_1483_2996# a_1805_2996# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7618 a_31070_9320# a_31800_9076# a_32008_9076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7619 a_5702_8272# a_5489_8272# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7620 a_25889_6047# a_25676_6047# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7621 a_11404_3580# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7622 a_30335_n6161# a_30863_n6157# a_31071_n6157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7623 a_120_n2222# a_649_n2313# a_857_n2313# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7624 a_38156_5982# a_39143_5548# a_39094_5738# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7625 vdd d2 a_2999_6357# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7626 vdd d2 a_23186_4132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7627 a_16671_n7630# a_16458_n7630# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7628 a_31590_n3158# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7629 vdd a_9135_n4085# a_8927_n4085# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7630 a_28127_n9621# a_28380_n9825# a_27987_n9110# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7631 a_25360_5698# a_25360_5241# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7632 a_38051_5275# a_38304_5262# a_37277_527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7633 a_26096_n6193# a_26827_n6503# a_27035_n6503# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7634 vdd a_3139_6868# a_2931_6868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7635 a_28014_n8182# a_28271_n8198# a_28020_n5782# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7636 a_6639_n9831# a_6426_n9831# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7637 a_12803_7642# a_12822_6362# a_12773_6552# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7638 a_11727_3001# a_11514_3001# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7639 gnd d0 a_24263_n8437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7640 a_25891_1635# a_25678_1635# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7641 a_10463_n8382# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7642 a_34039_n5671# a_34042_n4929# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7643 a_31071_n5054# a_30650_n5054# a_30335_n5058# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7644 a_648_1059# a_435_1059# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7645 a_5176_1951# a_5703_2203# a_5911_2203# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7646 vdd a_13173_n2087# a_12965_n2087# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7647 gnd a_23327_n4269# a_23119_n4269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7648 a_7944_n3022# a_8928_n3536# a_8883_n3332# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7649 gnd d0 a_9134_8322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7650 a_11713_505# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7651 a_20305_2807# a_20305_2578# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7652 a_1583_9090# a_1370_9090# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7653 vdd d3 a_3031_n3764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7654 a_30335_n5058# a_30336_n4601# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7655 a_14985_485# a_14876_485# a_9888_364# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7656 a_33105_n4070# a_34089_n4584# a_34044_n4380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7657 a_6851_n2110# a_6430_n2110# a_5912_n1800# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7658 a_1895_500# a_1682_500# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7659 a_20622_1594# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7660 vdd d1 a_8194_9115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7661 a_26098_3841# a_26828_3597# a_27036_3597# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7662 gnd a_8087_5276# a_7879_5276# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7663 a_15942_n6771# a_16672_n6527# a_16880_n6527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7664 a_34039_6251# a_34296_6061# a_33104_5764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7665 vdd a_28240_n9314# a_28032_n9314# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7666 a_431_n9480# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7667 a_24007_n8975# a_24264_n8991# a_23072_n8477# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7668 a_8876_n7378# a_8882_n6641# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7669 a_38159_6908# a_38412_6895# a_38019_6397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7670 a_7804_1999# a_7989_2497# a_7944_2510# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7671 a_21772_2453# a_21559_2453# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7672 a_15939_n9526# a_15518_n9526# a_15203_n9530# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7673 a_5910_4409# a_6641_4719# a_6849_4719# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7674 a_12807_n7977# a_12821_n9297# a_12776_n9093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7675 a_31070_7663# a_31801_7973# a_32009_7973# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7676 a_35920_n2889# a_35707_n2889# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7677 a_20302_n9924# a_20302_n9695# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7678 a_28018_7482# a_28271_7469# a_28020_5270# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7679 a_17973_n8542# a_18957_n9056# a_18908_n9040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7680 a_35921_n3443# a_35708_n3443# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7681 a_38158_1570# a_39145_1136# a_39096_1326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7682 a_6427_8028# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7683 a_15204_n7554# a_15204_n7324# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7684 a_26097_n6747# a_25676_n6747# a_25360_n6427# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7685 a_38016_n4891# a_38273_n4907# a_38051_n3587# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7686 a_30335_n6620# a_30864_n6711# a_31072_n6711# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7687 a_31070_7663# a_30649_7663# a_30334_7868# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7688 gnd a_14110_n2946# a_13902_n2946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7689 a_3826_n2737# a_3822_n2925# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7690 a_16673_3621# a_16460_3621# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7691 a_21040_8212# a_20619_8212# a_20303_8093# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7692 a_2748_1958# a_2933_2456# a_2884_2646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7693 a_31071_4354# a_30650_4354# a_30336_4102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7694 a_5175_n3366# a_5175_n3137# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7695 a_12805_3230# a_12824_1950# a_12775_2140# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7696 a_15519_6620# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7697 vdd d0 a_19165_n9056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7698 a_15205_5952# a_15734_6071# a_15942_6071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7699 a_119_3700# a_119_3470# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7700 a_31073_n4505# a_30652_n4505# a_30336_n4414# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7701 a_28129_5800# a_29113_6097# a_29064_6287# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7702 gnd a_35153_n10719# a_34945_n10719# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7703 gnd d5 a_2830_n10672# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7704 a_10885_n7833# a_11615_n7589# a_11823_n7589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7705 a_12774_4346# a_13031_4156# a_12809_3053# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7706 a_1481_n5908# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7707 a_10151_n1768# a_10679_n1764# a_10887_n1764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7708 a_2887_n6290# a_3140_n6494# a_2742_n7070# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7709 a_25361_3722# a_25361_3492# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7710 gnd d0 a_9136_3910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7711 vdd d0 a_39351_n5174# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7712 a_15522_n1805# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7713 gnd a_18226_n7643# a_18018_n7643# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7714 a_35705_n10061# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7715 a_2742_n7070# a_2999_n7086# a_2772_n8160# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7716 a_35393_n2249# a_35922_n2340# a_36130_n2340# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7717 a_38017_n2685# a_38207_n2109# a_38162_n1905# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7718 a_15523_n2359# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7719 a_35918_n10061# a_35705_n10061# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7720 a_31802_n5364# a_31589_n5364# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7721 a_5175_n4010# a_5175_n3553# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7722 gnd a_13172_2461# a_12964_2461# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7723 a_31729_n6978# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7724 a_12774_n4869# a_12964_n4293# a_12915_n4277# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7725 a_30862_6560# a_30649_6560# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7726 a_9875_n10838# a_9825_n10854# a_4778_n10717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7727 a_16781_5254# a_16568_5254# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7728 a_21040_n7809# a_20619_n7809# a_20303_n7489# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7729 a_38047_5452# a_38304_5262# a_37277_527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7730 a_21979_5762# a_21911_6273# a_21989_7389# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7731 a_35919_n8958# a_35706_n8958# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7732 a_15735_2762# a_15522_2762# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7733 gnd d0 a_4078_n5147# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7734 a_17971_n3215# a_18958_n2987# a_18913_n2783# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7735 a_10147_n9489# a_10148_n9032# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7736 vdd a_8198_n2123# a_7990_n2123# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7737 a_28020_3070# a_28273_3057# a_28016_5447# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7738 a_27034_8009# a_26613_8009# a_26095_7699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7739 a_25361_n4221# a_25890_n4541# a_26098_n4541# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7740 a_11841_n3701# a_11544_n4791# a_11825_n4280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7741 a_9987_364# a_9566_364# a_5053_480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7742 a_7801_n9129# a_8054_n9333# a_7832_n8013# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7743 a_12803_7642# a_12822_6362# a_12777_6375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7744 a_20834_3800# a_20621_3800# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7745 a_36967_n5935# a_36754_n5935# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7746 a_39095_n5712# a_39098_n4970# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7747 a_29063_7390# a_29320_7200# a_28128_6903# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7748 a_20833_n5603# a_20620_n5603# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7749 a_32961_2121# a_33151_1339# a_33106_1352# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7750 a_854_n5068# a_1585_n5378# a_1793_n5378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7751 a_9566_364# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7752 a_18911_7786# a_18907_7963# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7753 a_22928_n7051# a_23185_n7067# a_22958_n8141# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7754 a_10147_9449# a_10676_9339# a_10884_9339# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7755 a_6850_n3213# a_6783_n2621# a_6861_n3560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7756 vdd a_14110_n6809# a_13902_n6809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7757 a_11512_5213# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7758 a_27037_1391# a_26616_1391# a_26098_1081# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7759 a_31072_3251# a_30651_3251# a_30336_3456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7760 vdd d0 a_9134_8322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7761 gnd a_14107_n9564# a_13899_n9564# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7762 a_21039_7658# a_20618_7658# a_20303_7863# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7763 gnd d0 a_34294_6610# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7764 a_17859_n8206# a_17878_n7132# a_17829_n7116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7765 a_31073_n4505# a_31803_n4261# a_32011_n4261# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7766 a_39099_6115# a_39352_6102# a_38160_5805# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7767 a_3821_n8994# a_3824_n8252# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7768 a_11404_n4280# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7769 vdd a_8087_5276# a_7879_5276# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7770 a_3822_n5685# a_4079_n5701# a_2887_n5187# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7771 a_36646_n4302# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7772 a_17973_8030# a_18957_8327# a_18908_8517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7773 a_32025_n5894# a_31698_n8094# a_32025_n8094# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7774 gnd d0 a_14109_5526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7775 a_1585_n6481# a_1372_n6481# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7776 gnd a_19166_2258# a_18958_2258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7777 a_17969_n8730# a_18226_n8746# a_17828_n9322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7778 a_30333_9201# a_30333_8971# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7779 a_10678_n5627# a_10465_n5627# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7780 a_21882_n3677# a_21669_n3677# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7781 gnd a_8194_9115# a_7986_9115# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7782 a_117_n8611# a_117_n8381# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7783 a_36857_n7611# a_36644_n7611# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7784 gnd a_18116_n8222# a_17908_n8222# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7785 gnd d0 a_39350_9411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7786 a_16781_7454# a_16568_7454# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7787 a_38014_n9303# a_38204_n8727# a_38159_n8523# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7788 a_23071_n9580# a_23324_n9784# a_22931_n9069# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7789 a_25360_5054# a_25889_4944# a_26097_4944# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7790 a_21040_n6152# a_21771_n6462# a_21979_n6462# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7791 a_36127_n6198# a_35706_n6198# a_35391_n5745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7792 a_29067_n8828# a_29063_n9016# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7793 gnd a_30219_n10835# a_30011_n10835# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7794 a_26614_n6503# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7795 a_22964_n3541# a_23217_n3745# a_22960_n5929# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7796 a_38049_n7999# a_38302_n8203# a_38051_n5787# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7797 a_38158_1570# a_39145_1136# a_39100_1149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7798 a_30336_3686# a_30336_3456# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7799 a_27045_n5753# a_26936_n5930# a_27144_n5930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7800 a_11826_n2074# a_11405_n2074# a_10887_n1764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7801 a_2889_1366# a_3873_1663# a_3824_1853# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7802 gnd a_14109_8286# a_13901_8286# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7803 a_2887_n6290# a_3871_n6804# a_3822_n6788# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7804 a_24013_n1615# a_24009_n1803# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7805 gnd d0 a_29318_8852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7806 a_25358_9466# a_25358_9237# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7807 a_25362_n2244# a_25362_n2015# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7808 a_15521_n5668# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7809 a_2748_1958# a_2933_2456# a_2888_2469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7810 a_11512_7413# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7811 a_25891_n2335# a_25678_n2335# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7812 a_10148_8117# a_10677_8236# a_10885_8236# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7813 a_2745_n9088# a_2930_n9803# a_2885_n9599# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7814 a_854_8231# a_433_8231# a_117_8112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7815 a_18912_n7749# a_18908_n7937# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7816 a_30652_3805# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7817 a_118_n5302# a_647_n5622# a_855_n5622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7818 a_11614_9095# a_11401_9095# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7819 gnd d1 a_13171_4667# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7820 a_2774_n5948# a_2823_n3764# a_2778_n3560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7821 a_6847_n9831# a_6780_n9239# a_6864_n8149# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7822 a_15942_n6771# a_15521_n6771# a_15205_n6451# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7823 a_30863_n6157# a_30650_n6157# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7824 a_11755_n9203# a_11542_n9203# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7825 a_5175_n3553# a_5703_n4006# a_5911_n4006# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7826 gnd d1 a_18225_n9849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7827 a_15734_n4011# a_15521_n4011# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7828 gnd a_33357_n5377# a_33149_n5377# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7829 a_645_9334# a_432_9334# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7830 a_15941_4414# a_15520_4414# a_15205_4619# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7831 a_36643_9117# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7832 a_11824_n6486# a_11756_n6997# a_11834_n7936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7833 a_16459_n6527# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7834 a_37065_n7611# a_36998_n7019# a_37076_n7958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7835 a_15206_3059# a_15206_2872# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7836 a_8881_8335# a_8877_8512# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7837 a_30650_7114# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7838 a_15735_n4565# a_15522_n4565# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7839 vdd d1 a_38414_n3212# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7840 gnd d0 a_29322_n1860# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7841 a_37076_7435# a_36785_6319# a_37066_5808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7842 a_17975_3618# a_18959_3915# a_18910_4105# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7843 a_37083_n3723# a_36786_n4813# a_37066_n5405# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7844 a_30864_n2848# a_30651_n2848# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7845 gnd d2 a_23185_6338# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7846 a_10887_n3421# a_10466_n3421# a_10150_n3330# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7847 gnd d0 a_14111_1114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7848 a_5910_7169# a_5489_7169# a_5173_7279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7849 a_30334_6995# a_30334_6765# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7850 a_853_n7274# a_432_n7274# a_118_n6821# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7851 vdd a_13172_2461# a_12964_2461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7852 a_30648_8766# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7853 a_34037_n10083# a_34294_n10099# a_33102_n9585# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7854 a_10149_n6826# a_10149_n6639# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7855 a_24012_n3821# a_24265_n4025# a_23070_n4253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7856 vdd d1 a_38413_5792# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7857 a_7803_n4717# a_7988_n5432# a_7943_n5228# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7858 a_18908_n5177# a_19165_n5193# a_17970_n5421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7859 a_25361_3722# a_25890_3841# a_26098_3841# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7860 a_10885_7133# a_10464_7133# a_10148_7014# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7861 a_16783_3042# a_16570_3042# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7862 a_24011_4412# a_24264_4399# a_23069_4833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7863 gnd d0 a_4080_3869# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7864 a_25676_6047# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7865 vdd d0 a_14109_n7912# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7866 a_30651_n6711# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7867 a_21772_n4256# a_21559_n4256# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7868 a_15939_n9526# a_16670_n9836# a_16878_n9836# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7869 a_22930_2116# a_23187_1926# a_22960_3206# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7870 a_6643_1410# a_6430_1410# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7871 a_1793_4678# a_1372_4678# a_854_4368# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7872 a_38019_6397# a_38204_6895# a_38159_6908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7873 a_32119_5194# a_31698_5194# a_32025_5313# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7874 a_5704_n1800# a_5491_n1800# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7875 gnd a_14111_3874# a_13903_3874# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7876 a_36127_n7855# a_35706_n7855# a_35390_n7535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7877 a_38047_n5975# a_38304_n5991# a_37846_n10683# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7878 a_28014_7659# a_28033_6379# a_27988_6392# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7879 a_17973_n8542# a_18957_n9056# a_18912_n8852# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7880 a_21991_2977# a_21700_1861# a_21981_1350# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7881 a_11543_n6997# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7882 a_27045_n5753# a_26725_n3718# a_27052_n3718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7883 a_36997_8525# a_36784_8525# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7884 a_24009_2937# a_24266_2747# a_23074_2450# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7885 a_11514_3001# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7886 a_27989_n4698# a_28174_n5413# a_28129_n5209# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7887 a_11616_n6486# a_11403_n6486# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7888 a_649_1613# a_436_1613# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7889 vdd d0 a_34294_6610# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7890 a_34038_5697# a_34043_4971# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7891 a_10466_n1764# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7892 a_34042_8280# a_34295_8267# a_33103_7970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7893 a_16673_n3218# a_16460_n3218# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7894 a_34037_n10083# a_34040_n9341# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7895 a_435_1059# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7896 vdd d0 a_19167_2812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7897 gnd d0 a_24267_n2373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7898 a_2778_n3560# a_2792_n4880# a_2743_n4864# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7899 a_36644_8014# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7900 a_36126_6601# a_35705_6601# a_35391_6349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7901 vdd d0 a_14109_5526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7902 a_32991_5411# a_33040_3021# a_32991_3211# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7903 a_39098_8321# a_39094_8498# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7904 a_8878_3546# a_8883_2820# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7905 gnd a_9134_8322# a_8926_8322# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7906 a_3821_n6234# a_3826_n5497# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7907 a_35709_n2340# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7908 a_1370_9090# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7909 a_647_4922# a_434_4922# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7910 gnd d1 a_8196_4703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7911 a_35390_n7951# a_35918_n8404# a_36126_n8404# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7912 a_18910_8889# a_19163_8876# a_17968_9310# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7913 vdd d1 a_23326_n5372# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7914 a_35391_6162# a_35391_5933# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7915 gnd d4 a_3031_n5964# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7916 vdd a_8194_9115# a_7986_9115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7917 gnd d0 a_29319_n8478# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7918 a_6429_n3213# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7919 a_32008_9076# a_31941_8484# a_32025_7513# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7920 a_17829_6593# a_18086_6403# a_17859_7683# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7921 a_20305_n3077# a_20834_n3397# a_21042_n3397# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7922 vdd d0 a_39350_9411# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7923 a_855_n6725# a_434_n6725# a_118_n6405# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7924 vdd d2 a_38274_1972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7925 a_20831_6555# a_20618_6555# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7926 a_14710_n10722# a_17709_n10718# a_16989_n5954# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7927 gnd d2 a_3000_4151# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7928 gnd d0 a_4079_n2941# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7929 gnd d2 a_23187_1926# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7930 vdd a_28381_7993# a_28173_7993# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7931 a_18910_n4628# a_19167_n4644# a_17975_n4130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7932 a_29069_n1656# a_29065_n1844# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7933 gnd a_3140_4662# a_2932_4662# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7934 a_25677_n4541# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7935 a_2889_1366# a_3873_1663# a_3828_1676# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7936 vdd a_14109_8286# a_13901_8286# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7937 a_38161_n4111# a_39145_n4625# a_39100_n4421# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7938 a_30862_9320# a_30649_9320# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7939 a_16881_2518# a_16460_2518# a_15943_2762# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7940 a_1794_3575# a_1373_3575# a_856_3819# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7941 a_23068_n7562# a_24055_n7334# a_24010_n7130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7942 a_13858_n4399# a_14111_n4603# a_12919_n4089# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7943 a_39094_n7918# a_39097_n7176# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7944 a_29063_n9016# a_29320_n9032# a_28128_n8518# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7945 a_15732_7723# a_15519_7723# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7946 a_26097_n6747# a_26827_n6503# a_27035_n6503# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7947 a_22289_481# a_21868_481# a_22190_481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7948 a_118_n5718# a_118_n5531# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7949 a_17863_7506# a_17877_8609# a_17832_8622# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7950 a_38162_n1905# a_39146_n2419# a_39097_n2403# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7951 a_16460_3621# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7952 a_5176_1305# a_5178_1206# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7953 a_31588_6870# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7954 a_31730_n4772# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7955 a_36999_4113# a_36786_4113# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7956 vdd d0 a_34297_n4584# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7957 a_23069_n5356# a_24056_n5128# a_24007_n5112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7958 vdd a_29320_n6272# a_29112_n6272# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7959 vdd d0 a_34296_2198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7960 a_20621_n3397# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7961 a_34044_3868# a_34297_3855# a_33105_3558# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7962 vdd a_39350_n10140# a_39142_n10140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7963 vdd d0 a_14111_1114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7964 a_34849_466# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7965 gnd a_9136_3910# a_8928_3910# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7966 gnd a_9137_n2433# a_8929_n2433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7967 a_10148_7887# a_10676_7682# a_10884_7682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7968 a_21558_n6462# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7969 a_35392_3956# a_35392_3727# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7970 a_13856_8299# a_13852_8476# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7971 vdd a_13029_8568# a_12821_8568# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7972 a_23075_n1859# a_23328_n2063# a_22930_n2639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7973 a_1803_n5731# a_1694_n5908# a_1902_n5908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7974 a_10150_n4204# a_10150_n3974# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7975 a_12807_7465# a_12821_8568# a_12772_8758# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7976 a_17831_2181# a_18088_1991# a_17861_3271# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7977 a_32010_4664# a_31943_4072# a_32027_3101# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7978 vdd d0 a_39352_4999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7979 gnd a_24265_n2922# a_24057_n2922# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7980 a_17971_n3215# a_18228_n3231# a_17835_n2516# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7981 a_32960_4327# a_33150_3545# a_33101_3735# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7982 a_644_8780# a_431_8780# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7983 a_20833_2143# a_20620_2143# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7984 a_21667_7389# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7985 a_118_5219# a_118_5032# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7986 a_35709_1640# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7987 a_36644_n7611# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7988 gnd a_13171_n6499# a_12963_n6499# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7989 a_6850_2513# a_6783_1921# a_6861_3037# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7990 a_5175_4157# a_5702_4409# a_5910_4409# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7991 a_25360_n5094# a_25361_n4637# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7992 a_26096_7150# a_25675_7150# a_25359_7031# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7993 a_15939_n9526# a_15518_n9526# a_15204_n9073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7994 a_3820_7917# a_3825_7191# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7995 vdd d1 a_18228_n4334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X7996 a_21980_n3153# a_21559_n3153# a_21041_n2843# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7997 a_15522_2762# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7998 a_5174_4614# a_5175_4157# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X7999 a_37066_4705# a_36645_4705# a_36127_4395# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8000 a_435_n4519# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8001 gnd d0 a_4076_8830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8002 a_23073_n6271# a_24057_n6785# a_24012_n6581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8003 a_16880_n5424# a_16459_n5424# a_15942_n5668# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8004 a_30864_4908# a_30651_4908# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8005 a_10678_n3970# a_10465_n3970# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8006 a_20621_3800# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8007 a_6567_n9239# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8008 a_19317_288# a_29752_345# a_25239_461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8009 a_35921_n3443# a_35708_n3443# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8010 a_36785_n7019# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8011 a_15734_3311# a_15521_3311# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8012 a_7803_4205# a_7988_4703# a_7943_4716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8013 a_5173_8382# a_5173_8153# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8014 a_21771_4659# a_21558_4659# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8015 a_32991_5411# a_33040_3021# a_32995_3034# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8016 a_17865_3094# a_17879_4197# a_17834_4210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8017 vdd a_9134_8322# a_8926_8322# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8018 a_34037_n7323# a_34043_n6586# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8019 a_13853_n2930# a_13859_n2193# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8020 a_38159_n8523# a_39143_n9037# a_39094_n9021# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8021 a_38047_n3775# a_38066_n2701# a_38021_n2497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8022 gnd d0 a_9134_n5188# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8023 a_31899_486# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8024 a_15205_5952# a_15205_5722# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8025 a_5909_6615# a_5488_6615# a_5173_6820# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8026 a_10149_6327# a_10149_6140# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8027 gnd a_34294_6610# a_34086_6610# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8028 a_31073_n4505# a_30652_n4505# a_30336_n4185# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8029 a_12779_n2475# a_13032_n2679# a_12805_n3753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8030 gnd d0 a_39352_n2968# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8031 a_5703_6066# a_5490_6066# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8032 a_24012_n5478# a_24008_n5666# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8033 a_21989_7389# a_21880_7389# a_21994_5308# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8034 a_27984_n7092# a_28241_n7108# a_28014_n8182# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8035 a_36857_6911# a_36644_6911# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8036 vdd d2 a_3000_4151# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8037 a_10147_n9719# a_10676_n10039# a_10884_n10039# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8038 a_34041_n2362# a_34298_n2378# a_33106_n1864# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8039 a_119_2597# a_648_2716# a_856_2716# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8040 a_13852_4613# a_13858_3887# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8041 a_34042_n4929# a_34295_n5133# a_33100_n5361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8042 gnd a_9134_n9051# a_8926_n9051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8043 a_10150_3475# a_10678_3270# a_10886_3270# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8044 vdd a_3140_4662# a_2932_4662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8045 a_12917_n7398# a_13901_n7912# a_13856_n7708# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8046 vdd d2 a_33218_n2660# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8047 vdd a_8057_n2715# a_7849_n2715# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8048 a_16672_5827# a_16459_5827# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8049 a_16457_n9836# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8050 a_12914_n6483# a_13171_n6499# a_12773_n7075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8051 a_11824_n5383# a_11403_n5383# a_10885_n5073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8052 a_16890_n7977# a_16781_n8154# a_16895_n5954# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8053 gnd a_39352_n6831# a_39144_n6831# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8054 a_11933_5213# a_11926_505# a_12134_505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8055 a_12809_3053# a_12823_4156# a_12774_4346# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8056 a_119_3013# a_119_2826# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8057 a_38162_1393# a_39146_1690# a_39101_1703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8058 gnd a_24262_n9540# a_24054_n9540# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8059 gnd a_29321_n5723# a_29113_n5723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8060 a_31802_n5364# a_31589_n5364# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8061 a_3823_n3479# a_3826_n2737# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8062 gnd a_4078_n9010# a_3870_n9010# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8063 a_16670_9136# a_16457_9136# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8064 vdd d0 a_29319_n7375# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8065 a_8878_n4069# a_8883_n3332# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8066 a_10884_7682# a_11615_7992# a_11823_7992# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8067 a_37067_3602# a_36646_3602# a_36129_3846# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8068 a_32008_9076# a_31587_9076# a_31069_8766# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8069 a_37068_n2096# a_36647_n2096# a_36130_n2340# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8070 gnd d0 a_9135_6116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8071 a_29068_6110# a_29064_6287# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8072 gnd a_29318_8852# a_29110_8852# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8073 a_6848_6925# a_6427_6925# a_5909_6615# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8074 a_25360_n6656# a_25360_n6427# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8075 a_25361_n4450# a_25890_n4541# a_26098_n4541# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8076 gnd a_19167_n1884# a_18959_n1884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8077 vdd d0 a_9133_n10154# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8078 a_26098_n1781# a_25677_n1781# a_24985_n1506# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8079 a_36967_n5935# a_36754_n5935# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8080 a_20833_n5603# a_20620_n5603# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8081 a_9888_364# a_14663_485# a_14985_485# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8082 a_21770_n7565# a_21557_n7565# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8083 a_30334_n7910# a_30862_n8363# a_31070_n8363# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8084 a_29069_n3313# a_29065_n3501# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8085 a_11401_9095# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8086 a_17828_n9322# a_18085_n9338# a_17863_n8018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8087 a_26099_n2335# a_25678_n2335# a_25362_n2244# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8088 a_11758_n2585# a_11545_n2585# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8089 a_35705_n8404# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8090 a_32010_4664# a_31589_4664# a_31072_4908# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8091 a_30861_8766# a_30648_8766# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8092 a_24006_7898# a_24263_7708# a_23068_8142# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8093 a_35391_4830# a_35391_4600# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8094 a_2573_n10656# a_2823_n5964# a_2774_n5948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8095 gnd d0 a_9136_n4639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8096 a_432_9334# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8097 a_21978_7968# a_21910_8479# a_21994_7508# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8098 a_15734_4968# a_15521_4968# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8099 a_38049_n7999# a_38063_n9319# a_38018_n9115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8100 a_30862_n10020# a_30649_n10020# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8101 gnd d1 a_13170_n7602# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8102 vdd d1 a_8195_n7638# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8103 a_32960_4327# a_33150_3545# a_33105_3558# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8104 a_37175_5235# a_36754_5235# a_37081_5354# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8105 a_18915_1722# a_19168_1709# a_17976_1412# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8106 a_28018_7482# a_28032_8585# a_27983_8775# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8107 a_33100_n6464# a_34087_n6236# a_34042_n6032# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8108 vdd a_38413_5792# a_38205_5792# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8109 a_5909_n8418# a_5488_n8418# a_5173_n7965# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8110 a_36129_2743# a_35708_2743# a_35392_2853# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8111 a_31071_5457# a_30650_5457# a_30335_5662# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8112 a_27036_3597# a_26615_3597# a_26097_3287# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8113 vdd a_8054_n9333# a_7846_n9333# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8114 vdd d2 a_33215_n9278# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8115 a_5702_n5109# a_5489_n5109# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8116 a_26828_n3194# a_26615_n3194# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8117 a_16674_1415# a_16461_1415# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8118 a_21041_6006# a_20620_6006# a_20304_5887# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8119 a_3823_2956# a_3826_2225# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8120 a_20305_3910# a_20834_3800# a_21042_3800# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8121 a_18908_8517# a_18911_7786# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8122 a_31072_2148# a_30651_2148# a_30337_1896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8123 a_17829_n7116# a_18019_n6540# a_17974_n6336# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8124 a_21041_n6706# a_21771_n6462# a_21979_n6462# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8125 a_16570_3042# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8126 vdd a_38272_n7113# a_38064_n7113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8127 a_15206_n3371# a_15206_n3142# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8128 a_26614_n6503# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8129 a_39098_8321# a_39351_8308# a_38159_8011# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8130 gnd a_13170_7976# a_12962_7976# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8131 a_7800_n2699# a_7990_n2123# a_7945_n1919# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8132 a_6430_1410# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8133 a_26095_9356# a_26825_9112# a_27033_9112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8134 a_32009_7973# a_31588_7973# a_31071_8217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8135 vdd a_28271_7469# a_28063_7469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8136 a_21038_n9461# a_20617_n9461# a_20302_n9465# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8137 vdd a_4078_n6250# a_3870_n6250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8138 a_12912_9269# a_13899_8835# a_13850_9025# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8139 a_11755_8503# a_11542_8503# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8140 a_29068_n3862# a_29321_n4066# a_28126_n4294# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8141 a_29064_2424# a_29070_1698# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8142 gnd a_8055_n7127# a_7847_n7127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8143 a_39093_n7364# a_39099_n6627# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8144 a_6849_5822# a_6428_5822# a_5911_6066# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8145 a_36784_8525# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8146 a_30334_n8367# a_30334_n7910# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8147 a_27246_522# a_27137_522# a_25140_461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8148 a_25362_1745# a_25362_1516# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8149 gnd a_19164_n8502# a_18956_n8502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8150 a_20303_8509# a_20830_8761# a_21038_8761# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8151 vdd a_39350_n7380# a_39142_n7380# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8152 a_26095_n8399# a_25674_n8399# a_25359_n7946# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8153 a_436_1613# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8154 vdd a_34294_6610# a_34086_6610# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8155 a_16881_2518# a_16814_1926# a_16892_3042# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8156 a_5172_n9984# a_5172_n9755# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8157 a_118_n5531# a_647_n5622# a_855_n5622# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8158 a_38154_9291# a_39141_8857# a_39096_8870# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8159 a_30862_7663# a_30649_7663# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8160 vdd a_19167_2812# a_18959_2812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8161 vdd a_4080_3869# a_3872_3869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8162 a_11755_n9203# a_11542_n9203# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8163 a_30863_4354# a_30650_4354# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8164 vdd a_25122_n10714# a_24914_n10714# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8165 a_15735_3865# a_15522_3865# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8166 a_18911_9443# a_19164_9430# a_17972_9133# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8167 a_434_4922# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8168 gnd a_8196_4703# a_7988_4703# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8169 a_26094_n9502# a_26825_n9812# a_27033_n9812# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8170 a_1481_n5908# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8171 vdd d2 a_8056_n4921# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8172 a_35393_n1790# a_35921_n1786# a_36129_n1786# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8173 a_25360_4595# a_25361_4138# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8174 a_26936_n8130# a_26723_n8130# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8175 a_21980_3556# a_21912_4067# a_21996_3096# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8176 vdd d7 a_30219_n10835# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8177 gnd a_9133_n10154# a_8925_n10154# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8178 a_15735_n4565# a_15522_n4565# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8179 a_33105_n2967# a_33358_n3171# a_32965_n2456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8180 a_26829_n2091# a_26616_n2091# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8181 a_12809_3053# a_12823_4156# a_12778_4169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8182 vdd a_38274_1972# a_38066_1972# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8183 a_37083_n3723# a_36786_n4813# a_37067_n4302# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8184 a_35393_n2020# a_35922_n2340# a_36130_n2340# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8185 a_20303_8322# a_20303_8093# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8186 a_29064_5184# a_29321_4994# a_28129_4697# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8187 gnd d3 a_13060_n8181# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8188 a_10887_n3421# a_10466_n3421# a_10150_n3101# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8189 a_18913_n2783# a_19166_n2987# a_17971_n3215# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8190 a_24010_n2357# a_24013_n1615# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8191 a_32009_n8673# a_31588_n8673# a_31071_n8917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8192 a_432_n10034# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8193 a_20305_n4596# a_20832_n5049# a_21040_n5049# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8194 gnd d0 a_29323_n2414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8195 a_38018_8603# a_38271_8590# a_38049_7487# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8196 a_28020_3070# a_28034_4173# a_27985_4363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8197 a_5176_n2450# a_5176_n2263# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8198 a_20621_n1740# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8199 gnd a_23325_n7578# a_23117_n7578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8200 gnd d1 a_33358_n4274# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8201 a_15521_n4011# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8202 a_31073_1045# a_30652_1045# a_30337_1250# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8203 a_15940_6620# a_15519_6620# a_15204_6825# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8204 vdd d0 a_9135_6116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8205 a_8882_3369# a_8878_3546# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8206 a_21040_n7809# a_20619_n7809# a_20303_n7718# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8207 a_33103_n7379# a_34087_n7893# a_34042_n7689# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8208 vdd d1 a_28382_n5413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8209 a_20622_n2294# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8210 a_5909_n10075# a_5488_n10075# a_5172_n9755# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8211 a_5173_7050# a_5173_6820# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8212 a_24964_n10698# a_24914_n10714# a_24865_n10698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8213 a_15940_n10080# a_16670_n9836# a_16878_n9836# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8214 a_2885_n2066# a_3872_n1838# a_3823_n1822# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8215 a_39100_3909# a_39353_3896# a_38161_3599# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8216 a_31801_7973# a_31588_7973# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8217 a_1371_n7584# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8218 a_7939_n5416# a_8926_n5188# a_8877_n5172# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8219 a_11757_4091# a_11544_4091# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8220 gnd a_4080_1109# a_3872_1109# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8221 a_34044_2765# a_34040_2942# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8222 a_36786_4113# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8223 a_18913_6134# a_18909_6311# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8224 a_30336_n3955# a_30336_n3498# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8225 a_10884_9339# a_10463_9339# a_10147_9220# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8226 a_1792_n8687# a_1371_n8687# a_853_n8377# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8227 vdd a_34296_2198# a_34088_2198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8228 a_22964_5229# a_23007_7428# a_22962_7441# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8229 a_25361_2848# a_25890_2738# a_26098_2738# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8230 a_17970_6001# a_18227_5811# a_17829_6593# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8231 a_33099_7044# a_34086_6610# a_34037_6800# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8232 a_30864_3251# a_30651_3251# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8233 a_26095_n10056# a_25674_n10056# a_25358_n9736# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8234 gnd a_34296_n6790# a_34088_n6790# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8235 a_16568_n8154# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8236 a_32965_n2456# a_33150_n3171# a_33105_n2967# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8237 a_28018_7482# a_28032_8585# a_27987_8598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8238 a_18910_8889# a_18906_9066# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8239 a_30334_6995# a_30863_7114# a_31071_7114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8240 a_35390_n8408# a_35918_n8404# a_36126_n8404# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8241 gnd d0 a_9132_8871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8242 a_12809_5253# a_13062_5240# a_12035_505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8243 a_6864_n8149# a_6750_n8149# a_6864_n5949# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8244 a_7937_n9828# a_8194_n9844# a_7801_n9129# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8245 a_22958_n8141# a_22977_n7067# a_22928_n7051# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8246 a_28125_n5397# a_29112_n5169# a_29063_n5153# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8247 a_24008_5143# a_24265_4953# a_23073_4656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8248 a_6429_n3213# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8249 a_30336_2812# a_30336_2583# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8250 vdd d2 a_8055_6398# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8251 a_10148_n8616# a_10148_n8386# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8252 a_648_3819# a_435_3819# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8253 a_31071_n7814# a_30650_n7814# a_30334_n7723# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8254 a_26826_n8709# a_26613_n8709# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8255 vdd d0 a_34293_8816# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8256 vdd a_39352_4999# a_39144_4999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8257 a_10149_5911# a_10678_6030# a_10886_6030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8258 a_5913_n2354# a_6643_n2110# a_6851_n2110# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8259 a_431_8780# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8260 a_855_6025# a_434_6025# a_118_5906# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8261 a_20620_2143# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8262 a_119_2597# a_119_2367# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8263 a_35920_6052# a_35707_6052# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8264 a_10676_n7279# a_10463_n7279# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8265 vdd d4 a_13062_n5969# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8266 a_21039_6555# a_21770_6865# a_21978_6865# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8267 vdd d0 a_4077_n8456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8268 a_11615_6889# a_11402_6889# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8269 a_38159_n8523# a_38412_n8727# a_38014_n9303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8270 a_25358_n9506# a_25359_n9049# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8271 a_10149_n5077# a_10677_n5073# a_10885_n5073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8272 a_36125_8807# a_35704_8807# a_35390_8555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8273 a_25677_n4541# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8274 a_15520_n5114# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8275 a_22929_4322# a_23119_3540# a_23070_3730# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8276 a_13851_6819# a_14108_6629# a_12913_7063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8277 a_646_7128# a_433_7128# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8278 gnd a_28273_n5986# a_28065_n5986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8279 gnd d0 a_4080_n3495# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8280 vdd d0 a_14110_n2946# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8281 a_25361_2619# a_25361_2389# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8282 a_15942_2208# a_15521_2208# a_15206_2413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8283 gnd a_4076_8830# a_3868_8830# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8284 a_20302_8966# a_20303_8509# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8285 gnd a_23215_n8157# a_23007_n8157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8286 a_2778_n3560# a_3031_n3764# a_2774_n5948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8287 a_32991_3211# a_33010_1931# a_32965_1944# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8288 gnd d2 a_18086_6403# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8289 vdd a_3141_n4288# a_2933_n4288# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8290 a_12772_n9281# a_13029_n9297# a_12807_n7977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8291 a_35393_1291# a_35395_1192# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8292 a_30651_4908# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8293 a_5173_8382# a_5702_8272# a_5910_8272# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8294 a_35391_n5558# a_35920_n5649# a_36128_n5649# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8295 a_15521_n5668# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8296 a_36128_n2889# a_35707_n2889# a_35393_n2436# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8297 a_7944_n4125# a_8928_n4639# a_8879_n4623# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8298 vdd a_33359_n2068# a_33151_n2068# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8299 a_32995_n3546# a_33009_n4866# a_32960_n4850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8300 a_31803_3561# a_31590_3561# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8301 a_6639_9131# a_6426_9131# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8302 a_32020_n5717# a_31911_n5894# a_32119_n5894# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8303 a_27045_7430# a_26936_7430# a_27050_5349# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8304 gnd d2 a_2999_6357# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8305 a_15521_3311# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8306 a_12777_n6887# a_12962_n7602# a_12913_n7586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8307 a_30649_6560# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8308 a_36129_n3443# a_35708_n3443# a_35392_n3352# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8309 a_28126_n3191# a_28383_n3207# a_27990_n2492# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8310 a_18910_1345# a_15209_1211# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8311 a_6848_n8728# a_6780_n9239# a_6864_n8149# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8312 a_31730_n4772# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8313 a_18907_9620# a_19164_9430# a_17972_9133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8314 a_10885_8236# a_10464_8236# a_10148_8346# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8315 a_12917_6886# a_13170_6873# a_12777_6375# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8316 a_3824_7740# a_3820_7917# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8317 gnd a_13030_6362# a_12822_6362# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8318 a_22759_n10637# a_23009_n5945# a_22964_n5741# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8319 a_25362_1516# a_25891_1635# a_26099_1635# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8320 a_29066_n2398# a_29069_n1656# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8321 a_17972_1589# a_18229_1399# a_17831_2181# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8322 a_26828_2494# a_26615_2494# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8323 a_5490_6066# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8324 a_18908_n5177# a_18914_n4440# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8325 a_20304_n6156# a_20304_n5699# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8326 a_18911_6683# a_18907_6860# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8327 a_30864_n2848# a_30651_n2848# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8328 vdd a_14108_n10118# a_13900_n10118# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8329 a_15940_n10080# a_15519_n10080# a_15203_n9989# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8330 a_21558_n6462# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8331 a_28020_3070# a_28034_4173# a_27989_4186# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8332 a_28130_n4106# a_29114_n4620# a_29065_n4604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8333 a_22927_8734# a_23117_7952# a_23072_7965# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8334 a_36998_6319# a_36785_6319# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8335 a_38155_8188# a_38412_7998# a_38014_8780# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8336 a_13857_n2742# a_13853_n2930# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8337 a_12912_n9792# a_13899_n9564# a_13854_n9360# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8338 vdd a_19168_n2438# a_18960_n2438# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8339 a_31911_5194# a_31698_5194# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8340 vdd d0 a_34295_4404# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8341 a_31071_n7814# a_31801_n7570# a_32009_n7570# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8342 a_11402_n7589# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8343 a_5910_n8972# a_6640_n8728# a_6848_n8728# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8344 a_36644_n7611# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8345 a_857_n2313# a_436_n2313# a_120_n2222# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8346 a_36126_7704# a_35705_7704# a_35390_7909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8347 a_3821_n7891# a_3824_n7149# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8348 a_1583_n9790# a_1370_n9790# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8349 a_21041_2143# a_21772_2453# a_21980_2453# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8350 a_21557_7968# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8351 a_39097_n2403# a_39354_n2419# a_38162_n1905# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8352 gnd a_24266_n3476# a_24058_n3476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8353 a_39098_n4970# a_39351_n5174# a_38156_n5402# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8354 gnd a_9135_6116# a_8927_6116# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8355 gnd a_14112_n2397# a_13904_n2397# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8356 gnd d1 a_8197_2497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8357 vdd d0 a_4077_n10113# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8358 a_16880_n5424# a_16459_n5424# a_15941_n5114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8359 gnd d2 a_18088_1991# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8360 a_22960_3206# a_22979_1926# a_22934_1939# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8361 a_20303_n7718# a_20832_n7809# a_21040_n7809# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8362 a_27144_n5930# a_26723_n5930# a_27045_n5753# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8363 a_29064_n4050# a_29321_n4066# a_28126_n4294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8364 a_32009_6870# a_31942_6278# a_32020_7394# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8365 a_21038_n9461# a_21769_n9771# a_21977_n9771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8366 a_117_n7508# a_117_n7278# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8367 vdd d0 a_39351_7205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8368 vdd a_33356_n8686# a_33148_n8686# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8369 a_9776_n10838# a_10033_n10854# a_9875_n10838# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8370 vdd d0 a_24264_n6231# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8371 a_26612_n9812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8372 gnd d2 a_28241_n7108# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8373 a_33099_7044# a_34086_6610# a_34041_6623# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8374 a_20832_4349# a_20619_4349# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8375 a_7834_n3601# a_7848_n4921# a_7803_n4717# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8376 a_21913_1861# a_21700_1861# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8377 a_27047_3018# a_26938_3018# a_27045_5230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8378 a_29067_n7725# a_29063_n7913# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8379 a_16673_n3218# a_16460_n3218# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8380 a_35708_n1786# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8381 gnd d2 a_3001_1945# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8382 a_26095_9356# a_25674_9356# a_25358_9237# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8383 a_15943_3865# a_16673_3621# a_16881_3621# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8384 gnd a_3141_2456# a_2933_2456# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8385 a_30336_2583# a_30336_2353# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8386 a_18909_5208# a_19166_5018# a_17974_4721# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8387 a_15521_4968# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8388 a_12809_n5765# a_12852_n8181# a_12803_n8165# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8389 a_11542_n9203# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8390 vdd d4 a_8087_n6005# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8391 a_35709_n2340# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8392 gnd a_38411_9101# a_38203_9101# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8393 a_20619_n5049# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8394 a_12805_5430# a_13062_5240# a_12035_505# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8395 a_32012_1355# a_31944_1866# a_32022_2982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8396 a_35918_6601# a_35705_6601# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8397 a_1795_1369# a_1374_1369# a_857_1613# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8398 a_7800_2176# a_7990_1394# a_7941_1584# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8399 a_18995_288# d8 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8400 a_21880_n5889# a_21667_n5889# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8401 vdd d1 a_3140_n5391# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8402 a_15733_5517# a_15520_5517# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8403 a_10886_4927# a_11616_4683# a_11824_4683# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8404 a_38016_4368# a_38273_4178# a_38051_3075# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8405 a_20306_n1744# a_19886_n1571# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8406 a_17968_9310# a_18955_8876# a_18906_9066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8407 a_30861_n9466# a_30648_n9466# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8408 a_5174_n6862# a_5701_n7315# a_5909_n7315# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8409 a_10147_n9948# a_10147_n9719# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8410 a_33099_8147# a_33356_7957# a_32958_8739# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8411 a_17859_7683# a_17878_6403# a_17833_6416# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8412 a_31073_2702# a_30652_2702# a_30336_2583# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8413 a_28020_n3582# a_28034_n4902# a_27989_n4698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8414 a_16461_1415# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8415 a_22929_4322# a_23119_3540# a_23074_3553# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8416 a_16457_n9836# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8417 a_15733_n7874# a_15520_n7874# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8418 a_8881_7232# a_8877_7409# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8419 a_13857_4990# a_14110_4977# a_12918_4680# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8420 a_16882_n2115# a_16814_n2626# a_16892_n3565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8421 a_433_n5068# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8422 a_36128_3292# a_35707_3292# a_35392_3497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8423 a_30334_6765# a_30862_6560# a_31070_6560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8424 a_39100_n4421# a_39353_n4625# a_38161_n4111# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8425 a_24009_n4563# a_24266_n4579# a_23074_n4065# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8426 a_16895_5373# a_16781_5254# a_16989_5254# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8427 a_31700_n3682# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8428 a_29064_3527# a_29321_3337# a_28126_3771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8429 a_15205_6181# a_15205_5952# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8430 a_24010_n7130# a_24263_n7334# a_23068_n7562# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8431 a_38156_n6505# a_39143_n6277# a_39098_n6073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8432 vdd d2 a_23186_n4861# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8433 a_10149_5681# a_10677_5476# a_10885_5476# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8434 a_3826_n6600# a_4079_n6804# a_2887_n6290# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8435 a_10149_n5723# a_10149_n5536# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8436 vdd a_13030_6362# a_12822_6362# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8437 a_1808_5327# a_1694_5208# a_1902_5208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8438 a_35919_n5095# a_35706_n5095# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8439 a_38161_3599# a_39145_3896# a_39100_3909# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8440 a_21770_n7565# a_21557_n7565# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8441 a_32961_2121# a_33151_1339# a_33102_1529# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8442 a_26096_8253# a_25675_8253# a_25359_8363# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8443 a_30334_n8367# a_30862_n8363# a_31070_n8363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8444 a_116_9215# a_116_8985# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8445 a_645_6574# a_432_6574# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8446 a_33101_2632# a_34088_2198# a_34043_2211# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8447 vdd d0 a_19163_n9605# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8448 a_26099_n2335# a_25678_n2335# a_25362_n2015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8449 a_35389_9471# a_35918_9361# a_36126_9361# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8450 a_35705_n8404# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8451 a_2881_n9787# a_3138_n9803# a_2745_n9088# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8452 vdd d0 a_34295_n6236# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8453 vdd a_9134_n6291# a_8926_n6291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8454 a_30650_4354# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8455 a_30337_n2208# a_30866_n2299# a_31074_n2299# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8456 a_17828_8799# a_18018_8017# a_17973_8030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8457 a_15522_3865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8458 a_37066_5808# a_36645_5808# a_36128_6052# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8459 gnd d1 a_28381_6890# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8460 a_119_n2866# a_120_n2409# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8461 a_12917_6886# a_13901_7183# a_13852_7373# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8462 vdd a_39352_n4071# a_39144_n4071# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8463 a_28123_9286# a_28380_9096# a_27987_8598# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8464 vdd a_29321_n2963# a_29113_n2963# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8465 a_12604_n10661# a_12854_n5969# a_12809_n5765# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8466 a_2882_n8684# a_3869_n8456# a_3824_n8252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8467 a_11614_n9795# a_11401_n9795# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8468 a_27144_n5930# a_28072_n10694# a_24865_n10698# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8469 a_1810_n3696# a_1513_n4786# a_1793_n5378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8470 a_10464_n5073# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8471 a_25362_1932# a_25362_1745# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8472 a_1372_n6481# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8473 a_30863_n8917# a_30650_n8917# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8474 a_10884_7682# a_10463_7682# a_10148_7430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8475 a_23072_6862# a_24056_7159# a_24011_7172# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8476 a_24008_n6769# a_24011_n6027# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8477 a_12915_n3174# a_13902_n2946# a_13857_n2742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8478 gnd d0 a_9137_1704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8479 a_27033_9112# a_26966_8520# a_27050_7549# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8480 gnd d0 a_24265_n5682# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8481 a_2889_n1878# a_3142_n2082# a_2744_n2658# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8482 a_12776_8581# a_12961_9079# a_12916_9092# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8483 a_39099_n6627# a_39095_n6815# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8484 a_15735_1105# a_15522_1105# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8485 a_28126_2668# a_28383_2478# a_27990_1980# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8486 a_35707_n5649# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8487 gnd a_18228_n3231# a_18020_n3231# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8488 a_10885_n6176# a_10464_n6176# a_10149_n5723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8489 a_18913_n3886# a_18909_n4074# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8490 a_39098_7218# a_39094_7395# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8491 vdd a_9135_6116# a_8927_6116# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8492 a_16890_7454# a_16781_7454# a_16895_5373# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8493 a_15203_n9760# a_15732_n10080# a_15940_n10080# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8494 a_21910_n9179# a_21697_n9179# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8495 a_31698_n5894# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8496 a_435_n4519# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8497 a_38161_n3008# a_38414_n3212# a_38021_n2497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8498 a_25888_7150# a_25675_7150# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8499 gnd a_4077_n10113# a_3869_n10113# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8500 a_38155_7085# a_39142_6651# a_39093_6841# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8501 a_853_n10034# a_432_n10034# a_116_n9714# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8502 a_10678_n3970# a_10465_n3970# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8503 a_6567_n9239# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8504 a_1803_7408# a_1694_7408# a_1808_5327# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8505 a_21038_n9461# a_20617_n9461# a_20303_n9008# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8506 a_25361_n4637# a_25888_n5090# a_26096_n5090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8507 gnd a_4081_1663# a_3873_1663# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8508 vdd d0 a_9136_n1879# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8509 a_36858_4705# a_36645_4705# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8510 a_23068_n8665# a_24055_n8437# a_24010_n8233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8511 a_32010_n6467# a_31942_n6978# a_32020_n7917# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8512 a_18908_n7937# a_19165_n7953# a_17973_n7439# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8513 a_21996_n3677# a_21699_n4767# a_21979_n5359# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8514 a_6848_n7625# a_6427_n7625# a_5910_n7869# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8515 gnd d1 a_38414_n4315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8516 a_5489_5512# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8517 a_10151_1269# a_10679_1064# a_10887_1064# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8518 a_35389_n10157# a_39093_n10124# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8519 vdd a_3141_2456# a_2933_2456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8520 a_38159_n7420# a_39143_n7934# a_39098_n7730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8521 a_2885_9087# a_3138_9074# a_2745_8576# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8522 a_646_5471# a_433_5471# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8523 a_647_2162# a_434_2162# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8524 a_30651_3251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8525 a_18912_n6092# a_19165_n6296# a_17970_n6524# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8526 a_16671_6930# a_16458_6930# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8527 a_26095_n10056# a_26825_n9812# a_27033_n9812# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8528 a_21043_1594# a_20622_1594# a_20306_1475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8529 a_17859_7683# a_18116_7493# a_17865_5294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8530 a_37068_1396# a_36647_1396# a_36130_1640# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8531 a_35391_5703# a_35391_5246# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8532 a_31588_n7570# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8533 a_6859_n7972# a_6568_n7033# a_6849_n6522# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8534 gnd a_14109_n5152# a_13901_n5152# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8535 gnd d0 a_14109_n9015# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8536 a_38160_n5214# a_39144_n5728# a_39095_n5712# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8537 gnd a_9132_8871# a_8924_8871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8538 vdd d0 a_34295_n7893# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8539 a_6849_4719# a_6428_4719# a_5910_4409# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8540 vdd a_29318_n9581# a_29110_n9581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8541 vdd a_8055_6398# a_7847_6398# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8542 vdd a_34293_8816# a_34085_8816# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8543 a_435_3819# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8544 a_645_n7274# a_432_n7274# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8545 a_32009_n8673# a_31588_n8673# a_31070_n8363# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8546 a_10886_3270# a_10465_3270# a_10150_3018# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8547 a_11402_6889# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8548 a_2885_n9599# a_3869_n10113# a_116_n10130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8549 a_8882_n5538# a_8878_n5726# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8550 a_32011_2458# a_31590_2458# a_31073_2702# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8551 a_24007_5692# a_24264_5502# a_23069_5936# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8552 a_20619_n7809# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8553 a_27984_n7092# a_28174_n6516# a_28125_n6500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8554 gnd a_9135_n5742# a_8927_n5742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8555 a_25361_n3991# a_25889_n3987# a_26097_n3987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8556 a_433_7128# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8557 a_21556_n9771# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8558 a_20302_n9695# a_20831_n10015# a_21039_n10015# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8559 a_16892_3042# a_16783_3042# a_16890_5254# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8560 a_36859_n3199# a_36646_n3199# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8561 a_13856_7196# a_13852_7373# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8562 a_23073_n5168# a_23326_n5372# a_22933_n4657# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8563 a_35392_2853# a_35392_2624# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8564 a_30337_1896# a_30337_1709# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8565 a_27045_n7953# a_26754_n7014# a_27035_n6503# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8566 a_15207_1540# a_15207_1310# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8567 a_20305_3451# a_20305_2994# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8568 a_10150_n3101# a_10150_n2871# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8569 a_36859_3602# a_36646_3602# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8570 a_31590_3561# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8571 a_6426_9131# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8572 a_15942_6071# a_15521_6071# a_15205_5952# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8573 gnd a_13169_n9808# a_12961_n9808# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8574 a_1805_2996# a_1696_2996# a_1803_5208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8575 vdd d0 a_9133_n8497# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8576 a_5175_n4469# a_5704_n4560# a_5912_n4560# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8577 gnd d1 a_23326_n6475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8578 a_2889_n1878# a_3873_n2392# a_3824_n2376# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8579 a_28014_7659# a_28033_6379# a_27984_6569# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8580 gnd d1 a_23324_9055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8581 a_12917_6886# a_13901_7183# a_13856_7196# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8582 a_433_n7828# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8583 a_24009_n9336# a_24005_n9524# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8584 a_23071_n9580# a_24055_n10094# a_20302_n10111# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8585 a_24013_2760# a_24266_2747# a_23074_2450# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8586 vdd a_8197_n4329# a_7989_n4329# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8587 a_2747_n4676# a_2932_n5391# a_2887_n5187# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8588 a_26615_2494# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8589 a_28128_6903# a_29112_7200# a_29063_7390# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8590 a_5488_n7315# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8591 a_29064_n6810# a_29067_n6068# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8592 vdd a_38415_n2109# a_38207_n2109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8593 a_34037_n8426# a_34294_n8442# a_33099_n8670# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8594 a_38018_n9115# a_38271_n9319# a_38049_n7999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8595 a_32027_3101# a_31730_4072# a_32010_4664# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8596 a_27035_n5400# a_26614_n5400# a_26097_n5644# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8597 a_15944_n2359# a_15523_n2359# a_15207_n2039# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8598 a_3828_n2188# a_3824_n2376# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8599 vdd d0 a_39351_5548# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8600 a_11756_6297# a_11543_6297# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8601 gnd d1 a_18227_n5437# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8602 a_13856_4436# a_14109_4423# a_12914_4857# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8603 a_11826_n2074# a_11758_n2585# a_11836_n3524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8604 a_5173_7279# a_5173_7050# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8605 a_39093_7944# a_39098_7218# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8606 a_5909_n8418# a_5488_n8418# a_5173_n8422# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8607 a_5176_1305# a_5704_1100# a_5912_1100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8608 vdd d0 a_14109_n6255# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8609 a_16601_n2626# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8610 a_18914_1168# a_18910_1345# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8611 a_36785_6319# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8612 a_647_n6725# a_434_n6725# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8613 a_31071_n7814# a_30650_n7814# a_30334_n7494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8614 a_36967_5235# a_36754_5235# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8615 a_20304_6303# a_20831_6555# a_21039_6555# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8616 vdd a_34295_4404# a_34087_4404# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8617 a_25358_n10152# a_25358_n9965# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8618 a_15205_4849# a_15205_4619# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8619 a_10149_5224# a_10149_5037# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8620 a_38155_7085# a_39142_6651# a_39097_6664# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8621 a_30863_5457# a_30650_5457# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8622 a_34039_n5671# a_34296_n5687# a_33104_n5173# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8623 a_5176_1764# a_5176_1535# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8624 vdd a_4081_1663# a_3873_1663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8625 a_24009_1280# a_24266_1090# a_23071_1524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8626 a_30864_2148# a_30651_2148# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8627 a_117_8528# a_117_8341# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8628 a_18912_7237# a_19165_7224# a_17973_6927# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8629 a_15736_1659# a_15523_1659# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8630 gnd a_8197_2497# a_7989_2497# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8631 a_3825_8294# a_4078_8281# a_2886_7984# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8632 gnd d0 a_39353_2793# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8633 a_30333_9201# a_30862_9320# a_31070_9320# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8634 a_27033_9112# a_26612_9112# a_26094_8802# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8635 a_38015_n7097# a_38205_n6521# a_38156_n6505# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8636 a_17968_n9833# a_18955_n9605# a_18910_n9401# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8637 a_21042_n3397# a_21772_n3153# a_21980_n3153# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8638 vdd d2 a_8054_8604# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8639 a_31698_5194# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8640 vdd d0 a_14111_n3500# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8641 a_30653_n2299# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8642 a_25140_461# a_26924_522# a_27144_5230# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8643 a_2881_9264# a_3138_9074# a_2745_8576# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8644 a_5173_7923# a_5173_7466# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8645 a_15941_n5114# a_16672_n5424# a_16880_n5424# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8646 a_12805_n3753# a_13062_n3769# a_12805_n5953# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8647 vdd a_34296_n4030# a_34088_n4030# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8648 a_15204_7928# a_15732_7723# a_15940_7723# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8649 a_21700_1861# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8650 a_38019_6397# a_38272_6384# a_38045_7664# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8651 a_36129_n3443# a_35708_n3443# a_35392_n3123# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8652 vdd a_4079_n2941# a_3871_n2941# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8653 a_855_n6725# a_1585_n6481# a_1793_n6481# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8654 a_28016_3247# a_28035_1967# a_27986_2157# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8655 gnd d0 a_14108_n7358# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8656 a_21038_8761# a_20617_8761# a_20302_8966# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8657 a_22928_6528# a_23118_5746# a_23069_5936# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8658 a_11545_n2585# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8659 a_34040_4045# a_34043_3314# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8660 a_13850_9025# a_14107_8835# a_12912_9269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8661 a_16892_3042# a_16601_1926# a_16882_1415# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8662 gnd a_8196_n6535# a_7988_n6535# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8663 gnd d2 a_18085_8609# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8664 a_29068_5007# a_29064_5184# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8665 a_25359_n7759# a_25888_n7850# a_26096_n7850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8666 a_26096_n5090# a_25675_n5090# a_25361_n4637# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8667 a_11618_n2074# a_11405_n2074# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8668 vdd d3 a_18116_n8222# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8669 a_35705_6601# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8670 a_25360_n5553# a_25360_n5324# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8671 a_8880_1894# a_8883_1163# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8672 a_11617_2477# a_11404_2477# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8673 vdd a_38412_n8727# a_38204_n8727# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8674 a_17972_9133# a_18956_9430# a_18907_9620# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8675 vdd d5 a_12861_n10677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8676 a_31802_5767# a_31589_5767# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8677 vdd d8 a_20790_n10911# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8678 a_36646_2499# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8679 a_15520_5517# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8680 a_29067_5556# a_29320_5543# a_28125_5977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8681 a_5174_5073# a_5174_4844# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8682 a_26097_n5644# a_25676_n5644# a_25360_n5553# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8683 vdd a_13031_n4885# a_12823_n4885# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8684 a_11758_1885# a_11545_1885# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8685 a_6643_n2110# a_6430_n2110# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8686 gnd d0 a_9134_n7948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8687 a_20621_n1740# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8688 gnd a_13029_8568# a_12821_8568# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8689 a_31800_9076# a_31587_9076# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8690 a_13851_7922# a_13856_7196# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8691 a_13852_n7896# a_14109_n7912# a_12917_n7398# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8692 a_25675_n5090# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8693 a_7941_n2107# a_8928_n1879# a_8883_n1675# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8694 a_20306_1891# a_20833_2143# a_21041_2143# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8695 a_857_n2313# a_436_n2313# a_120_n1993# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8696 a_5175_2867# a_5704_2757# a_5912_2757# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8697 a_26827_4700# a_26614_4700# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8698 a_17971_3795# a_18228_3605# a_17830_4387# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8699 a_38157_2673# a_39144_2239# a_39099_2252# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8700 a_30865_1045# a_30652_1045# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8701 gnd d0 a_24264_8262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8702 a_3821_8471# a_3824_7740# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8703 a_7804_n2511# a_7989_n3226# a_7940_n3210# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8704 a_36955_527# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8705 a_2672_n10656# a_4936_n10733# a_4778_n10717# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8706 a_8880_n2417# a_8883_n1675# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8707 a_18914_2825# a_19167_2812# a_17975_2515# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8708 a_32965_n2456# a_33218_n2660# a_32991_n3734# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8709 vdd d1 a_23324_9055# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8710 a_21039_n10015# a_21769_n9771# a_21977_n9771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8711 a_17832_n9134# a_18017_n9849# a_17972_n9645# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8712 vdd d2 a_8056_4192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8713 a_18908_7414# a_18911_6683# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8714 a_26612_n9812# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8715 a_23071_9068# a_24055_9365# a_24006_9555# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8716 a_16890_n7977# a_16599_n7038# a_16880_n6527# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8717 a_432_6574# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8718 a_15943_n1805# a_15522_n1805# a_15207_n1809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8719 a_17830_n4910# a_18020_n4334# a_17975_n4130# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8720 a_12917_n8501# a_13901_n9015# a_13852_n8999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8721 a_29065_n4604# a_29322_n4620# a_28130_n4106# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8722 a_21040_4349# a_21771_4659# a_21979_4659# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8723 a_28127_n2088# a_29114_n1860# a_29069_n1656# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8724 a_38021_1985# a_38274_1972# a_38047_3252# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8725 vdd a_4076_n9559# a_3868_n9559# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8726 a_28129_4697# a_28382_4684# a_27989_4186# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8727 a_13854_n3484# a_13857_n2742# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8728 a_33104_5764# a_33357_5751# a_32959_6533# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8729 a_33100_n6464# a_33357_n6480# a_32959_n7056# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8730 a_34044_n3277# a_34040_n3465# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8731 a_35921_n1786# a_35708_n1786# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8732 a_13852_4613# a_14109_4423# a_12914_4857# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8733 a_11542_n9203# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8734 a_16813_n4832# a_16600_n4832# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8735 a_5911_4963# a_5490_4963# a_5174_4844# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8736 gnd d0 a_34294_n10099# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8737 gnd d2 a_18087_4197# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8738 a_29066_n8274# a_29319_n8478# a_28124_n8706# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8739 a_11617_n3177# a_11404_n3177# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8740 a_5174_6176# a_5703_6066# a_5911_6066# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8741 a_10883_n9485# a_10462_n9485# a_10148_n9032# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8742 a_17831_n2704# a_18021_n2128# a_17972_n2112# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8743 a_30334_n7264# a_30335_n6807# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8744 a_22081_481# a_21868_481# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8745 a_26826_n8709# a_26613_n8709# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8746 a_25676_n3987# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8747 a_31804_1355# a_31591_1355# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8748 gnd a_9137_1704# a_8929_1704# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8749 a_33098_9250# a_34085_8816# a_34040_8829# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8750 a_30861_n9466# a_30648_n9466# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8751 a_5173_n7319# a_5701_n7315# a_5909_n7315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8752 a_29069_1144# a_29322_1131# a_28127_1565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8753 a_15522_1105# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8754 a_12035_505# a_12854_5240# a_12805_5430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8755 a_15942_6071# a_16672_5827# a_16880_5827# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8756 a_6640_n8728# a_6427_n8728# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8757 a_6851_1410# a_6430_1410# a_5912_1100# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8758 a_18911_n8298# a_18907_n8486# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8759 a_18908_7414# a_19165_7224# a_17973_6927# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8760 a_10886_6030# a_10465_6030# a_10149_6140# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8761 a_30335_n6620# a_30335_n6391# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8762 a_35391_n5099# a_35919_n5095# a_36127_n5095# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8763 a_3821_8471# a_4078_8281# a_2886_7984# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8764 a_3819_n9543# a_3825_n8806# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8765 gnd a_13031_4156# a_12823_4156# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8766 a_21981_n2050# a_21560_n2050# a_21043_n2294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8767 a_15733_n7874# a_15520_n7874# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8768 a_12916_n9604# a_13900_n10118# a_13851_n10102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8769 a_5176_1535# a_5705_1654# a_5913_1654# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8770 a_17660_n10702# a_17910_n6010# a_17865_n5806# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8771 a_21978_6865# a_21557_6865# a_21040_7109# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8772 a_7938_n8725# a_8925_n8497# a_8880_n8293# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8773 a_25675_7150# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8774 gnd d0 a_4079_4972# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8775 a_5491_n4560# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8776 a_16881_n3218# a_16814_n2626# a_16892_n3565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8777 a_35917_8807# a_35704_8807# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8778 a_35391_n5329# a_35920_n5649# a_36128_n5649# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8779 vdd a_28382_n5413# a_28174_n5413# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8780 a_6642_2513# a_6429_2513# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8781 a_15939_8826# a_16670_9136# a_16878_9136# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8782 a_3822_6265# a_3825_5534# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8783 a_10885_n6176# a_11616_n6486# a_11824_n6486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8784 a_35392_n4455# a_35392_n4226# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8785 a_32991_n3734# a_33010_n2660# a_32965_n2456# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8786 gnd d0 a_24266_3850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8787 a_20303_7219# a_20303_6990# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8788 a_17829_6593# a_18019_5811# a_17970_6001# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8789 a_10885_7133# a_11615_6889# a_11823_6889# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8790 a_7941_n2107# a_8198_n2123# a_7800_n2699# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8791 a_10150_2831# a_10150_2602# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8792 a_38015_6574# a_38272_6384# a_38045_7664# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8793 gnd d1 a_33356_n7583# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8794 a_31072_4908# a_30651_4908# a_30335_4789# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8795 gnd d1 a_8195_n8741# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8796 a_22928_6528# a_23118_5746# a_23073_5759# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8797 a_32962_n9074# a_33215_n9278# a_32993_n7958# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8798 a_23075_n1859# a_24059_n2373# a_24014_n2169# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8799 a_29063_5733# a_29068_5007# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8800 a_8882_2266# a_8878_2443# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8801 a_433_5471# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8802 a_3825_n4943# a_3821_n5131# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8803 a_21040_n6152# a_20619_n6152# a_20304_n5699# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8804 a_34041_9383# a_34294_9370# a_33102_9073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8805 a_16811_8544# a_16598_8544# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8806 a_20306_1704# a_20306_1475# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8807 a_23073_4656# a_24057_4953# a_24008_5143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8808 a_434_2162# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8809 a_36127_5498# a_35706_5498# a_35391_5703# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8810 a_15940_n8423# a_15519_n8423# a_15204_n8427# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8811 a_29068_n6622# a_29321_n6826# a_28129_n6312# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8812 a_17972_9133# a_18956_9430# a_18911_9443# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8813 a_30333_8971# a_30861_8766# a_31069_8766# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8814 a_12777_6375# a_12962_6873# a_12913_7063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8815 a_28124_n8706# a_29111_n8478# a_29066_n8274# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8816 a_12914_n6483# a_13901_n6255# a_13856_n6051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8817 a_29063_5733# a_29320_5543# a_28125_5977# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8818 a_20833_n3946# a_20620_n3946# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8819 a_25887_n7296# a_25674_n7296# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8820 a_2774_3225# a_2793_1945# a_2748_1958# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8821 a_11542_8503# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8822 a_18913_5031# a_18909_5208# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8823 vdd a_39353_n4625# a_39145_n4625# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8824 a_30863_n8917# a_30650_n8917# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8825 a_30336_n2852# a_30337_n2395# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8826 a_39096_n1849# a_39353_n1865# a_38158_n2093# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8827 a_13854_2961# a_13857_2230# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8828 a_31070_n7260# a_31801_n7570# a_32009_n7570# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8829 vdd a_24263_n7334# a_24055_n7334# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8830 vdd d0 a_4079_n6804# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8831 a_27986_n2680# a_28243_n2696# a_28016_n3770# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8832 a_33100_4838# a_34087_4404# a_34042_4417# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8833 a_5909_n8418# a_6640_n8728# a_6848_n8728# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8834 a_22858_n10637# a_22808_n10653# a_22088_n5889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8835 a_20305_n4409# a_20834_n4500# a_21042_n4500# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8836 vdd d0 a_24264_8262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8837 a_1727_n2580# a_1514_n2580# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8838 vdd d5 a_7886_n10713# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8839 a_21559_n3153# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8840 gnd a_39350_n8483# a_39142_n8483# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8841 a_5174_n6216# a_5174_n5759# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8842 a_12919_n2986# a_13903_n3500# a_13858_n3296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8843 gnd d1 a_28380_9096# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8844 a_12916_9092# a_13900_9389# a_13851_9579# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8845 a_16459_n5424# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8846 a_24010_1834# a_24013_1103# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8847 vdd d1 a_18229_1399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8848 a_29069_2801# a_29322_2788# a_28130_2491# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8849 a_35918_7704# a_35705_7704# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8850 gnd a_39354_n2419# a_39146_n2419# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8851 a_38051_n5787# a_38094_n8203# a_38045_n8187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8852 gnd a_24264_n5128# a_24056_n5128# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8853 a_20303_n7489# a_20832_n7809# a_21040_n7809# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8854 a_27144_n5930# a_26723_n5930# a_27050_n5930# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8855 a_20304_5013# a_20304_4784# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8856 a_10148_n7513# a_10148_n7283# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8857 a_36125_n9507# a_35704_n9507# a_35389_n9511# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8858 gnd a_4080_n4598# a_3872_n4598# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8859 a_23071_9068# a_24055_9365# a_24010_9378# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8860 a_36127_8258# a_36857_8014# a_37065_8014# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8861 gnd a_28271_7469# a_28063_7469# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8862 gnd d0 a_39350_7754# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8863 a_21996_n3677# a_21699_n4767# a_21980_n4256# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8864 a_31073_3805# a_30652_3805# a_30336_3915# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8865 gnd a_28381_n8722# a_28173_n8722# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8866 a_6848_n7625# a_6427_n7625# a_5909_n7315# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8867 a_10887_2721# a_11617_2477# a_11825_2477# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8868 a_25675_n7850# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8869 a_28125_4874# a_28382_4684# a_27989_4186# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8870 a_17865_n5806# a_17908_n8222# a_17863_n8018# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8871 gnd a_23324_9055# a_23116_9055# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8872 a_33100_5941# a_33357_5751# a_32959_6533# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8873 vdd d0 a_9137_n2433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8874 a_17835_2004# a_18020_2502# a_17975_2515# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8875 vdd a_3139_n7597# a_2931_n7597# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8876 gnd d3 a_33246_n8162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8877 a_34039_3491# a_34044_2765# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8878 a_1587_n2069# a_1374_n2069# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8879 a_25887_9356# a_25674_9356# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8880 a_30334_7411# a_30862_7663# a_31070_7663# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8881 a_16813_4132# a_16600_4132# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8882 a_3823_1299# a_122_1165# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8883 a_35392_3040# a_35392_2853# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8884 vdd d0 a_24265_n2922# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8885 a_7942_n7434# a_8926_n7948# a_8877_n7932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8886 a_21772_n3153# a_21559_n3153# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8887 a_36129_1086# a_35708_1086# a_35393_1291# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8888 a_17974_4721# a_18958_5018# a_18913_5031# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8889 a_30335_4559# a_30863_4354# a_31071_4354# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8890 vdd d0 a_14110_2217# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8891 a_8883_3923# a_8879_4100# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8892 vdd d3 a_8085_7488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8893 gnd d1 a_28382_n6516# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8894 a_33103_n8482# a_34087_n8996# a_34038_n8980# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8895 a_29065_1321# a_29322_1131# a_28127_1565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8896 a_12035_505# a_12854_5240# a_12809_5253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8897 a_25889_n6747# a_25676_n6747# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8898 gnd a_18118_n3810# a_17910_n3810# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8899 a_5488_7718# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8900 vdd d7 a_10033_n10854# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8901 a_119_n3512# a_647_n3965# a_855_n3965# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8902 a_24006_n8421# a_24011_n7684# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8903 a_6859_n5772# a_6539_n3737# a_6866_n3737# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8904 a_34040_8829# a_34036_9006# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8905 a_28127_n9621# a_29111_n10135# a_25358_n10152# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8906 gnd d1 a_13172_n3190# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8907 vdd a_13031_4156# a_12823_4156# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8908 a_35920_3292# a_35707_3292# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8909 vdd a_24265_n6785# a_24057_n6785# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8910 a_3824_6637# a_3820_6814# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8911 a_36754_5235# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8912 a_645_n7274# a_432_n7274# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8913 a_20618_9315# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8914 a_645_7677# a_432_7677# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8915 a_39093_n8467# a_39350_n8483# a_38155_n8711# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8916 a_35708_2743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8917 a_26097_6047# a_25676_6047# a_25360_6157# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8918 a_30865_2702# a_30652_2702# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8919 a_30650_5457# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8920 a_646_4368# a_433_4368# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8921 a_11824_4683# a_11757_4091# a_11841_3120# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8922 a_1792_6884# a_1371_6884# a_854_7128# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8923 a_29062_n7359# a_29319_n7375# a_28124_n7603# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8924 a_35390_7265# a_35919_7155# a_36127_7155# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8925 vdd a_34294_n7339# a_34086_n7339# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8926 a_1724_n9198# a_1511_n9198# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8927 a_30651_2148# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8928 a_21556_n9771# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8929 a_15523_1659# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8930 a_28128_n7415# a_29112_n7929# a_29063_n7913# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8931 a_10680_1618# a_10467_1618# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8932 a_12918_4680# a_13902_4977# a_13853_5167# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8933 a_5176_n1804# a_4799_n1525# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8934 a_10887_n1764# a_10466_n1764# a_10151_n1768# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8935 gnd a_39353_2793# a_39145_2793# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8936 a_31942_n6978# a_31729_n6978# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8937 a_3823_n4582# a_4080_n4598# a_2888_n4084# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8938 a_24012_n3821# a_24008_n4009# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8939 vdd a_38274_n2701# a_38066_n2701# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8940 vdd a_8054_8604# a_7846_8604# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8941 vdd a_19166_n5747# a_18958_n5747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8942 a_31071_8217# a_31801_7973# a_32009_7973# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8943 a_16989_5254# a_16568_5254# a_16890_5254# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8944 a_8883_n3332# a_9136_n3536# a_7944_n3022# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8945 a_25360_5928# a_25360_5698# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8946 a_10147_n10135# a_14108_n10118# a_12916_n9604# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8947 a_37846_n10683# a_38096_n5991# a_38051_n5787# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8948 vdd d2 a_3000_n4880# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8949 a_34037_9560# a_34294_9370# a_33102_9073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8950 a_11757_n4791# a_11544_n4791# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8951 a_32960_n4850# a_33150_n4274# a_33101_n4258# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8952 a_21880_n8089# a_21667_n8089# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8953 a_855_n5622# a_434_n5622# a_118_n5531# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8954 a_7060_541# a_6951_541# a_4954_480# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8955 a_10887_1064# a_11618_1374# a_11826_1374# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8956 a_20305_n4409# a_20305_n4180# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8957 a_10885_5476# a_10464_5476# a_10149_5224# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8958 a_12809_n5765# a_13062_n5969# a_12604_n10661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8959 a_22934_n2451# a_23119_n3166# a_23070_n3150# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8960 gnd d0 a_39352_3342# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8961 a_27034_6906# a_26967_6314# a_27045_7430# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8962 a_39095_n5712# a_39352_n5728# a_38160_n5214# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8963 a_38157_n3196# a_39144_n2968# a_39099_n2764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8964 vdd a_29320_7200# a_29112_7200# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8965 a_1902_5208# a_1481_5208# a_1803_5208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8966 a_1803_n5731# a_1483_n3696# a_1805_n3519# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8967 a_33102_1529# a_33359_1339# a_32961_2121# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8968 a_5176_1951# a_5176_1764# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8969 gnd a_19166_n4090# a_18958_n4090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8970 a_25888_8253# a_25675_8253# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8971 a_27988_6392# a_28173_6890# a_28124_7080# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8972 a_32025_7513# a_31728_8484# a_32008_9076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8973 vdd d0 a_39352_n6831# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8974 a_22964_5229# a_23007_7428# a_22958_7618# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8975 a_5488_n7315# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8976 vdd d4 a_33248_n5950# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8977 vdd a_8087_n6005# a_7879_n6005# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8978 a_25358_n9965# a_25358_n9736# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8979 a_11404_2477# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8980 vdd a_3029_n8176# a_2821_n8176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8981 gnd d0 a_39349_n9586# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8982 a_30335_n5058# a_30863_n5054# a_31071_n5054# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8983 a_18910_n3525# a_18913_n2783# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8984 a_36858_5808# a_36645_5808# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8985 a_38156_4879# a_39143_4445# a_39094_4635# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8986 a_35706_n5095# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8987 a_15941_8277# a_15520_8277# a_15204_8158# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8988 gnd d0 a_29320_8303# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8989 vdd a_9135_n2982# a_8927_n2982# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8990 a_16601_n2626# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8991 a_16671_6930# a_16458_6930# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8992 a_26938_n3718# a_26725_n3718# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8993 a_35390_n7305# a_35391_n6848# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8994 a_647_n6725# a_434_n6725# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X8995 a_35707_n5649# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8996 a_20619_8212# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8997 a_8882_n2778# a_8878_n2966# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X8998 a_32011_n3158# a_31590_n3158# a_31073_n3402# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8999 a_22088_5189# a_21667_5189# a_21989_5189# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9000 a_2886_6881# a_3139_6868# a_2746_6370# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9001 a_647_3265# a_434_3265# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9002 a_6850_n4316# a_6429_n4316# a_5912_n4560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9003 a_28130_n4106# a_28383_n4310# a_27985_n4886# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9004 a_35391_5933# a_35920_6052# a_36128_6052# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9005 a_26614_4700# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9006 a_28127_9109# a_29111_9406# a_29062_9596# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9007 a_30652_1045# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9008 gnd a_24264_8262# a_24056_8262# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9009 a_21769_9071# a_21556_9071# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9010 a_32020_7394# a_31729_6278# a_32009_6870# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9011 vdd d3 a_28271_n8198# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9012 a_16895_5373# a_16568_7454# a_16895_7573# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9013 a_11839_n8113# a_11725_n8113# a_11839_n5913# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9014 vdd d0 a_39350_7754# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9015 a_38160_5805# a_38413_5792# a_38015_6574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9016 a_8878_n6829# a_8881_n6087# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9017 a_13855_6642# a_14108_6629# a_12913_7063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9018 gnd a_10033_n10854# a_9825_n10854# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9019 gnd d5 a_28072_n10694# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9020 a_27035_n5400# a_26968_n4808# a_27052_n3718# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9021 a_10884_n8382# a_10463_n8382# a_10148_n8386# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9022 vdd a_23324_9055# a_23116_9055# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9023 a_32119_n5894# a_33047_n10658# a_32889_n10642# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9024 gnd d4 a_23217_5216# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9025 a_33105_n2967# a_34089_n3481# a_34044_n3277# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9026 a_11822_9095# a_11401_9095# a_10883_8785# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9027 vdd a_23186_n4861# a_22978_n4861# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9028 a_1808_5327# a_1481_7408# a_1808_7527# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9029 vdd a_8056_4192# a_7848_4192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9030 a_26098_2738# a_26828_2494# a_27036_2494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9031 a_18908_5757# a_19165_5567# a_17970_6001# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9032 a_31073_3805# a_31803_3561# a_32011_3561# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9033 a_15942_n5668# a_16672_n5424# a_16880_n5424# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9034 a_27047_n3541# a_26756_n2602# a_27036_n3194# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9035 vdd a_14111_n1843# a_13903_n1843# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9036 a_36860_1396# a_36647_1396# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9037 a_10887_1064# a_10466_1064# a_10153_1170# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9038 a_24007_n7872# a_24264_n7888# a_23072_n7374# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9039 a_39098_n7730# a_39351_n7934# a_38159_n7420# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9040 a_35392_n3539# a_35920_n3992# a_36128_n3992# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9041 a_17091_546# a_17910_5281# a_17861_5471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9042 a_38154_n9814# a_39141_n9586# a_39096_n9382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9043 a_13852_n7896# a_13855_n7154# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9044 a_24008_3486# a_24265_3296# a_23070_3730# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9045 a_29062_n8462# a_29067_n7725# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9046 a_5910_n8972# a_5489_n8972# a_5173_n8881# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9047 vdd a_4080_n3495# a_3872_n3495# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9048 a_31588_n7570# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9049 vdd d0 a_24264_n8991# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9050 a_32993_7446# a_33246_7433# a_32995_5234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9051 a_22960_5406# a_23009_3016# a_22960_3206# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9052 a_27246_522# a_28065_5257# a_28020_5270# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9053 vdd a_18227_n6540# a_18019_n6540# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9054 a_17865_5294# a_17908_7493# a_17863_7506# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9055 a_1694_n8108# a_1481_n8108# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9056 a_31591_1355# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9057 a_26097_n5644# a_25676_n5644# a_25360_n5324# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9058 gnd d0 a_29322_3891# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9059 gnd a_34298_n2378# a_34090_n2378# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9060 a_5910_5512# a_5489_5512# a_5174_5260# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9061 vdd a_9132_n9600# a_8924_n9600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9062 a_23071_n2047# a_23328_n2063# a_22930_n2639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9063 a_30335_n5517# a_30864_n5608# a_31072_n5608# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9064 a_38156_n6505# a_38413_n6521# a_38015_n7097# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9065 a_22088_n5889# a_21667_n5889# a_21994_n5889# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9066 a_20619_n7809# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9067 gnd d1 a_23325_6849# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9068 a_31069_n9466# a_30648_n9466# a_30333_n9470# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9069 a_10675_8785# a_10462_8785# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9070 a_29068_n3862# a_29064_n4050# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9071 a_3827_2779# a_4080_2766# a_2888_2469# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9072 a_32025_5313# a_31911_5194# a_32119_5194# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9073 vdd d2 a_38273_n4907# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9074 a_26924_522# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9075 a_31073_n3402# a_30652_n3402# a_30336_n3311# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9076 a_35704_8807# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9077 a_26095_7699# a_26826_8009# a_27034_8009# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9078 a_19119_n829# d9 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9079 a_24009_1280# a_20308_1146# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9080 a_24013_3863# a_24009_4040# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9081 vdd d1 a_8197_3600# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9082 a_28129_4697# a_29113_4994# a_29064_5184# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9083 a_35390_n8867# a_35390_n8638# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9084 gnd a_24266_3850# a_24058_3850# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9085 a_7945_n1919# a_8929_n2433# a_8884_n2229# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9086 a_2887_n5187# a_3140_n5391# a_2747_n4676# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9087 a_38162_1393# a_38415_1380# a_38017_2162# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9088 vdd d0 a_39352_3342# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9089 a_5175_n4240# a_5704_n4560# a_5912_n4560# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9090 a_39099_n5524# a_39095_n5712# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9091 a_26096_5493# a_25675_5493# a_25360_5241# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9092 a_24010_6618# a_24006_6795# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9093 a_433_n7828# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9094 a_30335_n6807# a_30335_n6620# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9095 a_1902_n5908# a_1481_n5908# a_1803_n5731# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9096 a_1803_5208# a_1483_2996# a_1810_3115# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9097 gnd d1 a_3140_n6494# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9098 a_20305_4097# a_20832_4349# a_21040_4349# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9099 a_21980_2453# a_21913_1861# a_21991_2977# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9100 a_15943_n1805# a_15522_n1805# a_14830_n1530# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9101 vdd a_14108_n8461# a_13900_n8461# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9102 a_15204_n9073# a_15204_n8886# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9103 a_30335_6308# a_30335_6121# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9104 a_38159_n8523# a_39143_n9037# a_39098_n8833# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9105 a_20533_n10895# a_30011_n10835# a_24964_n10698# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9106 a_38156_4879# a_39143_4445# a_39098_4458# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9107 a_12779_n2475# a_12964_n3190# a_12915_n3174# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9108 a_15944_n2359# a_15523_n2359# a_15207_n2268# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9109 a_3823_1299# a_4080_1109# a_2885_1543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9110 a_16813_n4832# a_16600_n4832# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9111 a_18913_5031# a_19166_5018# a_17974_4721# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9112 a_35919_n7855# a_35706_n7855# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9113 a_3825_n8806# a_3821_n8994# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9114 a_3826_6088# a_4079_6075# a_2887_5778# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9115 a_28131_n1900# a_29115_n2414# a_29070_n2210# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9116 a_21880_5189# a_21667_5189# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9117 a_3820_n7337# a_4077_n7353# a_2882_n7581# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9118 a_37068_n2096# a_37000_n2607# a_37078_n3546# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9119 a_32995_3034# a_33248_3021# a_32991_5411# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9120 a_20834_2697# a_20621_2697# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9121 vdd a_9134_n9051# a_8926_n9051# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9122 a_15205_5722# a_15733_5517# a_15941_5517# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9123 a_18910_n9401# a_19163_n9605# a_17968_n9833# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9124 a_32889_n10642# a_35153_n10719# a_29962_n10819# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9125 a_5912_1100# a_5491_1100# a_5178_1206# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9126 vdd a_24264_8262# a_24056_8262# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9127 vdd d2 a_18086_n7132# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9128 a_7830_n5989# a_7879_n3805# a_7830_n3789# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9129 a_38020_4191# a_38273_4178# a_38051_3075# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9130 a_23068_n8665# a_23325_n8681# a_22927_n9257# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9131 vdd a_14110_n5706# a_13902_n5706# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9132 gnd d2 a_8054_n9333# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9133 a_21700_n2561# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9134 vdd d0 a_9134_7219# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9135 a_21039_6555# a_20618_6555# a_20303_6760# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9136 a_35705_7704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9137 a_6537_7449# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9138 vdd d4 a_23217_5216# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9139 a_36130_1640# a_35709_1640# a_35393_1521# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9140 a_21994_n8089# a_21697_n9179# a_21978_n8668# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9141 a_11404_n3177# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9142 a_36646_n3199# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9143 a_17973_6927# a_18957_7224# a_18908_7414# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9144 gnd d0 a_14109_4423# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9145 a_1585_n5378# a_1372_n5378# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9146 a_29068_3350# a_29321_3337# a_28126_3771# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9147 a_35390_8368# a_35390_8139# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9148 a_17091_546# a_17910_5281# a_17865_5294# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9149 a_11825_n4280# a_11404_n4280# a_10887_n4524# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9150 a_6850_3616# a_6429_3616# a_5911_3306# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9151 a_37175_5235# a_37168_527# a_35171_466# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9152 a_26098_1081# a_25677_1081# a_25364_1187# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9153 a_28016_n5970# a_28065_n3786# a_28016_n3770# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9154 a_5175_3741# a_5704_3860# a_5912_3860# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9155 a_32989_7623# a_33246_7433# a_32995_5234# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9156 a_25674_9356# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9157 a_16600_4132# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9158 a_25359_n7530# a_25888_n7850# a_26096_n7850# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9159 vdd d1 a_18226_n8746# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9160 a_15940_n8423# a_15519_n8423# a_15204_n7970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9161 a_22960_5406# a_23009_3016# a_22964_3029# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9162 a_32989_n8146# a_33008_n7072# a_32959_n7056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9163 a_6641_4719# a_6428_4719# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9164 a_15205_n6451# a_15734_n6771# a_15942_n6771# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9165 a_20305_2348# a_20306_1891# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9166 a_8883_n1675# a_9136_n1879# a_7941_n2107# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9167 gnd d0 a_24265_6056# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9168 a_10150_3934# a_10679_3824# a_10887_3824# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9169 a_20833_n3946# a_20620_n3946# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9170 a_17828_8799# a_18018_8017# a_17969_8207# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9171 gnd a_14109_7183# a_13901_7183# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9172 gnd d1 a_23324_n9784# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9173 a_2887_n5187# a_3871_n5701# a_3822_n5685# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9174 a_34040_n4568# a_34043_n3826# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9175 vdd a_19164_n10159# a_18956_n10159# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9176 a_15733_n6217# a_15520_n6217# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9177 a_852_n9480# a_1583_n9790# a_1791_n9790# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9178 a_27035_n6503# a_26614_n6503# a_26097_n6747# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9179 gnd d3 a_23217_n3745# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9180 gnd d3 a_38302_n8203# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9181 a_37065_n8714# a_36997_n9225# a_37081_n8135# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9182 a_20834_n4500# a_20621_n4500# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9183 a_3823_2956# a_4080_2766# a_2888_2469# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9184 a_647_4922# a_434_4922# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9185 a_432_7677# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9186 a_10148_7014# a_10677_7133# a_10885_7133# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9187 a_11512_n8113# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9188 gnd a_2999_n7086# a_2791_n7086# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9189 a_23072_6862# a_24056_7159# a_24007_7349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9190 a_26755_n4808# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9191 a_30652_2702# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9192 vdd a_13169_9079# a_12961_9079# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9193 a_433_4368# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9194 a_29064_n5707# a_29067_n4965# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9195 gnd a_33217_n4866# a_33009_n4866# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9196 a_12776_8581# a_12961_9079# a_12912_9269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9197 a_15942_n5668# a_15521_n5668# a_15205_n5348# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9198 a_30863_n5054# a_30650_n5054# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9199 a_15734_n2908# a_15521_n2908# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9200 a_28130_2491# a_28383_2478# a_27990_1980# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9201 a_33105_3558# a_33358_3545# a_32960_4327# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9202 a_20302_n9465# a_20303_n9008# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9203 a_38158_1570# a_38415_1380# a_38017_2162# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X9204 a_16459_n5424# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9205 a_5912_2757# a_5491_2757# a_5175_2638# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9206 a_8877_n6275# a_8882_n5538# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X9207 a_35707_3292# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
C0 a_5053_480# a_4954_480# 3.47fF
C1 a_16989_5254# a_17091_546# 8.08fF
C2 a_22088_5189# a_22190_481# 8.08fF
C3 a_6958_5249# a_7060_541# 8.08fF
C4 a_6958_n5949# a_7629_n10697# 8.08fF
C5 a_32119_5194# a_32221_486# 8.08fF
C6 vdd d3 2.11fF
C7 a_12703_n10661# a_9776_n10838# 3.47fF
C8 a_11933_n5913# a_12604_n10661# 8.08fF
C9 a_1902_n5908# a_2573_n10656# 8.08fF
C10 a_1902_5208# a_2004_500# 8.08fF
C11 a_11933_5213# a_12035_505# 8.08fF
C12 a_25239_461# a_25140_461# 3.47fF
C13 a_22088_n5889# a_22759_n10637# 8.08fF
C14 a_27144_5230# a_27246_522# 8.08fF
C15 a_16989_n5954# a_17660_n10702# 8.08fF
C16 vdd d0 16.89fF
C17 a_27144_n5930# a_27815_n10678# 8.08fF
C18 a_37175_5235# a_37277_527# 8.08fF
C19 vdd d1 8.45fF
C20 a_37175_n5935# a_37846_n10683# 8.08fF
C21 a_32889_n10642# a_29962_n10819# 3.47fF
C22 a_32119_n5894# a_32790_n10642# 8.08fF
C23 vdd d2 4.22fF
C24 a_20533_n10895# gnd 11.31fF
C25 a_34896_n10703# gnd 4.59fF
C26 a_29962_n10819# gnd 7.14fF
C27 d6 gnd 2.63fF
C28 d5 gnd 5.25fF
C29 a_32889_n10642# gnd 3.40fF
C30 a_24865_n10698# gnd 4.59fF
C31 a_24964_n10698# gnd 6.50fF
C32 a_9875_n10838# gnd 11.66fF
C33 a_22858_n10637# gnd 3.40fF
C34 a_14710_n10722# gnd 4.59fF
C35 a_9776_n10838# gnd 7.14fF
C36 a_12703_n10661# gnd 3.40fF
C37 a_4679_n10717# gnd 4.59fF
C38 a_4778_n10717# gnd 6.50fF
C39 a_2672_n10656# gnd 3.40fF
C40 a_35389_n10157# gnd 6.43fF
C41 d0 gnd 191.06fF
C42 a_35389_n9970# gnd 2.22fF
C43 a_30333_n10116# gnd 6.43fF
C44 a_39093_n10124# gnd 2.23fF
C45 a_25358_n10152# gnd 6.43fF
C46 a_30333_n9929# gnd 2.22fF
C47 a_25358_n9965# gnd 2.22fF
C48 a_20302_n10111# gnd 6.43fF
C49 a_35389_n9741# gnd 2.38fF
C50 a_34037_n10083# gnd 2.23fF
C51 a_38158_n9626# gnd 2.52fF
C52 a_36126_n10061# gnd 2.38fF
C53 a_29062_n10119# gnd 2.23fF
C54 a_30333_n9700# gnd 2.38fF
C55 d1 gnd 99.71fF
C56 a_15203_n10176# gnd 6.43fF
C57 a_15203_n9989# gnd 2.22fF
C58 a_10147_n10135# gnd 6.43fF
C59 a_20302_n9924# gnd 2.22fF
C60 a_18907_n10143# gnd 2.23fF
C61 a_25358_n9736# gnd 2.38fF
C62 a_33102_n9585# gnd 2.52fF
C63 a_31070_n10020# gnd 2.38fF
C64 a_24006_n10078# gnd 2.23fF
C65 a_28127_n9621# gnd 2.52fF
C66 a_26095_n10056# gnd 2.38fF
C67 a_20302_n9695# gnd 2.38fF
C68 a_5172_n10171# gnd 6.43fF
C69 a_10147_n9948# gnd 2.22fF
C70 a_5172_n9984# gnd 2.22fF
C71 a_116_n10130# gnd 6.43fF
C72 a_15203_n9760# gnd 2.38fF
C73 a_39092_n9570# gnd 2.28fF
C74 a_38154_n9814# gnd 2.18fF
C75 a_39096_n9382# gnd 2.38fF
C76 a_35389_n9511# gnd 2.23fF
C77 a_36125_n9507# gnd 2.52fF
C78 a_34036_n9529# gnd 2.28fF
C79 a_33098_n9773# gnd 2.18fF
C80 a_13851_n10102# gnd 2.23fF
C81 a_17972_n9645# gnd 2.52fF
C82 a_15940_n10080# gnd 2.38fF
C83 a_8876_n10138# gnd 2.23fF
C84 a_10147_n9719# gnd 2.38fF
C85 a_23071_n9580# gnd 2.52fF
C86 a_21039_n10015# gnd 2.38fF
C87 a_34040_n9341# gnd 2.38fF
C88 a_29061_n9565# gnd 2.28fF
C89 a_28123_n9809# gnd 2.18fF
C90 a_29065_n9377# gnd 2.38fF
C91 a_30333_n9470# gnd 2.23fF
C92 a_31069_n9466# gnd 2.52fF
C93 a_25358_n9506# gnd 2.23fF
C94 a_26094_n9502# gnd 2.52fF
C95 a_24005_n9524# gnd 2.28fF
C96 a_23067_n9768# gnd 2.18fF
C97 a_116_n9943# gnd 2.22fF
C98 a_5172_n9755# gnd 2.38fF
C99 a_12916_n9604# gnd 2.52fF
C100 a_10884_n10039# gnd 2.38fF
C101 a_3820_n10097# gnd 2.23fF
C102 a_7941_n9640# gnd 2.52fF
C103 a_5909_n10075# gnd 2.38fF
C104 a_116_n9714# gnd 2.38fF
C105 a_24009_n9336# gnd 2.38fF
C106 d2 gnd 50.39fF
C107 a_35390_n9054# gnd 2.49fF
C108 a_18906_n9589# gnd 2.28fF
C109 a_17968_n9833# gnd 2.18fF
C110 a_18910_n9401# gnd 2.38fF
C111 a_20302_n9465# gnd 2.23fF
C112 a_21038_n9461# gnd 2.52fF
C113 a_15203_n9530# gnd 2.23fF
C114 a_15939_n9526# gnd 2.52fF
C115 a_13850_n9548# gnd 2.28fF
C116 a_12912_n9792# gnd 2.18fF
C117 a_2885_n9599# gnd 2.52fF
C118 a_853_n10034# gnd 2.38fF
C119 a_13854_n9360# gnd 2.38fF
C120 a_8875_n9584# gnd 2.28fF
C121 a_7937_n9828# gnd 2.18fF
C122 a_8879_n9396# gnd 2.38fF
C123 a_30334_n9013# gnd 2.49fF
C124 a_25359_n9049# gnd 2.49fF
C125 a_10147_n9489# gnd 2.23fF
C126 a_10883_n9485# gnd 2.52fF
C127 a_5172_n9525# gnd 2.23fF
C128 a_5908_n9521# gnd 2.52fF
C129 a_3819_n9543# gnd 2.28fF
C130 a_2881_n9787# gnd 2.18fF
C131 a_3823_n9355# gnd 2.38fF
C132 a_39098_n8833# gnd 2.49fF
C133 a_35390_n8867# gnd 2.28fF
C134 a_34042_n8792# gnd 2.49fF
C135 a_39094_n9021# gnd 2.23fF
C136 a_20303_n9008# gnd 2.49fF
C137 a_15204_n9073# gnd 2.49fF
C138 a_29067_n8828# gnd 2.49fF
C139 a_30334_n8826# gnd 2.28fF
C140 a_25359_n8862# gnd 2.28fF
C141 a_116_n9484# gnd 2.23fF
C142 a_852_n9480# gnd 2.52fF
C143 a_24011_n8787# gnd 2.49fF
C144 a_35390_n8638# gnd 2.38fF
C145 a_34038_n8980# gnd 2.23fF
C146 a_38159_n8523# gnd 2.52fF
C147 a_36127_n8958# gnd 2.18fF
C148 a_29063_n9016# gnd 2.23fF
C149 a_30334_n8597# gnd 2.38fF
C150 a_10148_n9032# gnd 2.49fF
C151 a_5173_n9068# gnd 2.49fF
C152 a_18912_n8852# gnd 2.49fF
C153 a_15204_n8886# gnd 2.28fF
C154 a_13856_n8811# gnd 2.49fF
C155 a_20303_n8821# gnd 2.28fF
C156 a_18908_n9040# gnd 2.23fF
C157 a_25359_n8633# gnd 2.38fF
C158 a_33103_n8482# gnd 2.52fF
C159 a_31071_n8917# gnd 2.18fF
C160 a_24007_n8975# gnd 2.23fF
C161 a_28128_n8518# gnd 2.52fF
C162 a_26096_n8953# gnd 2.18fF
C163 a_20303_n8592# gnd 2.38fF
C164 a_117_n9027# gnd 2.49fF
C165 a_8881_n8847# gnd 2.49fF
C166 a_10148_n8845# gnd 2.28fF
C167 a_5173_n8881# gnd 2.28fF
C168 a_3825_n8806# gnd 2.49fF
C169 a_15204_n8657# gnd 2.38fF
C170 a_39093_n8467# gnd 2.28fF
C171 a_38155_n8711# gnd 2.45fF
C172 a_39097_n8279# gnd 2.38fF
C173 a_35390_n8408# gnd 2.23fF
C174 a_36126_n8404# gnd 2.52fF
C175 a_34037_n8426# gnd 2.28fF
C176 a_33099_n8670# gnd 2.45fF
C177 a_13852_n8999# gnd 2.23fF
C178 a_17973_n8542# gnd 2.52fF
C179 a_15941_n8977# gnd 2.18fF
C180 a_8877_n9035# gnd 2.23fF
C181 a_10148_n8616# gnd 2.38fF
C182 a_23072_n8477# gnd 2.52fF
C183 a_21040_n8912# gnd 2.18fF
C184 a_34041_n8238# gnd 2.38fF
C185 a_29062_n8462# gnd 2.28fF
C186 a_28124_n8706# gnd 2.45fF
C187 a_29066_n8274# gnd 2.38fF
C188 a_30334_n8367# gnd 2.23fF
C189 a_31070_n8363# gnd 2.52fF
C190 a_25359_n8403# gnd 2.23fF
C191 a_26095_n8399# gnd 2.52fF
C192 a_24006_n8421# gnd 2.28fF
C193 a_23068_n8665# gnd 2.45fF
C194 a_117_n8840# gnd 2.28fF
C195 a_5173_n8652# gnd 2.38fF
C196 a_12917_n8501# gnd 2.52fF
C197 a_10885_n8936# gnd 2.18fF
C198 a_3821_n8994# gnd 2.23fF
C199 a_7942_n8537# gnd 2.52fF
C200 a_5910_n8972# gnd 2.18fF
C201 a_117_n8611# gnd 2.38fF
C202 a_24010_n8233# gnd 2.38fF
C203 a_18907_n8486# gnd 2.28fF
C204 a_17969_n8730# gnd 2.45fF
C205 a_18911_n8298# gnd 2.38fF
C206 a_38049_n7999# gnd 2.28fF
C207 d3 gnd 22.51fF
C208 a_37081_n8135# gnd 2.04fF
C209 a_35390_n7951# gnd 2.49fF
C210 a_32993_n7958# gnd 2.28fF
C211 a_20303_n8362# gnd 2.23fF
C212 a_21039_n8358# gnd 2.52fF
C213 a_15204_n8427# gnd 2.23fF
C214 a_15940_n8423# gnd 2.52fF
C215 a_13851_n8445# gnd 2.28fF
C216 a_12913_n8689# gnd 2.45fF
C217 a_2886_n8496# gnd 2.52fF
C218 a_854_n8931# gnd 2.18fF
C219 a_13855_n8257# gnd 2.38fF
C220 a_8876_n8481# gnd 2.28fF
C221 a_7938_n8725# gnd 2.45fF
C222 a_8880_n8293# gnd 2.38fF
C223 a_28018_n7994# gnd 2.28fF
C224 a_32025_n8094# gnd 2.04fF
C225 a_30334_n7910# gnd 2.49fF
C226 a_27050_n8130# gnd 2.04fF
C227 a_25359_n7946# gnd 2.49fF
C228 a_22962_n7953# gnd 2.28fF
C229 a_10148_n8386# gnd 2.23fF
C230 a_10884_n8382# gnd 2.52fF
C231 a_5173_n8422# gnd 2.23fF
C232 a_5909_n8418# gnd 2.52fF
C233 a_3820_n8440# gnd 2.28fF
C234 a_2882_n8684# gnd 2.45fF
C235 a_3824_n8252# gnd 2.38fF
C236 a_17863_n8018# gnd 2.28fF
C237 a_39098_n7730# gnd 2.49fF
C238 a_35390_n7764# gnd 2.28fF
C239 a_34042_n7689# gnd 2.49fF
C240 a_39094_n7918# gnd 2.23fF
C241 a_21994_n8089# gnd 2.04fF
C242 a_20303_n7905# gnd 2.49fF
C243 a_16895_n8154# gnd 2.04fF
C244 a_15204_n7970# gnd 2.49fF
C245 a_12807_n7977# gnd 2.28fF
C246 a_117_n8381# gnd 2.23fF
C247 a_853_n8377# gnd 2.52fF
C248 a_7832_n8013# gnd 2.28fF
C249 a_29067_n7725# gnd 2.49fF
C250 a_30334_n7723# gnd 2.28fF
C251 a_25359_n7759# gnd 2.28fF
C252 a_24011_n7684# gnd 2.49fF
C253 a_35390_n7535# gnd 2.38fF
C254 a_34038_n7877# gnd 2.23fF
C255 a_38159_n7420# gnd 2.52fF
C256 a_36127_n7855# gnd 2.45fF
C257 a_29063_n7913# gnd 2.23fF
C258 a_30334_n7494# gnd 2.38fF
C259 a_11839_n8113# gnd 2.04fF
C260 a_10148_n7929# gnd 2.49fF
C261 a_6864_n8149# gnd 2.04fF
C262 a_5173_n7965# gnd 2.49fF
C263 a_2776_n7972# gnd 2.28fF
C264 a_18912_n7749# gnd 2.49fF
C265 a_15204_n7783# gnd 2.28fF
C266 a_13856_n7708# gnd 2.49fF
C267 a_20303_n7718# gnd 2.28fF
C268 a_18908_n7937# gnd 2.23fF
C269 a_25359_n7530# gnd 2.38fF
C270 a_33103_n7379# gnd 2.52fF
C271 a_31071_n7814# gnd 2.45fF
C272 a_24007_n7872# gnd 2.23fF
C273 a_28128_n7415# gnd 2.52fF
C274 a_26096_n7850# gnd 2.45fF
C275 a_20303_n7489# gnd 2.38fF
C276 a_1808_n8108# gnd 2.04fF
C277 a_117_n7924# gnd 2.49fF
C278 a_8881_n7744# gnd 2.49fF
C279 a_10148_n7742# gnd 2.28fF
C280 a_5173_n7778# gnd 2.28fF
C281 a_3825_n7703# gnd 2.49fF
C282 a_15204_n7554# gnd 2.38fF
C283 a_39093_n7364# gnd 2.28fF
C284 a_38155_n7608# gnd 2.18fF
C285 a_39097_n7176# gnd 2.38fF
C286 a_35390_n7305# gnd 2.23fF
C287 a_36126_n7301# gnd 2.52fF
C288 a_34037_n7323# gnd 2.28fF
C289 a_33099_n7567# gnd 2.18fF
C290 a_13852_n7896# gnd 2.23fF
C291 a_17973_n7439# gnd 2.52fF
C292 a_15941_n7874# gnd 2.45fF
C293 a_8877_n7932# gnd 2.23fF
C294 a_10148_n7513# gnd 2.38fF
C295 a_23072_n7374# gnd 2.52fF
C296 a_21040_n7809# gnd 2.45fF
C297 a_34041_n7135# gnd 2.38fF
C298 a_29062_n7359# gnd 2.28fF
C299 a_28124_n7603# gnd 2.18fF
C300 a_29066_n7171# gnd 2.38fF
C301 a_38045_n8187# gnd 2.45fF
C302 a_30334_n7264# gnd 2.23fF
C303 a_31070_n7260# gnd 2.52fF
C304 a_25359_n7300# gnd 2.23fF
C305 a_26095_n7296# gnd 2.52fF
C306 a_24006_n7318# gnd 2.28fF
C307 a_23068_n7562# gnd 2.18fF
C308 a_117_n7737# gnd 2.28fF
C309 a_5173_n7549# gnd 2.38fF
C310 a_12917_n7398# gnd 2.52fF
C311 a_10885_n7833# gnd 2.45fF
C312 a_3821_n7891# gnd 2.23fF
C313 a_7942_n7434# gnd 2.52fF
C314 a_5910_n7869# gnd 2.45fF
C315 a_117_n7508# gnd 2.38fF
C316 a_24010_n7130# gnd 2.38fF
C317 a_37076_n7958# gnd 2.34fF
C318 a_35391_n6848# gnd 2.49fF
C319 a_32989_n8146# gnd 2.45fF
C320 a_18907_n7383# gnd 2.28fF
C321 a_17969_n7627# gnd 2.18fF
C322 a_18911_n7195# gnd 2.38fF
C323 a_28014_n8182# gnd 2.45fF
C324 a_20303_n7259# gnd 2.23fF
C325 a_21039_n7255# gnd 2.52fF
C326 a_15204_n7324# gnd 2.23fF
C327 a_15940_n7320# gnd 2.52fF
C328 a_13851_n7342# gnd 2.28fF
C329 a_12913_n7586# gnd 2.18fF
C330 a_2886_n7393# gnd 2.52fF
C331 a_854_n7828# gnd 2.45fF
C332 a_13855_n7154# gnd 2.38fF
C333 a_8876_n7378# gnd 2.28fF
C334 a_7938_n7622# gnd 2.18fF
C335 a_8880_n7190# gnd 2.38fF
C336 a_32020_n7917# gnd 2.34fF
C337 a_30335_n6807# gnd 2.49fF
C338 a_27045_n7953# gnd 2.34fF
C339 a_25360_n6843# gnd 2.49fF
C340 a_22958_n8141# gnd 2.45fF
C341 a_17859_n8206# gnd 2.45fF
C342 a_10148_n7283# gnd 2.23fF
C343 a_10884_n7279# gnd 2.52fF
C344 a_5173_n7319# gnd 2.23fF
C345 a_5909_n7315# gnd 2.52fF
C346 a_3820_n7337# gnd 2.28fF
C347 a_2882_n7581# gnd 2.18fF
C348 a_3824_n7149# gnd 2.38fF
C349 a_39099_n6627# gnd 2.49fF
C350 a_35391_n6661# gnd 2.28fF
C351 a_34043_n6586# gnd 2.49fF
C352 a_39095_n6815# gnd 2.23fF
C353 a_21989_n7912# gnd 2.34fF
C354 a_20304_n6802# gnd 2.49fF
C355 a_16890_n7977# gnd 2.34fF
C356 a_15205_n6867# gnd 2.49fF
C357 a_12803_n8165# gnd 2.45fF
C358 a_29068_n6622# gnd 2.49fF
C359 a_30335_n6620# gnd 2.28fF
C360 a_25360_n6656# gnd 2.28fF
C361 a_7828_n8201# gnd 2.45fF
C362 a_117_n7278# gnd 2.23fF
C363 a_853_n7274# gnd 2.52fF
C364 a_24012_n6581# gnd 2.49fF
C365 a_35391_n6432# gnd 2.38fF
C366 a_34039_n6774# gnd 2.23fF
C367 a_38160_n6317# gnd 2.52fF
C368 a_36128_n6752# gnd 2.18fF
C369 a_29064_n6810# gnd 2.23fF
C370 a_30335_n6391# gnd 2.38fF
C371 a_11834_n7936# gnd 2.34fF
C372 a_10149_n6826# gnd 2.49fF
C373 a_6859_n7972# gnd 2.34fF
C374 a_5174_n6862# gnd 2.49fF
C375 a_2772_n8160# gnd 2.45fF
C376 a_18913_n6646# gnd 2.49fF
C377 a_15205_n6680# gnd 2.28fF
C378 a_13857_n6605# gnd 2.49fF
C379 a_20304_n6615# gnd 2.28fF
C380 a_18909_n6834# gnd 2.23fF
C381 a_25360_n6427# gnd 2.38fF
C382 a_33104_n6276# gnd 2.52fF
C383 a_31072_n6711# gnd 2.18fF
C384 a_24008_n6769# gnd 2.23fF
C385 a_28129_n6312# gnd 2.52fF
C386 a_26097_n6747# gnd 2.18fF
C387 a_20304_n6386# gnd 2.38fF
C388 a_1803_n7931# gnd 2.34fF
C389 a_118_n6821# gnd 2.49fF
C390 a_8882_n6641# gnd 2.49fF
C391 a_10149_n6639# gnd 2.28fF
C392 a_5174_n6675# gnd 2.28fF
C393 a_3826_n6600# gnd 2.49fF
C394 a_15205_n6451# gnd 2.38fF
C395 a_39094_n6261# gnd 2.28fF
C396 a_38156_n6505# gnd 2.45fF
C397 a_39098_n6073# gnd 2.38fF
C398 a_35391_n6202# gnd 2.23fF
C399 a_36127_n6198# gnd 2.52fF
C400 a_34038_n6220# gnd 2.28fF
C401 a_33100_n6464# gnd 2.45fF
C402 a_13853_n6793# gnd 2.23fF
C403 a_17974_n6336# gnd 2.52fF
C404 a_15942_n6771# gnd 2.18fF
C405 a_8878_n6829# gnd 2.23fF
C406 a_10149_n6410# gnd 2.38fF
C407 a_23073_n6271# gnd 2.52fF
C408 a_21041_n6706# gnd 2.18fF
C409 a_34042_n6032# gnd 2.38fF
C410 a_37846_n10683# gnd 5.48fF
C411 a_29063_n6256# gnd 2.28fF
C412 a_28125_n6500# gnd 2.45fF
C413 a_29067_n6068# gnd 2.38fF
C414 a_30335_n6161# gnd 2.23fF
C415 a_31071_n6157# gnd 2.52fF
C416 a_25360_n6197# gnd 2.23fF
C417 a_26096_n6193# gnd 2.52fF
C418 a_24007_n6215# gnd 2.28fF
C419 a_23069_n6459# gnd 2.45fF
C420 a_118_n6634# gnd 2.28fF
C421 a_5174_n6446# gnd 2.38fF
C422 a_12918_n6295# gnd 2.52fF
C423 a_10886_n6730# gnd 2.18fF
C424 a_3822_n6788# gnd 2.23fF
C425 a_7943_n6331# gnd 2.52fF
C426 a_5911_n6766# gnd 2.18fF
C427 a_118_n6405# gnd 2.38fF
C428 a_24011_n6027# gnd 2.38fF
C429 a_38051_n5787# gnd 3.68fF
C430 d4 gnd 11.80fF
C431 a_37081_n5935# gnd 3.32fF
C432 a_37175_n5935# gnd 6.48fF
C433 a_35391_n5745# gnd 2.50fF
C434 a_32790_n10642# gnd 5.48fF
C435 a_32995_n5746# gnd 3.68fF
C436 a_27815_n10678# gnd 5.48fF
C437 a_18908_n6280# gnd 2.28fF
C438 a_17970_n6524# gnd 2.45fF
C439 a_18912_n6092# gnd 2.38fF
C440 a_20304_n6156# gnd 2.23fF
C441 a_21040_n6152# gnd 2.52fF
C442 a_15205_n6221# gnd 2.23fF
C443 a_15941_n6217# gnd 2.52fF
C444 a_13852_n6239# gnd 2.28fF
C445 a_12914_n6483# gnd 2.45fF
C446 a_2887_n6290# gnd 2.52fF
C447 a_855_n6725# gnd 2.18fF
C448 a_13856_n6051# gnd 2.38fF
C449 a_28020_n5782# gnd 3.68fF
C450 a_32025_n5894# gnd 3.32fF
C451 a_32119_n5894# gnd 6.48fF
C452 a_27050_n5930# gnd 3.32fF
C453 a_27144_n5930# gnd 6.48fF
C454 a_39099_n5524# gnd 2.50fF
C455 a_30335_n5704# gnd 2.50fF
C456 a_35391_n5558# gnd 2.28fF
C457 a_25360_n5740# gnd 2.50fF
C458 a_22759_n10637# gnd 5.48fF
C459 a_22964_n5741# gnd 3.68fF
C460 a_17660_n10702# gnd 5.48fF
C461 a_8877_n6275# gnd 2.28fF
C462 a_7939_n6519# gnd 2.45fF
C463 a_8881_n6087# gnd 2.38fF
C464 a_10149_n6180# gnd 2.23fF
C465 a_10885_n6176# gnd 2.52fF
C466 a_5174_n6216# gnd 2.23fF
C467 a_5910_n6212# gnd 2.52fF
C468 a_3821_n6234# gnd 2.28fF
C469 a_2883_n6478# gnd 2.45fF
C470 a_3825_n6046# gnd 2.38fF
C471 a_17865_n5806# gnd 3.68fF
C472 a_16895_n5954# gnd 3.32fF
C473 a_16989_n5954# gnd 6.48fF
C474 a_21994_n5889# gnd 3.32fF
C475 a_22088_n5889# gnd 6.48fF
C476 a_34043_n5483# gnd 2.50fF
C477 a_39095_n5712# gnd 2.23fF
C478 a_29068_n5519# gnd 2.50fF
C479 a_30335_n5517# gnd 2.28fF
C480 a_20304_n5699# gnd 2.50fF
C481 a_25360_n5553# gnd 2.28fF
C482 a_15205_n5764# gnd 2.50fF
C483 a_12604_n10661# gnd 5.48fF
C484 a_12809_n5765# gnd 3.68fF
C485 a_7629_n10697# gnd 5.48fF
C486 a_118_n6175# gnd 2.23fF
C487 a_854_n6171# gnd 2.52fF
C488 a_7834_n5801# gnd 3.68fF
C489 a_11839_n5913# gnd 3.32fF
C490 a_11933_n5913# gnd 6.48fF
C491 a_6864_n5949# gnd 3.32fF
C492 a_6958_n5949# gnd 6.48fF
C493 a_24012_n5478# gnd 2.50fF
C494 a_35391_n5329# gnd 2.38fF
C495 a_34039_n5671# gnd 2.23fF
C496 a_38160_n5214# gnd 2.52fF
C497 a_36128_n5649# gnd 2.45fF
C498 a_29064_n5707# gnd 2.23fF
C499 a_30335_n5288# gnd 2.38fF
C500 a_18913_n5543# gnd 2.50fF
C501 a_10149_n5723# gnd 2.50fF
C502 a_15205_n5577# gnd 2.28fF
C503 a_5174_n5759# gnd 2.50fF
C504 a_2573_n10656# gnd 5.48fF
C505 a_2778_n5760# gnd 3.68fF
C506 a_1808_n5908# gnd 3.32fF
C507 a_1902_n5908# gnd 6.48fF
C508 a_13857_n5502# gnd 2.50fF
C509 a_20304_n5512# gnd 2.28fF
C510 a_18909_n5731# gnd 2.23fF
C511 a_25360_n5324# gnd 2.38fF
C512 a_33104_n5173# gnd 2.52fF
C513 a_31072_n5608# gnd 2.45fF
C514 a_24008_n5666# gnd 2.23fF
C515 a_28129_n5209# gnd 2.52fF
C516 a_26097_n5644# gnd 2.45fF
C517 a_20304_n5283# gnd 2.38fF
C518 a_8882_n5538# gnd 2.50fF
C519 a_10149_n5536# gnd 2.28fF
C520 a_118_n5718# gnd 2.50fF
C521 a_5174_n5572# gnd 2.28fF
C522 a_3826_n5497# gnd 2.50fF
C523 a_15205_n5348# gnd 2.38fF
C524 a_39094_n5158# gnd 2.28fF
C525 a_38156_n5402# gnd 2.18fF
C526 a_39098_n4970# gnd 2.38fF
C527 a_35391_n5099# gnd 2.23fF
C528 a_36127_n5095# gnd 2.52fF
C529 a_34038_n5117# gnd 2.28fF
C530 a_33100_n5361# gnd 2.18fF
C531 a_13853_n5690# gnd 2.23fF
C532 a_17974_n5233# gnd 2.52fF
C533 a_15942_n5668# gnd 2.45fF
C534 a_8878_n5726# gnd 2.23fF
C535 a_10149_n5307# gnd 2.38fF
C536 a_23073_n5168# gnd 2.52fF
C537 a_21041_n5603# gnd 2.45fF
C538 a_34042_n4929# gnd 2.38fF
C539 a_29063_n5153# gnd 2.28fF
C540 a_28125_n5397# gnd 2.18fF
C541 a_29067_n4965# gnd 2.38fF
C542 a_30335_n5058# gnd 2.23fF
C543 a_31071_n5054# gnd 2.52fF
C544 a_25360_n5094# gnd 2.23fF
C545 a_26096_n5090# gnd 2.52fF
C546 a_24007_n5112# gnd 2.28fF
C547 a_23069_n5356# gnd 2.18fF
C548 a_118_n5531# gnd 2.28fF
C549 a_5174_n5343# gnd 2.38fF
C550 a_12918_n5192# gnd 2.52fF
C551 a_10886_n5627# gnd 2.45fF
C552 a_3822_n5685# gnd 2.23fF
C553 a_7943_n5228# gnd 2.52fF
C554 a_5911_n5663# gnd 2.45fF
C555 a_118_n5302# gnd 2.38fF
C556 a_24011_n4924# gnd 2.38fF
C557 a_35392_n4642# gnd 2.49fF
C558 a_18908_n5177# gnd 2.28fF
C559 a_17970_n5421# gnd 2.18fF
C560 a_18912_n4989# gnd 2.38fF
C561 a_20304_n5053# gnd 2.23fF
C562 a_21040_n5049# gnd 2.52fF
C563 a_15205_n5118# gnd 2.23fF
C564 a_15941_n5114# gnd 2.52fF
C565 a_13852_n5136# gnd 2.28fF
C566 a_12914_n5380# gnd 2.18fF
C567 a_2887_n5187# gnd 2.52fF
C568 a_855_n5622# gnd 2.45fF
C569 a_13856_n4948# gnd 2.38fF
C570 a_8877_n5172# gnd 2.28fF
C571 a_7939_n5416# gnd 2.18fF
C572 a_8881_n4984# gnd 2.38fF
C573 a_30336_n4601# gnd 2.49fF
C574 a_25361_n4637# gnd 2.49fF
C575 a_10149_n5077# gnd 2.23fF
C576 a_10885_n5073# gnd 2.52fF
C577 a_5174_n5113# gnd 2.23fF
C578 a_5910_n5109# gnd 2.52fF
C579 a_3821_n5131# gnd 2.28fF
C580 a_2883_n5375# gnd 2.18fF
C581 a_3825_n4943# gnd 2.38fF
C582 a_39100_n4421# gnd 2.49fF
C583 a_35392_n4455# gnd 2.28fF
C584 a_34044_n4380# gnd 2.49fF
C585 a_39096_n4609# gnd 2.23fF
C586 a_20305_n4596# gnd 2.49fF
C587 a_15206_n4661# gnd 2.49fF
C588 a_29069_n4416# gnd 2.49fF
C589 a_30336_n4414# gnd 2.28fF
C590 a_25361_n4450# gnd 2.28fF
C591 a_118_n5072# gnd 2.23fF
C592 a_854_n5068# gnd 2.52fF
C593 a_24013_n4375# gnd 2.49fF
C594 a_35392_n4226# gnd 2.38fF
C595 a_34040_n4568# gnd 2.23fF
C596 a_38161_n4111# gnd 2.52fF
C597 a_36129_n4546# gnd 2.18fF
C598 a_29065_n4604# gnd 2.23fF
C599 a_30336_n4185# gnd 2.38fF
C600 a_10150_n4620# gnd 2.49fF
C601 a_5175_n4656# gnd 2.49fF
C602 a_18914_n4440# gnd 2.49fF
C603 a_15206_n4474# gnd 2.28fF
C604 a_13858_n4399# gnd 2.49fF
C605 a_20305_n4409# gnd 2.28fF
C606 a_18910_n4628# gnd 2.23fF
C607 a_25361_n4221# gnd 2.38fF
C608 a_33105_n4070# gnd 2.52fF
C609 a_31073_n4505# gnd 2.18fF
C610 a_24009_n4563# gnd 2.23fF
C611 a_28130_n4106# gnd 2.52fF
C612 a_26098_n4541# gnd 2.18fF
C613 a_20305_n4180# gnd 2.38fF
C614 a_119_n4615# gnd 2.49fF
C615 a_8883_n4435# gnd 2.49fF
C616 a_10150_n4433# gnd 2.28fF
C617 a_5175_n4469# gnd 2.28fF
C618 a_3827_n4394# gnd 2.49fF
C619 a_15206_n4245# gnd 2.38fF
C620 a_39095_n4055# gnd 2.28fF
C621 a_38157_n4299# gnd 2.45fF
C622 a_39099_n3867# gnd 2.38fF
C623 a_35392_n3996# gnd 2.23fF
C624 a_36128_n3992# gnd 2.52fF
C625 a_34039_n4014# gnd 2.28fF
C626 a_33101_n4258# gnd 2.45fF
C627 a_13854_n4587# gnd 2.23fF
C628 a_17975_n4130# gnd 2.52fF
C629 a_15943_n4565# gnd 2.18fF
C630 a_8879_n4623# gnd 2.23fF
C631 a_10150_n4204# gnd 2.38fF
C632 a_23074_n4065# gnd 2.52fF
C633 a_21042_n4500# gnd 2.18fF
C634 a_34043_n3826# gnd 2.38fF
C635 a_29064_n4050# gnd 2.28fF
C636 a_28126_n4294# gnd 2.45fF
C637 a_29068_n3862# gnd 2.38fF
C638 a_38047_n5975# gnd 3.32fF
C639 a_30336_n3955# gnd 2.23fF
C640 a_31072_n3951# gnd 2.52fF
C641 a_25361_n3991# gnd 2.23fF
C642 a_26097_n3987# gnd 2.52fF
C643 a_24008_n4009# gnd 2.28fF
C644 a_23070_n4253# gnd 2.45fF
C645 a_119_n4428# gnd 2.28fF
C646 a_5175_n4240# gnd 2.38fF
C647 a_12919_n4089# gnd 2.52fF
C648 a_10887_n4524# gnd 2.18fF
C649 a_3823_n4582# gnd 2.23fF
C650 a_7944_n4125# gnd 2.52fF
C651 a_5912_n4560# gnd 2.18fF
C652 a_119_n4199# gnd 2.38fF
C653 a_24012_n3821# gnd 2.38fF
C654 a_18909_n4074# gnd 2.28fF
C655 a_17971_n4318# gnd 2.45fF
C656 a_18913_n3886# gnd 2.38fF
C657 a_38051_n3587# gnd 2.34fF
C658 a_37083_n3723# gnd 2.45fF
C659 a_37076_n5758# gnd 3.68fF
C660 a_35392_n3539# gnd 2.49fF
C661 a_32991_n5934# gnd 3.32fF
C662 a_32995_n3546# gnd 2.34fF
C663 a_28016_n5970# gnd 3.32fF
C664 a_20305_n3950# gnd 2.23fF
C665 a_21041_n3946# gnd 2.52fF
C666 a_15206_n4015# gnd 2.23fF
C667 a_15942_n4011# gnd 2.52fF
C668 a_13853_n4033# gnd 2.28fF
C669 a_12915_n4277# gnd 2.45fF
C670 a_2888_n4084# gnd 2.52fF
C671 a_856_n4519# gnd 2.18fF
C672 a_13857_n3845# gnd 2.38fF
C673 a_8878_n4069# gnd 2.28fF
C674 a_7940_n4313# gnd 2.45fF
C675 a_8882_n3881# gnd 2.38fF
C676 a_28020_n3582# gnd 2.34fF
C677 a_32027_n3682# gnd 2.45fF
C678 a_32020_n5717# gnd 3.68fF
C679 a_30336_n3498# gnd 2.49fF
C680 a_27052_n3718# gnd 2.45fF
C681 a_27045_n5753# gnd 3.68fF
C682 a_25361_n3534# gnd 2.49fF
C683 a_22960_n5929# gnd 3.32fF
C684 a_22964_n3541# gnd 2.34fF
C685 a_17861_n5994# gnd 3.32fF
C686 a_10150_n3974# gnd 2.23fF
C687 a_10886_n3970# gnd 2.52fF
C688 a_5175_n4010# gnd 2.23fF
C689 a_5911_n4006# gnd 2.52fF
C690 a_3822_n4028# gnd 2.28fF
C691 a_2884_n4272# gnd 2.45fF
C692 a_3826_n3840# gnd 2.38fF
C693 a_17865_n3606# gnd 2.34fF
C694 a_39100_n3318# gnd 2.49fF
C695 a_35392_n3352# gnd 2.28fF
C696 a_34044_n3277# gnd 2.49fF
C697 a_39096_n3506# gnd 2.23fF
C698 a_21996_n3677# gnd 2.45fF
C699 a_21989_n5712# gnd 3.68fF
C700 a_20305_n3493# gnd 2.49fF
C701 a_16897_n3742# gnd 2.45fF
C702 a_16890_n5777# gnd 3.68fF
C703 a_15206_n3558# gnd 2.49fF
C704 a_12805_n5953# gnd 3.32fF
C705 a_12809_n3565# gnd 2.34fF
C706 a_7830_n5989# gnd 3.32fF
C707 a_119_n3969# gnd 2.23fF
C708 a_855_n3965# gnd 2.52fF
C709 a_7834_n3601# gnd 2.34fF
C710 a_29069_n3313# gnd 2.49fF
C711 a_30336_n3311# gnd 2.28fF
C712 a_25361_n3347# gnd 2.28fF
C713 a_24013_n3272# gnd 2.49fF
C714 a_35392_n3123# gnd 2.38fF
C715 a_34040_n3465# gnd 2.23fF
C716 a_38161_n3008# gnd 2.52fF
C717 a_36129_n3443# gnd 2.45fF
C718 a_29065_n3501# gnd 2.23fF
C719 a_30336_n3082# gnd 2.38fF
C720 a_11841_n3701# gnd 2.45fF
C721 a_11834_n5736# gnd 3.68fF
C722 a_10150_n3517# gnd 2.49fF
C723 a_6866_n3737# gnd 2.45fF
C724 a_6859_n5772# gnd 3.68fF
C725 a_5175_n3553# gnd 2.49fF
C726 a_2774_n5948# gnd 3.32fF
C727 a_2778_n3560# gnd 2.34fF
C728 a_18914_n3337# gnd 2.49fF
C729 a_15206_n3371# gnd 2.28fF
C730 a_13858_n3296# gnd 2.49fF
C731 a_20305_n3306# gnd 2.28fF
C732 a_18910_n3525# gnd 2.23fF
C733 a_25361_n3118# gnd 2.38fF
C734 a_33105_n2967# gnd 2.52fF
C735 a_31073_n3402# gnd 2.45fF
C736 a_24009_n3460# gnd 2.23fF
C737 a_28130_n3003# gnd 2.52fF
C738 a_26098_n3438# gnd 2.45fF
C739 a_20305_n3077# gnd 2.38fF
C740 a_1810_n3696# gnd 2.45fF
C741 a_1803_n5731# gnd 3.68fF
C742 a_119_n3512# gnd 2.49fF
C743 a_8883_n3332# gnd 2.49fF
C744 a_10150_n3330# gnd 2.28fF
C745 a_5175_n3366# gnd 2.28fF
C746 a_3827_n3291# gnd 2.49fF
C747 a_15206_n3142# gnd 2.38fF
C748 a_39095_n2952# gnd 2.28fF
C749 a_38157_n3196# gnd 2.18fF
C750 a_39099_n2764# gnd 2.38fF
C751 a_35392_n2893# gnd 2.23fF
C752 a_36128_n2889# gnd 2.52fF
C753 a_34039_n2911# gnd 2.28fF
C754 a_33101_n3155# gnd 2.18fF
C755 a_13854_n3484# gnd 2.23fF
C756 a_17975_n3027# gnd 2.52fF
C757 a_15943_n3462# gnd 2.45fF
C758 a_8879_n3520# gnd 2.23fF
C759 a_10150_n3101# gnd 2.38fF
C760 a_23074_n2962# gnd 2.52fF
C761 a_21042_n3397# gnd 2.45fF
C762 a_34043_n2723# gnd 2.38fF
C763 a_29064_n2947# gnd 2.28fF
C764 a_28126_n3191# gnd 2.18fF
C765 a_29068_n2759# gnd 2.38fF
C766 a_38047_n3775# gnd 2.04fF
C767 a_30336_n2852# gnd 2.23fF
C768 a_31072_n2848# gnd 2.52fF
C769 a_25361_n2888# gnd 2.23fF
C770 a_26097_n2884# gnd 2.52fF
C771 a_24008_n2906# gnd 2.28fF
C772 a_23070_n3150# gnd 2.18fF
C773 a_119_n3325# gnd 2.28fF
C774 a_5175_n3137# gnd 2.38fF
C775 a_12919_n2986# gnd 2.52fF
C776 a_10887_n3421# gnd 2.45fF
C777 a_3823_n3479# gnd 2.23fF
C778 a_7944_n3022# gnd 2.52fF
C779 a_5912_n3457# gnd 2.45fF
C780 a_119_n3096# gnd 2.38fF
C781 a_24012_n2718# gnd 2.38fF
C782 a_37078_n3546# gnd 2.28fF
C783 a_35393_n2436# gnd 2.49fF
C784 a_32991_n3734# gnd 2.04fF
C785 a_18909_n2971# gnd 2.28fF
C786 a_17971_n3215# gnd 2.18fF
C787 a_18913_n2783# gnd 2.38fF
C788 a_28016_n3770# gnd 2.04fF
C789 a_20305_n2847# gnd 2.23fF
C790 a_21041_n2843# gnd 2.52fF
C791 a_15206_n2912# gnd 2.23fF
C792 a_15942_n2908# gnd 2.52fF
C793 a_13853_n2930# gnd 2.28fF
C794 a_12915_n3174# gnd 2.18fF
C795 a_2888_n2981# gnd 2.52fF
C796 a_856_n3416# gnd 2.45fF
C797 a_13857_n2742# gnd 2.38fF
C798 a_8878_n2966# gnd 2.28fF
C799 a_7940_n3210# gnd 2.18fF
C800 a_8882_n2778# gnd 2.38fF
C801 a_32022_n3505# gnd 2.28fF
C802 a_30337_n2395# gnd 2.49fF
C803 a_27047_n3541# gnd 2.28fF
C804 a_25362_n2431# gnd 2.49fF
C805 a_22960_n3729# gnd 2.04fF
C806 a_17861_n3794# gnd 2.04fF
C807 a_10150_n2871# gnd 2.23fF
C808 a_10886_n2867# gnd 2.52fF
C809 a_5175_n2907# gnd 2.23fF
C810 a_5911_n2903# gnd 2.52fF
C811 a_3822_n2925# gnd 2.28fF
C812 a_2884_n3169# gnd 2.18fF
C813 a_3826_n2737# gnd 2.38fF
C814 a_39101_n2215# gnd 2.49fF
C815 a_35393_n2249# gnd 2.28fF
C816 a_34045_n2174# gnd 2.49fF
C817 a_39097_n2403# gnd 2.23fF
C818 a_21991_n3500# gnd 2.28fF
C819 a_20306_n2390# gnd 2.49fF
C820 a_16892_n3565# gnd 2.28fF
C821 a_15207_n2455# gnd 2.49fF
C822 a_12805_n3753# gnd 2.04fF
C823 a_29070_n2210# gnd 2.49fF
C824 a_30337_n2208# gnd 2.28fF
C825 a_25362_n2244# gnd 2.28fF
C826 a_7830_n3789# gnd 2.04fF
C827 a_119_n2866# gnd 2.23fF
C828 a_855_n2862# gnd 2.52fF
C829 a_24014_n2169# gnd 2.49fF
C830 a_35393_n2020# gnd 2.38fF
C831 a_34041_n2362# gnd 2.23fF
C832 a_38162_n1905# gnd 2.52fF
C833 a_36130_n2340# gnd 2.18fF
C834 a_29066_n2398# gnd 2.23fF
C835 a_30337_n1979# gnd 2.38fF
C836 a_11836_n3524# gnd 2.28fF
C837 a_10151_n2414# gnd 2.49fF
C838 a_6861_n3560# gnd 2.28fF
C839 a_5176_n2450# gnd 2.49fF
C840 a_2774_n3748# gnd 2.04fF
C841 a_18915_n2234# gnd 2.49fF
C842 a_15207_n2268# gnd 2.28fF
C843 a_13859_n2193# gnd 2.49fF
C844 a_20306_n2203# gnd 2.28fF
C845 a_18911_n2422# gnd 2.23fF
C846 a_25362_n2015# gnd 2.38fF
C847 a_33106_n1864# gnd 2.52fF
C848 a_31074_n2299# gnd 2.18fF
C849 a_24010_n2357# gnd 2.23fF
C850 a_28131_n1900# gnd 2.52fF
C851 a_26099_n2335# gnd 2.18fF
C852 a_20306_n1974# gnd 2.38fF
C853 a_1805_n3519# gnd 2.28fF
C854 a_120_n2409# gnd 2.49fF
C855 a_8884_n2229# gnd 2.49fF
C856 a_10151_n2227# gnd 2.28fF
C857 a_5176_n2263# gnd 2.28fF
C858 a_3828_n2188# gnd 2.49fF
C859 a_15207_n2039# gnd 2.38fF
C860 a_39096_n1849# gnd 2.22fF
C861 a_38158_n2093# gnd 2.38fF
C862 a_39100_n1661# gnd 2.38fF
C863 a_35393_n1790# gnd 2.23fF
C864 a_36129_n1786# gnd 2.52fF
C865 a_34040_n1808# gnd 2.22fF
C866 a_33102_n2052# gnd 2.38fF
C867 a_13855_n2381# gnd 2.23fF
C868 a_17976_n1924# gnd 2.52fF
C869 a_15944_n2359# gnd 2.18fF
C870 a_8880_n2417# gnd 2.23fF
C871 a_10151_n1998# gnd 2.38fF
C872 a_23075_n1859# gnd 2.52fF
C873 a_21043_n2294# gnd 2.18fF
C874 a_34044_n1620# gnd 2.38fF
C875 a_29065_n1844# gnd 2.22fF
C876 a_28127_n2088# gnd 2.38fF
C877 a_29069_n1656# gnd 2.38fF
C878 a_35016_n1511# gnd 2.98fF
C879 a_30337_n1749# gnd 2.23fF
C880 a_31073_n1745# gnd 2.52fF
C881 a_30041_n1547# gnd 2.82fF
C882 a_25362_n1785# gnd 2.23fF
C883 a_26098_n1781# gnd 2.52fF
C884 a_24009_n1803# gnd 2.22fF
C885 a_23071_n2047# gnd 2.38fF
C886 a_120_n2222# gnd 2.28fF
C887 a_5176_n2034# gnd 2.38fF
C888 a_12920_n1883# gnd 2.52fF
C889 a_10888_n2318# gnd 2.18fF
C890 a_3824_n2376# gnd 2.23fF
C891 a_7945_n1919# gnd 2.52fF
C892 a_5913_n2354# gnd 2.18fF
C893 a_120_n1993# gnd 2.38fF
C894 a_24013_n1615# gnd 2.38fF
C895 a_18910_n1868# gnd 2.22fF
C896 a_17972_n2112# gnd 2.38fF
C897 a_18914_n1680# gnd 2.38fF
C898 a_24985_n1506# gnd 2.98fF
C899 a_20306_n1744# gnd 2.23fF
C900 a_21042_n1740# gnd 2.52fF
C901 a_19886_n1571# gnd 2.97fF
C902 a_15207_n1809# gnd 2.23fF
C903 a_15943_n1805# gnd 2.52fF
C904 a_13854_n1827# gnd 2.22fF
C905 a_12916_n2071# gnd 2.38fF
C906 a_2889_n1878# gnd 2.52fF
C907 a_857_n2313# gnd 2.18fF
C908 a_13858_n1639# gnd 2.38fF
C909 a_8879_n1863# gnd 2.22fF
C910 a_7941_n2107# gnd 2.38fF
C911 a_8883_n1675# gnd 2.38fF
C912 a_14830_n1530# gnd 2.98fF
C913 a_10151_n1768# gnd 2.23fF
C914 a_10887_n1764# gnd 2.52fF
C915 a_9855_n1566# gnd 2.82fF
C916 a_5176_n1804# gnd 2.23fF
C917 a_5912_n1800# gnd 2.52fF
C918 a_3823_n1822# gnd 2.22fF
C919 a_2885_n2066# gnd 2.38fF
C920 a_3827_n1634# gnd 2.38fF
C921 a_4799_n1525# gnd 2.98fF
C922 a_120_n1763# gnd 2.75fF
C923 a_856_n1759# gnd 2.79fF
C924 a_19441_n829# gnd 12.08fF
C925 a_35171_466# gnd 3.40fF
C926 a_30074_345# gnd 6.50fF
C927 a_32320_486# gnd 4.59fF
C928 a_19317_288# gnd 11.66fF
C929 a_19416_288# gnd 2.27fF
C930 a_25140_461# gnd 3.40fF
C931 a_25239_461# gnd 7.14fF
C932 a_22289_481# gnd 4.59fF
C933 a_14985_485# gnd 3.40fF
C934 a_9888_364# gnd 6.50fF
C935 a_9987_364# gnd 11.31fF
C936 a_12134_505# gnd 4.59fF
C937 a_4954_480# gnd 3.40fF
C938 a_5053_480# gnd 7.14fF
C939 a_2103_500# gnd 4.59fF
C940 a_39096_1326# gnd 2.22fF
C941 a_35395_1192# gnd 6.43fF
C942 a_34040_1285# gnd 2.22fF
C943 a_30339_1151# gnd 6.43fF
C944 a_39100_1149# gnd 2.38fF
C945 a_35393_1291# gnd 2.23fF
C946 a_34044_1108# gnd 2.38fF
C947 a_38158_1570# gnd 2.38fF
C948 a_36129_1086# gnd 2.52fF
C949 a_29065_1321# gnd 2.22fF
C950 a_25364_1187# gnd 6.43fF
C951 a_24009_1280# gnd 2.22fF
C952 a_20308_1146# gnd 6.43fF
C953 a_30337_1250# gnd 2.23fF
C954 a_33102_1529# gnd 2.38fF
C955 a_31073_1045# gnd 2.52fF
C956 a_29069_1144# gnd 2.38fF
C957 a_25362_1286# gnd 2.23fF
C958 a_24013_1103# gnd 2.38fF
C959 a_35393_1521# gnd 2.38fF
C960 a_36130_1640# gnd 2.18fF
C961 a_28127_1565# gnd 2.38fF
C962 a_26098_1081# gnd 2.52fF
C963 a_20306_1245# gnd 2.23fF
C964 a_18910_1345# gnd 2.22fF
C965 a_15209_1211# gnd 6.43fF
C966 a_13854_1304# gnd 2.22fF
C967 a_10153_1170# gnd 6.43fF
C968 a_23071_1524# gnd 2.38fF
C969 a_21042_1040# gnd 2.52fF
C970 a_18914_1168# gnd 2.38fF
C971 a_35393_1750# gnd 2.28fF
C972 a_30337_1480# gnd 2.38fF
C973 a_31074_1599# gnd 2.18fF
C974 a_30337_1709# gnd 2.28fF
C975 a_38162_1393# gnd 2.52fF
C976 a_39097_1880# gnd 2.23fF
C977 a_33106_1352# gnd 2.52fF
C978 a_34041_1839# gnd 2.23fF
C979 a_25362_1516# gnd 2.38fF
C980 a_26099_1635# gnd 2.18fF
C981 a_15207_1310# gnd 2.23fF
C982 a_13858_1127# gnd 2.38fF
C983 a_17972_1589# gnd 2.38fF
C984 a_15943_1105# gnd 2.52fF
C985 a_8879_1340# gnd 2.22fF
C986 a_5178_1206# gnd 6.43fF
C987 a_3823_1299# gnd 2.22fF
C988 a_122_1165# gnd 6.43fF
C989 a_10151_1269# gnd 2.23fF
C990 a_12916_1548# gnd 2.38fF
C991 a_10887_1064# gnd 2.52fF
C992 a_8883_1163# gnd 2.38fF
C993 a_5176_1305# gnd 2.23fF
C994 a_3827_1122# gnd 2.38fF
C995 a_25362_1745# gnd 2.28fF
C996 a_20306_1475# gnd 2.38fF
C997 a_21043_1594# gnd 2.18fF
C998 a_20306_1704# gnd 2.28fF
C999 a_39101_1703# gnd 2.49fF
C1000 a_28131_1388# gnd 2.52fF
C1001 a_29066_1875# gnd 2.23fF
C1002 a_23075_1347# gnd 2.52fF
C1003 a_24010_1834# gnd 2.23fF
C1004 a_34045_1662# gnd 2.49fF
C1005 a_29070_1698# gnd 2.49fF
C1006 a_15207_1540# gnd 2.38fF
C1007 a_15944_1659# gnd 2.18fF
C1008 a_7941_1584# gnd 2.38fF
C1009 a_5912_1100# gnd 2.52fF
C1010 a_120_1264# gnd 2.23fF
C1011 a_2885_1543# gnd 2.38fF
C1012 a_856_1059# gnd 2.52fF
C1013 a_15207_1769# gnd 2.28fF
C1014 a_10151_1499# gnd 2.38fF
C1015 a_10888_1618# gnd 2.18fF
C1016 a_10151_1728# gnd 2.28fF
C1017 a_17976_1412# gnd 2.52fF
C1018 a_18911_1899# gnd 2.23fF
C1019 a_12920_1371# gnd 2.52fF
C1020 a_13855_1858# gnd 2.23fF
C1021 a_5176_1535# gnd 2.38fF
C1022 a_5913_1654# gnd 2.18fF
C1023 a_5176_1764# gnd 2.28fF
C1024 a_120_1494# gnd 2.38fF
C1025 a_857_1613# gnd 2.18fF
C1026 a_120_1723# gnd 2.28fF
C1027 a_24014_1657# gnd 2.49fF
C1028 a_39095_2429# gnd 2.28fF
C1029 a_35393_1937# gnd 2.49fF
C1030 a_34039_2388# gnd 2.28fF
C1031 a_30337_1896# gnd 2.49fF
C1032 a_39099_2252# gnd 2.38fF
C1033 a_35392_2394# gnd 2.23fF
C1034 a_34043_2211# gnd 2.38fF
C1035 a_38157_2673# gnd 2.18fF
C1036 a_36128_2189# gnd 2.52fF
C1037 a_29064_2424# gnd 2.28fF
C1038 a_25362_1932# gnd 2.49fF
C1039 a_18915_1722# gnd 2.49fF
C1040 a_7945_1407# gnd 2.52fF
C1041 a_8880_1894# gnd 2.23fF
C1042 a_2889_1366# gnd 2.52fF
C1043 a_3824_1853# gnd 2.23fF
C1044 a_13859_1681# gnd 2.49fF
C1045 a_24008_2383# gnd 2.28fF
C1046 a_20306_1891# gnd 2.49fF
C1047 a_8884_1717# gnd 2.49fF
C1048 a_3828_1676# gnd 2.49fF
C1049 a_30336_2353# gnd 2.23fF
C1050 a_33101_2632# gnd 2.18fF
C1051 a_31072_2148# gnd 2.52fF
C1052 a_29068_2247# gnd 2.38fF
C1053 a_25361_2389# gnd 2.23fF
C1054 a_24012_2206# gnd 2.38fF
C1055 a_35392_2624# gnd 2.38fF
C1056 a_36129_2743# gnd 2.45fF
C1057 a_28126_2668# gnd 2.18fF
C1058 a_26097_2184# gnd 2.52fF
C1059 a_20305_2348# gnd 2.23fF
C1060 a_18909_2448# gnd 2.28fF
C1061 a_15207_1956# gnd 2.49fF
C1062 a_13853_2407# gnd 2.28fF
C1063 a_10151_1915# gnd 2.49fF
C1064 a_23070_2627# gnd 2.18fF
C1065 a_21041_2143# gnd 2.52fF
C1066 a_18913_2271# gnd 2.38fF
C1067 a_35392_2853# gnd 2.28fF
C1068 a_30336_2583# gnd 2.38fF
C1069 a_31073_2702# gnd 2.45fF
C1070 a_30336_2812# gnd 2.28fF
C1071 a_38161_2496# gnd 2.52fF
C1072 a_39096_2983# gnd 2.23fF
C1073 a_33105_2455# gnd 2.52fF
C1074 a_34040_2942# gnd 2.23fF
C1075 a_25361_2619# gnd 2.38fF
C1076 a_26098_2738# gnd 2.45fF
C1077 a_15206_2413# gnd 2.23fF
C1078 a_13857_2230# gnd 2.38fF
C1079 a_17971_2692# gnd 2.18fF
C1080 a_15942_2208# gnd 2.52fF
C1081 a_8878_2443# gnd 2.28fF
C1082 a_5176_1951# gnd 2.49fF
C1083 a_3822_2402# gnd 2.28fF
C1084 a_120_1910# gnd 2.49fF
C1085 a_10150_2372# gnd 2.23fF
C1086 a_12915_2651# gnd 2.18fF
C1087 a_10886_2167# gnd 2.52fF
C1088 a_8882_2266# gnd 2.38fF
C1089 a_5175_2408# gnd 2.23fF
C1090 a_3826_2225# gnd 2.38fF
C1091 a_25361_2848# gnd 2.28fF
C1092 a_20305_2578# gnd 2.38fF
C1093 a_21042_2697# gnd 2.45fF
C1094 a_20305_2807# gnd 2.28fF
C1095 a_28130_2491# gnd 2.52fF
C1096 a_29065_2978# gnd 2.23fF
C1097 a_23074_2450# gnd 2.52fF
C1098 a_24009_2937# gnd 2.23fF
C1099 a_15206_2643# gnd 2.38fF
C1100 a_15943_2762# gnd 2.45fF
C1101 a_7940_2687# gnd 2.18fF
C1102 a_5911_2203# gnd 2.52fF
C1103 a_119_2367# gnd 2.23fF
C1104 a_2884_2646# gnd 2.18fF
C1105 a_855_2162# gnd 2.52fF
C1106 a_15206_2872# gnd 2.28fF
C1107 a_10150_2602# gnd 2.38fF
C1108 a_10887_2721# gnd 2.45fF
C1109 a_10150_2831# gnd 2.28fF
C1110 a_37078_3023# gnd 2.28fF
C1111 a_32022_2982# gnd 2.28fF
C1112 a_17975_2515# gnd 2.52fF
C1113 a_18910_3002# gnd 2.23fF
C1114 a_39100_2806# gnd 2.49fF
C1115 a_34044_2765# gnd 2.49fF
C1116 a_38047_3252# gnd 2.04fF
C1117 a_32991_3211# gnd 2.04fF
C1118 a_27047_3018# gnd 2.28fF
C1119 a_21991_2977# gnd 2.28fF
C1120 a_12919_2474# gnd 2.52fF
C1121 a_13854_2961# gnd 2.23fF
C1122 a_5175_2638# gnd 2.38fF
C1123 a_5912_2757# gnd 2.45fF
C1124 a_5175_2867# gnd 2.28fF
C1125 a_119_2597# gnd 2.38fF
C1126 a_856_2716# gnd 2.45fF
C1127 a_119_2826# gnd 2.28fF
C1128 a_29069_2801# gnd 2.49fF
C1129 a_39095_3532# gnd 2.28fF
C1130 a_35392_3040# gnd 2.49fF
C1131 a_24013_2760# gnd 2.49fF
C1132 a_28016_3247# gnd 2.04fF
C1133 a_7944_2510# gnd 2.52fF
C1134 a_8879_2997# gnd 2.23fF
C1135 a_2888_2469# gnd 2.52fF
C1136 a_3823_2956# gnd 2.23fF
C1137 a_22960_3206# gnd 2.04fF
C1138 a_16892_3042# gnd 2.28fF
C1139 a_11836_3001# gnd 2.28fF
C1140 a_34039_3491# gnd 2.28fF
C1141 a_30336_2999# gnd 2.49fF
C1142 a_39099_3355# gnd 2.38fF
C1143 a_35392_3497# gnd 2.23fF
C1144 a_34043_3314# gnd 2.38fF
C1145 a_38157_3776# gnd 2.45fF
C1146 a_36128_3292# gnd 2.52fF
C1147 a_29064_3527# gnd 2.28fF
C1148 a_25361_3035# gnd 2.49fF
C1149 a_18914_2825# gnd 2.49fF
C1150 a_24008_3486# gnd 2.28fF
C1151 a_20305_2994# gnd 2.49fF
C1152 a_13858_2784# gnd 2.49fF
C1153 a_17861_3271# gnd 2.04fF
C1154 a_12805_3230# gnd 2.04fF
C1155 a_6861_3037# gnd 2.28fF
C1156 a_1805_2996# gnd 2.28fF
C1157 a_8883_2820# gnd 2.49fF
C1158 a_30336_3456# gnd 2.23fF
C1159 a_33101_3735# gnd 2.45fF
C1160 a_31072_3251# gnd 2.52fF
C1161 a_29068_3350# gnd 2.38fF
C1162 a_25361_3492# gnd 2.23fF
C1163 a_24012_3309# gnd 2.38fF
C1164 a_35392_3727# gnd 2.38fF
C1165 a_36129_3846# gnd 2.18fF
C1166 a_28126_3771# gnd 2.45fF
C1167 a_26097_3287# gnd 2.52fF
C1168 a_20305_3451# gnd 2.23fF
C1169 a_18909_3551# gnd 2.28fF
C1170 a_15206_3059# gnd 2.49fF
C1171 a_3827_2779# gnd 2.49fF
C1172 a_7830_3266# gnd 2.04fF
C1173 a_2774_3225# gnd 2.04fF
C1174 a_13853_3510# gnd 2.28fF
C1175 a_10150_3018# gnd 2.49fF
C1176 a_23070_3730# gnd 2.45fF
C1177 a_21041_3246# gnd 2.52fF
C1178 a_18913_3374# gnd 2.38fF
C1179 a_35392_3956# gnd 2.28fF
C1180 a_30336_3686# gnd 2.38fF
C1181 a_31073_3805# gnd 2.18fF
C1182 a_30336_3915# gnd 2.28fF
C1183 a_38161_3599# gnd 2.52fF
C1184 a_39096_4086# gnd 2.23fF
C1185 a_33105_3558# gnd 2.52fF
C1186 a_34040_4045# gnd 2.23fF
C1187 a_25361_3722# gnd 2.38fF
C1188 a_26098_3841# gnd 2.18fF
C1189 a_15206_3516# gnd 2.23fF
C1190 a_13857_3333# gnd 2.38fF
C1191 a_17971_3795# gnd 2.45fF
C1192 a_15942_3311# gnd 2.52fF
C1193 a_8878_3546# gnd 2.28fF
C1194 a_5175_3054# gnd 2.49fF
C1195 a_3822_3505# gnd 2.28fF
C1196 a_119_3013# gnd 2.49fF
C1197 a_10150_3475# gnd 2.23fF
C1198 a_12915_3754# gnd 2.45fF
C1199 a_10886_3270# gnd 2.52fF
C1200 a_8882_3369# gnd 2.38fF
C1201 a_5175_3511# gnd 2.23fF
C1202 a_3826_3328# gnd 2.38fF
C1203 a_25361_3951# gnd 2.28fF
C1204 a_20305_3681# gnd 2.38fF
C1205 a_21042_3800# gnd 2.18fF
C1206 a_20305_3910# gnd 2.28fF
C1207 a_39100_3909# gnd 2.49fF
C1208 a_37083_3142# gnd 2.45fF
C1209 a_28130_3594# gnd 2.52fF
C1210 a_29065_4081# gnd 2.23fF
C1211 a_23074_3553# gnd 2.52fF
C1212 a_24009_4040# gnd 2.23fF
C1213 a_34044_3868# gnd 2.49fF
C1214 a_32027_3101# gnd 2.45fF
C1215 a_38051_3075# gnd 2.34fF
C1216 a_32995_3034# gnd 2.34fF
C1217 a_29069_3904# gnd 2.49fF
C1218 a_27052_3137# gnd 2.45fF
C1219 a_15206_3746# gnd 2.38fF
C1220 a_15943_3865# gnd 2.18fF
C1221 a_7940_3790# gnd 2.45fF
C1222 a_5911_3306# gnd 2.52fF
C1223 a_119_3470# gnd 2.23fF
C1224 a_2884_3749# gnd 2.45fF
C1225 a_855_3265# gnd 2.52fF
C1226 a_15206_3975# gnd 2.28fF
C1227 a_10150_3705# gnd 2.38fF
C1228 a_10887_3824# gnd 2.18fF
C1229 a_10150_3934# gnd 2.28fF
C1230 a_17975_3618# gnd 2.52fF
C1231 a_18910_4105# gnd 2.23fF
C1232 a_12919_3577# gnd 2.52fF
C1233 a_13854_4064# gnd 2.23fF
C1234 a_5175_3741# gnd 2.38fF
C1235 a_5912_3860# gnd 2.18fF
C1236 a_5175_3970# gnd 2.28fF
C1237 a_119_3700# gnd 2.38fF
C1238 a_856_3819# gnd 2.18fF
C1239 a_119_3929# gnd 2.28fF
C1240 a_24013_3863# gnd 2.49fF
C1241 a_21996_3096# gnd 2.45fF
C1242 a_39094_4635# gnd 2.28fF
C1243 a_35392_4143# gnd 2.49fF
C1244 a_28020_3070# gnd 2.34fF
C1245 a_22964_3029# gnd 2.34fF
C1246 a_34038_4594# gnd 2.28fF
C1247 a_30336_4102# gnd 2.49fF
C1248 a_39098_4458# gnd 2.38fF
C1249 a_35391_4600# gnd 2.23fF
C1250 a_34042_4417# gnd 2.38fF
C1251 a_38156_4879# gnd 2.18fF
C1252 a_36127_4395# gnd 2.52fF
C1253 a_29063_4630# gnd 2.28fF
C1254 a_25361_4138# gnd 2.49fF
C1255 a_18914_3928# gnd 2.49fF
C1256 a_16897_3161# gnd 2.45fF
C1257 a_7944_3613# gnd 2.52fF
C1258 a_8879_4100# gnd 2.23fF
C1259 a_2888_3572# gnd 2.52fF
C1260 a_3823_4059# gnd 2.23fF
C1261 a_13858_3887# gnd 2.49fF
C1262 a_11841_3120# gnd 2.45fF
C1263 a_24007_4589# gnd 2.28fF
C1264 a_20305_4097# gnd 2.49fF
C1265 a_17865_3094# gnd 2.34fF
C1266 a_12809_3053# gnd 2.34fF
C1267 a_8883_3923# gnd 2.49fF
C1268 a_6866_3156# gnd 2.45fF
C1269 a_3827_3882# gnd 2.49fF
C1270 a_1810_3115# gnd 2.45fF
C1271 a_30335_4559# gnd 2.23fF
C1272 a_33100_4838# gnd 2.18fF
C1273 a_31071_4354# gnd 2.52fF
C1274 a_29067_4453# gnd 2.38fF
C1275 a_25360_4595# gnd 2.23fF
C1276 a_24011_4412# gnd 2.38fF
C1277 a_35391_4830# gnd 2.38fF
C1278 a_36128_4949# gnd 2.45fF
C1279 a_28125_4874# gnd 2.18fF
C1280 a_26096_4390# gnd 2.52fF
C1281 a_20304_4554# gnd 2.23fF
C1282 a_18908_4654# gnd 2.28fF
C1283 a_15206_4162# gnd 2.49fF
C1284 a_7834_3089# gnd 2.34fF
C1285 a_2778_3048# gnd 2.34fF
C1286 a_13852_4613# gnd 2.28fF
C1287 a_10150_4121# gnd 2.49fF
C1288 a_23069_4833# gnd 2.18fF
C1289 a_21040_4349# gnd 2.52fF
C1290 a_18912_4477# gnd 2.38fF
C1291 a_35391_5059# gnd 2.28fF
C1292 a_30335_4789# gnd 2.38fF
C1293 a_31072_4908# gnd 2.45fF
C1294 a_30335_5018# gnd 2.28fF
C1295 a_38160_4702# gnd 2.52fF
C1296 a_39095_5189# gnd 2.23fF
C1297 a_33104_4661# gnd 2.52fF
C1298 a_34039_5148# gnd 2.23fF
C1299 a_25360_4825# gnd 2.38fF
C1300 a_26097_4944# gnd 2.45fF
C1301 a_15205_4619# gnd 2.23fF
C1302 a_13856_4436# gnd 2.38fF
C1303 a_17970_4898# gnd 2.18fF
C1304 a_15941_4414# gnd 2.52fF
C1305 a_8877_4649# gnd 2.28fF
C1306 a_5175_4157# gnd 2.49fF
C1307 a_3821_4608# gnd 2.28fF
C1308 a_119_4116# gnd 2.49fF
C1309 a_10149_4578# gnd 2.23fF
C1310 a_12914_4857# gnd 2.18fF
C1311 a_10885_4373# gnd 2.52fF
C1312 a_8881_4472# gnd 2.38fF
C1313 a_5174_4614# gnd 2.23fF
C1314 a_3825_4431# gnd 2.38fF
C1315 a_25360_5054# gnd 2.28fF
C1316 a_20304_4784# gnd 2.38fF
C1317 a_21041_4903# gnd 2.45fF
C1318 a_20304_5013# gnd 2.28fF
C1319 a_28129_4697# gnd 2.52fF
C1320 a_29064_5184# gnd 2.23fF
C1321 a_39099_5012# gnd 2.50fF
C1322 a_37277_527# gnd 6.48fF
C1323 a_37076_5235# gnd 3.68fF
C1324 a_37175_5235# gnd 5.48fF
C1325 a_34043_4971# gnd 2.50fF
C1326 a_38047_5452# gnd 3.32fF
C1327 a_32221_486# gnd 6.48fF
C1328 a_32020_5194# gnd 3.68fF
C1329 a_32119_5194# gnd 5.48fF
C1330 a_23073_4656# gnd 2.52fF
C1331 a_24008_5143# gnd 2.23fF
C1332 a_15205_4849# gnd 2.38fF
C1333 a_15942_4968# gnd 2.45fF
C1334 a_7939_4893# gnd 2.18fF
C1335 a_5910_4409# gnd 2.52fF
C1336 a_118_4573# gnd 2.23fF
C1337 a_2883_4852# gnd 2.18fF
C1338 a_854_4368# gnd 2.52fF
C1339 a_15205_5078# gnd 2.28fF
C1340 a_10149_4808# gnd 2.38fF
C1341 a_10886_4927# gnd 2.45fF
C1342 a_10149_5037# gnd 2.28fF
C1343 a_17974_4721# gnd 2.52fF
C1344 a_18909_5208# gnd 2.23fF
C1345 a_32991_5411# gnd 3.32fF
C1346 a_29068_5007# gnd 2.50fF
C1347 a_39094_5738# gnd 2.28fF
C1348 a_35391_5246# gnd 2.50fF
C1349 a_27246_522# gnd 6.48fF
C1350 a_27045_5230# gnd 3.68fF
C1351 a_27144_5230# gnd 5.48fF
C1352 a_24012_4966# gnd 2.50fF
C1353 a_28016_5447# gnd 3.32fF
C1354 a_22190_481# gnd 6.48fF
C1355 a_21989_5189# gnd 3.68fF
C1356 a_22088_5189# gnd 5.48fF
C1357 a_12918_4680# gnd 2.52fF
C1358 a_13853_5167# gnd 2.23fF
C1359 a_5174_4844# gnd 2.38fF
C1360 a_5911_4963# gnd 2.45fF
C1361 a_5174_5073# gnd 2.28fF
C1362 a_118_4803# gnd 2.38fF
C1363 a_855_4922# gnd 2.45fF
C1364 a_118_5032# gnd 2.28fF
C1365 a_7943_4716# gnd 2.52fF
C1366 a_8878_5203# gnd 2.23fF
C1367 a_22960_5406# gnd 3.32fF
C1368 a_34038_5697# gnd 2.28fF
C1369 a_30335_5205# gnd 2.50fF
C1370 a_39098_5561# gnd 2.38fF
C1371 a_35391_5703# gnd 2.23fF
C1372 a_34042_5520# gnd 2.38fF
C1373 a_38156_5982# gnd 2.45fF
C1374 a_36127_5498# gnd 2.52fF
C1375 a_29063_5733# gnd 2.28fF
C1376 a_25360_5241# gnd 2.50fF
C1377 a_18913_5031# gnd 2.50fF
C1378 a_24007_5692# gnd 2.28fF
C1379 a_20304_5200# gnd 2.50fF
C1380 a_17091_546# gnd 6.48fF
C1381 a_16890_5254# gnd 3.68fF
C1382 a_16989_5254# gnd 5.48fF
C1383 a_13857_4990# gnd 2.50fF
C1384 a_17861_5471# gnd 3.32fF
C1385 a_12035_505# gnd 6.48fF
C1386 a_11834_5213# gnd 3.68fF
C1387 a_11933_5213# gnd 5.48fF
C1388 a_2887_4675# gnd 2.52fF
C1389 a_3822_5162# gnd 2.23fF
C1390 a_12805_5430# gnd 3.32fF
C1391 a_8882_5026# gnd 2.50fF
C1392 a_30335_5662# gnd 2.23fF
C1393 a_33100_5941# gnd 2.45fF
C1394 a_31071_5457# gnd 2.52fF
C1395 a_29067_5556# gnd 2.38fF
C1396 a_25360_5698# gnd 2.23fF
C1397 a_24011_5515# gnd 2.38fF
C1398 a_35391_5933# gnd 2.38fF
C1399 a_36128_6052# gnd 2.18fF
C1400 a_28125_5977# gnd 2.45fF
C1401 a_26096_5493# gnd 2.52fF
C1402 a_20304_5657# gnd 2.23fF
C1403 a_18908_5757# gnd 2.28fF
C1404 a_15205_5265# gnd 2.50fF
C1405 a_7060_541# gnd 6.48fF
C1406 a_6859_5249# gnd 3.68fF
C1407 a_6958_5249# gnd 5.48fF
C1408 a_3826_4985# gnd 2.50fF
C1409 a_7830_5466# gnd 3.32fF
C1410 a_2004_500# gnd 6.48fF
C1411 a_1803_5208# gnd 3.68fF
C1412 a_1902_5208# gnd 5.48fF
C1413 a_2774_5425# gnd 3.32fF
C1414 a_13852_5716# gnd 2.28fF
C1415 a_10149_5224# gnd 2.50fF
C1416 a_23069_5936# gnd 2.45fF
C1417 a_21040_5452# gnd 2.52fF
C1418 a_18912_5580# gnd 2.38fF
C1419 a_35391_6162# gnd 2.28fF
C1420 a_30335_5892# gnd 2.38fF
C1421 a_31072_6011# gnd 2.18fF
C1422 a_30335_6121# gnd 2.28fF
C1423 a_38160_5805# gnd 2.52fF
C1424 a_39095_6292# gnd 2.23fF
C1425 a_33104_5764# gnd 2.52fF
C1426 a_34039_6251# gnd 2.23fF
C1427 a_25360_5928# gnd 2.38fF
C1428 a_26097_6047# gnd 2.18fF
C1429 a_15205_5722# gnd 2.23fF
C1430 a_13856_5539# gnd 2.38fF
C1431 a_17970_6001# gnd 2.45fF
C1432 a_15941_5517# gnd 2.52fF
C1433 a_8877_5752# gnd 2.28fF
C1434 a_5174_5260# gnd 2.50fF
C1435 a_3821_5711# gnd 2.28fF
C1436 a_118_5219# gnd 2.50fF
C1437 a_10149_5681# gnd 2.23fF
C1438 a_12914_5960# gnd 2.45fF
C1439 a_10885_5476# gnd 2.52fF
C1440 a_8881_5575# gnd 2.38fF
C1441 a_5174_5717# gnd 2.23fF
C1442 a_3825_5534# gnd 2.38fF
C1443 a_25360_6157# gnd 2.28fF
C1444 a_20304_5887# gnd 2.38fF
C1445 a_21041_6006# gnd 2.18fF
C1446 a_20304_6116# gnd 2.28fF
C1447 a_39099_6115# gnd 2.49fF
C1448 a_28129_5800# gnd 2.52fF
C1449 a_29064_6287# gnd 2.23fF
C1450 a_23073_5759# gnd 2.52fF
C1451 a_24008_6246# gnd 2.23fF
C1452 a_34043_6074# gnd 2.49fF
C1453 a_29068_6110# gnd 2.49fF
C1454 a_15205_5952# gnd 2.38fF
C1455 a_15942_6071# gnd 2.18fF
C1456 a_7939_5996# gnd 2.45fF
C1457 a_5910_5512# gnd 2.52fF
C1458 a_118_5676# gnd 2.23fF
C1459 a_2883_5955# gnd 2.45fF
C1460 a_854_5471# gnd 2.52fF
C1461 a_15205_6181# gnd 2.28fF
C1462 a_10149_5911# gnd 2.38fF
C1463 a_10886_6030# gnd 2.18fF
C1464 a_10149_6140# gnd 2.28fF
C1465 a_17974_5824# gnd 2.52fF
C1466 a_18909_6311# gnd 2.23fF
C1467 a_12918_5783# gnd 2.52fF
C1468 a_13853_6270# gnd 2.23fF
C1469 a_5174_5947# gnd 2.38fF
C1470 a_5911_6066# gnd 2.18fF
C1471 a_5174_6176# gnd 2.28fF
C1472 a_118_5906# gnd 2.38fF
C1473 a_855_6025# gnd 2.18fF
C1474 a_118_6135# gnd 2.28fF
C1475 a_24012_6069# gnd 2.49fF
C1476 a_39093_6841# gnd 2.28fF
C1477 a_35391_6349# gnd 2.49fF
C1478 a_34037_6800# gnd 2.28fF
C1479 a_30335_6308# gnd 2.49fF
C1480 a_39097_6664# gnd 2.38fF
C1481 a_35390_6806# gnd 2.23fF
C1482 a_34041_6623# gnd 2.38fF
C1483 a_38155_7085# gnd 2.18fF
C1484 a_36126_6601# gnd 2.52fF
C1485 a_29062_6836# gnd 2.28fF
C1486 a_25360_6344# gnd 2.49fF
C1487 a_18913_6134# gnd 2.49fF
C1488 a_7943_5819# gnd 2.52fF
C1489 a_8878_6306# gnd 2.23fF
C1490 a_2887_5778# gnd 2.52fF
C1491 a_3822_6265# gnd 2.23fF
C1492 a_13857_6093# gnd 2.49fF
C1493 a_24006_6795# gnd 2.28fF
C1494 a_20304_6303# gnd 2.49fF
C1495 a_8882_6129# gnd 2.49fF
C1496 a_3826_6088# gnd 2.49fF
C1497 a_30334_6765# gnd 2.23fF
C1498 a_33099_7044# gnd 2.18fF
C1499 a_31070_6560# gnd 2.52fF
C1500 a_29066_6659# gnd 2.38fF
C1501 a_25359_6801# gnd 2.23fF
C1502 a_24010_6618# gnd 2.38fF
C1503 a_35390_7036# gnd 2.38fF
C1504 a_36127_7155# gnd 2.45fF
C1505 a_28124_7080# gnd 2.18fF
C1506 a_26095_6596# gnd 2.52fF
C1507 a_20303_6760# gnd 2.23fF
C1508 a_18907_6860# gnd 2.28fF
C1509 a_15205_6368# gnd 2.49fF
C1510 a_13851_6819# gnd 2.28fF
C1511 a_10149_6327# gnd 2.49fF
C1512 a_23068_7039# gnd 2.18fF
C1513 a_21039_6555# gnd 2.52fF
C1514 a_18911_6683# gnd 2.38fF
C1515 a_35390_7265# gnd 2.28fF
C1516 a_30334_6995# gnd 2.38fF
C1517 a_31071_7114# gnd 2.45fF
C1518 a_30334_7224# gnd 2.28fF
C1519 a_38159_6908# gnd 2.52fF
C1520 a_39094_7395# gnd 2.23fF
C1521 a_33103_6867# gnd 2.52fF
C1522 a_34038_7354# gnd 2.23fF
C1523 a_25359_7031# gnd 2.38fF
C1524 a_26096_7150# gnd 2.45fF
C1525 a_15204_6825# gnd 2.23fF
C1526 a_13855_6642# gnd 2.38fF
C1527 a_17969_7104# gnd 2.18fF
C1528 a_15940_6620# gnd 2.52fF
C1529 a_8876_6855# gnd 2.28fF
C1530 a_5174_6363# gnd 2.49fF
C1531 a_3820_6814# gnd 2.28fF
C1532 a_118_6322# gnd 2.49fF
C1533 a_10148_6784# gnd 2.23fF
C1534 a_12913_7063# gnd 2.18fF
C1535 a_10884_6579# gnd 2.52fF
C1536 a_8880_6678# gnd 2.38fF
C1537 a_5173_6820# gnd 2.23fF
C1538 a_3824_6637# gnd 2.38fF
C1539 a_25359_7260# gnd 2.28fF
C1540 a_20303_6990# gnd 2.38fF
C1541 a_21040_7109# gnd 2.45fF
C1542 a_20303_7219# gnd 2.28fF
C1543 a_28128_6903# gnd 2.52fF
C1544 a_29063_7390# gnd 2.23fF
C1545 a_23072_6862# gnd 2.52fF
C1546 a_24007_7349# gnd 2.23fF
C1547 a_15204_7055# gnd 2.38fF
C1548 a_15941_7174# gnd 2.45fF
C1549 a_7938_7099# gnd 2.18fF
C1550 a_5909_6615# gnd 2.52fF
C1551 a_117_6779# gnd 2.23fF
C1552 a_2882_7058# gnd 2.18fF
C1553 a_853_6574# gnd 2.52fF
C1554 a_15204_7284# gnd 2.28fF
C1555 a_10148_7014# gnd 2.38fF
C1556 a_10885_7133# gnd 2.45fF
C1557 a_10148_7243# gnd 2.28fF
C1558 a_37076_7435# gnd 2.34fF
C1559 a_37081_5354# gnd 3.32fF
C1560 a_32020_7394# gnd 2.34fF
C1561 a_32025_5313# gnd 3.32fF
C1562 a_17973_6927# gnd 2.52fF
C1563 a_18908_7414# gnd 2.23fF
C1564 a_39098_7218# gnd 2.49fF
C1565 a_38051_5275# gnd 3.68fF
C1566 a_34042_7177# gnd 2.49fF
C1567 a_38045_7664# gnd 2.45fF
C1568 a_32995_5234# gnd 3.68fF
C1569 a_32989_7623# gnd 2.45fF
C1570 a_27045_7430# gnd 2.34fF
C1571 a_27050_5349# gnd 3.32fF
C1572 a_21989_7389# gnd 2.34fF
C1573 a_21994_5308# gnd 3.32fF
C1574 a_12917_6886# gnd 2.52fF
C1575 a_13852_7373# gnd 2.23fF
C1576 a_5173_7050# gnd 2.38fF
C1577 a_5910_7169# gnd 2.45fF
C1578 a_5173_7279# gnd 2.28fF
C1579 a_117_7009# gnd 2.38fF
C1580 a_854_7128# gnd 2.45fF
C1581 a_117_7238# gnd 2.28fF
C1582 a_29067_7213# gnd 2.49fF
C1583 a_39093_7944# gnd 2.28fF
C1584 a_35390_7452# gnd 2.49fF
C1585 a_28020_5270# gnd 3.68fF
C1586 a_24011_7172# gnd 2.49fF
C1587 a_28014_7659# gnd 2.45fF
C1588 a_22964_5229# gnd 3.68fF
C1589 a_7942_6922# gnd 2.52fF
C1590 a_8877_7409# gnd 2.23fF
C1591 a_2886_6881# gnd 2.52fF
C1592 a_3821_7368# gnd 2.23fF
C1593 a_22958_7618# gnd 2.45fF
C1594 a_16890_7454# gnd 2.34fF
C1595 a_16895_5373# gnd 3.32fF
C1596 a_11834_7413# gnd 2.34fF
C1597 a_11839_5332# gnd 3.32fF
C1598 a_34037_7903# gnd 2.28fF
C1599 a_30334_7411# gnd 2.49fF
C1600 a_39097_7767# gnd 2.38fF
C1601 a_35390_7909# gnd 2.23fF
C1602 a_34041_7726# gnd 2.38fF
C1603 a_38155_8188# gnd 2.45fF
C1604 a_36126_7704# gnd 2.52fF
C1605 a_29062_7939# gnd 2.28fF
C1606 a_25359_7447# gnd 2.49fF
C1607 a_18912_7237# gnd 2.49fF
C1608 a_24006_7898# gnd 2.28fF
C1609 a_20303_7406# gnd 2.49fF
C1610 a_17865_5294# gnd 3.68fF
C1611 a_13856_7196# gnd 2.49fF
C1612 a_17859_7683# gnd 2.45fF
C1613 a_12809_5253# gnd 3.68fF
C1614 a_12803_7642# gnd 2.45fF
C1615 a_6859_7449# gnd 2.34fF
C1616 a_6864_5368# gnd 3.32fF
C1617 a_1803_7408# gnd 2.34fF
C1618 a_1808_5327# gnd 3.32fF
C1619 a_8881_7232# gnd 2.49fF
C1620 a_30334_7868# gnd 2.23fF
C1621 a_33099_8147# gnd 2.45fF
C1622 a_31070_7663# gnd 2.52fF
C1623 a_29066_7762# gnd 2.38fF
C1624 a_25359_7904# gnd 2.23fF
C1625 a_24010_7721# gnd 2.38fF
C1626 a_35390_8139# gnd 2.38fF
C1627 a_36127_8258# gnd 2.18fF
C1628 a_28124_8183# gnd 2.45fF
C1629 a_26095_7699# gnd 2.52fF
C1630 a_20303_7863# gnd 2.23fF
C1631 a_18907_7963# gnd 2.28fF
C1632 a_15204_7471# gnd 2.49fF
C1633 a_7834_5289# gnd 3.68fF
C1634 a_3825_7191# gnd 2.49fF
C1635 a_7828_7678# gnd 2.45fF
C1636 a_2778_5248# gnd 3.68fF
C1637 a_2772_7637# gnd 2.45fF
C1638 a_13851_7922# gnd 2.28fF
C1639 a_10148_7430# gnd 2.49fF
C1640 a_23068_8142# gnd 2.45fF
C1641 a_21039_7658# gnd 2.52fF
C1642 a_18911_7786# gnd 2.38fF
C1643 a_35390_8368# gnd 2.28fF
C1644 a_30334_8098# gnd 2.38fF
C1645 a_31071_8217# gnd 2.18fF
C1646 a_30334_8327# gnd 2.28fF
C1647 a_38159_8011# gnd 2.52fF
C1648 a_39094_8498# gnd 2.23fF
C1649 a_33103_7970# gnd 2.52fF
C1650 a_34038_8457# gnd 2.23fF
C1651 a_25359_8134# gnd 2.38fF
C1652 a_26096_8253# gnd 2.18fF
C1653 a_15204_7928# gnd 2.23fF
C1654 a_13855_7745# gnd 2.38fF
C1655 a_17969_8207# gnd 2.45fF
C1656 a_15940_7723# gnd 2.52fF
C1657 a_8876_7958# gnd 2.28fF
C1658 a_5173_7466# gnd 2.49fF
C1659 a_3820_7917# gnd 2.28fF
C1660 a_117_7425# gnd 2.49fF
C1661 a_10148_7887# gnd 2.23fF
C1662 a_12913_8166# gnd 2.45fF
C1663 a_10884_7682# gnd 2.52fF
C1664 a_8880_7781# gnd 2.38fF
C1665 a_5173_7923# gnd 2.23fF
C1666 a_3824_7740# gnd 2.38fF
C1667 a_25359_8363# gnd 2.28fF
C1668 a_20303_8093# gnd 2.38fF
C1669 a_21040_8212# gnd 2.18fF
C1670 a_20303_8322# gnd 2.28fF
C1671 a_39098_8321# gnd 2.49fF
C1672 a_37081_7554# gnd 2.04fF
C1673 a_28128_8006# gnd 2.52fF
C1674 a_29063_8493# gnd 2.23fF
C1675 a_23072_7965# gnd 2.52fF
C1676 a_24007_8452# gnd 2.23fF
C1677 a_34042_8280# gnd 2.49fF
C1678 a_32025_7513# gnd 2.04fF
C1679 a_38049_7487# gnd 2.28fF
C1680 a_32993_7446# gnd 2.28fF
C1681 a_29067_8316# gnd 2.49fF
C1682 a_27050_7549# gnd 2.04fF
C1683 a_15204_8158# gnd 2.38fF
C1684 a_15941_8277# gnd 2.18fF
C1685 a_7938_8202# gnd 2.45fF
C1686 a_5909_7718# gnd 2.52fF
C1687 a_117_7882# gnd 2.23fF
C1688 a_2882_8161# gnd 2.45fF
C1689 a_853_7677# gnd 2.52fF
C1690 a_15204_8387# gnd 2.28fF
C1691 a_10148_8117# gnd 2.38fF
C1692 a_10885_8236# gnd 2.18fF
C1693 a_10148_8346# gnd 2.28fF
C1694 a_17973_8030# gnd 2.52fF
C1695 a_18908_8517# gnd 2.23fF
C1696 a_12917_7989# gnd 2.52fF
C1697 a_13852_8476# gnd 2.23fF
C1698 a_5173_8153# gnd 2.38fF
C1699 a_5910_8272# gnd 2.18fF
C1700 a_5173_8382# gnd 2.28fF
C1701 a_117_8112# gnd 2.38fF
C1702 a_854_8231# gnd 2.18fF
C1703 a_117_8341# gnd 2.28fF
C1704 a_24011_8275# gnd 2.49fF
C1705 a_21994_7508# gnd 2.04fF
C1706 a_39092_9047# gnd 2.28fF
C1707 a_35390_8555# gnd 2.49fF
C1708 a_28018_7482# gnd 2.28fF
C1709 a_22962_7441# gnd 2.28fF
C1710 a_34036_9006# gnd 2.28fF
C1711 a_30334_8514# gnd 2.49fF
C1712 a_39096_8870# gnd 2.38fF
C1713 a_35389_9012# gnd 2.23fF
C1714 a_34040_8829# gnd 2.38fF
C1715 a_38154_9291# gnd 2.18fF
C1716 a_36125_8807# gnd 2.52fF
C1717 a_29061_9042# gnd 2.28fF
C1718 a_25359_8550# gnd 2.49fF
C1719 a_18912_8340# gnd 2.49fF
C1720 a_16895_7573# gnd 2.04fF
C1721 a_7942_8025# gnd 2.52fF
C1722 a_8877_8512# gnd 2.23fF
C1723 a_2886_7984# gnd 2.52fF
C1724 a_3821_8471# gnd 2.23fF
C1725 a_13856_8299# gnd 2.49fF
C1726 a_11839_7532# gnd 2.04fF
C1727 a_24005_9001# gnd 2.28fF
C1728 a_20303_8509# gnd 2.49fF
C1729 a_17863_7506# gnd 2.28fF
C1730 a_12807_7465# gnd 2.28fF
C1731 a_8881_8335# gnd 2.49fF
C1732 a_6864_7568# gnd 2.04fF
C1733 a_3825_8294# gnd 2.49fF
C1734 a_1808_7527# gnd 2.04fF
C1735 a_30333_8971# gnd 2.23fF
C1736 a_33098_9250# gnd 2.18fF
C1737 a_31069_8766# gnd 2.52fF
C1738 a_29065_8865# gnd 2.38fF
C1739 a_25358_9007# gnd 2.23fF
C1740 a_24009_8824# gnd 2.38fF
C1741 a_35389_9242# gnd 2.38fF
C1742 a_36126_9361# gnd 2.38fF
C1743 a_28123_9286# gnd 2.18fF
C1744 a_26094_8802# gnd 2.52fF
C1745 a_20302_8966# gnd 2.23fF
C1746 a_18906_9066# gnd 2.28fF
C1747 a_15204_8574# gnd 2.49fF
C1748 a_7832_7501# gnd 2.28fF
C1749 a_2776_7460# gnd 2.28fF
C1750 a_13850_9025# gnd 2.28fF
C1751 a_10148_8533# gnd 2.49fF
C1752 a_23067_9245# gnd 2.18fF
C1753 a_21038_8761# gnd 2.52fF
C1754 a_18910_8889# gnd 2.38fF
C1755 a_35389_9471# gnd 2.22fF
C1756 a_30333_9201# gnd 2.38fF
C1757 a_31070_9320# gnd 2.38fF
C1758 a_30333_9430# gnd 2.22fF
C1759 a_39097_9424# gnd 14.14fF
C1760 a_38158_9114# gnd 2.52fF
C1761 a_39093_9601# gnd 2.23fF
C1762 a_33102_9073# gnd 2.52fF
C1763 a_34037_9560# gnd 2.23fF
C1764 a_25358_9237# gnd 2.38fF
C1765 a_26095_9356# gnd 2.38fF
C1766 a_15203_9031# gnd 2.23fF
C1767 a_13854_8848# gnd 2.38fF
C1768 a_17968_9310# gnd 2.18fF
C1769 a_15939_8826# gnd 2.52fF
C1770 a_8875_9061# gnd 2.28fF
C1771 a_5173_8569# gnd 2.49fF
C1772 a_3819_9020# gnd 2.28fF
C1773 a_117_8528# gnd 2.49fF
C1774 a_10147_8990# gnd 2.23fF
C1775 a_12912_9269# gnd 2.18fF
C1776 a_10883_8785# gnd 2.52fF
C1777 a_8879_8884# gnd 2.38fF
C1778 a_5172_9026# gnd 2.23fF
C1779 a_3823_8843# gnd 2.38fF
C1780 a_25358_9466# gnd 2.22fF
C1781 a_20302_9196# gnd 2.38fF
C1782 a_21039_9315# gnd 2.38fF
C1783 a_20302_9425# gnd 2.22fF
C1784 a_34041_9383# gnd 2.98fF
C1785 a_29066_9419# gnd 2.82fF
C1786 a_28127_9109# gnd 2.52fF
C1787 a_29062_9596# gnd 2.23fF
C1788 a_23071_9068# gnd 2.52fF
C1789 a_24006_9555# gnd 2.23fF
C1790 a_15203_9261# gnd 2.38fF
C1791 a_15940_9380# gnd 2.38fF
C1792 a_7937_9305# gnd 2.18fF
C1793 a_5908_8821# gnd 2.52fF
C1794 a_116_8985# gnd 2.23fF
C1795 a_2881_9264# gnd 2.18fF
C1796 a_852_8780# gnd 2.52fF
C1797 a_15203_9490# gnd 2.22fF
C1798 a_10147_9220# gnd 2.38fF
C1799 a_10884_9339# gnd 2.38fF
C1800 a_10147_9449# gnd 2.22fF
C1801 a_24010_9378# gnd 2.98fF
C1802 a_18911_9443# gnd 2.97fF
C1803 a_17972_9133# gnd 2.52fF
C1804 a_18907_9620# gnd 2.23fF
C1805 a_12916_9092# gnd 2.52fF
C1806 a_13851_9579# gnd 2.23fF
C1807 a_5172_9256# gnd 2.38fF
C1808 a_5909_9375# gnd 2.38fF
C1809 a_5172_9485# gnd 2.22fF
C1810 a_116_9215# gnd 2.38fF
C1811 a_853_9334# gnd 2.38fF
C1812 a_13855_9402# gnd 2.98fF
C1813 a_8880_9438# gnd 2.82fF
C1814 a_7941_9128# gnd 2.52fF
C1815 a_8876_9615# gnd 2.23fF
C1816 a_2885_9087# gnd 2.52fF
C1817 a_3820_9574# gnd 2.23fF
C1818 a_3824_9397# gnd 2.98fF
C1819 vdd gnd 1895.70fF
