* SPICE3 file created from 9bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 vdd a_84977_12190# a_84769_12190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1 a_16310_7830# a_16567_7640# a_15995_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2 a_26960_4731# a_26851_4731# a_27059_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3 a_46686_11577# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_23738_10733# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5 a_76951_10731# a_76530_10731# a_76122_10415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_62003_11530# a_63096_12192# a_63051_12205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7 a_48518_4733# a_54071_446# a_54279_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_82181_4855# a_82273_3220# a_82228_3233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9 a_49843_3418# a_50100_3228# a_49800_4863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X10 a_76120_4407# a_76741_4723# a_76949_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X11 a_63048_10183# a_63052_9238# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X12 gnd a_51549_8556# a_51341_8556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 gnd d1 a_73220_3993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X14 a_18869_6969# a_19962_7631# a_19917_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X15 vdd d1 a_83928_3987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X16 a_28389_12214# a_28642_12201# a_28347_10692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 a_57607_11571# a_57394_11571# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 gnd d2 a_50102_9236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 a_11936_4046# a_11723_4046# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 a_45196_12255# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X21 a_37987_7651# a_38240_7638# a_37668_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X22 a_1436_2605# a_2276_3280# a_2484_3280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X23 gnd d0 a_52595_3991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 gnd a_8414_5515# a_8206_5515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X25 a_11724_13021# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X26 a_40539_4177# a_41636_3983# a_41587_4173# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_61997_5699# a_62254_5509# a_60550_6379# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X28 a_61997_5699# a_63094_5505# a_63045_5695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_39097_12208# a_40589_12962# a_40540_13152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_41588_13148# a_41845_12958# a_40540_13152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X31 a_69983_4731# a_69770_4731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X32 gnd a_84720_13827# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X33 gnd a_28643_9234# a_28435_9234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X34 a_63051_12973# a_63047_13150# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X35 a_44568_4731# a_45408_4727# a_45616_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X36 a_66240_5570# a_65819_5570# a_65411_5678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X37 a_66242_13025# a_65821_13025# a_65413_13133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X38 gnd a_20173_8546# a_19965_8546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 vdd d1 a_30088_2546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X40 a_68780_11575# a_68359_11575# a_68686_11694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X41 a_9205_7148# a_9462_6958# a_8157_7152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X42 a_63049_6197# a_63302_6184# a_62001_5522# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X43 vdd a_30088_3993# a_29880_3993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X44 a_35933_5561# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X45 gnd d0 a_9465_9231# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X46 a_79392_5680# a_79022_7006# a_77996_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X47 gnd a_63305_9993# a_63097_9993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_40544_11528# a_41637_12190# a_41588_12380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_3554_11577# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X50 a_45615_7694# a_46854_7014# a_47011_5688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 gnd a_52594_5511# a_52386_5511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_35890_7006# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X53 gnd d3 a_17635_10675# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_1436_3284# a_1015_3284# a_607_3363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X55 a_3510_4047# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X56 gnd a_84977_13637# a_83676_12975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X57 a_36105_13014# a_35892_13014# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X58 a_67290_12253# a_66869_12253# a_66242_12257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X59 a_67083_9286# a_66870_9286# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 gnd d0 a_31135_6188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X61 a_606_7382# a_606_7127# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X62 a_608_11688# a_609_11074# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X63 a_32987_7119# a_32987_6578# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X64 a_76741_4044# a_76528_4044# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 a_65820_4729# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X66 vdd d3 a_71732_10679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X67 a_12146_10054# a_11725_10054# a_11317_9621# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X68 a_11048_446# a_15673_4727# a_15995_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X69 a_2064_12255# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X70 a_84718_7819# a_84722_6963# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X71 a_77789_3272# a_77576_3272# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_33817_4723# a_33396_4723# a_32988_4407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 a_14431_4041# a_14218_4041# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X74 a_22282_10816# a_22903_10737# a_23111_10737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X75 vdd a_51549_8556# a_51341_8556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X76 a_45195_4727# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X77 a_37214_8596# a_37001_8596# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 a_65413_12336# a_65413_11941# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X79 vdd a_8417_10003# a_8209_10003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X80 vdd d2 a_50102_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X81 a_23948_7692# a_23735_7692# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X82 a_76740_7690# a_76527_7690# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X83 a_51290_4185# a_52387_3991# a_52342_4004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X84 a_60557_9243# a_62049_9997# a_62004_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X85 vdd a_8414_5515# a_8206_5515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X86 a_19916_10862# a_19920_10006# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X87 gnd a_6968_3228# a_6760_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X88 a_59442_7830# a_60557_4667# a_60512_4680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X89 a_6672_4686# a_6925_4673# a_5602_7836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_19915_13829# a_20172_13639# a_18871_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X91 a_58881_8598# a_58460_8598# a_57813_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 vdd a_28643_9234# a_28435_9234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X93 a_56115_7688# a_55902_7688# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X94 a_55275_5566# a_54854_5566# a_54446_5674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X95 a_33816_7011# a_33395_7011# a_32987_7119# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X96 a_40543_4000# a_40796_3987# a_39096_3233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X97 a_3973_5569# a_3552_5569# a_3874_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X98 vdd a_20173_8546# a_19965_8546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X99 a_72962_7150# a_74059_6956# a_74010_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X100 a_32988_4802# a_32988_4407# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X101 a_65822_9290# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 a_63045_6374# a_63302_6184# a_62001_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X103 a_23736_3278# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X104 a_19915_11703# a_19920_10685# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X105 a_55278_10733# a_56118_10729# a_56326_10729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X106 a_48518_4733# a_48097_4733# a_48173_8604# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X107 a_30878_5699# a_31135_5509# a_29830_5703# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X108 vdd d0 a_9465_9231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X109 gnd a_71773_3226# a_71565_3226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 a_81115_7828# a_82230_4665# a_82181_4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_84718_5693# a_84975_5503# a_83670_5697# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X112 a_22280_3617# a_22901_4050# a_23109_4050# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X113 a_74015_4002# a_74011_4179# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X114 vdd a_52594_5511# a_52386_5511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X115 a_25549_11575# a_25185_10053# a_24159_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X116 a_6711_3418# a_8207_2548# a_8158_2738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 a_68357_5567# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 gnd a_30087_5513# a_29879_5513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X119 a_30880_11707# a_31137_11517# a_29832_11711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X120 vdd d3 a_17635_10675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X121 gnd a_19122_5509# a_18914_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X122 a_75744_444# a_75531_444# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X123 a_76119_7769# a_76119_7374# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X124 a_11316_12332# a_11937_12253# a_12145_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X125 a_9212_10012# a_9465_9999# a_8160_10193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X126 a_33611_8605# a_33398_8605# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X127 a_54855_4725# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X128 a_55070_10733# a_54857_10733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X129 a_46857_10055# a_46644_10055# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_21685_433# a_32399_444# a_27059_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X131 a_23950_13700# a_23737_13700# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X132 a_72968_12981# a_74061_13643# a_74012_13833# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X133 a_45197_10735# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X134 gnd d4 a_70664_7644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 gnd d0 a_9463_2544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_84719_4173# a_84976_3983# a_83671_4177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X137 a_76950_13698# a_76529_13698# a_76121_13382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X138 vdd a_60809_12197# a_60601_12197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X139 gnd a_39308_10673# a_39100_10673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X140 a_43741_8721# a_43738_8033# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X141 a_66033_4050# a_65820_4050# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X142 a_23109_3282# a_22688_3282# a_22280_2966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X143 a_11317_11068# a_11317_10812# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X144 a_76949_3276# a_76528_3276# a_76120_2960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X145 gnd a_83929_12962# a_83721_12962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X146 a_16314_7653# a_17427_10675# a_17378_10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X147 a_82230_9241# a_82483_9228# a_82183_10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X148 vdd d0 a_63303_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X149 vdd d0 a_31137_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X150 a_52339_13156# a_52343_12211# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X151 vdd d0 a_63302_6952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X152 a_82227_6200# a_83719_6954# a_83670_7144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 a_43739_3363# a_44360_3284# a_44568_3284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 vdd a_83928_3987# a_83720_3987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X155 gnd d0 a_20171_4664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 a_6668_4863# a_6925_4673# a_5602_7836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X157 vdd d1 a_83927_5507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X158 a_51289_5705# a_52386_5511# a_52337_5701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X159 a_11935_5566# a_11722_5566# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X160 a_43740_13135# a_44361_13027# a_44569_13027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X161 a_60556_12210# a_62048_12964# a_61999_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X162 a_63047_13150# a_63304_12960# a_61999_13154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X163 a_19920_9238# a_20173_9225# a_18872_8563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X164 gnd a_50102_9236# a_49894_9236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X165 a_12144_3278# a_11723_3278# a_11315_3357# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X166 a_11723_4046# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X167 a_40538_5697# a_41635_5503# a_41586_5693# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X168 a_77998_13694# a_77577_13694# a_76950_13019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X169 a_8161_6975# a_9254_7637# a_9209_7650# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X170 a_18865_7146# a_19962_6952# a_19913_7142# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X171 a_2485_13702# a_2064_13702# a_1437_13027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X172 a_69770_4731# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X173 vdd d0 a_63304_12192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X174 a_70411_7657# a_71524_10679# a_71479_10692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X175 a_1228_4052# a_1015_4052# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X176 a_22279_8031# a_22279_7775# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X177 vdd a_71773_3226# a_71565_3226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X178 a_56325_12249# a_57564_13016# a_57721_11690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X179 a_83673_10185# a_83930_9995# a_82230_9241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X180 a_32987_6578# a_32987_6322# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X181 a_12144_3278# a_12984_3274# a_13192_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X182 a_81115_7828# a_82230_4665# a_82185_4678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X183 a_84720_12380# a_84724_11524# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X184 a_1227_7698# a_1014_7698# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X185 a_19914_4175# a_19918_3230# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X186 vdd a_30087_5513# a_29879_5513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X187 gnd a_9465_9231# a_9257_9231# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_22690_10058# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X189 a_83675_4000# a_84768_4662# a_84719_4852# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X190 a_2486_9288# a_2065_9288# a_1438_9292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X191 a_23737_13700# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X192 a_17420_12387# a_17677_12197# a_17382_10688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X193 a_55278_9286# a_54857_9286# a_54449_8970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X194 a_72968_12981# a_74061_13643# a_74016_13656# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X195 a_84721_10181# a_84978_9991# a_83673_10185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X196 vdd d4 a_70664_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X197 vdd d0 a_9463_2544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X198 gnd a_6927_10681# a_6719_10681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 gnd a_31135_6188# a_30927_6188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X200 a_55905_10729# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X201 a_45410_9288# a_45197_9288# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X202 a_43741_8721# a_44362_8613# a_44570_8613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X203 a_44146_6251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X204 a_22901_3282# a_22688_3282# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X205 a_76740_5564# a_76527_5564# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 vdd a_39308_10673# a_39100_10673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X207 a_33611_10052# a_33398_10052# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X208 a_12146_8607# a_11725_8607# a_11317_8715# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X209 a_67289_4725# a_66868_4725# a_66241_4729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X210 a_43009_401# a_42796_401# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X211 a_22282_10166# a_22282_9625# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X212 a_76951_10052# a_76530_10052# a_76122_9619# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X213 a_26506_8602# a_26293_8602# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 a_55067_6245# a_54854_6245# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X215 a_77576_3272# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X216 a_18867_13154# a_19964_12960# a_19919_12973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X217 a_1437_12259# a_1016_12259# a_608_12338# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X218 a_16314_7653# a_17427_10675# a_17382_10688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X219 a_74014_6969# a_74010_7146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X220 a_29831_4183# a_30928_3989# a_30883_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X221 vdd d0 a_20171_4664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X222 vdd a_50102_9236# a_49894_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X223 a_23735_7692# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X224 a_51289_5705# a_52386_5511# a_52341_5524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X225 a_74012_12386# a_74269_12196# a_72968_11534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X226 a_19916_9415# a_20173_9225# a_18872_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X227 a_51294_2561# a_51547_2548# a_49843_3418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X228 a_76120_3611# a_76741_4044# a_76949_4044# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X229 a_11317_8970# a_11938_9286# a_12146_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X230 a_15541_8598# a_15328_8598# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X231 a_11724_13700# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X232 a_33818_13019# a_34658_13694# a_34866_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X233 a_34656_7686# a_34443_7686# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X234 a_51296_10016# a_52389_10678# a_52344_10691# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X235 a_63051_13652# a_63047_13829# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X236 a_65819_6249# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X237 a_40542_5520# a_40795_5507# a_39091_6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X238 a_19919_12973# a_20172_12960# a_18867_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X239 a_44146_7019# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_28388_3239# a_28641_3226# a_28341_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X241 a_8159_13160# a_9256_12966# a_9211_12979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X242 a_11317_10417# a_11938_10733# a_12146_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X243 a_70191_4731# a_69770_4731# a_70092_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X244 gnd a_31137_13643# a_30929_13643# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X245 a_3876_11577# a_3512_10055# a_2486_9288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_19918_2551# a_20171_2538# a_18866_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 gnd a_41845_11511# a_41637_11511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 a_29832_13158# a_30929_12964# a_30884_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X249 vdd d0 a_9465_10678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X250 a_47008_11577# a_46644_10055# a_45618_10735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X251 vdd a_9465_9231# a_9257_9231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X252 a_22280_5064# a_22900_5570# a_23108_5570# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X253 a_79394_11688# a_79024_13014# a_77998_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X254 a_52339_12388# a_52596_12198# a_51295_11536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X255 a_83675_4000# a_84768_4662# a_84723_4675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X256 a_34443_6239# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X257 a_57563_4041# a_57350_4041# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X258 a_72962_7150# a_73219_6960# a_71519_6206# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X259 a_34864_7686# a_36103_7006# a_36260_5680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 vdd a_6927_10681# a_6719_10681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X261 vdd a_38240_7638# a_38032_7638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X262 a_52337_7827# a_52594_7637# a_51293_6975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X263 a_61999_11707# a_62256_11517# a_60552_12387# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X264 gnd d4 a_48991_7646# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X265 a_76120_2705# a_76122_2606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X266 a_72965_10191# a_74062_9997# a_74017_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X267 a_2484_3280# a_3723_4047# a_3874_5569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X268 a_84724_12971# a_84977_12958# a_83672_13152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X269 a_84724_11524# a_84720_11701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X270 gnd a_9463_2544# a_9255_2544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X271 a_23949_4725# a_23736_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_44567_7698# a_44146_7698# a_43738_7382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X273 a_39051_10863# a_39143_9228# a_39094_9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 a_24159_9286# a_23738_9286# a_23111_8611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 a_1014_6251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X276 a_66032_5570# a_65819_5570# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X277 a_52344_10012# a_52340_10189# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X278 a_55276_2599# a_54855_2599# a_54449_2608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X279 a_65820_4050# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X280 a_65412_4413# a_66033_4729# a_66241_4729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X281 a_43739_2968# a_43739_2713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X282 vdd d0 a_52596_12966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X283 gnd d0 a_41846_9223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X284 a_66868_3278# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X285 a_33817_4044# a_33396_4044# a_32988_3611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X286 a_22282_10166# a_22903_10058# a_23111_10058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X287 vdd a_63303_3217# a_63095_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X288 a_9212_8565# a_9208_8742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X289 a_25395_7012# a_25182_7012# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 vdd a_63302_6952# a_63094_6952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X291 vdd a_83927_5507# a_83719_5507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X292 a_82187_10686# a_82440_10673# a_81119_7651# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X293 a_11722_5566# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X294 a_54446_5929# a_54446_5674# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X295 a_66034_12257# a_65821_12257# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X296 a_13191_7688# a_12770_7688# a_12143_7013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X297 vdd d1 a_62256_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X298 a_33816_7690# a_33395_7690# a_32987_7769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X299 a_28384_3416# a_28641_3226# a_28341_4861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X300 a_77788_6239# a_77575_6239# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X301 a_14430_7008# a_14217_7008# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X302 a_1227_5572# a_1014_5572# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X303 a_84721_10181# a_84725_9236# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X304 a_54446_6324# a_55067_6245# a_55275_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X305 vdd a_31137_13643# a_30929_13643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X306 a_14683_11571# a_15541_8598# a_15749_8598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X307 a_63046_2728# a_54449_2608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X308 a_34867_9280# a_36106_10047# a_36257_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X309 a_25554_11694# a_25184_13020# a_24158_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 a_82187_10686# a_82274_12195# a_82229_12208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X311 vdd a_41845_11511# a_41637_11511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X312 a_11317_2608# a_11936_2599# a_12144_2599# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X313 a_14433_10049# a_14220_10049# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X314 a_59446_7653# a_59699_7640# a_59127_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X315 a_15886_4727# a_15673_4727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X316 vdd a_40797_12962# a_40589_12962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X317 a_76122_10810# a_76743_10731# a_76951_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 a_57716_11571# a_57352_10049# a_56326_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X319 vdd d0 a_41845_13637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X320 a_1436_4052# a_2276_4727# a_2484_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X321 a_45196_13702# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X322 vdd d4 a_48991_7646# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X323 vdd a_9463_2544# a_9255_2544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X324 a_6715_3241# a_6968_3228# a_6668_4863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 vdd d1 a_51549_10003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X326 a_66241_3282# a_65820_3282# a_65412_3361# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X327 a_11316_13129# a_11316_12588# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X328 a_23951_9286# a_23738_9286# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X329 a_65414_8719# a_65411_8031# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X330 a_54855_4046# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X331 a_55070_10054# a_54857_10054# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X332 gnd d1 a_51547_3995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X333 a_72964_13158# a_74061_12964# a_74012_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X334 a_63049_7644# a_63302_7631# a_62001_6969# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X335 a_49800_4863# a_49892_3228# a_49843_3418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_11724_11574# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 gnd a_73222_10001# a_73014_10001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X338 vdd d0 a_41846_9223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X339 a_26293_8602# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 vdd d1 a_19122_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X341 a_74011_4179# a_74268_3989# a_72963_4183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X342 a_49849_9249# a_51341_10003# a_51292_10193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X343 a_29830_5703# a_30927_5509# a_30882_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X344 a_82183_10863# a_82440_10673# a_81119_7651# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X345 a_76120_5058# a_76740_5564# a_76948_5564# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X346 a_66242_11578# a_65821_11578# a_65414_11072# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X347 a_2486_9288# a_3725_10055# a_3876_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X348 a_17418_6379# a_17675_6189# a_17380_4680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X349 a_55275_5566# a_56115_6241# a_56323_6241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X350 a_49847_3241# a_50100_3228# a_49800_4863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X351 gnd d0 a_20171_3985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X352 gnd d0 a_31135_7635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X353 a_12145_11574# a_12985_12249# a_13193_12249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X354 a_22687_7017# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_23108_6249# a_22687_6249# a_22279_6328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X356 a_76119_5672# a_76120_5058# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X357 gnd d0 a_41844_2536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X358 a_8162_4008# a_8415_3995# a_6715_3241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X359 a_44148_12259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X360 a_59442_7830# a_59699_7640# a_59127_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X361 a_2064_13702# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X362 vdd a_31138_9997# a_30930_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X363 a_19915_12382# a_19919_11526# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X364 a_65412_3361# a_65412_2966# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X365 a_23108_6249# a_23948_6245# a_24156_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X366 a_55277_13021# a_54856_13021# a_54448_13129# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X367 a_1227_7019# a_1014_7019# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X368 a_62002_2555# a_63095_3217# a_63050_3230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X369 a_9210_3236# a_9463_3223# a_8162_2561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X370 a_11317_10417# a_11317_10162# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X371 a_79238_10047# a_79025_10047# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 a_19916_8736# a_19917_7644# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X373 a_61997_7146# a_63094_6952# a_63049_6965# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X374 a_44147_3284# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 gnd a_19125_9997# a_18917_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X376 a_57350_4041# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X377 a_83671_4177# a_83928_3987# a_82228_3233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X378 a_55068_3278# a_54855_3278# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X379 a_11936_3278# a_11723_3278# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X380 a_83671_4177# a_84768_3983# a_84719_4173# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X381 gnd d0 a_20172_12192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X382 a_35893_10047# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X383 a_32990_8968# a_32990_8713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X384 a_51295_12983# a_51548_12970# a_49848_12216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X385 a_46644_10055# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X386 a_63045_7821# a_63302_7631# a_62001_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X387 a_23736_4725# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 a_44568_2605# a_44147_2605# a_43741_2614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 a_22282_10816# a_22282_10421# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X390 a_25547_5567# a_25183_4045# a_24157_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X391 a_34657_4719# a_34444_4719# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 gnd a_73221_11521# a_73013_11521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X393 a_74014_7648# a_74010_7825# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X394 a_40544_12975# a_41637_13637# a_41592_13650# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X395 gnd d3 a_71732_10679# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X396 a_33816_5564# a_33395_5564# a_32988_5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 gnd a_41846_9223# a_41638_9223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X398 a_79394_11688# a_79280_11569# a_79488_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X399 a_84722_6195# a_84718_6372# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X400 a_25182_7012# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 vout a_42796_401# a_43118_401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X402 vdd d0 a_31135_7635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X403 a_79022_7006# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X404 a_11316_13779# a_11937_13700# a_12145_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X405 vdd d1 a_83930_8548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X406 vdd d0 a_41844_2536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X407 a_59442_7830# a_60557_4667# a_60508_4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X408 a_77575_6239# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X409 a_19919_13652# a_20172_13639# a_18871_12977# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 a_77999_10727# a_77578_10727# a_76951_10052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X411 gnd d0 a_74267_6188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X412 a_11314_7121# a_11935_7013# a_12143_7013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X413 a_47013_11696# a_46643_13022# a_45617_12255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X414 a_11316_12588# a_11316_12332# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X415 gnd d1 a_8416_11523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X416 a_44149_8613# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_24158_13700# a_23737_13700# a_23110_13704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X418 a_76950_12251# a_77790_12247# a_77998_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X419 a_11317_9621# a_11938_10054# a_12146_10054# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X420 a_54180_446# a_58805_4727# a_59127_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X421 a_68359_11575# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X422 gnd d1 a_40798_9995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X423 a_606_5935# a_1227_6251# a_1435_6251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X424 a_76741_3276# a_76528_3276# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X425 gnd a_31137_12964# a_30929_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X426 a_41592_12971# a_41588_13148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X427 gnd d3 a_50059_10681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_83677_8561# a_84770_9223# a_84721_9413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X429 a_11938_8607# a_11725_8607# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X430 a_76949_4723# a_76528_4723# a_76120_4407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 a_15673_4727# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X432 a_76121_13777# a_76742_13698# a_76950_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_56117_12249# a_55904_12249# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X434 a_9206_3413# a_9463_3223# a_8162_2561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X435 a_72964_13158# a_73221_12968# a_71521_12214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X436 a_43739_4810# a_44360_4731# a_44568_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X437 a_47011_5688# a_46897_5569# a_47105_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X438 a_57721_11690# a_57607_11571# a_57815_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X439 a_3512_10055# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X440 a_76122_9363# a_76743_9284# a_76951_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 a_56116_3274# a_55903_3274# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X442 a_12144_4725# a_11723_4725# a_11315_4804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X443 a_33818_13698# a_33397_13698# a_32989_13777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X444 a_12772_12249# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X445 a_5178_4733# a_4965_4733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X446 a_52338_2734# a_43741_2614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X447 a_43118_401# a_64495_433# a_54279_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X448 a_1230_10739# a_1017_10739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X449 a_32987_7769# a_33608_7690# a_33816_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X450 a_64495_433# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X451 a_32988_5058# a_32988_4802# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X452 vdd d2 a_82482_12195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X453 a_30884_11530# a_31137_11517# a_29832_11711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X454 a_67291_9286# a_66870_9286# a_66243_9290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X455 a_29835_4006# a_30088_3993# a_28388_3239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X456 a_68529_13020# a_68316_13020# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X457 a_76948_7011# a_76527_7011# a_76119_7119# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X458 a_54854_5566# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X459 a_63051_11526# a_63047_11703# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X460 a_65412_2966# a_65412_2711# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X461 gnd a_51547_3995# a_51339_3995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X462 a_11315_2962# a_11315_2707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X463 a_12144_4725# a_12984_4721# a_13192_4721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X464 vdd d0 a_74269_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X465 a_40544_11528# a_40797_11515# a_39093_12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X466 vdd a_73221_11521# a_73013_11521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X467 a_606_7127# a_1227_7019# a_1435_7019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_76529_12251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X469 a_14262_11571# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X470 a_74010_5699# a_74267_5509# a_72962_5703# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X471 vdd a_41846_9223# a_41638_9223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X472 vdd a_19122_6956# a_18914_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X473 a_52341_6971# a_52337_7148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X474 vdd a_20171_2538# a_19963_2538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X475 gnd a_73220_2546# a_73012_2546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 a_37422_8596# a_37001_8596# a_36356_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X477 vdd a_83930_9995# a_83722_9995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X478 a_76119_8025# a_76119_7769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X479 gnd d1 a_62254_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 vdd d2 a_39348_6187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X481 a_65412_3617# a_66033_4050# a_66241_4050# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X482 a_45615_6247# a_45194_6247# a_44567_5572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X483 gnd d0 a_20170_5505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X484 a_34866_13694# a_36105_13014# a_36262_11688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X485 gnd d0 a_63303_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X486 a_32990_11066# a_32990_10810# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X487 a_65822_10737# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X488 a_76743_8605# a_76530_8605# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X489 gnd a_31135_7635# a_30927_7635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X490 a_80478_4725# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X491 a_18867_13154# a_19124_12964# a_17424_12210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X492 a_14432_13016# a_14219_13016# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X493 vdd d1 a_8416_11523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X494 a_44570_8613# a_44149_8613# a_43741_8721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X495 a_67083_10733# a_66870_10733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 gnd a_41844_2536# a_41636_2536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X497 a_28389_12214# a_29881_12968# a_29836_12981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X498 a_8161_6975# a_9254_7637# a_9205_7827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X499 a_70411_7657# a_71524_10679# a_71475_10869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X500 a_55067_7692# a_54854_7692# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X501 a_76529_13019# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X502 vdd d3 a_50059_10681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X503 a_83677_8561# a_84770_9223# a_84725_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X504 a_70411_7657# a_70664_7644# a_70092_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X505 a_84723_3996# a_84719_4173# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X506 a_1437_13706# a_1016_13706# a_608_13785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X507 a_76951_9284# a_76530_9284# a_76122_9363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X508 vdd d1 a_73219_6960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X509 a_76743_10731# a_76530_10731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X510 vdd a_62257_9997# a_62049_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X511 a_45197_9288# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X512 a_3509_7014# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X513 a_40538_7144# a_41635_6950# a_41590_6963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X514 vdd d0 a_52594_6958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X515 a_22688_3282# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X516 a_76122_10160# a_76743_10052# a_76951_10052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X517 a_41588_11701# a_41593_10683# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X518 a_57352_10049# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X519 a_83670_5697# a_83927_5507# a_82223_6377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X520 a_83670_5697# a_84767_5503# a_84718_5693# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_76122_10160# a_76122_9619# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X522 a_11723_3278# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X523 a_13193_13696# a_12772_13696# a_12145_13021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X524 a_43740_11943# a_44361_12259# a_44569_12259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X525 a_33608_6243# a_33395_6243# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X526 a_77577_12247# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_12983_7688# a_12770_7688# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_40540_11705# a_40797_11515# a_39093_12385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X529 a_15328_8598# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X530 a_76120_2705# a_76741_2597# a_76949_2597# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X531 a_55276_3278# a_56116_3274# a_56324_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X532 vdd a_73220_2546# a_73012_2546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X533 a_22280_2966# a_22901_3282# a_23109_3282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X534 a_33819_8605# a_34659_9280# a_34867_9280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X535 a_63049_6965# a_63302_6952# a_61997_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X536 a_43739_3619# a_43739_3363# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X537 a_2485_13702# a_3724_13022# a_3881_11696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 a_76951_10052# a_77791_10727# a_77999_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X539 a_71517_12391# a_71774_12201# a_71479_10692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X540 vdd d2 a_71772_6193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X541 a_33816_7690# a_34656_7686# a_34864_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 a_56118_10729# a_55905_10729# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X543 a_2484_3280# a_2063_3280# a_1436_2605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X544 a_52337_5701# a_52342_4683# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X545 a_57714_5563# a_57605_5563# a_57813_5563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X546 vdd a_31135_7635# a_30927_7635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X547 a_36260_5680# a_35890_7006# a_34864_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X548 a_30880_13154# a_30884_12209# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X549 gnd a_74270_10676# a_74062_10676# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X550 a_1017_9292# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X551 a_29833_8744# a_30930_8550# a_30881_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 vdd a_41844_2536# a_41636_2536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X553 a_19916_10183# a_20173_9993# a_18868_10187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X554 a_54857_9286# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X555 gnd d0 a_31135_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X556 gnd a_74267_6188# a_74059_6188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_63046_3407# a_63050_2551# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X558 a_51296_10016# a_52389_10678# a_52340_10868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 a_70407_7834# a_70664_7644# a_70092_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X560 a_66033_3282# a_65820_3282# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X561 a_32721_444# a_37346_4725# a_37668_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X562 gnd a_28598_4671# a_28390_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_33818_11572# a_33397_11572# a_32990_11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X564 a_77791_9280# a_77578_9280# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X565 gnd a_17635_10675# a_17427_10675# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X566 a_11725_8607# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X567 a_69638_8602# a_69425_8602# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X568 a_66868_4725# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X569 a_25552_5686# a_25438_5567# a_25646_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 gnd d0 a_84978_10670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X571 a_34657_3272# a_34444_3272# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X572 a_71520_3239# a_73012_3993# a_72967_4006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X573 a_55277_13700# a_54856_13700# a_54448_13779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X574 a_35892_13014# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X575 gnd a_62256_12964# a_62048_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X576 a_9210_4004# a_9206_4181# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X577 gnd d0 a_9465_10678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X578 a_40538_7144# a_40795_6954# a_39095_6200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X579 a_66034_13704# a_65821_13704# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X580 a_54449_8970# a_55070_9286# a_55278_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X581 a_77788_7686# a_77575_7686# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X582 a_72966_5526# a_74059_6188# a_74014_6201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X583 vdd a_71732_10679# a_71524_10679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X584 vdd a_50100_3228# a_49892_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X585 a_41587_2726# a_32990_2606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X586 a_22902_11578# a_22689_11578# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X587 a_606_7777# a_606_7382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X588 a_62003_11530# a_62256_11517# a_60552_12387# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X589 gnd a_38240_7638# a_38032_7638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X590 a_52341_7650# a_52594_7637# a_51293_6975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X591 a_23111_10737# a_23951_10733# a_24159_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X592 gnd d2 a_50099_6195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X593 vdd d2 a_60807_6189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X594 vdd d1 a_8415_2548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X595 gnd a_63304_12192# a_63096_12192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X596 a_44568_2605# a_45408_3280# a_45616_3280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X597 a_44362_9292# a_44149_9292# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X598 a_65412_5064# a_66032_5570# a_66240_5570# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X599 gnd a_62254_6956# a_62046_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X600 vdd a_39348_6187# a_39140_6187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X601 a_32990_10810# a_33611_10731# a_33819_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X602 a_11938_10733# a_11725_10733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X603 vdd a_74270_10676# a_74062_10676# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X604 a_29833_8744# a_30930_8550# a_30885_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X605 gnd a_63303_3217# a_63095_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 a_607_3363# a_1228_3284# a_1436_3284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X607 a_11316_13129# a_11937_13021# a_12145_13021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X608 a_1437_11580# a_1016_11580# a_609_11074# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X609 a_76530_8605# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X610 a_26960_4731# a_27324_7644# a_27275_7834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X611 a_54446_5674# a_54447_5060# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X612 a_68681_11575# a_68317_10053# a_67291_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X613 gnd d0 a_9462_6190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X614 vdd a_28598_4671# a_28390_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X615 a_12145_12253# a_11724_12253# a_11316_11937# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X616 a_41592_13650# a_41588_13827# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X617 a_3511_13022# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X618 vdd a_17635_10675# a_17427_10675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X619 a_77578_10727# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X620 vdd d0 a_84978_10670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X621 a_76742_13698# a_76529_13698# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X622 a_23109_4050# a_22688_4050# a_22280_3617# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X623 a_1015_2605# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X624 a_54855_2599# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X625 a_76949_4044# a_76528_4044# a_76120_3611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 gnd d0 a_84978_9223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_46642_4047# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X628 a_19913_5695# a_19918_4677# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X629 a_68527_7012# a_68314_7012# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X630 a_33817_3276# a_33396_3276# a_32988_3355# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X631 a_43739_4160# a_44360_4052# a_44568_4052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X632 a_71515_6383# a_73011_5513# a_72962_5703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X633 a_41593_9236# a_41846_9223# a_40545_8561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_14582_5563# a_14218_4041# a_13192_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X635 a_33818_13019# a_33397_13019# a_32989_13127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X636 vdd a_84977_12958# a_84769_12958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X637 a_12144_4046# a_11723_4046# a_11315_4154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X638 a_12145_13021# a_12985_13696# a_13193_13696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X639 gnd d0 a_41845_13637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X640 a_23108_7696# a_22687_7696# a_22279_7775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X641 a_56323_7688# a_55902_7688# a_55275_7013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X642 a_63050_2551# a_63046_2728# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X643 vdd a_9464_12966# a_9256_12966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X644 a_61999_13154# a_63096_12960# a_63051_12973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X645 a_1230_10060# a_1017_10060# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X646 a_32990_9619# a_32990_9363# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X647 a_12770_7688# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X648 a_76948_7690# a_76527_7690# a_76119_7769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X649 a_33395_6243# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X650 a_44148_13706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X651 a_43738_7382# a_44359_7698# a_44567_7698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X652 a_54279_446# a_64708_433# a_43118_401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_23111_8611# a_23951_9286# a_24159_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X654 a_2275_7694# a_2062_7694# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X655 a_54449_2608# a_55068_2599# a_55276_2599# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X656 a_52341_7650# a_52337_7827# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X657 a_609_8721# a_1230_8613# a_1438_8613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X658 a_32989_13127# a_32989_12586# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X659 gnd a_20172_11513# a_19964_11513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X660 a_59018_4727# a_58805_4727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X661 a_25438_5567# a_25225_5567# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 a_34866_12247# a_34445_12247# a_33818_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X663 a_44147_4731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_30885_10010# a_30881_10187# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X665 gnd d1 a_62257_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X666 a_9211_12211# a_9464_12198# a_8163_11536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X667 a_45617_12255# a_45196_12255# a_44569_11580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X668 a_82185_4678# a_82438_4665# a_81115_7828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X669 a_26960_4731# a_27324_7644# a_27279_7657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X670 a_55068_4725# a_54855_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 a_11936_4725# a_11723_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X672 a_22281_12336# a_22281_11941# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X673 a_5041_8604# a_4620_8604# a_3973_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X674 a_74017_8563# a_74270_8550# a_72965_8744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_44359_5572# a_44146_5572# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X676 a_32988_4407# a_32988_4152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X677 gnd d1 a_30089_11521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X678 a_65822_10058# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 gnd a_31135_6956# a_30927_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X680 a_44360_2605# a_44147_2605# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X681 a_55277_11574# a_54856_11574# a_54449_11068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X682 a_84723_4675# a_84719_4852# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X683 a_33819_8605# a_33398_8605# a_32990_8713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X684 a_65820_3282# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X685 a_8157_7152# a_9254_6958# a_9205_7148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X686 vdd d0 a_84978_9223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X687 a_55067_7013# a_54854_7013# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X688 a_60555_3235# a_62047_3989# a_61998_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 a_1437_13027# a_1016_13027# a_608_13135# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X690 a_57351_13016# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X691 a_69425_8602# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X692 a_71515_6383# a_73011_5513# a_72966_5526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X693 a_3975_11577# a_3554_11577# a_3881_11696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X694 a_76743_10052# a_76530_10052# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X695 a_41589_9413# a_41846_9223# a_40545_8561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X696 a_10939_446# a_10726_446# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X697 a_65414_11072# a_66034_11578# a_66242_11578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X698 a_76122_10810# a_76122_10415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X699 a_77575_7686# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X700 a_62002_2555# a_63095_3217# a_63046_3407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_44361_11580# a_44148_11580# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X702 gnd d0 a_74267_7635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 a_32990_10415# a_32990_10160# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X704 a_51292_10193# a_51549_10003# a_49849_9249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X705 a_65819_7017# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X706 a_49806_10694# a_49893_12203# a_49848_12216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X707 gnd d0 a_84976_2536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 a_3874_5569# a_3765_5569# a_3973_5569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X709 a_82227_6200# a_82480_6187# a_82185_4678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X710 vdd a_82482_12195# a_82274_12195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X711 a_22687_6249# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X712 a_65412_3617# a_65412_3361# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X713 gnd d4 a_5859_7646# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 a_18869_6969# a_19122_6956# a_17422_6202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X715 a_2485_12255# a_2064_12255# a_1437_12259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X716 a_19917_6197# a_20170_6184# a_18869_5522# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X717 vdd a_60807_6189# a_60599_6189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X718 a_607_2713# a_609_2614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X719 a_41591_2549# a_41844_2536# a_40539_2730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X720 a_36255_5561# a_35891_4039# a_34865_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X721 a_76741_4723# a_76528_4723# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X722 vdd a_20172_11513# a_19964_11513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X723 a_12146_10733# a_11725_10733# a_11317_10812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X724 vdd a_8415_2548# a_8207_2548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X725 a_1435_7698# a_1014_7698# a_606_7382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X726 a_22279_7125# a_22279_6584# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X727 a_54449_10812# a_55070_10733# a_55278_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 a_1017_10060# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X729 vdd d1 a_62257_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X730 a_74010_7825# a_74014_6969# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X731 a_66240_6249# a_67080_6245# a_67288_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X732 a_56116_4721# a_55903_4721# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X733 a_12772_13696# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X734 a_32989_13777# a_33610_13698# a_33818_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X735 a_82181_4855# a_82438_4665# a_81115_7828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X736 a_40544_12975# a_41637_13637# a_41588_13827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X737 a_71475_10869# a_71567_9234# a_71518_9424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 vdd d0 a_20172_13639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X739 a_1438_9292# a_2278_9288# a_2486_9288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 a_74013_8740# a_74270_8550# a_72965_8744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X741 a_84720_12380# a_84977_12190# a_83676_11528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X742 a_65411_8031# a_66035_8611# a_66243_8611# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X743 a_19915_13829# a_19919_12973# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X744 a_67290_13700# a_66869_13700# a_66242_13704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X745 a_9207_13156# a_9211_12211# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X746 vdd d1 a_30089_11521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X747 vdd d2 a_39351_9228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X748 a_64817_433# a_75531_444# a_70191_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X749 a_33610_12251# a_33397_12251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X750 gnd d1 a_83930_9995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_8164_10016# a_8417_10003# a_6717_9249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X752 gnd a_74270_9997# a_74062_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X753 a_3879_5688# a_3509_7014# a_2483_6247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X754 gnd a_9462_6190# a_9254_6190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X755 a_23737_12253# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X756 a_18868_8740# a_19965_8546# a_19916_8736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X757 gnd d0 a_31138_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X758 a_76950_12251# a_76529_12251# a_76121_11935# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X759 gnd d1 a_83930_8548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X760 a_51292_10193# a_52389_9999# a_52340_10189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X761 a_2483_6247# a_2062_6247# a_1435_6251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X762 a_44570_10739# a_44149_10739# a_43741_10818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X763 a_68679_5567# a_68315_4045# a_67289_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X764 a_77789_4719# a_77576_4719# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X765 a_23108_5570# a_22687_5570# a_22280_5064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X766 a_45618_9288# a_45197_9288# a_44570_9292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X767 gnd d1 a_40796_2540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X768 a_76948_5564# a_76527_5564# a_76120_5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X769 a_32989_12586# a_32989_12330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X770 a_33397_11572# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X771 a_34867_9280# a_34446_9280# a_33819_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X772 gnd a_84978_9223# a_84770_9223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 vdd d0 a_31137_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X774 a_47008_11577# a_46899_11577# a_47107_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X775 a_79278_5561# a_79065_5561# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_41588_12380# a_41592_11524# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X777 a_44148_11580# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X778 gnd d0 a_84978_9991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X779 a_68314_7012# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X780 a_43738_5680# a_44359_5572# a_44567_5572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X781 a_34864_7686# a_34443_7686# a_33816_7011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_19918_3230# a_19914_3407# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X783 a_12143_5566# a_11722_5566# a_11314_5674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X784 gnd d0 a_9465_9999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X785 vdd d0 a_74267_7635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X786 a_66034_13025# a_65821_13025# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X787 vdd d0 a_41846_9991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X788 a_33610_13019# a_33397_13019# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 vdd d0 a_84976_2536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X790 a_13194_10729# a_12773_10729# a_12146_10054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X791 a_45618_10735# a_45197_10735# a_44570_10739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X792 a_15749_8598# a_15328_8598# a_14683_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X793 vdd d4 a_5859_7646# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X794 a_54446_7121# a_55067_7013# a_55275_7013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 vdd a_52596_12966# a_52388_12966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X796 a_83673_8738# a_83930_8548# a_82226_9418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X797 a_19913_6374# a_20170_6184# a_18869_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X798 a_41587_2726# a_41844_2536# a_40539_2730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X799 vdd d3 a_17633_4667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X800 a_11314_5929# a_11935_6245# a_12143_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X801 a_2062_7694# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X802 a_52341_6971# a_52594_6958# a_51289_7152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X803 a_33611_9284# a_33398_9284# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X804 gnd a_28641_3226# a_28433_3226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X805 a_19920_10685# a_19916_10862# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X806 a_69846_8602# a_69983_4731# a_70191_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 a_58805_4727# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X808 a_25225_5567# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X809 a_71475_10869# a_71567_9234# a_71522_9247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X810 gnd a_20171_2538# a_19963_2538# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X811 vdd d0 a_63304_12960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X812 gnd a_62257_8550# a_62049_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 gnd d2 a_60809_12197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X814 a_32990_10160# a_33611_10052# a_33819_10052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X815 gnd d2 a_60810_9230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X816 a_52337_6380# a_52341_5524# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X817 a_63051_13652# a_65413_13783# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X818 a_43740_13390# a_44361_13706# a_44569_13706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X819 a_11723_4725# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X820 vdd d1 a_51546_6962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X821 a_11938_10054# a_11725_10054# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X822 a_18868_8740# a_19965_8546# a_19920_8559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X823 vdd d0 a_31138_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X824 a_66870_9286# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X825 a_1228_4731# a_1015_4731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X826 a_55276_4725# a_56116_4721# a_56324_4721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X827 a_54857_10733# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X828 a_68317_10053# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X829 vdd d1 a_40796_2540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X830 a_52338_4181# a_52342_3236# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X831 a_606_5680# a_607_5066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X832 a_60550_6379# a_62046_5509# a_61997_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 a_22281_12336# a_22902_12257# a_23110_12257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X834 gnd a_51548_11523# a_51340_11523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X835 a_49806_10694# a_50059_10681# a_48738_7659# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X836 vdd a_84978_9223# a_84770_9223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X837 a_23949_3278# a_23736_3278# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X838 vdd d1 a_19123_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X839 a_23109_4729# a_22688_4729# a_22280_4413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X840 a_28383_6383# a_29879_5513# a_29830_5703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 a_39095_6200# a_40587_6954# a_40538_7144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X842 a_22279_6584# a_22279_6328# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X843 vdd d0 a_20171_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X844 vdd d0 a_20170_6952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X845 a_63045_7142# a_63049_6197# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X846 a_34658_13694# a_34445_13694# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X847 a_30878_5699# a_30883_4681# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X848 a_37001_8596# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X849 a_47105_5569# a_47965_8604# a_48173_8604# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X850 a_82230_9241# a_83722_9995# a_83673_10185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 a_39053_4678# a_39140_6187# a_39091_6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X852 gnd d0 a_52595_3223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 a_40543_2553# a_41636_3215# a_41587_3405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X854 a_29833_10191# a_30090_10001# a_28390_9247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X855 a_8157_7152# a_8414_6962# a_6714_6208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X856 gnd a_74267_7635# a_74059_7635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 gnd d0 a_41845_12958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_23108_7017# a_22687_7017# a_22279_7125# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X859 gnd d0 a_41843_6182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 a_41587_3405# a_41591_2549# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X861 a_8159_11713# a_9256_11519# a_9211_11532# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X862 gnd a_84976_2536# a_84768_2536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 a_12143_7692# a_12983_7688# a_13191_7688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X864 a_44148_13027# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X865 a_72969_8567# a_74062_9229# a_74017_9242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X866 a_43738_6586# a_44359_7019# a_44567_7019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X867 vdd a_28641_3226# a_28433_3226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X868 a_6716_12216# a_8208_12970# a_8163_12983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X869 a_74012_13154# a_74269_12964# a_72964_13158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X870 a_55277_12253# a_56117_12249# a_56325_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 a_14587_5682# a_14217_7008# a_13191_7688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X872 a_46686_11577# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X873 a_29832_11711# a_30929_11517# a_30884_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X874 a_41592_11524# a_41588_11701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X875 a_76951_10731# a_76530_10731# a_76122_10810# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X876 a_609_10168# a_1230_10060# a_1438_10060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X877 a_1436_2605# a_1015_2605# a_609_2614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X878 vdd a_62257_8550# a_62049_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X879 a_54180_446# a_54071_446# a_54279_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X880 vdd d2 a_60810_9230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X881 a_83670_7144# a_84767_6950# a_84722_6963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X882 a_9212_10012# a_9208_10189# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X883 a_40541_10185# a_41638_9991# a_41593_10004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X884 a_12146_9286# a_11725_9286# a_11317_8970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X885 a_22900_7696# a_22687_7696# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X886 a_44147_4052# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 a_67290_12253# a_68529_13020# a_68686_11694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X888 a_72963_2736# a_74060_2542# a_74011_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X889 a_55068_4046# a_54855_4046# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X890 gnd d0 a_20172_12960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 a_60552_12387# a_60809_12197# a_60514_10688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X892 a_57607_11571# a_57394_11571# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X893 a_11936_4046# a_11723_4046# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X894 a_45196_12255# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X895 a_49847_3241# a_51339_3995# a_51294_4008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X896 gnd a_31138_8550# a_30930_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X897 a_44146_7698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X898 a_44567_6251# a_44146_6251# a_43738_5935# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 a_33609_2597# a_33396_2597# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X900 a_34444_3272# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X901 a_83676_12975# a_83929_12962# a_82229_12208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X902 vdd a_51548_11523# a_51340_11523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X903 a_49802_10871# a_50059_10681# a_48738_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X904 a_79025_10047# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X905 a_84725_9236# a_84721_9413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X906 a_28383_6383# a_29879_5513# a_29834_5526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X907 a_8160_8746# a_9257_8552# a_9208_8742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 a_65412_2966# a_66033_3282# a_66241_3282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X909 a_77576_4719# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 a_44568_4052# a_45408_4727# a_45616_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X911 a_76951_8605# a_77791_9280# a_77999_9280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X912 gnd a_40796_2540# a_40588_2540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X913 a_52341_5524# a_52337_5701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X914 vdd d0 a_52596_11519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X915 a_60514_10688# a_60601_12197# a_60552_12387# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X916 a_19913_6374# a_19917_5518# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X917 a_25184_13020# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X918 a_76948_7690# a_77788_7686# a_77996_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X919 vdd d0 a_52595_3223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X920 a_40543_2553# a_41636_3215# a_41591_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X921 a_79065_5561# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 a_35933_5561# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X923 vdd a_74267_7635# a_74059_7635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X924 a_79392_5680# a_79022_7006# a_77996_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X925 a_13191_6241# a_12770_6241# a_12143_5566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X926 a_71515_6383# a_71772_6193# a_71477_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X927 a_607_4810# a_1228_4731# a_1436_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X928 vdd d1 a_62256_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X929 a_13194_10729# a_14433_10049# a_14584_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X930 a_35890_7006# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X931 a_45615_6247# a_46854_7014# a_47011_5688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X932 vdd d0 a_41843_6182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X933 a_12145_13700# a_11724_13700# a_11316_13384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X934 vdd a_84976_2536# a_84768_2536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X935 gnd d0 a_74267_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X936 a_45410_10735# a_45197_10735# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X937 gnd a_71732_10679# a_71524_10679# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X938 gnd a_50100_3228# a_49892_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X939 a_27059_4731# a_26638_4731# a_26960_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X940 a_36105_13014# a_35892_13014# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X941 a_22689_12257# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 vdd d3 a_28600_10679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X943 a_18872_8563# a_19125_8550# a_17421_9420# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X944 a_82224_3410# a_83720_2540# a_83671_2730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_84723_2549# a_84719_2726# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X946 a_43740_11688# a_44361_11580# a_44569_11580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X947 a_67080_7692# a_66867_7692# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X948 a_29837_10014# a_30930_10676# a_30881_10866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X949 a_76741_4044# a_76528_4044# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X950 a_11048_446# a_15673_4727# a_15749_8598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X951 a_1017_10739# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_12146_10054# a_11725_10054# a_11317_10162# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X953 gnd d1 a_8415_2548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X954 a_9206_4181# a_9463_3991# a_8158_4185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X955 a_68684_5686# a_68570_5567# a_68778_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X956 a_52343_12979# a_52339_13156# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X957 a_77789_3272# a_77576_3272# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X958 a_14431_4041# a_14218_4041# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X959 a_33817_4723# a_33396_4723# a_32988_4802# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X960 a_22282_10421# a_22903_10737# a_23111_10737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X961 gnd d3 a_82440_10673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X962 a_54449_10162# a_55070_10054# a_55278_10054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X963 a_29830_7150# a_30087_6960# a_28387_6206# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X964 a_6674_10694# a_6927_10681# a_5606_7659# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_84721_10860# a_84725_10004# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X966 a_33398_9284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X967 a_40540_13152# a_41637_12958# a_41588_13148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_72963_2736# a_74060_2542# a_74015_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X969 a_606_8033# a_606_7777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X970 vdd a_51546_6962# a_51338_6962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X971 vdd a_31138_8550# a_30930_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X972 a_55904_12249# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 vdd a_63304_13639# a_63096_13639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X974 a_49842_6385# a_51338_5515# a_51289_5705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_74013_10187# a_74017_9242# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X976 a_8160_8746# a_9257_8552# a_9212_8565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X977 a_12144_2599# a_11723_2599# a_11317_2608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X978 a_3973_5569# a_3552_5569# a_3879_5688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X979 vdd a_40796_2540# a_40588_2540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X980 a_17422_6202# a_18914_6956# a_18865_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X981 a_70191_4731# a_75744_444# a_64817_433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_23736_3278# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X983 a_19918_3998# a_19914_4175# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X984 vdd d1 a_19122_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X985 a_44570_10060# a_44149_10060# a_43741_10168# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X986 gnd d1 a_30087_6960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X987 a_60550_6379# a_60807_6189# a_60512_4680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X988 gnd d2 a_17676_3222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X989 vdd a_19123_3989# a_18915_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X990 a_34866_13694# a_34445_13694# a_33818_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X991 a_54448_13779# a_54448_13384# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X992 a_55278_10054# a_56118_10729# a_56326_10729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X993 a_22282_9369# a_22282_8974# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X994 a_9211_13658# a_9464_13645# a_8163_12983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_45617_13702# a_45196_13702# a_44569_13027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X996 a_11315_3357# a_11936_3278# a_12144_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X997 vdd d0 a_9462_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X998 a_76120_2960# a_76120_2705# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X999 a_68357_5567# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1000 a_75744_444# a_75531_444# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1001 gnd a_41843_6182# a_41635_6182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1002 a_11316_11937# a_11937_12253# a_12145_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1003 a_41592_11524# a_41845_11511# a_40540_11705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1004 a_46857_10055# a_46644_10055# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1005 a_18868_8740# a_19125_8550# a_17421_9420# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1006 a_82224_3410# a_83720_2540# a_83675_2553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1007 a_29837_10014# a_30930_10676# a_30885_10689# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1008 a_76121_12330# a_76121_11935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1009 a_52344_8565# a_52597_8552# a_51292_8746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 vdd d3 a_82440_10673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1011 a_66240_7696# a_65819_7696# a_65411_7380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1012 a_18870_4002# a_19963_4664# a_19914_4854# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1013 a_6670_10871# a_6927_10681# a_5606_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1014 a_9209_5524# a_9462_5511# a_8157_5705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 a_22688_4050# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 a_44146_5572# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1017 a_66870_10733# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1018 a_84725_9236# a_84978_9223# a_83677_8561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1019 a_76949_3276# a_76528_3276# a_76120_3355# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1020 a_22901_2603# a_22688_2603# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1021 a_62002_2555# a_62255_2542# a_60551_3412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1022 gnd a_52597_9231# a_52389_9231# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1023 a_55067_5566# a_54854_5566# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1024 a_68316_13020# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1025 a_43741_10168# a_43741_9627# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1026 a_11723_4046# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1027 a_11935_5566# a_11722_5566# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1028 a_43740_12594# a_44361_13027# a_44569_13027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1029 a_76527_6243# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 a_22687_7696# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1031 a_55902_7688# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1032 a_33608_7011# a_33395_7011# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_49842_6385# a_51338_5515# a_51293_5528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1034 a_2485_13702# a_2064_13702# a_1437_13706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1035 gnd a_41846_10670# a_41638_10670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1036 a_19917_7644# a_20170_7631# a_18869_6969# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1037 a_1228_4052# a_1015_4052# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1038 a_66243_8611# a_67083_9286# a_67291_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1039 a_11317_8715# a_11938_8607# a_12146_8607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_33396_2597# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1041 vdd d2 a_17676_3222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1042 a_84719_4852# a_84723_3996# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1043 a_52340_8742# a_52341_7650# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1044 a_28345_4684# a_28432_6193# a_28387_6206# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1045 a_54857_10054# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1046 a_36356_11569# a_37214_8596# a_37422_8596# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1047 a_12144_2599# a_12984_3274# a_13192_3274# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1048 a_9207_13835# a_9464_13645# a_8163_12983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1049 vdd a_60765_4667# a_60557_4667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1050 vdd d0 a_31135_6188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1051 a_55275_7013# a_56115_7688# a_56323_7688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1052 vdd a_30089_12968# a_29881_12968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1053 vdd a_41843_6182# a_41635_6182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1054 gnd d1 a_51548_12970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1055 a_41588_11701# a_41845_11511# a_40540_11705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1056 gnd a_74267_6956# a_74059_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1057 a_22282_8974# a_22282_8719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1058 a_2483_7694# a_2062_7694# a_1435_7698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1059 a_52340_8742# a_52597_8552# a_51292_8746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1060 a_55275_7692# a_54854_7692# a_54446_7376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 a_55905_10729# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1062 a_43738_8033# a_44362_8613# a_44570_8613# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1063 a_609_10818# a_1230_10739# a_1438_10739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1064 vdd d0 a_31136_4668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1065 a_18870_4002# a_19963_4664# a_19918_4677# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1066 a_76740_5564# a_76527_5564# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1067 a_76121_12330# a_76742_12251# a_76950_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1068 a_9205_5701# a_9462_5511# a_8157_5705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1069 a_30881_9419# a_31138_9229# a_29837_8567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1070 a_77576_3272# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1071 gnd a_8415_2548# a_8207_2548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1072 a_55069_12253# a_54856_12253# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1073 a_76951_10052# a_76530_10052# a_76122_10160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1074 a_84721_9413# a_84978_9223# a_83677_8561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1075 a_26506_8602# a_26293_8602# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1076 a_61998_2732# a_62255_2542# a_60551_3412# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1077 a_1230_9292# a_1017_9292# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1078 vdd a_52597_9231# a_52389_9231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1079 a_40539_4177# a_40796_3987# a_39096_3233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1080 a_23111_10737# a_22690_10737# a_22282_10421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1081 a_74014_6201# a_74010_6378# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1082 gnd d0 a_20172_13639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 vdd a_41846_10670# a_41638_10670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1084 a_76121_11935# a_76121_11680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1085 a_19913_7821# a_20170_7631# a_18869_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1086 a_19919_12205# a_19915_12382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1087 gnd d2 a_39351_9228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1088 a_11314_7376# a_11935_7692# a_12143_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1089 a_80554_8596# a_80133_8596# a_79488_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1090 a_65819_6249# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1091 a_30883_2555# a_31136_2542# a_29831_2736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1092 vdd d0 a_74269_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1093 a_44146_7019# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1094 a_84723_2549# a_84976_2536# a_83671_2730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1095 a_79387_5561# a_79023_4039# a_77997_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1096 a_36356_11569# a_35935_11569# a_36257_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1097 a_70191_4731# a_69770_4731# a_69846_8602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1098 a_66034_11578# a_65821_11578# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1099 gnd a_52595_2544# a_52387_2544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1100 a_45616_4727# a_46855_4047# a_47006_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1101 a_35891_4039# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1102 vdd a_19122_5509# a_18914_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1103 gnd a_63304_12960# a_63096_12960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 vdd d1 a_73221_12968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1105 a_3876_11577# a_3512_10055# a_2486_10735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1106 a_54449_8715# a_54446_8027# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1107 a_30878_6378# a_30882_5522# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1108 a_34659_10727# a_34446_10727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_9208_10189# a_9465_9999# a_8160_10193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1110 a_6714_6208# a_8206_6962# a_8157_7152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1111 a_34445_13694# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1112 a_14681_5563# a_14260_5563# a_14582_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1113 gnd d0 a_31137_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 a_28386_9424# a_29882_8554# a_29833_8744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1115 vdd a_9462_7637# a_9254_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1116 a_34443_6239# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1117 a_19915_12382# a_20172_12192# a_18871_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1118 a_11938_9286# a_11725_9286# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1119 a_51296_8569# a_52389_9231# a_52340_9421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1120 a_18867_11707# a_19124_11517# a_17420_12387# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1121 a_607_4160# a_1228_4052# a_1436_4052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1122 a_63051_11526# a_63304_11513# a_61999_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1123 a_34864_6239# a_36103_7006# a_36260_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1124 a_22280_5064# a_22280_4808# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1125 a_12145_13021# a_11724_13021# a_11316_12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1126 a_30879_4179# a_30883_3234# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1127 gnd d2 a_71774_12201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 a_14683_11571# a_14262_11571# a_14584_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1129 a_23949_4725# a_23736_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1130 a_22281_13783# a_22902_13704# a_23110_13704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1131 a_83677_8561# a_83930_8548# a_82226_9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1132 a_606_7382# a_1227_7698# a_1435_7698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1133 a_6672_4686# a_6759_6195# a_6714_6208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1134 gnd d3 a_17633_4667# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1135 a_52343_13658# a_52339_13835# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1136 a_41586_7140# a_41590_6195# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1137 a_21784_433# a_21363_433# a_21685_433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1138 a_45616_3280# a_45195_3280# a_44568_2605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1139 a_1014_6251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1140 gnd d1 a_83928_2540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1141 a_29833_10191# a_30930_9997# a_30881_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1142 a_21363_433# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 a_66241_2603# a_65820_2603# a_65414_2612# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1144 gnd a_17678_9230# a_17470_9230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1145 a_77999_9280# a_77578_9280# a_76951_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1146 a_63052_8559# a_63305_8546# a_62000_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1147 a_22687_5570# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1148 a_24156_7692# a_23735_7692# a_23108_7017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1149 a_33817_4044# a_33396_4044# a_32988_4152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1150 a_8162_4008# a_9255_4670# a_9206_4860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1151 a_22282_9625# a_22903_10058# a_23111_10058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1152 a_77996_7686# a_77575_7686# a_76948_7011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1153 vdd d1 a_19124_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1154 a_25395_7012# a_25182_7012# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1155 a_12983_6241# a_12770_6241# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1156 a_54447_3357# a_54447_2962# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1157 a_11722_5566# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1158 a_33395_7011# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1159 a_30879_2732# a_31136_2542# a_29831_2736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1160 a_84719_2726# a_84976_2536# a_83671_2730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1161 a_39055_10686# a_39142_12195# a_39097_12208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1162 a_19918_4677# a_19914_4854# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1163 a_1227_5572# a_1014_5572# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1164 a_77790_13694# a_77577_13694# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1165 a_25648_11575# a_26506_8602# a_26714_8602# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1166 a_17380_4680# a_17467_6189# a_17418_6379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1167 a_54446_5929# a_55067_6245# a_55275_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1168 vdd a_52595_2544# a_52387_2544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1169 a_17376_4857# a_17633_4667# a_16310_7830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1170 a_76529_13698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1171 a_2278_10735# a_2065_10735# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1172 a_76743_9284# a_76530_9284# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1173 gnd a_30088_2546# a_29880_2546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1174 a_1014_7019# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1175 a_48097_4733# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1176 a_44570_9292# a_44149_9292# a_43741_8976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1177 a_17421_9420# a_18917_8550# a_18868_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1178 gnd d2 a_17677_12197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1179 a_18867_11707# a_19964_11513# a_19915_11703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 a_56118_9282# a_55905_9282# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1181 a_15886_4727# a_15673_4727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1182 a_76122_10415# a_76743_10731# a_76951_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1183 a_28386_9424# a_29882_8554# a_29837_8567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1184 gnd d0 a_20171_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1185 vdd d0 a_63302_5505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1186 a_9211_12979# a_9464_12966# a_8159_13160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1187 a_57716_11571# a_57352_10049# a_56326_10729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1188 a_51296_8569# a_52389_9231# a_52344_9244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1189 vdd a_31135_6188# a_30927_6188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1190 a_46856_13022# a_46643_13022# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1191 a_63047_11703# a_63304_11513# a_61999_11707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1192 a_25227_11575# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1193 a_45196_13702# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1194 a_77998_12247# a_77577_12247# a_76950_11572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1195 a_60557_9243# a_60810_9230# a_60510_10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 a_8161_5528# a_9254_6190# a_9209_6203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1197 a_60554_6202# a_62046_6956# a_62001_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1198 a_8159_11713# a_9256_11519# a_9207_11709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1199 a_83673_10185# a_84770_9991# a_84725_10004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1200 vdd d1 a_83928_2540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1201 vdd d0 a_63303_3985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1202 a_30882_5522# a_30878_5699# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1203 a_72969_8567# a_74062_9229# a_74013_9419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1204 a_11936_2599# a_11723_2599# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1205 a_51290_2738# a_52387_2544# a_52338_2734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1206 vdd a_31136_4668# a_30928_4668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1207 a_13194_9282# a_12773_9282# a_12146_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1208 vdd a_17678_9230# a_17470_9230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1209 a_63048_8736# a_63305_8546# a_62000_8740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1210 a_11724_11574# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1211 a_22688_4729# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1212 a_29832_11711# a_30929_11517# a_30880_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1213 a_26293_8602# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1214 a_18866_4179# a_19963_3985# a_19914_4175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 a_8162_4008# a_9255_4670# a_9210_4683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1216 a_54448_11682# a_54449_11068# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1217 a_9205_7827# a_9209_6971# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1218 a_51293_6975# a_51546_6962# a_49846_6208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1219 a_40538_5697# a_40795_5507# a_39091_6377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1220 a_74013_10866# a_74017_10010# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1221 a_83675_2553# a_84768_3215# a_84719_3405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1222 a_43741_10818# a_43741_10423# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1223 a_22279_7775# a_22900_7696# a_23108_7696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1224 vdd d0 a_41843_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1225 a_66242_11578# a_65821_11578# a_65413_11686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1226 a_71479_10692# a_71566_12201# a_71517_12391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1227 a_72968_11534# a_74061_12196# a_74016_12209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1228 vdd d0 a_20173_9993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1229 a_72966_5526# a_73219_5513# a_71515_6383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1230 a_22689_13704# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1231 gnd d0 a_84975_6182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1232 a_22687_7017# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1233 a_41590_6195# a_41843_6182# a_40542_5520# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1234 vdd a_30088_2546# a_29880_2546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1235 gnd a_41846_9991# a_41638_9991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1236 a_19917_6965# a_20170_6952# a_18865_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1237 a_17421_9420# a_18917_8550# a_18872_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1238 a_68572_11575# a_68359_11575# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1239 a_74012_11707# a_74017_10689# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1240 a_18867_11707# a_19964_11513# a_19919_11526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1241 a_84721_9413# a_84725_8557# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1242 a_63052_8559# a_63048_8736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1243 a_49845_9426# a_51341_8556# a_51292_8746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1244 a_24156_7692# a_25395_7012# a_25552_5686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1245 a_30885_10689# a_31138_10676# a_29837_10014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1246 a_17424_12210# a_18916_12964# a_18871_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1247 gnd d0 a_52596_11519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_66032_7696# a_65819_7696# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 a_2484_4727# a_2063_4727# a_1436_4052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1250 a_23108_5570# a_23948_6245# a_24156_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1251 a_74011_2732# a_65414_2612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1252 a_76120_3611# a_76120_3355# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1253 a_52342_4683# a_52595_4670# a_51294_4008# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1254 a_65821_12257# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1255 a_60553_9420# a_60810_9230# a_60510_10865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1256 a_79238_10047# a_79025_10047# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1257 a_11725_9286# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1258 a_76741_2597# a_76528_2597# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1259 a_606_5680# a_1227_5572# a_1435_5572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1260 a_45407_7694# a_45194_7694# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1261 a_67082_12253# a_66869_12253# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1262 gnd d1 a_62256_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_11314_7376# a_11314_7121# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1264 a_55068_3278# a_54855_3278# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1265 gnd a_39350_12195# a_39142_12195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1266 gnd a_74270_8550# a_74062_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1267 a_46644_10055# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1268 a_51290_2738# a_52387_2544# a_52342_2557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1269 a_23736_4725# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1270 a_17382_10688# a_17469_12197# a_17420_12387# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1271 a_14220_10049# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1272 a_44568_2605# a_44147_2605# a_43739_2713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1273 a_76742_12251# a_76529_12251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1274 gnd d3 a_28600_10679# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 gnd a_83928_2540# a_83720_2540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1276 a_34657_4719# a_34444_4719# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1277 a_12985_13696# a_12772_13696# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1278 gnd a_40797_11515# a_40589_11515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1279 a_83675_2553# a_84768_3215# a_84723_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1280 a_11315_4804# a_11936_4725# a_12144_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1281 a_33816_5564# a_33395_5564# a_32987_5672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1282 a_79389_11569# a_79280_11569# a_79488_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1283 a_25182_7012# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1284 a_56323_6241# a_55902_6241# a_55275_5566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1285 a_72962_5703# a_73219_5513# a_71515_6383# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1286 a_72962_5703# a_74059_5509# a_74010_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1287 a_76529_11572# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1288 a_76122_9363# a_76122_8968# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1289 vout a_42796_401# a_21784_433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1290 vdd d0 a_84975_6182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1291 vdd a_9464_11519# a_9256_11519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1292 a_23111_10058# a_22690_10058# a_22282_9625# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1293 a_79022_7006# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1294 a_12770_6241# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1295 a_52337_6380# a_52594_6190# a_51293_5528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1296 a_41586_6372# a_41843_6182# a_40542_5520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1297 a_3881_11696# a_3511_13022# a_2485_12255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1298 vdd a_8416_12970# a_8208_12970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1299 a_77999_10727# a_77578_10727# a_76951_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1300 a_32399_444# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1301 gnd d3 a_71730_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1302 a_47013_11696# a_46643_13022# a_45617_13702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1303 a_71522_9247# a_73014_10001# a_72969_10014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1304 a_11314_6580# a_11935_7013# a_12143_7013# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1305 gnd a_63304_13639# a_63096_13639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1306 a_52339_13156# a_52596_12966# a_51291_13160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1307 a_76530_9284# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1308 a_44149_8613# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1309 a_49845_9426# a_51341_8556# a_51296_8569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1310 a_76950_11572# a_77790_12247# a_77998_12247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1311 gnd a_82480_6187# a_82272_6187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1312 a_30881_10866# a_31138_10676# a_29837_10014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1313 a_34659_9280# a_34446_9280# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1314 a_54180_446# a_58805_4727# a_58881_8598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1315 gnd a_20170_6184# a_19962_6184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 a_76949_4723# a_76528_4723# a_76120_4802# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1317 a_56117_12249# a_55904_12249# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1318 a_25398_10053# a_25185_10053# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1319 a_52338_4860# a_52595_4670# a_51294_4008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1320 a_15673_4727# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1321 vdd a_63302_5505# a_63094_5505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1322 a_57716_11571# a_57607_11571# a_57815_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1323 a_43739_4415# a_44360_4731# a_44568_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1324 a_47006_5569# a_46897_5569# a_47105_5569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1325 gnd a_6969_12203# a_6761_12203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1326 gnd a_74269_12196# a_74061_12196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1327 a_76951_8605# a_76530_8605# a_76119_8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 a_5178_4733# a_4965_4733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1329 a_609_8721# a_606_8033# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1330 a_32987_7769# a_32987_7374# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1331 a_76119_7769# a_76740_7690# a_76948_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1332 a_1015_3284# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1333 vdd a_74270_8550# a_74062_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1334 gnd d0 a_9462_7637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1335 a_51295_11536# a_52388_12198# a_52339_12388# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1336 vdd a_31137_12196# a_30929_12196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1337 a_22282_9625# a_22282_9369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1338 a_71477_4684# a_71564_6193# a_71515_6383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1339 a_52343_13658# a_54448_13779# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1340 a_30881_8740# a_30882_7648# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1341 a_82223_6377# a_83719_5507# a_83670_5697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1342 a_29831_2736# a_30928_2542# a_30879_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1343 vdd a_83928_2540# a_83720_2540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1344 vdd a_63303_3985# a_63095_3985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1345 a_25396_4045# a_25183_4045# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1346 a_12144_4046# a_12984_4721# a_13192_4721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1347 a_22281_13133# a_22902_13025# a_23110_13025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1348 gnd d0 a_84977_12190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1349 a_44570_9292# a_45410_9288# a_45618_9288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1350 a_11723_2599# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1351 vdd a_40797_11515# a_40589_11515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1352 a_606_6586# a_1227_7019# a_1435_7019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1353 a_14262_11571# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1354 a_25554_11694# a_25440_11575# a_25648_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1355 a_18865_5699# a_19962_5505# a_19913_5695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1356 gnd d0 a_9464_12198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1357 a_609_10168# a_609_9627# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1358 a_17423_3235# a_17676_3222# a_17376_4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1359 vdd d0 a_41845_12190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1360 a_6670_10871# a_6762_9236# a_6713_9426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1361 a_54447_3357# a_55068_3278# a_55276_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1362 a_30884_12977# a_30880_13154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1363 vdd a_41843_7629# a_41635_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1364 a_22280_2711# a_22901_2603# a_23109_2603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1365 a_8158_4185# a_9255_3991# a_9206_4181# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1366 a_45615_6247# a_45194_6247# a_44567_6251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1367 a_34866_12247# a_36105_13014# a_36262_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1368 gnd a_84975_6182# a_84767_6182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1369 a_65822_10737# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1370 gnd d0 a_41843_6950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1371 vdd d3 a_71730_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1372 a_14432_13016# a_14219_13016# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1373 a_81115_7828# a_81372_7638# a_80800_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1374 a_22280_4413# a_22280_4158# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1375 a_23110_12257# a_23950_12253# a_24158_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1376 a_67083_10733# a_66870_10733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1377 a_74015_4681# a_74011_4858# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1378 a_57721_11690# a_57351_13016# a_56325_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1379 a_19920_9238# a_19916_9415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1380 a_1435_6251# a_1014_6251# a_606_5935# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1381 a_71521_12214# a_73013_12968# a_72964_13158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1382 a_76529_13019# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1383 vdd a_20170_6184# a_19962_6184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1384 a_55069_13700# a_54856_13700# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1385 vdd a_19125_9997# a_18917_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1386 a_1017_8613# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 a_44360_3284# a_44147_3284# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 a_36260_5680# a_36146_5561# a_36354_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1389 a_32989_12330# a_33610_12251# a_33818_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 vdd d2 a_82483_9228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1391 a_76743_10731# a_76530_10731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1392 a_33819_9284# a_33398_9284# a_32990_8968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1393 a_3509_7014# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1394 a_66033_2603# a_65820_2603# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1395 a_11937_12253# a_11724_12253# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1396 a_34446_10727# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1397 a_76122_9619# a_76743_10052# a_76951_10052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1398 gnd a_60765_4667# a_60557_4667# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1399 a_45194_7694# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1400 a_60508_4857# a_60600_3222# a_60551_3412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1401 a_63050_4677# a_63303_4664# a_62002_4002# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1402 a_65819_7696# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1403 a_65413_13133# a_65413_12592# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1404 a_32989_13382# a_32989_13127# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1405 a_33608_6243# a_33395_6243# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1406 a_77577_12247# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1407 a_54449_8715# a_55070_8607# a_55278_8607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1408 a_29831_2736# a_30928_2542# a_30883_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1409 a_76528_2597# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1410 a_49848_12216# a_51340_12970# a_51291_13160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1411 vdd d1 a_73220_3993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1412 a_84720_13148# a_84977_12958# a_83672_13152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1413 a_1229_12259# a_1016_12259# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1414 a_28385_12391# a_28642_12201# a_28347_10692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1415 a_82229_12208# a_82482_12195# a_82187_10686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1416 a_55276_2599# a_56116_3274# a_56324_3274# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1417 a_17419_3412# a_17676_3222# a_17376_4857# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1418 a_43738_6330# a_43738_5935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1419 a_49846_6208# a_50099_6195# a_49804_4686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1420 gnd d0 a_31136_4668# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1421 a_5041_8604# a_5178_4733# a_5386_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1422 a_2485_12255# a_3724_13022# a_3881_11696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1423 a_6670_10871# a_6762_9236# a_6717_9249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1424 vdd d0 a_52595_3991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1425 a_72968_11534# a_73221_11521# a_71517_12391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 a_30885_9242# a_31138_9229# a_29837_8567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1427 a_34443_7686# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1428 a_61997_5699# a_63094_5505# a_63049_5518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1429 vdd d0 a_74267_6188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1430 a_84720_13148# a_84724_12203# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1431 vdd a_84975_6182# a_84767_6182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1432 gnd d1 a_8417_10003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1433 a_44362_8613# a_44149_8613# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1434 a_39095_6200# a_39348_6187# a_39053_4678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1435 a_19919_13652# a_22281_13783# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1436 vdd a_52596_11519# a_52388_11519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1437 a_22689_13025# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1438 a_83676_11528# a_84769_12190# a_84720_12380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1439 a_65414_9369# a_66035_9290# a_66243_9290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1440 a_23109_3282# a_23949_3278# a_24157_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1441 a_77791_10727# a_77578_10727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1442 a_9208_10189# a_9212_9244# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1443 a_33818_11572# a_33397_11572# a_32989_11680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1444 vdd a_63305_9993# a_63097_9993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1445 a_54854_7692# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1446 a_61998_4179# a_63095_3985# a_63050_3998# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1447 vdd d0 a_74268_4668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1448 a_32721_444# a_37346_4725# a_37422_8596# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1449 a_40544_11528# a_41637_12190# a_41592_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1450 gnd d0 a_74269_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1451 a_79237_13014# a_79024_13014# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1452 a_52342_3236# a_52338_3413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1453 gnd a_19124_12964# a_18916_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1454 a_69638_8602# a_69425_8602# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1455 a_12986_9282# a_12773_9282# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1456 a_25547_5567# a_25438_5567# a_25646_5567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1457 a_35892_13014# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1458 a_30885_10010# a_31138_9997# a_29833_10191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1459 gnd d4 a_27532_7644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1460 a_60508_4857# a_60600_3222# a_60555_3235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1461 a_63046_4854# a_63303_4664# a_62002_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1462 a_46643_13022# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1463 a_52342_4004# a_52595_3991# a_51290_4185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1464 a_33610_13698# a_33397_13698# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1465 a_607_2968# a_607_2713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1466 gnd a_50101_12203# a_49893_12203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 gnd d2 a_28643_9234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1468 gnd a_9462_7637# a_9254_7637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 a_23737_13700# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1470 a_18871_11530# a_19124_11517# a_17420_12387# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1471 a_40545_10008# a_40798_9995# a_39098_9241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1472 a_54446_7376# a_55067_7692# a_55275_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1473 a_22279_7380# a_22279_7125# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1474 gnd a_20173_10672# a_19965_10672# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1475 a_32988_2705# a_32990_2606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1476 a_33817_2597# a_33396_2597# a_32990_2606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1477 a_74015_2555# a_74268_2542# a_72963_2736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_25183_4045# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1479 a_28385_12391# a_29881_11521# a_29832_11711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1480 a_23111_10058# a_23951_10733# a_24159_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1481 gnd a_73219_6960# a_73011_6960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1482 a_79023_4039# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1483 gnd d1 a_73219_5513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1484 a_36146_5561# a_35933_5561# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1485 a_52339_13835# a_52343_12979# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1486 a_72964_11711# a_73221_11521# a_71517_12391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1487 a_36103_7006# a_35890_7006# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1488 a_42796_401# d8 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1489 a_57813_5563# a_57392_5563# a_57714_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1490 gnd d0 a_52594_5511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1491 a_11315_4154# a_11936_4046# a_12144_4046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1492 a_32990_10415# a_33611_10731# a_33819_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1493 a_37668_4725# a_38032_7638# a_37987_7651# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1494 a_32987_6322# a_33608_6243# a_33816_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1495 a_11938_10733# a_11725_10733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1496 a_57719_5682# a_57349_7008# a_56323_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1497 gnd a_41843_6950# a_41635_6950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1498 a_11316_12588# a_11937_13021# a_12145_13021# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1499 a_68681_11575# a_68317_10053# a_67291_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1500 a_12143_6245# a_12983_6241# a_13191_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1501 gnd d1 a_40797_12962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1502 a_36257_11569# a_35893_10047# a_34867_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1503 a_12145_12253# a_11724_12253# a_11316_12332# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1504 a_74012_11707# a_74269_11517# a_72964_11711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1505 a_72969_8567# a_73222_8554# a_71518_9424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1506 a_43739_4160# a_43739_3619# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1507 a_43738_5935# a_43738_5680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1508 a_74012_12386# a_74016_11530# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1509 a_19914_4854# a_19918_3998# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1510 a_3511_13022# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1511 a_43740_12338# a_43740_11943# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1512 a_54448_12332# a_55069_12253# a_55277_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1513 a_54446_7121# a_54446_6580# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1514 a_17380_4680# a_17633_4667# a_16310_7830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1515 a_65819_5570# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1516 vdd d4 a_27532_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1517 a_83675_2553# a_83928_2540# a_82224_3410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1518 a_54447_3613# a_54447_3357# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1519 a_67288_7692# a_66867_7692# a_66240_7017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1520 a_65820_2603# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1521 a_76949_4044# a_76528_4044# a_76120_4152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1522 a_68527_7012# a_68314_7012# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1523 a_43739_3619# a_44360_4052# a_44568_4052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1524 vdd d2 a_28643_9234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1525 a_14582_5563# a_14218_4041# a_13192_4721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1526 a_63045_5695# a_63050_4677# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1527 vdd a_20173_10672# a_19965_10672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1528 a_76527_7011# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1529 a_74011_2732# a_74268_2542# a_72963_2736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1530 a_52344_10691# a_52340_10868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1531 gnd d0 a_9462_6958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1532 a_28385_12391# a_29881_11521# a_29836_11534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1533 a_33395_6243# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1534 gnd d1 a_62255_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1535 a_41593_8557# a_41589_8734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1536 a_64817_433# a_64708_433# a_43118_401# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1537 gnd d2 a_71773_3226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1538 vdd d1 a_73219_5513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1539 a_609_10818# a_609_10423# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1540 a_84725_10004# a_84721_10181# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1541 a_606_8033# a_1230_8613# a_1438_8613# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1542 a_23108_7017# a_23948_7692# a_24156_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1543 a_59018_4727# a_58805_4727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1544 gnd a_31136_4668# a_30928_4668# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1545 vdd d0 a_52594_5511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1546 a_40538_5697# a_41635_5503# a_41590_5516# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1547 a_30884_13656# a_30880_13833# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1548 a_25438_5567# a_25225_5567# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1549 a_65821_13704# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1550 a_12986_10729# a_12773_10729# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1551 a_44147_4731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1552 vdd a_74267_6188# a_74059_6188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1553 a_9211_12979# a_9207_13156# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1554 a_9209_6203# a_9205_6380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1555 a_67082_13700# a_66869_13700# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1556 a_45617_12255# a_45196_12255# a_44569_12259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1557 a_41589_10860# a_41593_10004# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1558 a_55068_4725# a_54855_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1559 a_13193_12249# a_12772_12249# a_12145_11574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1560 gnd d0 a_41843_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1561 a_5041_8604# a_4620_8604# a_3975_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1562 a_72965_8744# a_73222_8554# a_71518_9424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1563 a_32987_5672# a_32988_5058# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1564 a_65822_10058# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1565 a_5386_4733# a_10939_446# a_11147_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1566 a_55277_11574# a_54856_11574# a_54448_11682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1567 a_74017_10689# a_74270_10676# a_72969_10014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1568 a_40539_4177# a_41636_3983# a_41591_3996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1569 a_39097_12208# a_40589_12962# a_40544_12975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1570 a_28388_3239# a_29880_3993# a_29831_4183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 vdd a_74268_4668# a_74060_4668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1572 a_74017_9242# a_74013_9419# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1573 a_83671_2730# a_83928_2540# a_82224_3410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1574 a_25554_11694# a_25184_13020# a_24158_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1575 a_33610_11572# a_33397_11572# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1576 a_56326_9282# a_55905_9282# a_55278_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1577 a_69425_8602# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1578 a_33816_6243# a_34656_6239# a_34864_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1579 a_57351_13016# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1580 a_55069_13021# a_54856_13021# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1581 a_12773_9282# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1582 a_33609_3276# a_33396_3276# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1583 a_41591_3228# a_41587_3405# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1584 a_11316_13779# a_11316_13384# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1585 a_76743_10052# a_76530_10052# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1586 gnd a_27532_7644# a_27324_7644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 vdd d0 a_84975_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1588 a_10939_446# a_10726_446# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1589 a_65411_7775# a_66032_7696# a_66240_7696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_41586_7819# a_41843_7629# a_40542_6967# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1591 a_62004_10010# a_62257_9997# a_60557_9243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1592 a_74016_11530# a_74012_11707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1593 a_43740_11943# a_43740_11688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1594 gnd d2 a_60808_3222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_63050_3998# a_63303_3985# a_61998_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1596 a_54856_12253# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1597 a_1438_10739# a_2278_10735# a_2486_10735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1598 a_65819_7017# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1599 a_34444_4719# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1600 a_84722_6195# a_84975_6182# a_83674_5520# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1601 a_65411_6328# a_65411_5933# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1602 vdd d2 a_71773_3226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1603 a_76950_13019# a_77790_13694# a_77998_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1604 gnd a_52594_6190# a_52386_6190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1605 gnd a_39349_3220# a_39141_3220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_36255_5561# a_35891_4039# a_34865_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1607 a_36148_11569# a_35935_11569# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1608 gnd a_20170_7631# a_19962_7631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1609 a_74015_2555# a_74011_2732# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1610 a_56117_13696# a_55904_13696# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1611 a_67288_7692# a_68527_7012# a_68684_5686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1612 a_82183_10863# a_82275_9228# a_82230_9241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1613 a_54446_6580# a_54446_6324# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1614 a_54449_10417# a_55070_10733# a_55278_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1615 a_66240_5570# a_67080_6245# a_67288_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1616 gnd d0 a_31136_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1617 a_11314_5674# a_11935_5566# a_12143_5566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1618 gnd a_74269_13643# a_74061_13643# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1619 a_63047_13150# a_63051_12205# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1620 gnd d3 a_50057_4673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1621 a_1015_4731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1622 gnd a_84977_11511# a_84769_11511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1623 a_51295_12983# a_52388_13645# a_52339_13835# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1624 gnd a_9464_11519# a_9256_11519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1625 a_61999_11707# a_63096_11513# a_63047_11703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1626 a_74013_10866# a_74270_10676# a_72969_10014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1627 a_1435_7698# a_2275_7694# a_2483_7694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1628 a_68530_10053# a_68317_10053# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1629 a_3879_5688# a_3509_7014# a_2483_7694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1630 a_19917_6197# a_19913_6374# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1631 gnd d3 a_39306_4665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1632 a_76950_12251# a_76529_12251# a_76121_12330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1633 gnd d0 a_9464_13645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1634 a_77789_4719# a_77576_4719# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1635 a_72962_7150# a_74059_6956# a_74014_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1636 vdd a_27532_7644# a_27324_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1637 a_54447_4804# a_55068_4725# a_55276_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1638 a_76948_5564# a_76527_5564# a_76119_5672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1639 gnd a_71774_12201# a_71566_12201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1640 a_8164_10016# a_9257_10678# a_9212_10691# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1641 a_79278_5561# a_79065_5561# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1642 a_43739_5066# a_44359_5572# a_44567_5572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1643 a_45615_7694# a_45194_7694# a_44567_7698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1644 a_68314_7012# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1645 a_55902_6241# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1646 vdd d2 a_60808_3222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1647 a_23110_13704# a_23950_13700# a_24158_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1648 a_1438_9292# a_1017_9292# a_609_9371# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1649 a_84718_6372# a_84975_6182# a_83674_5520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1650 a_33610_13019# a_33397_13019# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1651 a_79488_11569# a_80346_8596# a_80554_8596# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1652 gnd a_9462_6958# a_9254_6958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1653 a_13194_10729# a_12773_10729# a_12146_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1654 gnd d1 a_62254_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1655 a_76950_13019# a_76529_13019# a_76121_12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1656 gnd a_20173_9993# a_19965_9993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 a_54446_6580# a_55067_7013# a_55275_7013# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1658 vdd a_39349_3220# a_39141_3220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1659 gnd a_62255_3989# a_62047_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1660 vdd a_20170_7631# a_19962_7631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1661 a_9207_12388# a_9464_12198# a_8163_11536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1662 a_80691_4725# a_80478_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1663 a_71477_4684# a_71730_4671# a_70407_7834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1664 a_44360_4731# a_44147_4731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1665 a_32612_444# a_32399_444# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1666 a_58805_4727# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1667 vdd d3 a_50057_4673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1668 a_11937_13700# a_11724_13700# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1669 vdd a_74269_13643# a_74061_13643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1670 a_32987_8025# a_32987_7769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1671 a_49843_3418# a_51339_2548# a_51294_2561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1672 a_70092_4731# a_69983_4731# a_70191_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1673 a_25225_5567# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1674 a_68686_11694# a_68316_13020# a_67290_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1675 vdd a_84977_11511# a_84769_11511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1676 a_51295_12983# a_52388_13645# a_52343_13658# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1677 gnd d1 a_30090_10001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1678 a_32990_9619# a_33611_10052# a_33819_10052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1679 gnd a_6970_9236# a_6762_9236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1680 a_65412_4158# a_65412_3617# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1681 a_65411_5933# a_65411_5678# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1682 vdd a_83929_12962# a_83721_12962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1683 a_61999_11707# a_63096_11513# a_63051_11526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1684 gnd a_41843_7629# a_41635_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1685 a_82227_6200# a_83719_6954# a_83674_6967# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1686 a_14587_5682# a_14473_5563# a_14681_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1687 a_11316_13384# a_11937_13700# a_12145_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1688 vdd d0 a_74270_9229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1689 a_48738_7659# a_48991_7646# a_48419_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1690 a_60555_3235# a_62047_3989# a_62002_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1691 a_43739_4810# a_43739_4415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1692 a_11314_5929# a_11314_5674# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1693 a_77577_13694# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1694 a_11938_10054# a_11725_10054# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1695 vdd d3 a_39306_4665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1696 vdd d0 a_84977_13637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1697 a_60556_12210# a_62048_12964# a_62003_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1698 gnd a_17677_12197# a_17469_12197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1699 vdd d0 a_52597_10678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1700 a_2275_6247# a_2062_6247# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1701 a_71516_3416# a_73012_2546# a_72963_2736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1702 a_18870_2555# a_19963_3217# a_19918_3230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1703 a_1229_13706# a_1016_13706# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1704 vdd d0 a_9464_13645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1705 a_23738_9286# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1706 a_81119_7651# a_81372_7638# a_80800_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1707 a_18865_7146# a_19962_6952# a_19917_6965# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1708 a_51293_5528# a_52386_6190# a_52337_6380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1709 a_68528_4045# a_68315_4045# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1710 a_1016_12259# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_55276_4046# a_56116_4721# a_56324_4721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1712 a_54857_10733# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1713 a_19916_9415# a_19920_8559# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1714 gnd a_71775_9234# a_71567_9234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_23109_4729# a_22688_4729# a_22280_4808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1716 a_22281_11941# a_22902_12257# a_23110_12257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1717 a_33396_3276# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1718 gnd d2 a_82483_9228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 a_6713_9426# a_8209_8556# a_8160_8746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1720 vdd a_84975_7629# a_84767_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1721 a_65412_2711# a_66033_2603# a_66241_2603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1722 a_82223_6377# a_82480_6187# a_82185_4678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1723 a_44569_12259# a_44148_12259# a_43740_11943# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1724 vdd d1 a_51547_3995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1725 a_607_3619# a_607_3363# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1726 gnd d0 a_84975_6950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1727 gnd a_60808_3222# a_60600_3222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1728 a_23109_4729# a_23949_4725# a_24157_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1729 a_63049_5518# a_63302_5505# a_61997_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1730 vdd a_73222_10001# a_73014_10001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1731 a_84722_6963# a_84718_7140# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1732 gnd d0 a_9465_8552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 a_41590_6963# a_41843_6950# a_40538_7144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1734 a_71473_4861# a_71730_4671# a_70407_7834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1735 a_49849_9249# a_51341_10003# a_51296_10016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1736 a_30883_3234# a_30879_3411# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1737 a_55277_11574# a_56117_12249# a_56325_12249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1738 a_24159_10733# a_25398_10053# a_25549_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1739 a_63052_10006# a_63048_10183# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1740 a_15995_4727# a_16359_7640# a_16310_7830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1741 a_79392_5680# a_79278_5561# a_79486_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1742 a_1436_2605# a_1015_2605# a_607_2713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1743 a_9211_13658# a_9207_13835# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1744 gnd d0 a_31135_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1745 vdd a_6970_9236# a_6762_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1746 a_77996_7686# a_79235_7006# a_79392_5680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1747 gnd a_31136_3989# a_30928_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1748 gnd a_50057_4673# a_49849_4673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1749 vdd a_74270_9997# a_74062_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1750 a_43741_9371# a_44362_9292# a_44570_9292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1751 a_65821_13025# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1752 a_48734_7836# a_48991_7646# a_48419_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1753 a_44147_4052# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1754 a_8158_4185# a_8415_3995# a_6715_3241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1755 a_51292_10193# a_52389_9999# a_52344_10012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1756 a_11317_9365# a_11317_8970# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1757 a_12143_7692# a_11722_7692# a_11314_7376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1758 a_55068_4046# a_54855_4046# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1759 a_33398_8605# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1760 a_80346_8596# a_80133_8596# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1761 a_71516_3416# a_73012_2546# a_72967_2559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1762 gnd a_52596_11519# a_52388_11519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1763 gnd a_39306_4665# a_39098_4665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1764 a_44567_6251# a_44146_6251# a_43738_6330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1765 a_44362_10060# a_44149_10060# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_74017_10010# a_74270_9997# a_72965_10191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_12146_9286# a_12986_9282# a_13194_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1768 vdd a_71775_9234# a_71567_9234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1769 a_34444_3272# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1770 a_19915_13150# a_20172_12960# a_18867_13154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1771 a_79025_10047# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1772 a_77576_4719# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1773 vdd d0 a_9465_9999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1774 a_32990_8968# a_33611_9284# a_33819_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1775 a_76119_7374# a_76119_7119# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1776 a_60514_10688# a_60767_10675# a_59446_7653# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1777 a_52338_3413# a_52342_2557# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1778 gnd d0 a_74268_4668# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1779 vdd d0 a_20172_12192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1780 a_6713_9426# a_8209_8556# a_8164_8569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1781 a_48173_8604# a_47752_8604# a_47105_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1782 vdd d1 a_19124_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1783 gnd d0 a_63304_11513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1784 a_41593_10683# a_41846_10670# a_40545_10008# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1785 a_79065_5561# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1786 a_18870_4002# a_19123_3989# a_17423_3235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1787 a_83676_12975# a_84769_13637# gnd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1788 a_13191_6241# a_12770_6241# a_12143_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1789 vdd a_60808_3222# a_60600_3222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1790 a_607_4415# a_1228_4731# a_1436_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1791 a_63045_6374# a_63049_5518# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1792 gnd a_41845_12190# a_41637_12190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1793 gnd d1 a_51546_5515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1794 a_13194_9282# a_14433_10049# a_14584_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1795 vdd d0 a_9465_8552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1796 a_11147_446# a_10726_446# a_11048_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1797 a_44567_7019# a_44146_7019# a_43738_6586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1798 a_66241_3282# a_67081_3278# a_67289_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1799 gnd a_62254_5509# a_62046_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1800 a_45410_10735# a_45197_10735# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1801 a_27059_4731# a_26638_4731# a_26714_8602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1802 a_54448_13779# a_55069_13700# a_55277_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1803 a_22689_12257# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1804 a_15995_4727# a_16359_7640# a_16314_7653# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1805 a_63046_4175# a_63050_3230# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1806 vdd d2 a_60809_12197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1807 a_77578_9280# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1808 a_11316_11682# a_11937_11574# a_12145_11574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1809 a_55070_9286# a_54857_9286# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1810 gnd a_20170_6952# a_19962_6952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1811 vdd a_50057_4673# a_49849_4673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1812 a_68679_5567# a_68570_5567# a_68778_5567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1813 a_1017_10739# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1814 a_52343_12211# a_52339_12388# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1815 a_34864_6239# a_34443_6239# a_33816_5564# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1816 a_3874_5569# a_3510_4047# a_2484_3280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 gnd d1 a_83929_12962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1818 a_54449_9621# a_55070_10054# a_55278_10054# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1819 a_51296_8569# a_51549_8556# a_49845_9426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1820 a_41586_5693# a_41591_4675# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1821 a_8163_12983# a_8416_12970# a_6716_12216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1822 gnd a_74269_12964# a_74061_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1823 a_11316_11682# a_11317_11068# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1824 a_79067_11569# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1825 a_2484_3280# a_2063_3280# a_1436_3284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1826 a_37668_4725# a_38032_7638# a_37983_7828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1827 a_1015_4052# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1828 a_60550_6379# a_62046_5509# a_62001_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1829 a_8161_5528# a_8414_5515# a_6710_6385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1830 a_51291_13160# a_52388_12966# a_52339_13156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_608_12338# a_608_11943# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1832 vdd d1 a_40798_9995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1833 vdd a_39306_4665# a_39098_4665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1834 a_76949_2597# a_76528_2597# a_76122_2606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1835 a_55904_12249# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1836 a_28390_9247# a_28643_9234# a_28343_10869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1837 a_608_12338# a_1229_12259# a_1437_12259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1838 gnd a_51549_10003# a_51341_10003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1839 a_54449_8970# a_54449_8715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1840 a_2062_6247# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1841 vdd d0 a_63303_2538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1842 a_68315_4045# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1843 a_45616_4727# a_45195_4727# a_44568_4052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1844 a_9210_4683# a_9206_4860# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1845 a_6712_12393# a_8208_11523# a_8159_11713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1846 a_74016_11530# a_74269_11517# a_72964_11711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1847 a_22903_10737# a_22690_10737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1848 a_1014_7698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1849 a_39053_4678# a_39140_6187# a_39095_6200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1850 a_60510_10865# a_60767_10675# a_59446_7653# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1851 a_19920_8559# a_20173_8546# a_18868_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1852 a_75853_444# a_75744_444# a_64817_433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1853 gnd d0 a_9464_12966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 a_41589_10860# a_41846_10670# a_40545_10008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1855 a_8157_7152# a_9254_6958# a_9209_6971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1856 a_23110_12257# a_22689_12257# a_22281_11941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1857 vdd d0 a_63304_11513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1858 a_29831_4183# a_30088_3993# a_28388_3239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1859 a_25648_11575# a_25227_11575# a_25549_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1860 a_79235_7006# a_79022_7006# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1861 a_54447_4154# a_55068_4046# a_55276_4046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1862 a_45617_13702# a_45196_13702# a_44569_13706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1863 a_57394_11571# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1864 a_47011_5688# a_46641_7014# a_45615_6247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1865 a_11315_2962# a_11936_3278# a_12144_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1866 vdd d1 a_51546_5515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1867 vdd a_51547_3995# a_51339_3995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1868 gnd a_84975_6950# a_84767_6950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1869 a_32990_2606# a_33609_2597# a_33817_2597# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1870 a_1228_3284# a_1015_3284# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1871 gnd a_9465_8552# a_9257_8552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1872 a_45618_10735# a_46857_10055# a_47008_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1873 a_37983_7828# a_39098_4665# a_39049_4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1874 a_34658_12247# a_34445_12247# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1875 a_17420_12387# a_18916_11517# a_18871_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1876 a_44360_4052# a_44147_4052# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1877 a_33609_4723# a_33396_4723# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1878 vdd d0 a_20170_5505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1879 a_72964_13158# a_74061_12964# a_74016_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1880 a_51292_8746# a_51549_8556# a_49845_9426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1881 gnd a_31135_5509# a_30927_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1882 a_11937_13021# a_11724_13021# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1883 a_65412_4808# a_65412_4413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1884 a_30880_13833# a_30884_12977# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1885 a_66870_10733# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1886 a_66867_7692# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1887 a_22901_2603# a_22688_2603# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1888 a_44146_5572# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1889 a_5602_7836# a_6717_4673# a_6668_4863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1890 a_8157_5705# a_8414_5515# a_6710_6385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1891 a_58673_8598# a_58460_8598# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1892 a_28386_9424# a_28643_9234# a_28343_10869# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1893 a_55067_5566# a_54854_5566# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1894 a_54856_13700# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1895 a_1437_11580# a_1016_11580# a_608_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1896 a_80133_8596# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1897 a_54447_5060# a_54447_4804# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1898 a_33608_7011# a_33395_7011# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1899 a_76527_6243# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1900 a_39096_3233# a_40588_3987# a_40539_4177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 a_60514_10688# a_60601_12197# a_60556_12210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1902 a_1230_8613# a_1017_8613# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1903 vdd d0 a_20171_3985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1904 a_3765_5569# a_3552_5569# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1905 a_6712_12393# a_8208_11523# a_8163_11536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1906 a_19916_8736# a_20173_8546# a_18868_8740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1907 a_56325_13696# a_55904_13696# a_55277_13021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1908 a_11314_8027# a_11938_8607# a_12146_8607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1909 a_1229_13027# a_1016_13027# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 gnd d0 a_31138_10676# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1911 a_82229_12208# a_83721_12962# a_83672_13152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1912 a_54857_10054# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1913 a_71520_3239# a_71773_3226# a_71473_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1914 gnd a_74268_4668# a_74060_4668# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1915 a_3767_11577# a_3554_11577# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1916 a_63052_10685# a_63305_10672# a_62004_10010# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1917 a_66240_7017# a_67080_7692# a_67288_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1918 a_83670_5697# a_84767_5503# a_84722_5516# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1919 a_22900_6249# a_22687_6249# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 a_23109_4050# a_22688_4050# a_22280_4158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1921 a_608_11943# a_608_11688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1922 a_29834_5526# a_30087_5513# a_28383_6383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1923 a_18869_5522# a_19122_5509# a_17418_6379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1924 gnd d0 a_84975_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1925 a_84722_7642# a_84718_7819# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1926 gnd a_51546_5515# a_51338_5515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1927 vdd a_9465_8552# a_9257_8552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1928 a_37983_7828# a_39098_4665# a_39053_4678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1929 a_32989_13777# a_32989_13382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1930 a_41590_7642# a_41843_7629# a_40542_6967# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1931 a_2277_12255# a_2064_12255# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1932 a_14584_11571# a_14220_10049# a_13194_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1933 a_83671_4177# a_84768_3983# a_84723_3996# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1934 a_52339_11709# a_52596_11519# a_51291_11713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1935 a_14217_7008# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1936 a_30885_10689# a_30881_10866# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1937 a_49802_10871# a_49894_9236# a_49845_9426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1938 a_9211_13658# a_11316_13779# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1939 a_51291_13160# a_51548_12970# a_49848_12216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1940 gnd d1 a_8414_6962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1941 a_76121_11935# a_76742_12251# a_76950_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1942 a_609_10423# a_1230_10739# a_1438_10739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1943 a_55905_9282# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1944 a_52337_7148# a_52594_6958# a_51289_7152# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1945 a_76948_6243# a_77788_6239# a_77996_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1946 a_55069_12253# a_54856_12253# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1947 a_82183_10863# a_82275_9228# a_82226_9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 a_72967_4006# a_73220_3993# a_71520_3239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1949 a_5602_7836# a_6717_4673# a_6672_4686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1950 a_44568_3284# a_44147_3284# a_43739_2968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1951 a_49849_9249# a_50102_9236# a_49802_10871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1952 a_23111_10737# a_22690_10737# a_22282_10816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1953 a_84718_7819# a_84975_7629# a_83674_6967# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1954 a_1014_5572# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1955 a_79024_13014# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1956 a_65414_10816# a_66035_10737# a_66243_10737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1957 vdd a_52594_7637# a_52386_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1958 gnd d1 a_19123_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1959 a_18872_10010# a_19965_10672# a_19916_10862# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1960 a_23111_9290# a_22690_9290# a_22282_9369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1961 gnd d0 a_41846_8544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1962 a_60555_3235# a_60808_3222# a_60508_4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1963 a_44362_10739# a_44149_10739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1964 vdd a_63303_2538# a_63095_2538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1965 vdd d0 a_31138_10676# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1966 a_67080_6245# a_66867_6245# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 a_36356_11569# a_35935_11569# a_36262_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1968 a_71516_3416# a_71773_3226# a_71473_4861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1969 a_13192_3274# a_12771_3274# a_12144_2599# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1970 a_79387_5561# a_79023_4039# a_77997_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1971 a_76121_13127# a_76742_13019# a_76950_13019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_63048_10862# a_63305_10672# a_62004_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1973 a_66034_11578# a_65821_11578# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1974 a_45616_3280# a_46855_4047# a_47006_5569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1975 a_35891_4039# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1976 a_47107_11577# a_46686_11577# a_47008_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1977 gnd d0 a_9463_4670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1978 a_29830_5703# a_30087_5513# a_28383_6383# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1979 a_13193_13696# a_14432_13016# a_14589_11690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1980 a_9212_9244# a_9465_9231# a_8164_8569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1981 gnd d0 a_74268_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1982 a_54446_5674# a_55067_5566# a_55275_5566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1983 a_29836_12981# a_30089_12968# a_28389_12214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1984 vdd a_31137_12964# a_30929_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1985 a_66243_10737# a_67083_10733# a_67291_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1986 a_44149_9292# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1987 a_34659_10727# a_34446_10727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1988 a_41593_10004# a_41846_9991# a_40541_10185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1989 a_32987_7119# a_33608_7011# a_33816_7011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1990 vdd a_51546_5515# a_51338_5515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1991 a_14681_5563# a_14260_5563# a_14587_5682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1992 a_8164_10016# a_9257_10678# a_9208_10868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1993 a_2278_9288# a_2065_9288# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1994 vdd d2 a_50099_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1995 a_607_3619# a_1228_4052# a_1436_4052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1996 gnd d2 a_28642_12201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1997 a_22279_7775# a_22279_7380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1998 vdd a_63304_12192# a_63096_12192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1999 a_30882_6201# a_31135_6188# a_29834_5526# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 gnd d3 a_28598_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2001 a_11935_7692# a_11722_7692# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2002 a_48173_8604# a_48310_4733# a_48518_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2003 a_1016_13706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2004 a_12145_13021# a_11724_13021# a_11316_13129# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2005 vdd d0 a_41845_12958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2006 a_49802_10871# a_49894_9236# a_49849_9249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2007 a_64708_433# a_64495_433# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2008 a_22281_13133# a_22281_12592# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2009 a_22281_13388# a_22902_13704# a_23110_13704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2010 a_54448_13129# a_55069_13021# a_55277_13021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2011 a_14683_11571# a_14262_11571# a_14589_11690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2012 gnd a_59699_7640# a_59491_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2013 a_30884_12209# a_31137_12196# a_29836_11534# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2014 a_63048_8736# a_63049_7644# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2015 a_21784_433# a_21363_433# a_11147_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2016 a_80554_8596# a_80691_4725# a_75853_444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2017 a_33396_4723# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2018 a_21363_433# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2019 a_66241_2603# a_65820_2603# a_65412_2711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2020 a_1017_10060# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2021 a_49845_9426# a_50102_9236# a_49802_10871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2022 vdd d0 a_9462_6190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2023 a_44569_13706# a_44148_13706# a_43740_13390# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2024 a_47965_8604# a_47752_8604# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2025 a_49843_3418# a_51339_2548# a_51290_2738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2026 a_33398_10731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2027 a_58460_8598# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2028 vdd d1 a_62254_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2029 a_41588_13148# a_41592_12203# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2030 vdd d0 a_41846_8544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2031 vdd d1 a_19123_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2032 gnd d1 a_30088_3993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2033 a_17423_3235# a_18915_3989# a_18866_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2034 gnd a_30089_11521# a_29881_11521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2035 a_18872_10010# a_19965_10672# a_19920_10685# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2036 a_12983_6241# a_12770_6241# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2037 a_60551_3412# a_60808_3222# a_60508_4857# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2038 a_39091_6377# a_40587_5507# a_40538_5697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2039 a_33395_7011# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2040 a_11314_5674# a_11315_5060# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2041 a_3552_5569# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2042 gnd d0 a_74270_9229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2043 a_28341_4861# a_28433_3226# a_28384_3416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2044 a_55277_13021# a_56117_13696# a_56325_13696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2045 gnd d0 a_84977_13637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2046 gnd d0 a_52597_10678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2047 a_25646_5567# a_26506_8602# a_26714_8602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2048 vdd d0 a_9463_4670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2049 a_2278_10735# a_2065_10735# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2050 a_9212_9244# a_9208_9421# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2051 gnd d2 a_28640_6193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2052 a_66240_6249# a_65819_6249# a_65411_5933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2053 gnd d0 a_31136_3221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2054 a_18870_2555# a_19963_3217# a_19914_3407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2055 a_48097_4733# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2056 a_22903_10058# a_22690_10058# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2057 a_9208_9421# a_9465_9231# a_8164_8569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2058 a_1014_7019# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2059 a_23108_5570# a_22687_5570# a_22279_5678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2060 a_76740_7690# a_76527_7690# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2061 a_44148_11580# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2062 a_46856_13022# a_46643_13022# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2063 gnd a_84975_7629# a_84767_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2064 a_25227_11575# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2065 a_52337_7148# a_52341_6203# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2066 vdd d3 a_28598_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2067 a_77998_12247# a_77577_12247# a_76950_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2068 a_51293_6975# a_52386_7637# a_52341_7650# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2069 a_56323_7688# a_57562_7008# a_57719_5682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2070 a_9210_2557# a_9463_2544# a_8158_2738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2071 vdd a_59699_7640# a_59491_7640# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2072 a_61998_2732# a_63095_2538# a_63050_2551# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2073 gnd d1 a_51549_8556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2074 a_44359_7698# a_44146_7698# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2075 a_6716_12216# a_6969_12203# a_6674_10694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2076 gnd a_8414_6962# a_8206_6962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2077 a_9210_2557# a_9206_2734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2078 a_55068_2599# a_54855_2599# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2079 a_30879_3411# a_30883_2555# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2080 gnd d1 a_73221_11521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2081 vdd a_9465_10678# a_9257_10678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2082 a_76528_3276# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2083 a_33609_4044# a_33396_4044# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2084 a_22688_4729# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2085 a_9207_13835# a_9211_12979# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2086 a_63045_7142# a_63302_6952# a_61997_7146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2087 a_41586_6372# a_41590_5516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2088 a_63046_3407# a_63303_3217# a_62002_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2089 a_19918_4677# a_20171_4664# a_18870_4002# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2090 a_28347_10692# a_28434_12201# a_28385_12391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2091 vdd a_30089_11521# a_29881_11521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2092 gnd d0 a_63305_9225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2093 a_46854_7014# a_46641_7014# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2094 a_28341_4861# a_28433_3226# a_28388_3239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2095 a_40540_13152# a_41637_12958# a_41592_12971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2096 a_33608_7690# a_33395_7690# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2097 a_66241_4729# a_67081_4725# a_67289_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2098 gnd a_41846_8544# a_41638_8544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2099 a_84722_6963# a_84975_6950# a_83670_7144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2100 a_55275_6245# a_54854_6245# a_54446_5929# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2101 gnd a_19123_2542# a_18915_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2102 a_22689_13704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2103 a_54856_13021# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2104 a_54449_9621# a_54449_9365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2105 a_41587_4173# a_41591_3228# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2106 vdd d0 a_31136_3221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2107 vdd d0 a_31135_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2108 a_68572_11575# a_68359_11575# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2109 gnd a_9463_4670# a_9255_4670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2110 gnd d0 a_31138_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2111 a_24156_6245# a_25395_7012# a_25552_5686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2112 gnd d0 a_74267_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2113 gnd a_74268_3989# a_74060_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2114 a_65413_13388# a_65413_13133# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2115 a_63052_10006# a_63305_9993# a_62000_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2116 a_65412_2711# a_65414_2612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2117 a_2484_4727# a_2063_4727# a_1436_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2118 a_76119_6322# a_76119_5927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2119 a_65821_12257# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2120 gnd d1 a_19124_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2121 a_2065_9288# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2122 a_607_5066# a_1227_5572# a_1435_5572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2123 vdd a_62256_12964# a_62048_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2124 a_35935_11569# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2125 a_83673_8738# a_84770_8544# a_84721_8734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2126 a_55904_13696# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2127 gnd a_17675_6189# a_17467_6189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2128 a_9206_2734# a_9463_2544# a_8158_2738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2129 a_608_13785# a_1229_13706# a_1437_13706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2130 a_83676_12975# a_84769_13637# a_84720_13827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2131 a_67082_12253# a_66869_12253# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2132 vdd d1 a_51549_8556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2133 a_76122_11066# a_76122_10810# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2134 a_29833_10191# a_30930_9997# a_30885_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2135 a_11722_7692# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2136 a_54447_4409# a_54447_4154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2137 a_9212_10691# a_9208_10868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2138 gnd d2 a_6967_6195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2139 vdd d1 a_73221_11521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2140 a_14220_10049# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2141 a_55278_9286# a_56118_9282# a_56326_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2142 a_76742_12251# a_76529_12251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2143 a_23110_13704# a_22689_13704# a_22281_13388# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2144 a_57714_5563# a_57350_4041# a_56324_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2145 a_609_9627# a_1230_10060# a_1438_10060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2146 a_34445_12247# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2147 vdd d1 a_83930_9995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2148 a_19914_4854# a_20171_4664# a_18870_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2149 vdd a_41845_13637# a_41637_13637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2150 a_41593_10004# a_41589_10181# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2151 vdd d0 a_63305_9225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2152 a_47752_8604# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2153 vdd a_9462_6190# a_9254_6190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2154 a_11315_4409# a_11936_4725# a_12144_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2155 a_8160_10193# a_8417_10003# a_6717_9249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2156 a_33397_13698# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2157 vdd a_62254_6956# a_62046_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2158 a_17380_4680# a_17467_6189# a_17422_6202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2159 a_56323_6241# a_55902_6241# a_55275_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2160 a_76529_11572# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2161 a_17418_6379# a_18914_5509# a_18865_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2162 a_23111_10058# a_22690_10058# a_22282_10166# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2163 vdd a_41846_8544# a_41638_8544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2164 vdd a_19123_2542# a_18915_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2165 a_84722_5516# a_84718_5693# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2166 a_12770_6241# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2167 a_52338_4860# a_52342_4004# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2168 vdd d2 a_17677_12197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2169 a_32989_11680# a_32990_11066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2170 a_65414_10166# a_66035_10058# a_66243_10058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2171 gnd a_30087_6960# a_29879_6960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2172 a_3881_11696# a_3511_13022# a_2485_13702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2173 a_32399_444# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2174 a_6715_3241# a_8207_3995# a_8158_4185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2175 a_68570_5567# a_68357_5567# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2176 a_18868_10187# a_19965_9993# a_19916_10183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2177 vdd d0 a_84978_9991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2178 a_76742_13019# a_76529_13019# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2179 gnd d1 a_40795_6954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2180 gnd d0 a_63303_2538# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2181 vdd a_9463_4670# a_9255_4670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2182 a_56326_10729# a_55905_10729# a_55278_10054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2183 gnd a_31136_3221# a_30928_3221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2184 a_24156_6245# a_23735_6245# a_23108_5570# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2185 a_8162_2561# a_9255_3223# a_9206_3413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2186 gnd d0 a_9463_3991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2187 a_25398_10053# a_25185_10053# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2188 a_77996_6239# a_77575_6239# a_76948_5564# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2189 a_32988_2960# a_32988_2705# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2190 a_83673_8738# a_84770_8544# a_84725_8557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2191 a_76951_8605# a_76530_8605# a_76122_8713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2192 a_8160_10193# a_9257_9999# a_9208_10189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2193 a_29837_8567# a_30090_8554# a_28386_9424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2194 a_12145_13700# a_11724_13700# a_11316_13779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2195 a_77790_12247# a_77577_12247# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2196 a_1016_13027# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2197 a_22903_9290# a_22690_9290# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2198 a_40543_2553# a_40796_2540# a_39092_3410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 a_25396_4045# a_25183_4045# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2200 a_39055_10686# a_39308_10673# a_37987_7651# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2201 a_76120_4152# a_76120_3611# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2202 a_76119_5927# a_76119_5672# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2203 a_22281_12592# a_22902_13025# a_23110_13025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2204 a_43741_11074# a_44361_11580# a_44569_11580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2205 a_12984_3274# a_12771_3274# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2206 gnd d0 a_41844_4662# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2207 a_33396_4044# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2208 a_33608_5564# a_33395_5564# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2209 a_25549_11575# a_25440_11575# a_25648_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2210 a_17420_12387# a_18916_11517# a_18867_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2211 vdd a_52597_10678# a_52389_10678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2212 a_44567_7698# a_45407_7694# a_45615_7694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2213 a_54447_2962# a_55068_3278# a_55276_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2214 a_44569_13027# a_44148_13027# a_43740_12594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2215 gnd a_63305_9225# a_63097_9225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2216 a_30884_12209# a_30880_12386# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2217 a_609_9371# a_1230_9292# a_1438_9292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2218 a_22282_2612# a_22901_2603# a_23109_2603# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2219 gnd a_20172_12192# a_19964_12192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2220 a_33398_10052# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2221 a_2277_13702# a_2064_13702# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2222 gnd d0 a_74270_10676# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2223 a_57815_11571# a_58673_8598# a_58881_8598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2224 a_33395_7690# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2225 a_33817_3276# a_34657_3272# a_34865_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2226 a_22279_5678# a_22280_5064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2227 a_23110_11578# a_23950_12253# a_24158_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2228 a_29834_5526# a_30927_6188# a_30878_6378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2229 vdd a_31135_6956# a_30927_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2230 vdd a_31136_3221# a_30928_3221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2231 a_57721_11690# a_57351_13016# a_56325_13696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2232 gnd d0 a_84977_12958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2233 gnd d0 a_52597_9999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2234 a_82230_9241# a_83722_9995# a_83677_10008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2235 a_1435_6251# a_1014_6251# a_606_6330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2236 a_41592_13650# a_43740_13785# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2237 a_8162_2561# a_9255_3223# a_9210_3236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2238 a_1017_8613# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2239 gnd a_71730_4671# a_71522_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2240 a_44568_4731# a_44147_4731# a_43739_4415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2241 gnd a_74267_5509# a_74059_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2242 a_47105_5569# a_46684_5569# a_47006_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2243 a_36255_5561# a_36146_5561# a_36354_5561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2244 a_32989_11935# a_33610_12251# a_33818_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2245 a_75853_444# a_80478_4725# a_80800_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_22279_6328# a_22900_6249# a_23108_6249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2247 gnd d1 a_62257_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2248 a_66033_2603# a_65820_2603# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2249 a_11937_12253# a_11724_12253# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2250 a_34446_10727# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2251 a_29833_8744# a_30090_8554# a_28386_9424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2252 a_33816_7690# a_33395_7690# a_32987_7374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2253 a_17382_10688# a_17469_12197# a_17424_12210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2254 a_67083_9286# a_66870_9286# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2255 gnd a_8416_11523# a_8208_11523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2256 a_40539_2730# a_40796_2540# a_39092_3410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2257 a_75531_444# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2258 a_51294_4008# a_51547_3995# a_49847_3241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2259 a_13192_4721# a_12771_4721# a_12144_4046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2260 a_39051_10863# a_39308_10673# a_37987_7651# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2261 a_54446_8027# a_55070_8607# a_55278_8607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2262 a_1435_7019# a_1014_7019# a_606_6586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2263 gnd a_6967_6195# a_6759_6195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2264 a_39097_12208# a_39350_12195# a_39055_10686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2265 a_52343_11532# a_52596_11519# a_51291_11713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_63048_10862# a_63052_10006# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2267 gnd a_40798_9995# a_40590_9995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2268 vdd d0 a_41844_4662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2269 a_72962_5703# a_74059_5509# a_74014_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2270 a_1229_12259# a_1016_12259# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2271 a_18865_7146# a_19122_6956# a_17422_6202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2272 a_32989_13127# a_33610_13019# a_33818_13019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2273 a_37214_8596# a_37001_8596# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2274 a_66032_6249# a_65819_6249# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2275 a_52342_3236# a_52595_3223# a_51294_2561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2276 a_5287_4733# a_5178_4733# a_5386_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2277 vdd a_63305_9225# a_63097_9225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2278 a_22688_4050# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2279 a_30884_13656# a_32989_13777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2280 a_58881_8598# a_58460_8598# a_57815_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2281 a_45407_6247# a_45194_6247# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2282 a_19918_3998# a_20171_3985# a_18866_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2283 vdd d0 a_74270_10676# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2284 gnd a_71772_6193# a_71564_6193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2285 a_30882_7648# a_31135_7635# a_29834_6973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2286 vdd a_82480_6187# a_82272_6187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2287 a_68316_13020# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2288 a_63047_11703# a_63052_10685# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2289 a_84722_7642# a_84975_7629# a_83674_6967# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2290 a_44362_8613# a_44149_8613# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2291 a_24157_4725# a_25396_4045# a_25547_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2292 gnd d2 a_82480_6187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2293 gnd a_52594_7637# a_52386_7637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2294 a_57349_7008# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2295 a_22689_13025# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2296 a_23109_2603# a_23949_3278# a_24157_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2297 a_30884_13656# a_31137_13643# a_29836_12981# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2298 a_70092_4731# a_70456_7644# a_70407_7834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2299 a_77791_10727# a_77578_10727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2300 a_3725_10055# a_3512_10055# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2301 a_41589_8734# a_41590_7642# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2302 gnd a_40795_6954# a_40587_6954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2303 gnd a_63303_2538# a_63095_2538# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2304 vdd a_71730_4671# a_71522_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2305 a_12985_12249# a_12772_12249# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2306 a_79237_13014# a_79024_13014# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2307 vdd d4 a_38240_7638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2308 a_51295_11536# a_52388_12198# a_52343_12211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2309 a_12145_11574# a_11724_11574# a_11317_11068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2310 gnd a_9463_3991# a_9255_3991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2311 a_76121_13127# a_76121_12586# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2312 a_62004_8563# a_63097_9225# a_63048_9415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2313 a_82223_6377# a_83719_5507# a_83674_5520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2314 a_46643_13022# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2315 vdd a_8416_11523# a_8208_11523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2316 a_60552_12387# a_62048_11517# a_62003_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2317 a_66243_9290# a_65822_9290# a_65414_9369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2318 gnd d0 a_84978_8544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2319 a_608_13135# a_1229_13027# a_1437_13027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2320 a_83672_13152# a_84769_12958# a_84720_13148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2321 vdd d0 a_9464_12198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2322 a_76950_13698# a_76529_13698# a_76121_13777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2323 a_22690_9290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2324 a_41593_8557# a_41846_8544# a_40541_8738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2325 a_65411_8031# a_65411_7775# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2326 a_56324_3274# a_55903_3274# a_55276_2599# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2327 a_23109_3282# a_22688_3282# a_22280_3361# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2328 a_25183_4045# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2329 a_76530_10731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2330 a_79023_4039# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2331 a_52338_3413# a_52595_3223# a_51294_2561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2332 a_12771_3274# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2333 gnd a_41844_4662# a_41636_4662# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2334 a_33395_5564# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2335 a_36146_5561# a_35933_5561# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2336 a_23110_13025# a_22689_13025# a_22281_12592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2337 a_43739_2968# a_44360_3284# a_44568_3284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2338 a_42796_401# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2339 a_81119_7651# a_82232_10673# a_82183_10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2340 a_36103_7006# a_35890_7006# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2341 a_2276_3280# a_2063_3280# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2342 a_11315_3613# a_11936_4046# a_12144_4046# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2343 a_57813_5563# a_57392_5563# a_57719_5682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2344 a_77998_13694# a_77577_13694# a_76950_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2345 a_30878_7825# a_31135_7635# a_29834_6973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2346 a_30878_7146# a_30882_6201# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2347 a_76119_6322# a_76740_6243# a_76948_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2348 a_32987_5927# a_33608_6243# a_33816_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2349 a_1437_12259# a_2277_12255# a_2485_12255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2350 a_57719_5682# a_57349_7008# a_56323_7688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2351 a_74014_6201# a_74267_6188# a_72966_5526# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2352 a_26638_4731# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2353 a_23951_10733# a_23738_10733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2354 a_30880_13833# a_31137_13643# a_29836_12981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2355 a_70092_4731# a_70456_7644# a_70411_7657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2356 a_12143_5566# a_12983_6241# a_13191_6241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2357 a_36257_11569# a_35893_10047# a_34867_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2358 a_37559_4725# a_37346_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2359 a_25397_13020# a_25184_13020# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2360 a_76122_10415# a_76122_10160# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2361 a_17378_10865# a_17470_9230# a_17421_9420# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2362 a_43739_3363# a_43739_2968# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2363 a_77999_10727# a_79238_10047# a_79389_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2364 gnd d4 a_59699_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2365 a_76528_4723# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2366 a_54448_11937# a_55069_12253# a_55277_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2367 a_84724_11524# a_84977_11511# a_83672_11705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2368 a_23111_8611# a_22690_8611# a_22279_8031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2369 a_57565_10049# a_57352_10049# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2370 a_9208_9421# a_9212_8565# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2371 a_54446_6324# a_54446_5929# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2372 a_62004_8563# a_63097_9225# a_63052_9238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2373 a_65820_2603# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2374 a_55278_9286# a_54857_9286# a_54449_9365# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2375 a_39095_6200# a_40587_6954# a_40542_6967# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2376 vdd d0 a_84978_8544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2377 a_76527_7011# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2378 a_41589_8734# a_41846_8544# a_40541_8738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2379 a_51293_6975# a_52386_7637# a_52337_7827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2380 vdd a_41844_4662# a_41636_4662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2381 gnd d0 a_74268_3221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2382 a_61998_2732# a_63095_2538# a_63046_2728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2383 a_19919_12973# a_19915_13150# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2384 a_72969_10014# a_73222_10001# a_71522_9247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2385 gnd a_84978_10670# a_84770_10670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2386 a_28387_6206# a_28640_6193# a_28345_4684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2387 a_63050_3230# a_63046_3407# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2388 a_45616_3280# a_45195_3280# a_44568_3284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2389 a_22900_7017# a_22687_7017# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2390 a_62001_6969# a_62254_6956# a_60554_6202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2391 a_39091_6377# a_39348_6187# a_39053_4678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2392 gnd d0 a_41844_3983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2393 a_81119_7651# a_82232_10673# a_82187_10686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2394 gnd a_9465_10678# a_9257_10678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2395 a_12986_10729# a_12773_10729# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2396 a_44570_10739# a_45410_10735# a_45618_10735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 a_62004_10010# a_63097_10672# a_63048_10862# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2398 a_22687_5570# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2399 a_65821_13704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2400 a_76121_12586# a_76121_12330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2401 a_19917_5518# a_20170_5505# a_18865_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2402 a_45194_6247# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2403 a_63050_3230# a_63303_3217# a_62002_2555# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2404 a_9211_12211# a_9207_12388# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2405 a_1436_3284# a_1015_3284# a_607_2968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2406 a_13193_12249# a_12772_12249# a_12145_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2407 a_54279_446# a_53858_446# a_54180_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2408 gnd d0 a_74270_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2409 a_17378_10865# a_17470_9230# a_17425_9243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2410 a_11048_446# a_10939_446# a_11147_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2411 vdd d0 a_20172_12960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2412 vdd d4 a_59699_7640# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2413 a_84720_11701# a_84977_11511# a_83672_11705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2414 a_30881_10187# a_31138_9997# a_29833_10191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2415 vdd d1 a_40798_8548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2416 a_83672_13152# a_83929_12962# a_82229_12208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2417 a_33610_11572# a_33397_11572# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2418 a_23948_7692# a_23735_7692# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2419 a_55069_13021# a_54856_13021# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2420 a_33816_5564# a_34656_6239# a_34864_6239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2421 a_76950_11572# a_76529_11572# a_76122_11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2422 a_40545_8561# a_41638_9223# a_41589_9413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2423 gnd d0 a_52597_9231# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2424 a_33609_3276# a_33396_3276# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2425 a_32988_3611# a_32988_3355# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2426 a_44568_4052# a_44147_4052# a_43739_3619# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2427 a_11725_10733# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2428 a_18872_10010# a_19125_9997# a_17425_9243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2429 a_52344_8565# a_52340_8742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2430 a_30879_4858# a_30883_4002# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2431 a_56115_7688# a_55902_7688# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2432 a_28390_9247# a_29882_10001# a_29833_10191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2433 gnd a_84978_8544# a_84770_8544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2434 a_44567_7698# a_44146_7698# a_43738_7777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2435 a_49848_12216# a_50101_12203# a_49806_10694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2436 a_1438_10060# a_2278_10735# a_2486_10735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2437 a_66243_10737# a_65822_10737# a_65414_10421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2438 a_41586_7819# a_41590_6963# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2439 a_54856_12253# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2440 a_24159_9286# a_23738_9286# a_23111_9290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2441 a_54854_6245# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2442 vdd d0 a_74268_3221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2443 a_34865_3272# a_34444_3272# a_33817_2597# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2444 a_34444_4719# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2445 a_39098_9241# a_40590_9995# a_40541_10185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2446 vdd d0 a_74267_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2447 a_55276_2599# a_54855_2599# a_54447_2707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2448 a_54447_4154# a_54447_3613# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2449 vdd a_84978_10670# a_84770_10670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2450 a_1438_8613# a_1017_8613# a_606_8033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2451 a_74010_5699# a_74015_4681# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2452 a_48734_7836# a_49849_4673# a_49800_4863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2453 a_36148_11569# a_35935_11569# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2454 vdd d3 a_60765_4667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2455 a_62004_10010# a_63097_10672# a_63052_10685# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2456 a_67288_6245# a_68527_7012# a_68684_5686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2457 gnd d1 a_8416_12970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2458 a_79488_11569# a_79067_11569# a_79389_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 a_46897_5569# a_46684_5569# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2460 a_13191_7688# a_12770_7688# a_12143_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2461 a_2063_3280# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2462 a_11315_5060# a_11935_5566# a_12143_5566# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2463 gnd a_41845_13637# a_41637_13637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2464 a_72965_8744# a_74062_8550# a_74013_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2465 a_54449_10162# a_54449_9621# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2466 a_32990_9363# a_32990_8968# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2467 a_4833_8604# a_4620_8604# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2468 a_1015_4731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2469 a_14681_5563# a_15541_8598# a_15749_8598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2470 a_30882_6969# a_31135_6956# a_29830_7150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2471 a_34446_9280# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2472 a_68530_10053# a_68317_10053# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2473 gnd a_52594_6958# a_52386_6958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2474 vdd d1 a_51547_2548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2475 a_12984_4721# a_12771_4721# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2476 a_30884_12977# a_31137_12964# a_29832_13158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2477 a_72964_11711# a_74061_11517# a_74016_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2478 a_6714_6208# a_6967_6195# a_6672_4686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2479 a_63049_6197# a_63045_6374# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2480 gnd a_28642_12201# a_28434_12201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2481 vdd a_28600_10679# a_28392_10679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2482 a_40545_8561# a_41638_9223# a_41593_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2483 vdd d0 a_52597_9231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2484 a_71521_12214# a_73013_12968# a_72968_12981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2485 a_57815_11571# a_57394_11571# a_57716_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2486 a_17422_6202# a_18914_6956# a_18869_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2487 vdd d1 a_30087_6960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2488 a_54447_4409# a_55068_4725# a_55276_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2489 a_40544_12975# a_40797_12962# a_39097_12208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2490 vdd d2 a_71774_12201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2491 a_49804_4686# a_49891_6195# a_49842_6385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2492 vdd d1 a_62255_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2493 a_22281_11686# a_22902_11578# a_23110_11578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2494 vdd a_84978_8544# a_84770_8544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2495 a_55902_6241# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2496 vdd d0 a_20171_2538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2497 gnd a_73220_3993# a_73012_3993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2498 gnd d1 a_73220_2546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2499 a_29834_6973# a_30927_7635# a_30878_7825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2500 a_82185_4678# a_82272_6187# a_82223_6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2501 a_40539_2730# a_41636_2536# a_41587_2726# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2502 gnd d0 a_52595_2544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2503 a_36104_4039# a_35891_4039# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2504 a_76950_13019# a_76529_13019# a_76121_13127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2505 a_39093_12385# a_40589_11515# a_40540_11705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2506 gnd d1 a_83927_6954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2507 a_8158_2738# a_8415_2548# a_6711_3418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2508 a_48734_7836# a_49849_4673# a_49804_4686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2509 a_22282_8974# a_22903_9290# a_23111_9290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2510 gnd a_74268_3221# a_74060_3221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2511 a_32988_3355# a_33609_3276# a_33817_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2512 a_1227_7698# a_1014_7698# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2513 a_66240_7017# a_65819_7017# a_65411_6584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2514 a_80691_4725# a_80478_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2515 a_44360_4731# a_44147_4731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2516 gnd d1 a_8417_8556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2517 a_41592_12203# a_41845_12190# a_40544_11528# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2518 a_76530_10052# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2519 a_67288_6245# a_66867_6245# a_66240_5570# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2520 gnd a_41844_3983# a_41636_3983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2521 gnd d0 a_41843_5503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2522 a_65413_11941# a_65413_11686# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2523 a_32612_444# a_32399_444# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2524 a_72965_8744# a_74062_8550# a_74017_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2525 a_2486_9288# a_2065_9288# a_1438_8613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2526 a_36262_11688# a_35892_13014# a_34866_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2527 gnd a_52597_10678# a_52389_10678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2528 a_63047_12382# a_63051_11526# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2529 a_9209_6203# a_9462_6190# a_8161_5528# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2530 a_21784_433# a_43009_401# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2531 a_14582_5563# a_14473_5563# a_14681_5563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2532 vref a_608_13785# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2533 a_45410_9288# a_45197_9288# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2534 a_3722_7014# a_3509_7014# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2535 a_11315_3357# a_11315_2962# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2536 gnd d4 a_16567_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2537 a_22901_3282# a_22688_3282# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2538 a_66035_9290# a_65822_9290# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2539 vdd a_82483_9228# a_82275_9228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2540 vdd a_40798_8548# a_40590_8548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2541 a_2275_6247# a_2062_6247# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2542 a_1229_13706# a_1016_13706# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2543 gnd d0 a_63305_10672# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2544 a_68528_4045# a_68315_4045# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2545 a_1016_12259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2546 gnd d2 a_17678_9230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2547 gnd d0 a_84976_4662# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 a_62000_10187# a_62257_9997# a_60557_9243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2549 a_34659_9280# a_34446_9280# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2550 a_23735_7692# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2551 a_44147_3284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2552 a_76528_4044# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2553 vdd a_20172_13639# a_19964_13639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2554 a_41591_4675# a_41844_4662# a_40543_4000# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2555 a_44567_5572# a_44146_5572# a_43739_5066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2556 a_11317_9365# a_11938_9286# a_12146_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2557 a_15541_8598# a_15328_8598# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2558 a_33396_3276# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2559 a_14218_4041# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2560 a_33818_13698# a_34658_13694# a_34866_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2561 a_34656_7686# a_34443_7686# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2562 a_65414_2612# a_66033_2603# a_66241_2603# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2563 vdd d1 a_73220_2546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2564 a_32990_8713# a_33611_8605# a_33819_8605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2565 a_606_6330# a_606_5935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2566 a_44569_12259# a_44148_12259# a_43740_12338# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2567 a_29834_6973# a_30927_7635# a_30882_7648# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2568 a_76527_7690# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2569 a_55275_7013# a_54854_7013# a_54446_6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2570 a_76949_3276# a_77789_3272# a_77997_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2571 a_40539_2730# a_41636_2536# a_41591_2549# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2572 vdd d0 a_52595_2544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2573 a_23109_4050# a_23949_4725# a_24157_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2574 vdd d1 a_51548_12970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2575 a_39093_12385# a_40589_11515# a_40544_11528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2576 a_82226_9418# a_83722_8548# a_83677_8561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2577 a_63050_3998# a_63046_4175# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2578 a_19919_13652# a_19915_13829# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2579 a_22902_12257# a_22689_12257# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2580 vdd a_74268_3221# a_74060_3221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2581 vdd d0 a_31136_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2582 a_51289_7152# a_52386_6958# a_52337_7148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2583 vdd a_74267_6956# a_74059_6956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2584 vdd d1 a_8417_8556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2585 a_24159_9286# a_25398_10053# a_25549_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2586 a_79387_5561# a_79278_5561# a_79486_5561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2587 a_71479_10692# a_71566_12201# a_71521_12214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2588 vdd a_31137_11517# a_30929_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2589 gnd a_84978_9991# a_84770_9991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2590 a_22903_8611# a_22690_8611# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2591 a_62004_8563# a_62257_8550# a_60553_9420# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2592 a_22689_11578# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2593 a_77996_6239# a_79235_7006# a_79392_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2594 a_65411_6328# a_66032_6249# a_66240_6249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2595 a_46684_5569# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2596 gnd a_9465_9999# a_9257_9999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2597 a_62000_10187# a_63097_9993# a_63048_10183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2598 a_65821_13025# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2599 vdd a_41846_9991# a_41638_9991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2600 a_4620_8604# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2601 a_76948_7690# a_76527_7690# a_76119_7374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2602 a_55070_8607# a_54857_8607# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2603 a_54448_13384# a_54448_13129# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2604 vdd d4 a_16567_7640# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2605 a_43741_11074# a_43741_10818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2606 a_33398_8605# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2607 a_56324_4721# a_55903_4721# a_55276_4046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2608 vdd d0 a_63305_10672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2609 vdd d2 a_17678_9230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2610 vdd d0 a_84976_4662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2611 a_76121_13382# a_76742_13698# a_76950_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2612 vdd a_51547_2548# a_51339_2548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2613 a_12771_4721# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2614 a_17382_10688# a_17635_10675# a_16314_7653# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2615 vdd d2 a_50100_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2616 a_41587_4852# a_41844_4662# a_40543_4000# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2617 a_76122_8968# a_76743_9284# a_76951_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2618 a_55069_13700# a_54856_13700# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2619 a_65413_13783# a_65413_13388# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2620 a_62003_12977# a_62256_12964# a_60556_12210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2621 vdd a_63304_12960# a_63096_12960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2622 a_48173_8604# a_47752_8604# a_47107_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2623 gnd d4 a_38240_7638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2624 vdd d1 a_62254_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2625 vdd a_39350_12195# a_39142_12195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2626 vdd a_62255_3989# a_62047_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2627 a_1437_13706# a_2277_13702# a_2485_13702# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2628 a_6714_6208# a_8206_6962# a_8161_6975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2629 a_71475_10869# a_71732_10679# a_70411_7657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2630 a_11725_10054# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2631 a_74014_7648# a_74267_7635# a_72966_6973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2632 gnd a_83929_11515# a_83721_11515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2633 a_30881_9419# a_30885_8563# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2634 a_1435_6251# a_2275_6247# a_2483_6247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2635 gnd a_20171_4664# a_19963_4664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2636 a_67289_4725# a_68528_4045# a_68679_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2637 a_54447_4804# a_54447_4409# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2638 a_60552_12387# a_62048_11517# a_61999_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2639 a_11147_446# a_10726_446# a_5386_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2640 gnd d0 a_31137_12196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2641 a_66243_10058# a_65822_10058# a_65414_9625# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2642 a_44567_7019# a_44146_7019# a_43738_7127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2643 gnd d0 a_63302_6184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2644 a_66241_2603# a_67081_3278# a_67289_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2645 a_11315_2707# a_11936_2599# a_12144_2599# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2646 a_24159_10733# a_23738_10733# a_23111_10058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2647 vdd d0 a_9462_6958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2648 gnd a_83927_6954# a_83719_6954# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2649 a_1228_2605# a_1015_2605# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2650 a_63051_12205# a_63304_12192# a_62003_11530# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2651 gnd a_8417_8556# a_8209_8556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2652 a_62000_8740# a_62257_8550# a_60553_9420# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2653 gnd a_41843_5503# a_41635_5503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2654 a_11317_11068# a_11937_11574# a_12145_11574# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2655 a_33819_10731# a_33398_10731# a_32990_10415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2656 a_607_4160# a_607_3619# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2657 a_606_5935# a_606_5680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2658 vdd a_17677_12197# a_17469_12197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2659 a_54449_10812# a_54449_10417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2660 a_41589_10181# a_41593_9236# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2661 a_34864_6239# a_34443_6239# a_33816_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2662 a_3874_5569# a_3510_4047# a_2484_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2663 a_1229_11580# a_1016_11580# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2664 a_79067_11569# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2665 a_39094_9418# a_39351_9228# a_39051_10863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2666 gnd a_41845_12958# a_41637_12958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2667 a_66241_3282# a_65820_3282# a_65412_2966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2668 a_1015_4052# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2669 a_23951_9286# a_23738_9286# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2670 a_30885_8563# a_31138_8550# a_29833_8744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2671 a_71519_6206# a_73011_6960# a_72962_7150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2672 a_44359_6251# a_44146_6251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2673 gnd a_16567_7640# a_16359_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2674 a_65822_9290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2675 a_84725_8557# a_84978_8544# a_83673_8738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2676 a_608_11943# a_1229_12259# a_1437_12259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2677 a_17378_10865# a_17635_10675# a_16314_7653# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2678 a_2062_6247# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2679 a_68315_4045# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2680 gnd a_52597_8552# a_52389_8552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2681 a_45616_4727# a_45195_4727# a_44568_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2682 vdd a_6969_12203# a_6761_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2683 a_22903_10737# a_22690_10737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2684 a_45197_9288# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2685 a_55903_3274# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2686 a_82228_3233# a_82481_3220# a_82181_4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2687 gnd a_84976_4662# a_84768_4662# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 vdd a_74269_12196# a_74061_12196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2689 a_22688_3282# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2690 a_76527_5564# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2691 a_23110_12257# a_22689_12257# a_22281_12336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2692 a_25648_11575# a_25227_11575# a_25554_11694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2693 a_79235_7006# a_79022_7006# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2694 a_56324_4721# a_57563_4041# a_57714_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_52340_10868# a_52597_10678# a_51296_10016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2696 a_22282_8719# a_22279_8031# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2697 a_74010_7825# a_74267_7635# a_72966_6973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2698 a_71477_4684# a_71564_6193# a_71519_6206# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2699 a_54447_3613# a_55068_4046# a_55276_4046# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2700 a_1436_4731# a_1015_4731# a_607_4415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2701 a_13193_13696# a_12772_13696# a_12145_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2702 vdd a_83929_11515# a_83721_11515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2703 a_43738_7127# a_43738_6586# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2704 vdd a_20171_4664# a_19963_4664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2705 a_22281_13388# a_22281_13133# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2706 gnd a_20172_12960# a_19964_12960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2707 a_65413_12336# a_66034_12257# a_66242_12257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2708 a_57394_11571# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2709 a_68686_11694# a_68572_11575# a_68780_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2710 a_12983_7688# a_12770_7688# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2711 a_47011_5688# a_46641_7014# a_45615_7694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2712 a_9207_13156# a_9464_12966# a_8159_13160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2713 a_18871_11530# a_19964_12192# a_19915_12382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2714 a_44361_12259# a_44148_12259# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2715 vdd d0 a_84977_12190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2716 a_15328_8598# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2717 a_76122_2606# a_76741_2597# a_76949_2597# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2718 a_46899_11577# a_46686_11577# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2719 vdd d0 a_63302_6184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2720 a_29830_7150# a_30927_6956# a_30878_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2721 vdd d0 a_31135_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2722 a_18865_5699# a_19962_5505# a_19917_5518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2723 vdd a_31136_3989# a_30928_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2724 a_45618_9288# a_46857_10055# a_47008_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2725 vdd a_8417_8556# a_8209_8556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2726 a_74010_6378# a_74014_5522# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2727 a_84720_13827# a_84724_12971# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2728 a_19919_11526# a_20172_11513# a_18867_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2729 a_8158_4185# a_9255_3991# a_9210_4004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2730 a_68778_5567# a_68357_5567# a_68679_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2731 a_74012_13154# a_74016_12209# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2732 a_66242_12257# a_67082_12253# a_67290_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2733 a_66243_8611# a_65822_8611# a_65411_8031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2734 a_33816_7011# a_34656_7686# a_34864_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2735 a_44360_4052# a_44147_4052# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2736 a_34658_12247# a_34445_12247# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2737 a_33609_4723# a_33396_4723# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2738 a_22690_8611# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2739 a_8163_11536# a_9256_12198# a_9207_12388# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2740 a_45409_12255# a_45196_12255# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2741 a_30885_8563# a_30881_8740# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2742 a_22279_7125# a_22900_7017# a_23108_7017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2743 a_11937_13021# a_11724_13021# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2744 vdd a_62256_11517# a_62048_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2745 a_52342_4004# a_52338_4181# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2746 a_51289_7152# a_51546_6962# a_49846_6208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2747 a_18866_4179# a_19963_3985# a_19918_3998# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2748 a_76121_11680# a_76742_11572# a_76950_11572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2749 a_74013_10187# a_74270_9997# a_72965_10191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2750 a_54857_9286# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2751 a_74011_4179# a_74015_3234# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2752 gnd a_52597_9999# a_52389_9999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2753 a_30881_8740# a_31138_8550# a_29833_8744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2754 a_13191_7688# a_14430_7008# a_14587_5682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2755 a_29836_11534# a_30929_12196# a_30880_12386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2756 a_84721_8734# a_84978_8544# a_83673_8738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2757 vdd a_16567_7640# a_16359_7640# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2758 a_54446_7771# a_54446_7376# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2759 a_55069_11574# a_54856_11574# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 a_84719_2726# a_76122_2606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2761 a_22280_3361# a_22280_2966# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2762 a_3765_5569# a_3552_5569# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2763 a_1230_8613# a_1017_8613# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2764 gnd a_30090_8554# a_29882_8554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2765 vdd a_52597_8552# a_52389_8552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2766 a_82224_3410# a_82481_3220# a_82181_4855# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2767 vdd a_84976_4662# a_84768_4662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2768 a_18866_4179# a_19123_3989# a_17423_3235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2769 gnd d1 a_40798_8548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2770 a_19914_3407# a_20171_3217# a_18870_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2771 a_1229_13027# a_1016_13027# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2772 a_48738_7659# a_49851_10681# a_49802_10871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2773 gnd d0 a_63305_9993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 a_19913_7142# a_20170_6952# a_18865_7146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2775 a_66032_7017# a_65819_7017# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2776 gnd d0 a_84976_3983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2777 a_33397_12251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2778 a_3767_11577# a_3554_11577# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2779 gnd d0 a_20173_9225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2780 a_65819_5570# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2781 a_22900_6249# a_22687_6249# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2782 a_41591_3996# a_41844_3983# a_40539_4177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2783 vdd a_62254_5509# a_62046_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2784 a_12143_6245# a_11722_6245# a_11314_5929# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2785 a_63050_4677# a_63046_4854# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2786 a_84725_10683# a_84721_10860# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2787 a_72967_4006# a_74060_4668# a_74015_4681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2788 a_24158_13700# a_25397_13020# a_25554_11694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2789 gnd d0 a_52596_12198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2790 a_82225_12385# a_82482_12195# a_82187_10686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2791 a_49842_6385# a_50099_6195# a_49804_4686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2792 a_14584_11571# a_14220_10049# a_13194_10729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2793 a_2277_12255# a_2064_12255# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2794 a_14217_7008# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2795 gnd a_63302_6184# a_63094_6184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2796 a_77997_4719# a_79236_4039# a_79387_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2797 a_19915_11703# a_20172_11513# a_18867_11707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2798 vdd a_9462_6958# a_9254_6958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2799 a_41590_6195# a_41586_6372# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2800 a_56326_10729# a_57565_10049# a_57716_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2801 a_51292_8746# a_52389_8552# a_52340_8742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2802 a_54071_446# a_53858_446# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2803 a_55278_10733# a_54857_10733# a_54449_10417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2804 vdd d1 a_8417_10003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2805 a_8157_5705# a_9254_5511# a_9205_5701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2806 a_76948_5564# a_77788_6239# a_77996_6239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2807 a_33818_13698# a_33397_13698# a_32989_13382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2808 a_60551_3412# a_62047_2542# a_61998_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2809 gnd d3 a_60765_4667# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2810 a_43740_13135# a_43740_12594# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2811 a_83676_11528# a_84769_12190# a_84724_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2812 a_607_2968# a_1228_3284# a_1436_3284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2813 a_67291_9286# a_66870_9286# a_66243_8611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2814 a_43738_6586# a_43738_6330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2815 a_67082_13700# a_66869_13700# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2816 a_3975_11577# a_4833_8604# a_5041_8604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2817 a_1014_5572# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2818 a_6717_9249# a_8209_10003# a_8160_10193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2819 a_39049_4855# a_39141_3220# a_39092_3410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2820 a_74014_5522# a_74010_5699# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2821 a_79024_13014# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2822 a_65414_10421# a_66035_10737# a_66243_10737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2823 vdd a_30090_8554# a_29882_8554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2824 a_15749_8598# a_15886_4727# a_11048_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2825 a_77997_3272# a_77576_3272# a_76949_2597# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2826 a_32988_4802# a_33609_4723# a_33817_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2827 a_76742_13698# a_76529_13698# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2828 a_66869_12253# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2829 a_44362_10739# a_44149_10739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2830 a_19919_11526# a_19915_11703# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2831 a_48738_7659# a_49851_10681# a_49806_10694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2832 a_67080_6245# a_66867_6245# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2833 a_37422_8596# a_37001_8596# a_36354_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2834 a_9206_2734# a_609_2614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2835 a_54855_2599# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2836 a_13192_3274# a_12771_3274# a_12144_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2837 a_52338_4181# a_52595_3991# a_51290_4185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2838 a_76121_12586# a_76742_13019# a_76950_13019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2839 vdd d0 a_20173_9225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2840 gnd d1 a_51547_2548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2841 vdd a_50101_12203# a_49893_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2842 a_47107_11577# a_46686_11577# a_47013_11696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2843 a_72964_11711# a_74061_11517# a_74012_11707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2844 a_60512_4680# a_60599_6189# a_60550_6379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2845 a_60508_4857# a_60765_4667# a_59442_7830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2846 a_13193_12249# a_14432_13016# a_14589_11690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2847 gnd a_28600_10679# a_28392_10679# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2848 a_40541_10185# a_40798_9995# a_39098_9241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2849 a_56323_7688# a_55902_7688# a_55275_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2850 a_27275_7834# a_28390_4671# a_28341_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2851 a_54447_5060# a_55067_5566# a_55275_5566# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2852 a_66243_10058# a_67083_10733# a_67291_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2853 a_25440_11575# a_25227_11575# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2854 a_33819_10731# a_34659_10727# a_34867_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2855 a_32987_6578# a_33608_7011# a_33816_7011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2856 a_76119_7119# a_76740_7011# a_76948_7011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 a_22280_2966# a_22280_2711# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2858 gnd a_73221_12968# a_73013_12968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2859 a_12770_7688# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2860 a_10726_446# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2861 a_74014_6969# a_74267_6956# a_72962_7150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2862 vdd a_63302_6184# a_63094_6184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2863 gnd a_20171_3985# a_19963_3985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2864 a_2275_7694# a_2062_7694# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2865 a_55067_7692# a_54854_7692# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2866 a_9209_6971# a_9205_7148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2867 gnd d0 a_20171_2538# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2868 a_48419_4733# a_48310_4733# a_48518_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2869 vdd a_31135_5509# a_30927_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2870 gnd d3 a_39308_10673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2871 a_74017_10010# a_74013_10187# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2872 a_51292_8746# a_52389_8552# a_52344_8565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2873 a_1016_13706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2874 a_43741_10423# a_43741_10168# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2875 a_76951_9284# a_76530_9284# a_76122_8968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2876 a_64708_433# a_64495_433# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2877 a_54448_12588# a_55069_13021# a_55277_13021# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2878 a_607_4810# a_607_4415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2879 a_8157_5705# a_9254_5511# a_9209_5524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2880 a_79389_11569# a_79025_10047# a_77999_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2881 a_8162_2561# a_8415_2548# a_6711_3418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2882 a_60551_3412# a_62047_2542# a_62002_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2883 a_80800_4725# a_80691_4725# a_75853_444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2884 a_33396_4723# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2885 a_39096_3233# a_40588_3987# a_40543_4000# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2886 a_44569_13706# a_44148_13706# a_43740_13785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2887 a_65413_11686# a_65414_11072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2888 a_33819_10052# a_33398_10052# a_32990_9619# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2889 a_47965_8604# a_47752_8604# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2890 gnd a_51548_12970# a_51340_12970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2891 a_33398_10731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2892 a_28387_6206# a_29879_6960# a_29830_7150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2893 a_39049_4855# a_39141_3220# a_39096_3233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2894 a_41591_3996# a_41587_4173# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2895 a_22902_13704# a_22689_13704# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2896 a_2483_7694# a_3722_7014# a_3879_5688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2897 a_54447_2707# a_54449_2608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2898 a_3552_5569# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2899 a_41588_13827# a_41845_13637# a_40544_12975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2900 vdd d0 a_41843_6950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2901 a_62001_5522# a_63094_6184# a_63045_6374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2902 a_83671_2730# a_84768_2536# a_84719_2726# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2903 a_22280_3361# a_22901_3282# a_23109_3282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2904 a_79236_4039# a_79023_4039# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2905 a_5287_4733# a_5651_7646# a_5602_7836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2906 a_47006_5569# a_46642_4047# a_45616_3280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2907 a_18865_5699# a_19122_5509# a_17418_6379# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2908 a_51295_11536# a_51548_11523# a_49844_12393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2909 gnd a_82483_9228# a_82275_9228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2910 gnd a_40798_8548# a_40590_8548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2911 a_83674_6967# a_83927_6954# a_82227_6200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2912 a_65411_7125# a_65411_6584# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2913 a_66240_6249# a_65819_6249# a_65411_6328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2914 gnd a_84976_3983# a_84768_3983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2915 gnd d0 a_84975_5503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2916 a_22903_10058# a_22690_10058# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2917 a_27275_7834# a_28390_4671# a_28345_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2918 a_52341_5524# a_52594_5511# a_51289_5705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2919 gnd a_20173_9225# a_19965_9225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2920 a_11314_7121# a_11314_6580# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2921 a_66867_6245# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2922 a_41590_5516# a_41843_5503# a_40538_5697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2923 a_14473_5563# a_14260_5563# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2924 a_43740_12594# a_43740_12338# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2925 a_9205_7827# a_9462_7637# a_8161_6975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2926 a_11315_3613# a_11315_3357# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2927 gnd a_20172_13639# a_19964_13639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_1436_4052# a_1015_4052# a_607_3619# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 a_45617_13702# a_46856_13022# a_47013_11696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2930 gnd d3 a_6927_10681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2931 a_1017_9292# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2932 a_33817_4723# a_34657_4719# a_34865_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2933 a_23110_13025# a_23950_13700# a_24158_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2934 vdd d3 a_39308_10673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2935 a_66033_3282# a_65820_3282# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2936 gnd d2 a_39350_12195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2937 a_56325_12249# a_55904_12249# a_55277_11574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2938 vdd a_83930_8548# a_83722_8548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2939 a_56323_6241# a_57562_7008# a_57719_5682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2940 a_65821_11578# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2941 a_82226_9418# a_83722_8548# a_83673_8738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2942 a_1435_7698# a_1014_7698# a_606_7777# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2943 a_45408_3280# a_45195_3280# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2944 a_63047_13829# a_63051_12973# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2945 a_1438_10060# a_1017_10060# a_609_9627# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2946 a_9205_5701# a_9210_4683# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2947 a_32989_13382# a_33610_13698# a_33818_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2948 a_17425_9243# a_17678_9230# a_17378_10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2949 a_49848_12216# a_51340_12970# a_51295_12983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2950 a_19917_6965# a_19913_7142# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2951 a_84723_4675# a_84976_4662# a_83675_4000# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2952 a_19916_10183# a_19920_9238# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2953 a_1438_8613# a_2278_9288# a_2486_9288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2954 a_54449_9365# a_55070_9286# a_55278_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2955 a_76528_3276# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2956 a_33609_4044# a_33396_4044# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2957 a_11937_13700# a_11724_13700# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2958 gnd a_31137_11517# a_30929_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2959 a_77788_7686# a_77575_7686# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2960 gnd a_52595_4670# a_52387_4670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2961 a_22282_8719# a_22903_8611# a_23111_8611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2962 a_68686_11694# a_68316_13020# a_67290_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2963 a_76742_11572# a_76529_11572# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2964 a_609_11074# a_609_10818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2965 a_28388_3239# a_29880_3993# a_29835_4006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2966 a_43741_9371# a_43741_8976# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2967 a_74013_8740# a_74014_7648# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2968 a_46854_7014# a_46641_7014# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2969 a_83671_2730# a_84768_2536# a_84723_2549# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2970 a_66241_4050# a_67081_4725# a_67289_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2971 gnd d0 a_31137_13643# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2972 gnd d0 a_63302_7631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2973 a_62001_5522# a_63094_6184# a_63049_6197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2974 a_54856_13021# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2975 a_5287_4733# a_5651_7646# a_5606_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2976 a_54854_7013# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2977 a_55275_6245# a_54854_6245# a_54446_6324# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2978 a_51291_11713# a_51548_11523# a_49844_12393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2979 a_26714_8602# a_26293_8602# a_25646_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2980 a_29835_2559# a_30088_2546# a_28384_3416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2981 vdd d0 a_74268_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2982 a_16310_7830# a_17425_4667# a_17380_4680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2983 a_54448_12332# a_54448_11937# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2984 gnd d0 a_41845_11511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2985 vdd a_20173_9225# a_19965_9225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2986 a_44362_9292# a_44149_9292# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2987 a_32987_7374# a_32987_7119# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2988 a_52337_5701# a_52594_5511# a_51289_5705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2989 gnd a_51547_2548# a_51339_2548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2990 gnd d2 a_50100_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2991 a_66035_8611# a_65822_8611# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2992 a_34864_7686# a_34443_7686# a_33816_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2993 a_30878_6378# a_31135_6188# a_29834_5526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2994 vdd a_19124_12964# a_18916_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2995 a_1016_11580# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2996 vdd d3 a_6927_10681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2997 gnd a_28640_6193# a_28432_6193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2998 a_14589_11690# a_14219_13016# a_13193_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2999 gnd d2 a_6969_12203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3000 gnd d0 a_74269_12196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 a_60510_10865# a_60602_9230# a_60553_9420# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3002 a_67291_10733# a_66870_10733# a_66243_10058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3003 vdd a_52594_6190# a_52386_6190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3004 gnd d1 a_8415_3995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3005 a_35935_11569# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3006 a_63052_10685# a_63048_10862# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3007 a_71479_10692# a_71732_10679# a_70411_7657# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3008 gnd a_20170_5505# a_19962_5505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3009 a_63052_9238# a_63048_9415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3010 a_2062_7694# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3011 a_608_13390# a_1229_13706# a_1437_13706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3012 a_33611_9284# a_33398_9284# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3013 a_2065_10735# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3014 a_44569_11580# a_44148_11580# a_43741_11074# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3015 a_55903_4721# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3016 a_30879_4858# a_31136_4668# a_29835_4006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3017 a_17421_9420# a_17678_9230# a_17378_10865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3018 gnd d0 a_9463_3223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3019 a_84719_4852# a_84976_4662# a_83675_4000# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3020 a_57714_5563# a_57350_4041# a_56324_4721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3021 a_17423_3235# a_18915_3989# a_18870_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3022 a_23110_13704# a_22689_13704# a_22281_13783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3023 a_55278_10054# a_54857_10054# a_54449_9621# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3024 a_49846_6208# a_51338_6962# a_51289_7152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3025 vdd a_73219_6960# a_73011_6960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3026 a_65411_6584# a_65411_6328# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3027 vdd a_52595_4670# a_52387_4670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3028 a_34445_12247# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3029 a_39091_6377# a_40587_5507# a_40542_5520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3030 a_12145_13700# a_12985_13696# a_13193_13696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3031 a_65413_13783# a_66034_13704# a_66242_13704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3032 a_5606_7659# a_6719_10681# a_6670_10871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3033 gnd a_30090_10001# a_29882_10001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3034 a_11314_6580# a_11314_6324# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3035 a_47752_8604# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3036 a_23108_7696# a_22687_7696# a_22279_7380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3037 a_67081_3278# a_66868_3278# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3038 a_44361_13706# a_44148_13706# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3039 vdd d0 a_31137_13643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3040 vdd d0 a_63302_7631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3041 a_39098_9241# a_39351_9228# a_39051_10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3042 a_43738_7777# a_44359_7698# a_44567_7698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3043 a_11935_6245# a_11722_6245# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3044 a_63047_13829# a_63304_13639# a_62003_12977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3045 vdd d0 a_41845_11511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3046 a_23111_9290# a_23951_9286# a_24159_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3047 a_40542_5520# a_41635_6182# a_41586_6372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3048 gnd d0 a_52594_6190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3049 a_84719_3405# a_84723_2549# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3050 a_29831_2736# a_30088_2546# a_28384_3416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3051 a_76122_8713# a_76119_8025# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3052 a_54447_2707# a_55068_2599# a_55276_2599# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3053 a_65414_9625# a_66035_10058# a_66243_10058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3054 vdd a_41843_6950# a_41635_6950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3055 a_76121_13382# a_76121_13127# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3056 vdd d1 a_40797_12962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3057 vdd a_71774_12201# a_71566_12201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3058 a_32988_4152# a_33609_4044# a_33817_4044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3059 a_68570_5567# a_68357_5567# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3060 a_66242_13704# a_67082_13700# a_67290_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3061 a_44362_10060# a_44149_10060# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3062 a_34658_13694# a_34445_13694# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3063 a_76742_13019# a_76529_13019# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3064 a_25552_5686# a_25182_7012# a_24156_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3065 a_56326_10729# a_55905_10729# a_55278_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3066 gnd a_84975_5503# a_84767_5503# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3067 a_8163_12983# a_9256_13645# a_9207_13835# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3068 a_45409_13702# a_45196_13702# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3069 a_43741_8976# a_43741_8721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3070 a_24156_6245# a_23735_6245# a_23108_6249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3071 a_30883_4002# a_30879_4179# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3072 a_2276_4727# a_2063_4727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3073 a_14260_5563# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3074 a_60510_10865# a_60602_9230# a_60557_9243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3075 a_51294_4008# a_52387_4670# a_52338_4860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3076 a_77996_6239# a_77575_6239# a_76948_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3077 a_32987_7374# a_33608_7690# a_33816_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3078 a_1435_5572# a_1014_5572# a_607_5066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3079 vdd a_20173_9993# a_19965_9993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3080 a_29836_12981# a_30929_13643# a_30880_13833# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3081 a_54448_11937# a_54448_11682# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3082 a_32989_11680# a_33610_11572# a_33818_11572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3083 a_52344_10691# a_52597_10678# a_51296_10016# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3084 a_9209_7650# a_9205_7827# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3085 a_12143_7013# a_12983_7688# a_13191_7688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3086 a_40540_11705# a_41637_11511# a_41588_11701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3087 a_65820_3282# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3088 a_22901_4050# a_22688_4050# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3089 a_77790_12247# a_77577_12247# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3090 a_11937_11574# a_11724_11574# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3091 gnd d1 a_73222_10001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3092 vdd d0 a_9463_3223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3093 a_54448_13384# a_55069_13700# a_55277_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3094 a_45195_3280# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3095 a_1016_13027# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3096 vdd d1 a_30090_10001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3097 a_77578_9280# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3098 a_22900_7696# a_22687_7696# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3099 a_76120_3355# a_76120_2960# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3100 a_76740_6243# a_76527_6243# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3101 a_6674_10694# a_6761_12203# a_6712_12393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3102 a_5606_7659# a_6719_10681# a_6674_10694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3103 a_12146_9286# a_11725_9286# a_11317_9365# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3104 a_12984_3274# a_12771_3274# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3105 a_33608_5564# a_33395_5564# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3106 a_84724_12203# a_84720_12380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3107 a_33396_4044# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3108 a_18871_12977# a_19964_13639# a_19919_13652# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3109 a_77575_7686# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3110 a_56115_6241# a_55902_6241# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3111 a_41591_4675# a_41587_4852# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3112 a_44569_13027# a_44148_13027# a_43740_13135# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3113 a_51293_5528# a_52386_6190# a_52341_6203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3114 gnd d0 a_52596_13645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3115 gnd a_62256_11517# a_62048_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3116 a_33398_10052# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3117 a_40542_5520# a_41635_6182# a_41590_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3118 a_11317_10162# a_11317_9621# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3119 a_2277_13702# a_2064_13702# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3120 vdd d0 a_31138_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3121 gnd a_63302_7631# a_63094_7631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3122 a_22902_13025# a_22689_13025# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3123 a_44149_10060# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3124 a_33817_2597# a_34657_3272# a_34865_3272# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3125 vdd a_74268_3989# a_74060_3989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3126 vdd d0 a_74267_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3127 a_8163_12983# a_9256_13645# a_9211_13658# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3128 a_76948_7011# a_77788_7686# a_77996_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3129 gnd a_50099_6195# a_49891_6195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3130 a_43739_5066# a_43739_4810# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3131 a_12772_13696# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3132 gnd d1 a_19125_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3133 a_65822_8611# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3134 vdd a_17675_6189# a_17467_6189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3135 a_51294_4008# a_52387_4670# a_52342_4683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3136 a_63045_5695# a_63302_5505# a_61997_5699# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3137 a_608_11688# a_1229_11580# a_1437_11580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3138 a_65411_7125# a_66032_7017# a_66240_7017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3139 a_19918_3230# a_20171_3217# a_18870_2555# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3140 a_75853_444# a_80478_4725# a_80554_8596# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3141 a_44568_4731# a_44147_4731# a_43739_4810# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3142 a_47105_5569# a_46684_5569# a_47011_5688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3143 a_29836_12981# a_30929_13643# a_30884_13656# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3144 a_67291_10733# a_68530_10053# a_68681_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3145 a_54446_8027# a_54446_7771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3146 a_22279_5933# a_22900_6249# a_23108_6249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3147 a_22280_3617# a_22280_3361# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3148 a_29832_13158# a_30089_12968# a_28389_12214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3149 a_23950_12253# a_23737_12253# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3150 a_40540_11705# a_41637_11511# a_41592_11524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3151 gnd d2 a_50101_12203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3152 gnd a_8415_3995# a_8207_3995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3153 a_63046_4854# a_63050_3998# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3154 a_66869_13700# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3155 a_67080_7692# a_66867_7692# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3156 a_75531_444# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3157 a_63046_4175# a_63303_3985# a_61998_4179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3158 a_72967_4006# a_74060_4668# a_74011_4858# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3159 a_608_13135# a_608_12594# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3160 a_1438_10739# a_1017_10739# a_609_10423# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3161 gnd d2 a_71775_9234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3162 a_13192_4721# a_12771_4721# a_12144_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3163 a_45618_9288# a_45197_9288# a_44570_8613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3164 a_19917_7644# a_19913_7821# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3165 a_1435_7019# a_1014_7019# a_606_7127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3166 gnd a_9463_3223# a_9255_3223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3167 a_25185_10053# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3168 a_65414_9369# a_65414_8974# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3169 a_17376_4857# a_17468_3222# a_17419_3412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3170 a_46855_4047# a_46642_4047# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3171 a_17418_6379# a_18914_5509# a_18869_5522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3172 gnd d1 a_30089_12968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3173 a_32989_12586# a_33610_13019# a_33818_13019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3174 a_30882_6969# a_30878_7146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3175 a_66032_6249# a_65819_6249# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3176 a_55276_3278# a_54855_3278# a_54447_2962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3177 a_84723_3996# a_84976_3983# a_83671_4177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3178 a_23109_2603# a_22688_2603# a_22282_2612# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3179 vdd d0 a_52596_13645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3180 a_22281_11941# a_22281_11686# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3181 gnd a_52595_3991# a_52387_3991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3182 a_15749_8598# a_15328_8598# a_14681_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3183 a_45407_6247# a_45194_6247# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3184 vdd a_63302_7631# a_63094_7631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3185 a_43739_2713# a_44360_2605# a_44568_2605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3186 a_84725_10683# a_84978_10670# a_83677_10008# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3187 a_11722_6245# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3188 a_54856_13700# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3189 a_80800_4725# a_81164_7638# a_81119_7651# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3190 a_12144_2599# a_11723_2599# a_11315_2707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3191 a_24157_3278# a_25396_4045# a_25547_5567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3192 a_34865_4719# a_34444_4719# a_33817_4044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3193 gnd d0 a_31137_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3194 a_57349_7008# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3195 gnd d0 a_63302_6952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3196 gnd a_84977_12190# a_84769_12190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3197 a_1227_6251# a_1014_6251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3198 a_32987_5672# a_33608_5564# a_33816_5564# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3199 a_63051_12973# a_63304_12960# a_61999_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3200 a_36354_5561# a_35933_5561# a_36255_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3201 a_3725_10055# a_3512_10055# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3202 gnd a_9464_12198# a_9256_12198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3203 a_44569_12259# a_45409_12255# a_45617_12255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3204 a_62003_11530# a_63096_12192# a_63047_12382# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3205 a_12985_12249# a_12772_12249# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3206 vdd a_41845_12190# a_41637_12190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3207 a_8160_10193# a_9257_9999# a_9212_10012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3208 a_52340_10868# a_52344_10012# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3209 a_2063_4727# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3210 a_12145_11574# a_11724_11574# a_11316_11682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3211 a_60512_4680# a_60765_4667# a_59442_7830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3212 a_54448_11682# a_55069_11574# a_55277_11574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3213 a_609_10423# a_609_10168# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3214 a_66241_4050# a_65820_4050# a_65412_3617# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3215 a_66870_9286# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3216 a_58881_8598# a_59018_4727# a_54180_446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3217 a_22900_5570# a_22687_5570# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3218 a_62001_6969# a_63094_7631# a_63045_7821# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3219 a_14475_11571# a_14262_11571# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3220 vdd d2 a_71775_9234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3221 a_55278_8607# a_54857_8607# a_54446_8027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3222 a_608_12594# a_1229_13027# a_1437_13027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3223 vdd a_9463_3223# a_9255_3223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3224 a_52339_11709# a_52344_10691# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3225 a_17425_9243# a_18917_9997# a_18868_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3226 a_66240_7696# a_65819_7696# a_65411_7775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3227 a_9205_6380# a_9209_5524# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3228 a_56324_3274# a_55903_3274# a_55276_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3229 a_17376_4857# a_17468_3222# a_17423_3235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3230 a_76530_10731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3231 a_5386_4733# a_4965_4733# a_5287_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3232 a_37001_8596# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3233 a_12771_3274# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3234 a_33395_5564# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3235 a_23110_13025# a_22689_13025# a_22281_13133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3236 a_11724_12253# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3237 a_37987_7651# a_39100_10673# a_39051_10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3238 a_66035_10737# a_65822_10737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3239 gnd a_30088_3993# a_29880_3993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3240 vdd a_51549_10003# a_51341_10003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3241 a_29834_5526# a_30927_6188# a_30882_6201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3242 a_65413_13133# a_66034_13025# a_66242_13025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3243 a_55902_7688# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3244 a_48310_4733# a_48097_4733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3245 a_84721_10860# a_84978_10670# a_83677_10008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3246 gnd d1 a_40796_3987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3247 a_9206_4181# a_9210_3236# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3248 a_76119_5927# a_76740_6243# a_76948_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3249 a_18867_13154# a_19964_12960# a_19915_13150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3250 a_66242_12257# a_65821_12257# a_65413_11941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3251 vdd d0 a_52597_9999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3252 a_44361_13027# a_44148_13027# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3253 a_1437_11580# a_2277_12255# a_2485_12255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3254 a_19914_2728# a_11317_2608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3255 a_24157_3278# a_23736_3278# a_23109_2603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3256 a_26638_4731# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3257 vdd a_74267_5509# a_74059_5509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3258 a_23951_10733# a_23738_10733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3259 a_11316_13384# a_11316_13129# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3260 a_65414_8974# a_65414_8719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3261 vdd d1 a_62257_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3262 a_36354_5561# a_37214_8596# a_37422_8596# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3263 a_37559_4725# a_37346_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3264 gnd d0 a_41844_3215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3265 a_41592_13650# a_41845_13637# a_40544_12975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3266 a_608_12594# a_608_12338# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3267 a_77999_9280# a_79238_10047# a_79389_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3268 gnd a_5859_7646# a_5651_7646# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3269 a_29835_4006# a_30928_4668# a_30883_4681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3270 a_76528_4723# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3271 a_23111_8611# a_22690_8611# a_22282_8719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3272 a_44567_6251# a_45407_6247# a_45615_6247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3273 a_57565_10049# a_57352_10049# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3274 a_8159_13160# a_9256_12966# a_9207_13156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3275 a_22281_13783# a_22281_13388# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3276 gnd a_8417_10003# a_8209_10003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3277 a_43741_10168# a_44362_10060# a_44570_10060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3278 a_51290_4185# a_52387_3991# a_52338_4181# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3279 a_9209_7650# a_9462_7637# a_8161_6975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3280 a_62001_6969# a_63094_7631# a_63049_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3281 a_29832_13158# a_30929_12964# a_30880_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3282 a_44146_7698# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3283 a_52344_10012# a_52597_9999# a_51292_10193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3284 a_55275_7692# a_54854_7692# a_54446_7771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3285 gnd a_70664_7644# a_70456_7644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3286 a_22901_4729# a_22688_4729# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3287 vdd a_39351_9228# a_39143_9228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3288 a_33609_2597# a_33396_2597# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3289 vdd d0 a_84975_6950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3290 a_65412_3361# a_66033_3282# a_66241_3282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3291 a_72966_6973# a_73219_6960# a_71519_6206# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3292 gnd a_83930_8548# a_83722_8548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3293 a_41586_7140# a_41843_6950# a_40538_7144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3294 a_37987_7651# a_39100_10673# a_39055_10686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3295 a_63051_12205# a_63047_12382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3296 a_11147_446# a_21576_433# a_21784_433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3297 a_54856_11574# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3298 a_22900_7017# a_22687_7017# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3299 a_46641_7014# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3300 gnd a_82481_3220# a_82273_3220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3301 a_84722_5516# a_84975_5503# a_83670_5697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3302 a_57605_5563# a_57392_5563# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3303 vdd d2 a_82480_6187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3304 gnd d0 a_74269_13643# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3305 a_44570_10060# a_45410_10735# a_45618_10735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3306 a_12146_10733# a_12986_10729# a_13194_10729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3307 a_33816_6243# a_33395_6243# a_32987_5927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3308 a_12143_7013# a_11722_7013# a_11314_6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3309 a_57562_7008# a_57349_7008# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3310 a_45194_6247# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3311 a_11317_10812# a_11317_10417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3312 a_41593_9236# a_41589_9413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3313 a_39094_9418# a_40590_8548# a_40545_8561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3314 a_76949_4723# a_77789_4719# a_77997_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3315 a_54279_446# a_53858_446# a_48518_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3316 a_44149_10739# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3317 a_9209_5524# a_9205_5701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3318 gnd d0 a_52596_12966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3319 a_65412_5064# a_65412_4808# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3320 a_71518_9424# a_73014_8554# a_72965_8744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3321 gnd a_63302_6952# a_63094_6952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3322 a_11315_5060# a_11315_4804# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3323 vdd d0 a_41844_3215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3324 vdd a_5859_7646# a_5651_7646# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3325 a_16310_7830# a_17425_4667# a_17376_4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3326 gnd d1 a_62256_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3327 a_84718_7140# a_84722_6195# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3328 a_34445_13694# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3329 a_43741_9627# a_43741_9371# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3330 a_1436_3284# a_2276_3280# a_2484_3280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3331 gnd d3 a_82438_4665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3332 a_33398_9284# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3333 gnd d0 a_74270_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3334 gnd a_52596_12198# a_52388_12198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3335 a_11938_9286# a_11725_9286# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3336 a_32987_6322# a_32987_5927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3337 a_67081_4725# a_66868_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3338 a_76950_11572# a_76529_11572# a_76121_11680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3339 a_44568_4052# a_44147_4052# a_43739_4160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3340 a_11725_10733# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3341 vdd a_70664_7644# a_70456_7644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3342 a_41591_2549# a_41587_2726# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3343 a_66240_5570# a_65819_5570# a_65412_5064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3344 gnd a_60810_9230# a_60602_9230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3345 a_37422_8596# a_37559_4725# a_32721_444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3346 gnd a_40797_12962# a_40589_12962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3347 gnd d0 a_63304_12192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3348 gnd a_50059_10681# a_49851_10681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3349 a_63048_9415# a_63052_8559# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3350 a_69846_8602# a_69425_8602# a_68778_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3351 a_66243_10737# a_65822_10737# a_65414_10816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3352 a_34866_13694# a_34445_13694# a_33818_13019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3353 a_54854_6245# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3354 a_34865_3272# a_34444_3272# a_33817_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3355 a_72963_4183# a_73220_3993# a_71520_3239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3356 a_72963_4183# a_74060_3989# a_74011_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3357 a_30882_7648# a_30878_7825# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3358 a_1438_8613# a_1017_8613# a_609_8721# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3359 a_83677_10008# a_83930_9995# a_82230_9241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3360 a_24156_7692# a_23735_7692# a_23108_7696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3361 vdd a_82481_3220# a_82273_3220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3362 a_43739_4415# a_43739_4160# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3363 a_30883_4681# a_31136_4668# a_29835_4006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3364 vdd d0 a_74269_13643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3365 a_77996_7686# a_77575_7686# a_76948_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3366 a_41588_13827# a_41592_12971# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3367 a_68780_11575# a_69638_8602# a_69846_8602# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3368 a_74010_6378# a_74267_6188# a_72966_5526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3369 a_79488_11569# a_79067_11569# a_79394_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3370 vdd a_20170_6952# a_19962_6952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3371 vdd a_20171_3217# a_19963_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3372 a_26851_4731# a_26638_4731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3373 a_46897_5569# a_46684_5569# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3374 a_9207_11709# a_9464_11519# a_8159_11713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3375 gnd d1 a_40795_5507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3376 vdd d1 a_83929_12962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3377 a_4833_8604# a_4620_8604# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3378 gnd a_40796_3987# a_40588_3987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3379 gnd d1 a_19122_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3380 a_77790_13694# a_77577_13694# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3381 a_3724_13022# a_3511_13022# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3382 a_8159_13160# a_8416_12970# a_6716_12216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3383 vdd a_74269_12964# a_74061_12964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3384 a_71518_9424# a_73014_8554# a_72969_8567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3385 gnd d0 a_20170_6184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3386 a_74015_3234# a_74011_3411# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3387 a_76743_9284# a_76530_9284# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3388 a_84725_10004# a_84978_9991# a_83673_10185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3389 a_63051_13652# a_63304_13639# a_62003_12977# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3390 a_51291_13160# a_52388_12966# a_52343_12979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3391 a_44570_9292# a_44149_9292# a_43741_9371# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3392 a_74011_4858# a_74268_4668# a_72967_4006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3393 a_41589_10181# a_41846_9991# a_40541_10185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3394 a_56118_9282# a_55905_9282# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3395 gnd a_41844_3215# a_41636_3215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3396 vdd d3 a_82438_4665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3397 vdd d0 a_74270_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3398 a_12984_4721# a_12771_4721# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3399 a_19917_5518# a_19913_5695# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3400 a_12773_10729# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3401 vdd d0 a_84977_12958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3402 vdd d2 a_28642_12201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3403 a_57815_11571# a_57394_11571# a_57721_11690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3404 a_52337_7827# a_52341_6971# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3405 a_14219_13016# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3406 a_27279_7657# a_27532_7644# a_26960_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3407 a_18866_2732# a_19963_2538# a_19918_2551# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3408 vdd d0 a_9464_12966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3409 a_74016_12209# a_74269_12196# a_72968_11534# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3410 a_82228_3233# a_83720_3987# a_83671_4177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3411 vdd a_60810_9230# a_60602_9230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3412 a_40542_6967# a_41635_7629# a_41590_7642# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3413 vdd d0 a_52594_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3414 a_66241_4729# a_65820_4729# a_65412_4413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3415 a_22687_7696# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3416 a_22282_11072# a_22902_11578# a_23110_11578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3417 a_44147_2605# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3418 a_30880_12386# a_31137_12196# a_29836_11534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3419 vdd a_50059_10681# a_49851_10681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3420 a_33396_2597# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3421 a_66243_9290# a_67083_9286# a_67291_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3422 a_83674_5520# a_84767_6182# a_84718_6372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3423 a_61997_7146# a_63094_6952# a_63045_7142# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3424 vdd a_84975_6950# a_84767_6950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3425 a_11936_2599# a_11723_2599# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3426 a_22280_4158# a_22901_4050# a_23109_4050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3427 gnd d0 a_20172_11513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3428 a_41593_10683# a_41589_10860# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3429 a_39096_3233# a_39349_3220# a_39049_4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3430 a_36104_4039# a_35891_4039# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3431 a_76120_3355# a_76741_3276# a_76949_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3432 a_32988_4152# a_32988_3611# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3433 a_32987_5927# a_32987_5672# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3434 a_66240_7017# a_65819_7017# a_65411_7125# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3435 a_68684_5686# a_68314_7012# a_67288_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3436 a_32988_2960# a_33609_3276# a_33817_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3437 a_13192_4721# a_14431_4041# a_14582_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3438 a_83676_11528# a_83929_11515# a_82225_12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3439 a_76530_10052# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3440 a_55275_7692# a_56115_7688# a_56323_7688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3441 a_67288_6245# a_66867_6245# a_66240_6249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3442 vdd d1 a_30088_3993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3443 a_22279_7380# a_22900_7696# a_23108_7696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3444 a_57392_5563# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3445 vdd d0 a_74270_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3446 a_23950_13700# a_23737_13700# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3447 a_66035_10058# a_65822_10058# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3448 a_18871_12977# a_19964_13639# a_19915_13829# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3449 a_36262_11688# a_35892_13014# a_34866_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3450 vdd d0 a_20170_6184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3451 a_41587_4852# a_41591_3996# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3452 a_28345_4684# a_28598_4671# a_27275_7834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3453 a_9208_8742# a_9209_7650# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3454 vdd d2 a_28640_6193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3455 a_77998_13694# a_79237_13014# a_79394_11688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3456 a_2483_7694# a_2062_7694# a_1435_7019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3457 a_76119_7119# a_76119_6578# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3458 a_43118_401# a_43009_401# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3459 a_66033_4050# a_65820_4050# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3460 a_24158_12253# a_23737_12253# a_23110_11578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3461 a_3722_7014# a_3509_7014# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3462 vdd a_41844_3215# a_41636_3215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3463 a_57564_13016# a_57351_13016# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3464 a_27059_4731# a_32612_444# a_21685_433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3465 a_25646_5567# a_25225_5567# a_25547_5567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3466 a_18868_10187# a_19125_9997# a_17425_9243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3467 a_32990_10160# a_32990_9619# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3468 a_33818_12251# a_33397_12251# a_32989_11935# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3469 a_43738_7382# a_43738_7127# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3470 a_41592_12971# a_41845_12958# a_40540_13152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3471 a_27275_7834# a_27532_7644# a_26960_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3472 a_66032_7696# a_65819_7696# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3473 gnd a_82438_4665# a_82230_4665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3474 a_55276_4725# a_54855_4725# a_54447_4409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3475 a_1230_9292# a_1017_9292# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3476 a_76528_4044# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3477 a_11725_9286# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3478 a_76741_2597# a_76528_2597# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3479 a_82229_12208# a_83721_12962# a_83676_12975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3480 a_45407_7694# a_45194_7694# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3481 a_44567_5572# a_44146_5572# a_43738_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3482 a_43741_10818# a_44362_10739# a_44570_10739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3483 a_14218_4041# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3484 a_32987_8025# a_33611_8605# a_33819_8605# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3485 a_76122_8713# a_76743_8605# a_76951_8605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3486 a_6712_12393# a_6969_12203# a_6674_10694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3487 a_80554_8596# a_80133_8596# a_79486_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3488 a_11314_7771# a_11935_7692# a_12143_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3489 a_76120_4802# a_76120_4407# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3490 a_83674_5520# a_84767_6182# a_84722_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3491 a_9209_6971# a_9462_6958# a_8157_7152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3492 vdd d0 a_20172_11513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3493 a_55275_7013# a_54854_7013# a_54446_7121# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3494 a_76949_2597# a_77789_3272# a_77997_3272# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3495 a_39092_3410# a_39349_3220# a_39049_4855# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3496 a_62002_4002# a_62255_3989# a_60555_3235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3497 a_22902_12257# a_22689_12257# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3498 a_52339_12388# a_52343_11532# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3499 a_70407_7834# a_71522_4671# a_71473_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3500 gnd a_9464_13645# a_9256_13645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3501 a_12985_13696# a_12772_13696# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3502 a_44569_13706# a_45409_13702# a_45617_13702# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3503 a_83672_13152# a_84769_12958# a_84724_12971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3504 a_28347_10692# a_28434_12201# a_28389_12214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3505 a_83672_11705# a_83929_11515# a_82225_12385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3506 a_82187_10686# a_82274_12195# a_82225_12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3507 a_23948_6245# a_23735_6245# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3508 a_19913_7821# a_19917_6965# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3509 a_5606_7659# a_5859_7646# a_5287_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3510 vdd d1 a_8414_6962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3511 a_71517_12391# a_73013_11521# a_72964_11711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3512 gnd d1 a_30087_5513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3513 a_22689_11578# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3514 a_22903_8611# a_22690_8611# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3515 a_65411_5933# a_66032_6249# a_66240_6249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3516 a_53858_446# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3517 a_28341_4861# a_28598_4671# a_27275_7834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3518 a_46684_5569# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3519 gnd d0 a_74269_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3520 a_79280_11569# a_79067_11569# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3521 gnd a_40795_5507# a_40587_5507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3522 a_4620_8604# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3523 a_48419_4733# a_48783_7646# a_48734_7836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3524 a_22281_11686# a_22282_11072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3525 a_55070_8607# a_54857_8607# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3526 gnd a_19122_6956# a_18914_6956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3527 a_34865_4719# a_36104_4039# a_36255_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3528 a_29837_8567# a_30930_9229# a_30885_9242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3529 a_76530_9284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3530 a_19914_3407# a_19918_2551# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3531 gnd d1 a_51549_10003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3532 a_65414_9625# a_65414_9369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3533 a_11317_8715# a_11314_8027# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3534 a_606_7777# a_1227_7698# a_1435_7698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3535 a_63048_10183# a_63305_9993# a_62000_10187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3536 a_80800_4725# a_81164_7638# a_81115_7828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3537 a_56324_4721# a_55903_4721# a_55276_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3538 vdd a_82438_4665# a_82230_4665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3539 a_12771_4721# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3540 a_71522_9247# a_71775_9234# a_71475_10869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3541 a_11724_13700# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3542 a_18871_12977# a_19124_12964# a_17424_12210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3543 a_82185_4678# a_82272_6187# a_82227_6200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3544 a_28343_10869# a_28600_10679# a_27279_7657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3545 a_54855_3278# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3546 a_1015_3284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3547 a_1437_13027# a_2277_13702# a_2485_13702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3548 a_66242_13704# a_65821_13704# a_65413_13388# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3549 gnd d1 a_73219_6960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3550 vdd d2 a_6967_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3551 a_22688_2603# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3552 a_11725_10054# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3553 a_11935_7013# a_11722_7013# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3554 a_24157_4725# a_23736_4725# a_23109_4050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3555 vdd a_84977_13637# a_84769_13637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3556 a_19920_10685# a_20173_10672# a_18872_10010# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3557 a_1435_5572# a_2275_6247# a_2483_6247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3558 a_77997_4719# a_77576_4719# a_76949_4044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3559 a_23110_11578# a_22689_11578# a_22282_11072# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3560 a_40538_7144# a_41635_6950# a_41586_7140# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3561 a_76119_6578# a_76119_6322# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3562 a_67289_3278# a_68528_4045# a_68679_5567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3563 a_70407_7834# a_71522_4671# a_71477_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3564 vdd a_9464_13645# a_9256_13645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3565 a_76529_13698# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3566 a_44570_8613# a_45410_9288# a_45618_9288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3567 a_11723_2599# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3568 a_65412_4413# a_65412_4158# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3569 a_22279_5678# a_22900_5570# a_23108_5570# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3570 a_62003_12977# a_63096_13639# a_63051_13652# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3571 a_43740_13390# a_43740_13135# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3572 a_74016_12977# a_74012_13154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3573 a_24159_10733# a_23738_10733# a_23111_10737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3574 a_66243_10058# a_65822_10058# a_65414_10166# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3575 a_11315_4409# a_11315_4154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3576 a_79486_5561# a_79065_5561# a_79387_5561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3577 a_71517_12391# a_73013_11521# a_72968_11534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3578 a_5602_7836# a_5859_7646# a_5287_4733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3579 a_1228_2605# a_1015_2605# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3580 vdd d1 a_30087_5513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3581 a_30883_4002# a_31136_3989# a_29831_4183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3582 a_49804_4686# a_50057_4673# a_48734_7836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3583 a_33819_10731# a_33398_10731# a_32990_10810# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3584 a_607_3363# a_607_2968# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3585 a_48419_4733# a_48783_7646# a_48738_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3586 a_6715_3241# a_8207_3995# a_8162_4008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3587 a_18868_10187# a_19965_9993# a_19920_10006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3588 gnd d2 a_17675_6189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3589 a_21576_433# a_21363_433# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3590 a_37346_4725# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3591 a_52343_11532# a_52339_11709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3592 a_66032_5570# a_65819_5570# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3593 a_36106_10047# a_35893_10047# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3594 gnd d1 a_19125_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3595 a_65820_4050# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3596 a_39053_4678# a_39306_4665# a_37983_7828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3597 a_44359_6251# a_44146_6251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3598 a_76121_13777# a_76121_13382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3599 gnd d1 a_51548_11523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3600 vdd d0 a_9463_3991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3601 a_55277_12253# a_54856_12253# a_54448_11937# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3602 a_13194_9282# a_12773_9282# a_12146_8607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3603 a_71518_9424# a_71775_9234# a_71475_10869# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3604 a_54857_8607# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3605 a_44360_3284# a_44147_3284# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3606 a_11316_12332# a_11316_11937# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3607 a_33819_9284# a_33398_9284# a_32990_9363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3608 a_76740_7011# a_76527_7011# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3609 a_55903_3274# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3610 a_76527_5564# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3611 a_4965_4733# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3612 a_29835_4006# a_30928_4668# a_30879_4858# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3613 a_45194_7694# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3614 a_65414_11072# a_65414_10816# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3615 a_19918_2551# a_19914_2728# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3616 a_56324_3274# a_57563_4041# a_57714_5563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3617 a_1436_4731# a_1015_4731# a_607_4810# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3618 a_30881_10866# a_30885_10010# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3619 gnd d1 a_83928_3987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3620 a_65413_11941# a_66034_12257# a_66242_12257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3621 a_19916_10862# a_20173_10672# a_18872_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3622 a_36262_11688# a_36148_11569# a_36356_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3623 a_68681_11575# a_68572_11575# a_68780_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3624 a_62001_5522# a_62254_5509# a_60550_6379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3625 a_44361_12259# a_44148_12259# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3626 a_44359_7019# a_44146_7019# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3627 a_67289_3278# a_66868_3278# a_66241_2603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3628 a_22280_4808# a_22901_4729# a_23109_4729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3629 a_46899_11577# a_46686_11577# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3630 gnd a_39351_9228# a_39143_9228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3631 a_40542_6967# a_40795_6954# a_39095_6200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3632 vdd a_9465_9999# a_9257_9999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3633 a_52340_10189# a_52344_9244# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3634 gnd d0 a_84976_3215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3635 a_34867_10727# a_34446_10727# a_33819_10052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3636 a_23735_6245# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3637 a_41591_3228# a_41844_3215# a_40543_2553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3638 gnd a_52596_13645# a_52388_13645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3639 vdd a_20172_12192# a_19964_12192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3640 a_30880_11707# a_30885_10689# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3641 a_66243_8611# a_65822_8611# a_65414_8719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3642 a_49800_4863# a_50057_4673# a_48734_7836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3643 a_68778_5567# a_68357_5567# a_68684_5686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3644 a_66242_11578# a_67082_12253# a_67290_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3645 vdd a_8414_6962# a_8206_6962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3646 a_33818_12251# a_34658_12247# a_34866_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3647 vdd a_19124_11517# a_18916_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3648 gnd a_63304_11513# a_63096_11513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3649 a_34656_6239# a_34443_6239# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3650 a_3723_4047# a_3510_4047# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3651 a_22690_8611# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3652 a_22279_6584# a_22900_7017# a_23108_7017# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3653 a_45409_12255# a_45196_12255# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3654 a_54447_2962# a_54447_2707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3655 a_2276_3280# a_2063_3280# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3656 a_6710_6385# a_8206_5515# a_8157_5705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3657 a_74013_9419# a_74270_9229# a_72969_8567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3658 vdd d1 a_19125_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3659 a_14589_11690# a_14475_11571# a_14683_11571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3660 a_76122_11066# a_76742_11572# a_76950_11572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3661 a_13191_6241# a_14430_7008# a_14587_5682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3662 a_66033_4729# a_65820_4729# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3663 a_39049_4855# a_39306_4665# a_37983_7828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3664 vdd d1 a_51548_11523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3665 a_28343_10869# a_28435_9234# a_28386_9424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3666 a_41589_9413# a_41593_8557# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3667 a_39094_9418# a_40590_8548# a_40541_8738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3668 gnd d2 a_82482_12195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3669 a_55069_11574# a_54856_11574# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3670 a_65411_7380# a_65411_7125# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3671 a_607_2713# a_1228_2605# a_1436_2605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3672 a_32990_10810# a_32990_10415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3673 a_72969_10014# a_74062_10676# a_74013_10866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3674 a_54854_7692# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3675 a_45408_4727# a_45195_4727# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3676 a_18872_8563# a_19965_9225# a_19916_9415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3677 a_84718_7140# a_84975_6950# a_83670_7144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3678 gnd d0 a_9462_5511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3679 a_25397_13020# a_25184_13020# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3680 vdd a_52594_6958# a_52386_6958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3681 gnd d1 a_62255_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3682 a_66032_7017# a_65819_7017# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3683 a_3881_11696# a_3767_11577# a_3975_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3684 gnd a_83930_9995# a_83722_9995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3685 a_55276_4046# a_54855_4046# a_54447_3613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3686 a_33397_12251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3687 a_76948_6243# a_76527_6243# a_76119_5927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3688 gnd d2 a_39349_3220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3689 a_51290_4185# a_51547_3995# a_49847_3241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3690 a_60557_9243# a_62049_9997# a_62000_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3691 vdd a_6967_6195# a_6759_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3692 a_43738_6330# a_44359_6251# a_44567_6251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3693 a_39093_12385# a_39350_12195# a_39055_10686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3694 vdd a_40798_9995# a_40590_9995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3695 gnd d0 a_20170_7631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3696 a_33817_2597# a_33396_2597# a_32988_2705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3697 a_11722_7013# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3698 a_12143_6245# a_11722_6245# a_11314_6324# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3699 a_2486_10735# a_2065_10735# a_1438_10060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3700 a_9212_8565# a_9465_8552# a_8160_8746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3701 a_11316_11937# a_11316_11682# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3702 vdd d0 a_84976_3215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3703 a_22690_10737# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3704 a_77997_3272# a_79236_4039# a_79387_5561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3705 a_41587_3405# a_41844_3215# a_40543_2553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3706 vdd a_52596_13645# a_52388_13645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3707 a_56326_9282# a_57565_10049# a_57716_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3708 gnd a_9464_12966# a_9256_12966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3709 a_61999_13154# a_63096_12960# a_63047_13150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3710 a_54071_446# a_53858_446# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3711 vdd a_63304_11513# a_63096_11513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3712 a_30878_7825# a_30882_6969# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3713 vdd a_71772_6193# a_71564_6193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3714 a_30882_5522# a_31135_5509# a_29830_5703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3715 a_55278_10733# a_54857_10733# a_54449_10812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3716 a_74016_13656# a_74269_13643# a_72968_12981# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3717 a_33397_13019# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3718 a_6710_6385# a_8206_5515# a_8161_5528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3719 a_41592_12203# a_41588_12380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3720 a_33611_10731# a_33398_10731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3721 gnd a_20171_3217# a_19963_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3722 a_26714_8602# a_26851_4731# a_27059_4731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3723 vdd d0 a_63304_13639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3724 a_23738_10733# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3725 a_28343_10869# a_28435_9234# a_28390_9247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3726 a_9211_11532# a_9464_11519# a_8159_11713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3727 a_72969_10014# a_74062_10676# a_74017_10689# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3728 a_3973_5569# a_4833_8604# a_5041_8604# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3729 gnd a_19125_8550# a_18917_8550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3730 a_18872_8563# a_19965_9225# a_19920_9238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3731 vdd d0 a_31138_9229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3732 a_74011_3411# a_74015_2555# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3733 vdd a_9463_3991# a_9255_3991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3734 a_15995_4727# a_15886_4727# a_11048_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3735 vdd d0 a_9462_5511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3736 a_77997_3272# a_77576_3272# a_76949_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3737 vdd d1 a_62255_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3738 a_76120_4802# a_76741_4723# a_76949_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3739 a_84725_8557# a_84721_8734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3740 a_32988_4407# a_33609_4723# a_33817_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3741 a_66869_12253# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3742 vdd a_30087_6960# a_29879_6960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3743 gnd a_60809_12197# a_60601_12197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3744 a_67288_7692# a_66867_7692# a_66240_7696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3745 a_71473_4861# a_71565_3226# a_71516_3416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3746 a_74015_4681# a_74268_4668# a_72967_4006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3747 a_11724_13021# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3748 vdd d1 a_40795_6954# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3749 a_71521_12214# a_71774_12201# a_71479_10692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3750 vdd d2 a_39349_3220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3751 vdd d0 a_20170_7631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3752 gnd d2 a_71772_6193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3753 a_69983_4731# a_69770_4731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3754 a_33819_10052# a_34659_10727# a_34867_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3755 a_76119_6578# a_76740_7011# a_76948_7011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3756 a_52341_6203# a_52337_6380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3757 a_18866_2732# a_19963_2538# a_19914_2728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3758 gnd d0 a_31136_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3759 gnd a_83928_3987# a_83720_3987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3760 gnd d1 a_83927_5507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3761 a_51293_5528# a_51546_5515# a_49842_6385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3762 a_66242_13025# a_65821_13025# a_65413_12592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3763 a_25440_11575# a_25227_11575# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3764 a_9208_8742# a_9465_8552# a_8160_8746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3765 a_24158_13700# a_23737_13700# a_23110_13025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3766 a_40542_6967# a_41635_7629# a_41586_7819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3767 gnd d0 a_52594_7637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3768 a_10726_446# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3769 a_68780_11575# a_68359_11575# a_68681_11575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3770 a_74016_13656# a_74012_13833# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3771 a_19920_10006# a_20173_9993# a_18868_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3772 a_8163_11536# a_9256_12198# a_9211_12211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3773 gnd a_31138_10676# a_30930_10676# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3774 gnd d2 a_6970_9236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3775 gnd a_84976_3215# a_84768_3215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3776 a_3554_11577# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3777 a_51289_7152# a_52386_6958# a_52341_6971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3778 a_74012_13833# a_74269_13643# a_72968_12981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3779 vdd a_52597_9999# a_52389_9999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3780 a_79389_11569# a_79025_10047# a_77999_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3781 a_68529_13020# a_68316_13020# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3782 a_71520_3239# a_73012_3993# a_72963_4183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3783 a_3510_4047# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3784 a_67290_12253# a_66869_12253# a_66242_11578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3785 gnd d3 a_60767_10675# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3786 a_84723_3228# a_84719_3405# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3787 a_33819_10052# a_33398_10052# a_32990_10160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3788 a_76122_8968# a_76122_8713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3789 a_83674_6967# a_84767_7629# a_84722_7642# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3790 a_2063_3280# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3791 gnd d0 a_41846_10670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3792 vdd a_19125_8550# a_18917_8550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3793 a_65819_7696# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3794 gnd d1 a_30090_8554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3795 a_65820_4729# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3796 a_2064_12255# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3797 a_17424_12210# a_17677_12197# a_17382_10688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3798 a_72967_2559# a_74060_3221# a_74011_3411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3799 a_76528_2597# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3800 a_22902_13704# a_22689_13704# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3801 a_63046_2728# a_63303_2538# a_61998_2732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3802 a_65412_4158# a_66033_4050# a_66241_4050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3803 a_45195_4727# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3804 a_2483_6247# a_3722_7014# a_3879_5688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3805 a_79236_4039# a_79023_4039# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3806 a_34446_9280# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3807 gnd d0 a_63305_8546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3808 a_71473_4861# a_71565_3226# a_71520_3239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3809 gnd a_9462_5511# a_9254_5511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3810 gnd a_62255_2542# a_62047_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3811 a_47006_5569# a_46642_4047# a_45616_4727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3812 a_34443_7686# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3813 a_8164_8569# a_9257_9231# a_9208_9421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3814 a_65411_7380# a_66032_7696# a_66240_7696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3815 a_55275_5566# a_54854_5566# a_54447_5060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3816 vdd d0 a_52596_12198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3817 a_33816_7011# a_33395_7011# a_32987_6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3818 a_11314_6324# a_11314_5929# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3819 a_66867_6245# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3820 vdd d0 a_31136_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3821 a_29831_4183# a_30928_3989# a_30879_4179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3822 a_51289_5705# a_51546_5515# a_49842_6385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3823 a_14473_5563# a_14260_5563# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3824 a_9208_10868# a_9212_10012# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3825 a_1436_4052# a_1015_4052# a_607_4160# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3826 a_45617_12255# a_46856_13022# a_47013_11696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3827 a_72965_10191# a_73222_10001# a_71522_9247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3828 a_48518_4733# a_48097_4733# a_48419_4733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3829 a_33817_4044# a_34657_4719# a_34865_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3830 a_28383_6383# a_28640_6193# a_28345_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3831 vdd a_31138_10676# a_30930_10676# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3832 vdd d2 a_6970_9236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3833 vdd a_84976_3215# a_84768_3215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3834 a_56325_12249# a_55904_12249# a_55277_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3835 a_65821_11578# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3836 a_25549_11575# a_25185_10053# a_24159_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3837 a_76121_11680# a_76122_11066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3838 a_19913_5695# a_20170_5505# a_18865_5699# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3839 a_9207_11709# a_9212_10691# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3840 a_12986_9282# a_12773_9282# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3841 vdd d3 a_60767_10675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3842 a_33611_8605# a_33398_8605# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3843 gnd a_52596_12966# a_52388_12966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3844 a_55070_10733# a_54857_10733# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3845 a_54855_4725# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3846 a_76120_5058# a_76120_4802# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3847 vdd d0 a_41846_10670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3848 a_21685_433# a_32399_444# a_32721_444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3849 a_33610_13698# a_33397_13698# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3850 a_52343_12211# a_52596_12198# a_51295_11536# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3851 a_45197_10735# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3852 a_22279_8031# a_22903_8611# a_23111_8611# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3853 a_63049_6965# a_63045_7142# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3854 a_65414_10421# a_65414_10166# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3855 vdd d1 a_30090_8554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3856 a_1435_7019# a_2275_7694# a_2483_7694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3857 a_76742_11572# a_76529_11572# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3858 a_54446_7771# a_55067_7692# a_55275_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3859 a_72967_2559# a_74060_3221# a_74015_3234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3860 a_33819_9284# a_34659_9280# a_34867_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3861 gnd a_48991_7646# a_48783_7646# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3862 a_9210_3236# a_9206_3413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3863 a_19914_4175# a_20171_3985# a_18866_4179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3864 vdd a_41845_12958# a_41637_12958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3865 vdd d0 a_63305_8546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3866 vdd a_9462_5511# a_9254_5511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3867 gnd d0 a_63304_12960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3868 vdd a_31138_9229# a_30930_9229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3869 a_60512_4680# a_60599_6189# a_60554_6202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3870 a_72965_10191# a_74062_9997# a_74013_10187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3871 a_29837_8567# a_30930_9229# a_30881_9419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3872 a_54854_7013# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3873 vdd a_62255_2542# a_62047_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3874 gnd a_82440_10673# a_82232_10673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3875 a_26714_8602# a_26293_8602# a_25648_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3876 gnd d1 a_51546_6962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3877 a_8164_8569# a_9257_9231# a_9212_9244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3878 a_12144_3278# a_11723_3278# a_11315_2962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3879 a_59446_7653# a_60559_10675# a_60510_10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3880 a_28390_9247# a_29882_10001# a_29837_10014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3881 vdd a_40795_6954# a_40587_6954# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3882 a_40545_10008# a_41638_10670# a_41589_10860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3883 a_66035_8611# a_65822_8611# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3884 a_69770_4731# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3885 a_49844_12393# a_50101_12203# a_49806_10694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3886 gnd a_83927_5507# a_83719_5507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3887 a_14589_11690# a_14219_13016# a_13193_13696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3888 a_39098_9241# a_40590_9995# a_40545_10008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3889 a_79486_5561# a_80346_8596# a_80554_8596# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3890 gnd a_31136_2542# a_30928_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3891 a_608_13390# a_608_13135# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3892 a_28347_10692# a_28600_10679# a_27279_7657# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3893 a_67291_10733# a_66870_10733# a_66243_10737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3894 a_77791_9280# a_77578_9280# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3895 gnd d0 a_20170_6952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3896 a_56325_13696# a_57564_13016# a_57721_11690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3897 a_72968_12981# a_73221_12968# a_71521_12214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3898 a_8158_2738# a_9255_2544# a_9206_2734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3899 a_55277_13700# a_54856_13700# a_54448_13384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3900 gnd a_84977_13637# a_84769_13637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3901 a_40541_8738# a_40798_8548# a_39094_9418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3902 a_65413_12592# a_65413_12336# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3903 a_2065_10735# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3904 a_8161_6975# a_8414_6962# a_6714_6208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3905 a_62003_12977# a_63096_13639# a_63047_13829# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3906 a_22690_10058# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3907 a_11315_4154# a_11315_3613# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3908 a_55903_4721# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3909 a_30880_12386# a_30884_11530# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3910 a_52344_9244# a_52597_9231# a_51296_8569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3911 a_55278_10054# a_54857_10054# a_54449_10162# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3912 a_6716_12216# a_8208_12970# a_8159_13160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3913 a_65413_13388# a_66034_13704# a_66242_13704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3914 a_74016_12977# a_74269_12964# a_72964_13158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3915 vdd a_48991_7646# a_48783_7646# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3916 a_44146_6251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3917 a_33611_10052# a_33398_10052# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3918 a_12146_8607# a_11725_8607# a_11314_8027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3919 a_67081_3278# a_66868_3278# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3920 a_67289_4725# a_66868_4725# a_66241_4050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3921 a_44361_13706# a_44148_13706# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3922 a_6710_6385# a_6967_6195# a_6672_4686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3923 a_43009_401# a_42796_401# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3924 a_83670_7144# a_84767_6950# a_84718_7140# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3925 a_55067_6245# a_54854_6245# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3926 a_18870_2555# a_19123_2542# a_17419_3412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3927 a_1437_12259# a_1016_12259# a_608_11943# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3928 a_49806_10694# a_49893_12203# a_49844_12393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3929 a_30881_10187# a_30885_9242# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3930 a_51296_10016# a_51549_10003# a_49849_9249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3931 a_23738_9286# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3932 a_11935_6245# a_11722_6245# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3933 a_44568_3284# a_45408_3280# a_45616_3280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3934 a_65411_5678# a_66032_5570# a_66240_5570# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3935 vdd a_28642_12201# a_28434_12201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3936 gnd a_82482_12195# a_82274_12195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3937 vdd a_82440_10673# a_82232_10673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3938 gnd a_63305_8546# a_63097_8546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3939 a_606_7127# a_606_6586# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3940 a_49804_4686# a_49891_6195# a_49846_6208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3941 a_59446_7653# a_60559_10675# a_60514_10688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3942 a_23108_7696# a_23948_7692# a_24156_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3943 a_76120_4152# a_76741_4044# a_76949_4044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3944 a_32988_3611# a_33609_4044# a_33817_4044# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3945 a_9210_4683# a_9463_4670# a_8162_4008# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3946 a_40545_10008# a_41638_10670# a_41593_10683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3947 a_25552_5686# a_25182_7012# a_24156_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3948 vdd a_73220_3993# a_73012_3993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3949 a_74015_4002# a_74268_3989# a_72963_4183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3950 a_49844_12393# a_51340_11523# a_51291_11713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3951 a_45409_13702# a_45196_13702# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3952 a_2276_4727# a_2063_4727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3953 a_29830_5703# a_30927_5509# a_30878_5699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3954 a_28389_12214# a_29881_12968# a_29832_13158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3955 vdd a_31136_2542# a_30928_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3956 a_14260_5563# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3957 a_32989_12330# a_32989_11935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3958 a_76119_7374# a_76740_7690# a_76948_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3959 a_11317_10812# a_11938_10733# a_12146_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3960 a_1435_5572# a_1014_5572# a_606_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3961 a_74016_13656# a_76121_13777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3962 a_84724_12203# a_84977_12190# a_83676_11528# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3963 a_23111_9290# a_22690_9290# a_22282_8974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3964 a_54449_9365# a_54449_8970# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3965 a_8158_2738# a_9255_2544# a_9210_2557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3966 a_17422_6202# a_17675_6189# a_17380_4680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3967 vdd a_17633_4667# a_17425_4667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3968 a_32990_11066# a_33610_11572# a_33818_11572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3969 a_41588_12380# a_41845_12190# a_40544_11528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3970 gnd d0 a_52594_6958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3971 vdd d0 a_41843_5503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3972 a_79394_11688# a_79024_13014# a_77998_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3973 a_47008_11577# a_46644_10055# a_45618_9288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3974 a_11937_11574# a_11724_11574# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3975 a_56326_9282# a_55905_9282# a_55278_8607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3976 a_57563_4041# a_57350_4041# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3977 gnd a_31138_9997# a_30930_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3978 a_12773_9282# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3979 a_52340_9421# a_52597_9231# a_51296_8569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3980 a_43741_8976# a_44362_9292# a_44570_9292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3981 a_76740_6243# a_76527_6243# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3982 a_1230_10060# a_1017_10060# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3983 a_9205_6380# a_9462_6190# a_8161_5528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3984 a_2484_4727# a_3723_4047# a_3874_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3985 gnd a_19124_11517# a_18916_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3986 a_12143_7692# a_11722_7692# a_11314_7771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3987 a_61997_7146# a_62254_6956# a_60554_6202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3988 a_56115_6241# a_55902_6241# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3989 vdd d0 a_41844_3983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3990 a_80346_8596# a_80133_8596# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3991 a_18866_2732# a_19123_2542# a_17419_3412# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3992 a_1229_11580# a_1016_11580# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3993 gnd d0 a_41846_9991# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3994 a_83675_4000# a_83928_3987# a_82228_3233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3995 a_65412_4808# a_66033_4729# a_66241_4729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3996 a_76950_13698# a_77790_13694# a_77998_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3997 a_74017_9242# a_74270_9229# a_72969_8567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3998 vdd a_63305_8546# a_63097_8546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3999 a_29834_6973# a_30087_6960# a_28387_6206# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4000 a_52342_2557# a_52595_2544# a_51290_2738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4001 a_30884_11530# a_30880_11707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4002 a_12146_8607# a_12986_9282# a_13194_9282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4003 a_66868_3278# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4004 a_22902_13025# a_22689_13025# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4005 a_6668_4863# a_6760_3228# a_6715_3241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4006 a_56117_13696# a_55904_13696# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4007 gnd a_51546_6962# a_51338_6962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4008 a_30883_3234# a_31136_3221# a_29835_2559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4009 a_9206_4860# a_9463_4670# a_8162_4008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4010 a_43738_7777# a_43738_7382# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4011 a_49844_12393# a_51340_11523# a_51295_11536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4012 a_84723_3228# a_84976_3215# a_83675_2553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4013 a_74010_7146# a_74014_6201# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4014 a_66034_12257# a_65821_12257# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4015 gnd a_52595_3223# a_52387_3223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4016 gnd a_73219_5513# a_73011_5513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4017 a_77788_6239# a_77575_6239# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4018 a_65822_8611# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4019 a_14430_7008# a_14217_7008# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4020 a_65411_6584# a_66032_7017# a_66240_7017# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4021 a_67291_9286# a_68530_10053# a_68681_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4022 a_22279_6328# a_22279_5933# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4023 a_84718_5693# a_84723_4675# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4024 a_19915_13150# a_19919_12205# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4025 a_34867_10727# a_36106_10047# a_36257_11569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4026 vdd d4 a_81372_7638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4027 vdd a_74269_11517# a_74061_11517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4028 a_23950_12253# a_23737_12253# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4029 a_14433_10049# a_14220_10049# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4030 vdd a_73221_12968# a_73013_12968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4031 a_51291_11713# a_52388_11519# a_52343_11532# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4032 vdd a_84978_9991# a_84770_9991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4033 a_62000_8740# a_63097_8546# a_63048_8736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4034 a_606_6586# a_606_6330# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4035 a_39092_3410# a_40588_2540# a_40539_2730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4036 a_52342_4683# a_52338_4860# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4037 gnd d1 a_40797_11515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4038 a_1438_10739# a_1017_10739# a_609_10818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4039 a_62000_10187# a_63097_9993# a_63052_10006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4040 a_1436_4731# a_2276_4727# a_2484_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4041 a_32989_11935# a_32989_11680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4042 a_44361_11580# a_44148_11580# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4043 a_46855_4047# a_46642_4047# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4044 a_25185_10053# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4045 a_45615_7694# a_45194_7694# a_44567_7019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4046 a_63049_7644# a_63045_7821# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4047 vdd d0 a_9464_11519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4048 gnd d0 a_63303_4664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4049 a_76122_9619# a_76122_9363# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4050 a_30882_6201# a_30878_6378# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4051 a_55276_3278# a_54855_3278# a_54447_3357# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4052 a_54855_4046# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4053 a_55070_10054# a_54857_10054# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4054 a_1438_9292# a_1017_9292# a_609_8976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4055 a_63052_9238# a_63305_9225# a_62004_8563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4056 a_23109_2603# a_22688_2603# a_22280_2711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4057 vdd d1 a_8416_12970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4058 a_27279_7657# a_28392_10679# a_28347_10692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4059 a_29837_10014# a_30090_10001# a_28390_9247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4060 a_52338_2734# a_52595_2544# a_51290_2738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4061 a_76949_2597# a_76528_2597# a_76120_2705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4062 gnd d0 a_63304_13639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4063 a_65414_8974# a_66035_9290# a_66243_9290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4064 a_11722_6245# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4065 a_43741_2614# a_44360_2605# a_44568_2605# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4066 a_30879_3411# a_31136_3221# a_29835_2559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4067 a_34865_4719# a_34444_4719# a_33817_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4068 a_30878_7146# a_31135_6956# a_29830_7150# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4069 a_84719_3405# a_84976_3215# a_83675_2553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4070 a_1227_6251# a_1014_6251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4071 a_76119_5672# a_76740_5564# a_76948_5564# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4072 a_32988_5058# a_33608_5564# a_33816_5564# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4073 gnd d0 a_31138_9229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4074 a_55275_6245# a_56115_6241# a_56323_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4075 vdd a_52595_3223# a_52387_3223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4076 vdd a_73219_5513# a_73011_5513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4077 a_36354_5561# a_35933_5561# a_36260_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4078 a_2486_10735# a_3725_10055# a_3876_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4079 a_74014_5522# a_74267_5509# a_72962_5703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4080 a_67290_13700# a_66869_13700# a_66242_13025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4081 a_30880_13154# a_31137_12964# a_29832_13158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4082 a_12145_12253# a_12985_12249# a_13193_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4083 a_44569_11580# a_45409_12255# a_45617_12255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4084 a_23108_6249# a_22687_6249# a_22279_5933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4085 a_2063_4727# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4086 a_40541_10185# a_41638_9991# a_41589_10181# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4087 gnd d2 a_39348_6187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4088 a_76120_4407# a_76120_4152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4089 a_33608_7690# a_33395_7690# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4090 a_77577_13694# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4091 vdd d0 a_31137_12196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4092 a_2064_13702# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4093 a_44148_12259# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4094 a_54449_11068# a_55069_11574# a_55277_11574# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4095 a_40540_13152# a_40797_12962# a_39097_12208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4096 a_63047_12382# a_63304_12192# a_62003_11530# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4097 a_24158_12253# a_25397_13020# a_25554_11694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4098 a_62000_8740# a_63097_8546# a_63052_8559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4099 a_49847_3241# a_51339_3995# a_51290_4185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4100 a_59127_4727# a_59018_4727# a_54180_446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4101 vdd a_41843_5503# a_41635_5503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4102 vdd d1 a_40797_11515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4103 a_34867_9280# a_34446_9280# a_33819_8605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4104 a_39092_3410# a_40588_2540# a_40543_2553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4105 a_43740_13785# a_43740_13390# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4106 a_74012_13833# a_74016_12977# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4107 a_55277_13021# a_54856_13021# a_54448_12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4108 a_14475_11571# a_14262_11571# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4109 a_55278_8607# a_54857_8607# a_54449_8715# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4110 a_1227_7019# a_1014_7019# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4111 a_11315_4804# a_11315_4409# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4112 gnd a_84977_12958# a_84769_12958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4113 a_57350_4041# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4114 a_9207_12388# a_9211_11532# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4115 a_28384_3416# a_29880_2546# a_29831_2736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4116 a_22280_4158# a_22280_3617# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4117 a_22279_5933# a_22279_5678# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4118 vdd d1 a_83927_6954# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4119 vdd d0 a_63303_4664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4120 a_5386_4733# a_4965_4733# a_5041_8604# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4121 a_35893_10047# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4122 a_63048_9415# a_63305_9225# a_62004_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4123 a_66867_7692# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4124 a_51294_2561# a_52387_3223# a_52338_3413# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4125 a_11936_3278# a_11723_3278# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4126 a_74011_4858# a_74015_4002# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4127 gnd a_62257_9997# a_62049_9997# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4128 a_11724_12253# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4129 a_58673_8598# a_58460_8598# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4130 a_66035_10737# a_65822_10737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4131 vdd a_41844_3983# a_41636_3983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4132 a_80133_8596# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4133 a_71519_6206# a_71772_6193# a_71477_4684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4134 gnd d0 a_74268_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4135 a_65413_12592# a_66034_13025# a_66242_13025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4136 a_29836_11534# a_30089_11521# a_28385_12391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4137 a_48310_4733# a_48097_4733# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4138 a_83674_5520# a_83927_5507# a_82223_6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4139 a_83674_6967# a_84767_7629# a_84718_7819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4140 a_25547_5567# a_25183_4045# a_24157_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4141 a_44361_13027# a_44148_13027# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4142 a_66242_12257# a_65821_12257# a_65413_12336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4143 a_54449_11068# a_54449_10812# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4144 a_56325_13696# a_55904_13696# a_55277_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4145 vdd d1 a_19125_9997# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4146 a_24157_3278# a_23736_3278# a_23109_3282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4147 a_63050_2551# a_63303_2538# a_61998_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4148 gnd a_17676_3222# a_17468_3222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4149 a_6717_9249# a_6970_9236# a_6670_10871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4150 a_9210_4004# a_9463_3991# a_8158_4185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4151 a_18871_11530# a_19964_12192# a_19919_12205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4152 a_19920_10006# a_19916_10183# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4153 a_44567_5572# a_45407_6247# a_45615_6247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4154 a_43739_2713# a_43741_2614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4155 a_77575_6239# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4156 a_52343_13658# a_52596_13645# a_51295_12983# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4157 a_41590_6963# a_41586_7140# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4158 a_74017_10689# a_74013_10866# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4159 vdd a_81372_7638# a_81164_7638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4160 a_11317_10162# a_11938_10054# a_12146_10054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4161 gnd d1 a_73222_8554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4162 a_68359_11575# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4163 a_606_6330# a_1227_6251# a_1435_6251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4164 a_11938_8607# a_11725_8607# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4165 a_76741_3276# a_76528_3276# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4166 a_22901_4729# a_22688_4729# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4167 a_40541_8738# a_41638_8544# a_41589_8734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4168 gnd d0 a_52597_8552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4169 a_17419_3412# a_18915_2542# a_18866_2732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4170 a_3512_10055# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4171 a_609_9371# a_609_8976# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4172 a_56116_3274# a_55903_3274# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4173 a_32990_9363# a_33611_9284# a_33819_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4174 a_28384_3416# a_29880_2546# a_29835_2559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4175 a_12144_4725# a_11723_4725# a_11315_4409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4176 a_12772_12249# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4177 a_9208_10868# a_9465_10678# a_8164_10016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4178 a_43118_401# a_64495_433# a_64817_433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4179 a_1230_10739# a_1017_10739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4180 a_51294_2561# a_52387_3223# a_52342_3236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4181 a_64495_433# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4182 a_44568_3284# a_44147_3284# a_43739_3363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4183 a_29836_11534# a_30929_12196# a_30884_12209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4184 a_54856_11574# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4185 a_76948_7011# a_76527_7011# a_76119_6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4186 a_21685_433# a_21576_433# a_21784_433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4187 gnd a_63303_4664# a_63095_4664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4188 a_54854_5566# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4189 a_46641_7014# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4190 vdd d0 a_74268_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4191 a_57605_5563# a_57392_5563# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4192 a_29832_11711# a_30089_11521# a_28385_12391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4193 a_33816_6243# a_33395_6243# a_32987_6322# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4194 a_12146_10054# a_12986_10729# a_13194_10729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4195 a_12143_7013# a_11722_7013# a_11314_7121# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4196 a_57562_7008# a_57349_7008# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4197 a_76529_12251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4198 a_65414_10166# a_65414_9625# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4199 a_72966_5526# a_74059_6188# a_74010_6378# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4200 a_76949_4044# a_77789_4719# a_77997_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4201 vdd a_9464_12198# a_9256_12198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4202 vdd d0 a_63305_9993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4203 a_22903_9290# a_22690_9290# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4204 a_65411_7775# a_65411_7380# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4205 a_9211_11532# a_9207_11709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4206 a_44149_10739# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4207 vdd a_17676_3222# a_17468_3222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4208 a_11314_7771# a_11314_7376# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4209 a_9206_3413# a_9210_2557# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4210 a_83677_10008# a_84770_10670# a_84721_10860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4211 a_6713_9426# a_6970_9236# a_6670_10871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4212 gnd d1 a_19124_12964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4213 a_19920_8559# a_19916_8736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4214 gnd a_31138_9229# a_30930_9229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4215 a_55070_9286# a_54857_9286# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4216 gnd d2 a_60807_6189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4217 vdd d2 a_6968_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4218 a_52339_13835# a_52596_13645# a_51295_12983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4219 a_67290_13700# a_68529_13020# a_68686_11694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4220 a_44149_9292# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4221 a_76743_8605# a_76530_8605# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4222 a_80478_4725# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4223 a_30879_2732# a_22282_2612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4224 a_44570_8613# a_44149_8613# a_43738_8033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4225 gnd a_39348_6187# a_39140_6187# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4226 vdd d1 a_73222_8554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4227 a_33395_7690# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4228 a_67081_4725# a_66868_4725# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4229 a_61999_13154# a_62256_12964# a_60556_12210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4230 gnd d0 a_20173_10672# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4231 a_22282_11072# a_22282_10816# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4232 a_17425_9243# a_18917_9997# a_18872_10010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4233 a_11935_7692# a_11722_7692# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4234 a_1437_13706# a_1016_13706# a_608_13390# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4235 a_76951_9284# a_77791_9280# a_77999_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4236 a_17419_3412# a_18915_2542# a_18870_2555# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4237 a_37668_4725# a_37559_4725# a_32721_444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4238 a_40541_8738# a_41638_8544# a_41593_8557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4239 vdd d0 a_52597_8552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4240 a_25184_13020# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4241 vdd a_74270_9229# a_74062_9229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4242 a_1014_7698# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4243 a_69846_8602# a_69425_8602# a_68780_11575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4244 a_40545_8561# a_40798_8548# a_39094_9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4245 a_45408_3280# a_45195_3280# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4246 a_1438_10060# a_1017_10060# a_609_10168# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4247 a_57352_10049# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4248 a_52344_9244# a_52340_9421# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4249 a_28345_4684# a_28432_6193# a_28383_6383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4250 a_29835_2559# a_30928_3221# a_30879_3411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4251 vdd d1 a_40796_3987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4252 vdd a_63303_4664# a_63095_4664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4253 a_60554_6202# a_62046_6956# a_61997_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4254 vdd a_83927_6954# a_83719_6954# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4255 a_43738_5680# a_43739_5066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4256 a_43740_12338# a_44361_12259# a_44569_12259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4257 a_11723_3278# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4258 a_6717_9249# a_8209_10003# a_8164_10016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4259 a_58460_8598# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4260 a_68778_5567# a_69638_8602# a_69846_8602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4261 a_18869_5522# a_19962_6184# a_19913_6374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4262 gnd d0 a_63303_3985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4263 a_11317_8970# a_11317_8715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4264 a_32988_2705# a_33609_2597# a_33817_2597# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4265 a_1228_3284# a_1015_3284# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4266 a_26851_4731# a_26638_4731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4267 gnd a_74268_2542# a_74060_2542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4268 a_609_8976# a_609_8721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4269 a_3724_13022# a_3511_13022# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4270 a_76951_10731# a_77791_10727# a_77999_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4271 a_83677_10008# a_84770_10670# a_84725_10683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4272 a_32990_8713# a_32987_8025# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4273 a_71519_6206# a_73011_6960# a_72966_6973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4274 a_56118_10729# a_55905_10729# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4275 a_36260_5680# a_35890_7006# a_34864_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4276 a_57719_5682# a_57605_5563# a_57813_5563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4277 a_37983_7828# a_38240_7638# a_37668_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4278 a_52342_2557# a_52338_2734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4279 a_12773_10729# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4280 a_52340_10189# a_52597_9999# a_51292_10193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4281 a_62002_4002# a_63095_4664# a_63046_4854# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4282 vdd d0 a_20173_10672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4283 a_63049_5518# a_63045_5695# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4284 a_84718_6372# a_84722_5516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4285 a_14219_13016# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4286 a_1016_11580# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4287 gnd a_73222_8554# a_73014_8554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4288 a_66241_4729# a_65820_4729# a_65412_4808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4289 a_44570_10060# a_44149_10060# a_43741_9627# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4290 a_17424_12210# a_18916_12964# a_18867_13154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4291 a_11725_8607# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4292 a_44359_7698# a_44146_7698# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4293 a_44147_2605# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4294 a_66868_4725# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4295 vdd a_20172_12960# a_19964_12960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4296 gnd a_17633_4667# a_17425_4667# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4297 a_34657_3272# a_34444_3272# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4298 gnd a_60767_10675# a_60559_10675# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4299 a_55068_2599# a_54855_2599# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4300 a_84719_4173# a_84723_3228# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4301 a_22280_4808# a_22280_4413# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4302 a_66240_7696# a_67080_7692# a_67288_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4303 a_29835_2559# a_30928_3221# a_30883_3234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4304 a_66034_13704# a_65821_13704# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4305 a_44569_11580# a_44148_11580# a_43740_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4306 a_29830_7150# a_30927_6956# a_30882_6969# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4307 gnd d2 a_82481_3220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4308 gnd d3 a_6925_4673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4309 a_68684_5686# a_68314_7012# a_67288_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4310 a_76120_2960# a_76741_3276# a_76949_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4311 a_32988_3355# a_32988_2960# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4312 a_13192_3274# a_14431_4041# a_14582_5563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4313 a_84720_13827# a_84977_13637# a_83676_12975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4314 a_54448_13129# a_54448_12588# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4315 a_18869_5522# a_19962_6184# a_19917_6197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4316 a_22902_11578# a_22689_11578# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4317 vdd a_74268_2542# a_74060_2542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4318 a_57392_5563# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4319 vdd d1 a_30089_12968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4320 a_74013_9419# a_74017_8563# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4321 a_607_5066# a_607_4810# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4322 a_19919_12205# a_20172_12192# a_18871_11530# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4323 a_66035_10058# a_65822_10058# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4324 a_59127_4727# a_59491_7640# a_59442_7830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4325 a_66243_9290# a_65822_9290# a_65414_8974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4326 a_22690_9290# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4327 vdd d0 a_84975_5503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4328 a_77998_12247# a_79237_13014# a_79394_11688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4329 a_24158_12253# a_23737_12253# a_23110_12257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4330 a_30883_4681# a_30879_4858# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4331 vdd a_52596_12198# a_52388_12198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4332 a_41586_5693# a_41843_5503# a_40538_5697# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4333 a_25646_5567# a_25225_5567# a_25552_5686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4334 a_57564_13016# a_57351_13016# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4335 a_6672_4686# a_6759_6195# a_6710_6385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4336 a_11315_2707# a_11317_2608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4337 a_32721_444# a_32612_444# a_21685_433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4338 a_43740_11688# a_43741_11074# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4339 a_55905_9282# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4340 gnd a_60807_6189# a_60599_6189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4341 vdd a_6968_3228# a_6760_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4342 a_66242_13025# a_67082_13700# a_67290_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4343 a_41590_7642# a_41586_7819# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4344 a_6668_4863# a_6760_3228# a_6711_3418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4345 a_62002_4002# a_63095_4664# a_63050_4677# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4346 gnd a_8416_12970# a_8208_12970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4347 a_33818_12251# a_33397_12251# a_32989_12330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4348 a_76530_8605# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4349 a_55276_4725# a_54855_4725# a_54447_4804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4350 a_52343_12979# a_52596_12966# a_51291_13160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4351 vdd d2 a_39350_12195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4352 vdd d0 a_84976_3983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4353 a_43741_10423# a_44362_10739# a_44570_10739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4354 vdd a_73222_8554# a_73014_8554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4355 a_72963_4183# a_74060_3989# a_74015_4002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4356 a_77578_10727# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4357 a_76119_8025# a_76743_8605# a_76951_8605# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4358 a_11722_7692# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4359 a_41587_4173# a_41844_3983# a_40539_4177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4360 gnd d1 a_83929_11515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4361 gnd d4 a_81372_7638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4362 a_8163_11536# a_8416_11523# a_6712_12393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4363 gnd a_74269_11517# a_74061_11517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4364 a_43738_8033# a_43738_7777# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4365 vdd a_60767_10675# a_60559_10675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4366 a_55278_8607# a_56118_9282# a_56326_9282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4367 a_1015_2605# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4368 a_54449_10417# a_54449_10162# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4369 vdd d2 a_82481_3220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4370 a_46642_4047# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4371 a_22901_4050# a_22688_4050# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4372 a_39055_10686# a_39142_12195# a_39093_12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4373 a_51291_11713# a_52388_11519# a_52339_11709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4374 a_6711_3418# a_8207_2548# a_8162_2561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4375 vdd d3 a_6925_4673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4376 a_74015_3234# a_74268_3221# a_72967_2559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4377 a_33817_3276# a_33396_3276# a_32988_2960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4378 a_44569_13027# a_45409_13702# a_45617_13702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4379 a_45195_3280# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4380 a_12144_4046# a_11723_4046# a_11315_3613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4381 a_33818_13019# a_33397_13019# a_32989_12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4382 vdd a_40796_3987# a_40588_3987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4383 vdd d1 a_40795_5507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4384 a_23948_6245# a_23735_6245# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4385 a_33397_13698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4386 gnd d0 a_84977_11511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4387 a_59127_4727# a_59491_7640# a_59446_7653# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4388 a_44148_13706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4389 a_2278_9288# a_2065_9288# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4390 a_63045_7821# a_63049_6965# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4391 gnd a_63303_3985# a_63095_3985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4392 gnd d0 a_63302_5505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4393 gnd d0 a_9464_11519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4394 a_65414_10816# a_65414_10421# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4395 a_53858_446# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4396 a_79280_11569# a_79067_11569# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4397 a_27279_7657# a_28392_10679# a_28343_10869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4398 a_8161_5528# a_9254_6190# a_9205_6380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4399 a_34865_3272# a_36104_4039# a_36255_5561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4400 a_34866_12247# a_34445_12247# a_33818_11572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4401 a_44149_10060# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4402 a_82226_9418# a_82483_9228# a_82183_10863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4403 a_83673_10185# a_84770_9991# a_84721_10181# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4404 vdd a_28640_6193# a_28432_6193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4405 a_82228_3233# a_83720_3987# a_83675_4000# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4406 vdd d2 a_6969_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4407 a_74017_8563# a_74013_8740# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4408 a_11936_4725# a_11723_4725# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4409 vdd d0 a_74269_12196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4410 vdd d1 a_8415_3995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4411 gnd d0 a_52595_4670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4412 a_40543_4000# a_41636_4662# a_41587_4852# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4413 a_44359_5572# a_44146_5572# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4414 vdd a_20170_5505# a_19962_5505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4415 a_54448_12588# a_54448_12332# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4416 a_44360_2605# a_44147_2605# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4417 a_609_11074# a_1229_11580# a_1437_11580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4418 vdd d1 a_83929_11515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4419 a_33819_8605# a_33398_8605# a_32987_8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4420 a_608_13785# a_608_13390# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4421 a_54855_3278# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4422 a_66242_13704# a_65821_13704# a_65413_13783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4423 a_84724_12971# a_84720_13148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4424 a_8159_11713# a_8416_11523# a_6712_12393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4425 gnd d0 a_20173_9993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4426 a_22688_2603# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4427 a_72968_11534# a_74061_12196# a_74012_12386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4428 a_55067_7013# a_54854_7013# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4429 a_55277_13700# a_56117_13696# a_56325_13696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4430 a_11935_7013# a_11722_7013# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4431 a_24157_4725# a_23736_4725# a_23109_4729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4432 a_1437_13027# a_1016_13027# a_608_12594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4433 a_23110_11578# a_22689_11578# a_22281_11686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4434 a_77997_4719# a_77576_4719# a_76949_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4435 a_66869_13700# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4436 a_74010_7146# a_74267_6956# a_72962_7150# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4437 a_74011_3411# a_74268_3221# a_72967_2559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4438 a_65411_5678# a_65412_5064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4439 a_3975_11577# a_3554_11577# a_3876_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4440 gnd a_63305_10672# a_63097_10672# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4441 vdd a_30090_10001# a_29882_10001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4442 vdd a_20171_3985# a_19963_3985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4443 a_65413_11686# a_66034_11578# a_66242_11578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4444 a_74016_12209# a_74012_12386# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4445 gnd a_6925_4673# a_6717_4673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4446 a_79486_5561# a_79065_5561# a_79392_5680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4447 vdd d0 a_84977_11511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4448 a_44567_7019# a_45407_7694# a_45615_7694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4449 a_54446_7376# a_54446_7121# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4450 gnd d1 a_19123_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4451 a_60553_9420# a_62049_8550# a_62000_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4452 a_609_8976# a_1230_9292# a_1438_9292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4453 gnd d2 a_28641_3226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4454 a_3879_5688# a_3765_5569# a_3973_5569# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4455 a_82225_12385# a_83721_11515# a_83672_11705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4456 vdd d0 a_52594_6190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4457 a_57813_5563# a_58673_8598# a_58881_8598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4458 a_22687_6249# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4459 a_2485_12255# a_2064_12255# a_1437_11580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4460 a_76741_4723# a_76528_4723# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4461 a_12146_10733# a_11725_10733# a_11317_10417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4462 a_21576_433# a_21363_433# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4463 a_37346_4725# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4464 vdd a_51548_12970# a_51340_12970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4465 a_22282_10421# a_22282_10166# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4466 a_28387_6206# a_29879_6960# a_29834_6973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4467 vdd a_84975_5503# a_84767_5503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4468 a_36106_10047# a_35893_10047# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4469 a_77999_9280# a_77578_9280# a_76951_8605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4470 a_56116_4721# a_55903_4721# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4471 a_51290_2738# a_51547_2548# a_49843_3418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4472 a_54857_8607# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4473 a_55277_12253# a_54856_12253# a_54448_12332# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4474 a_83672_11705# a_84769_11511# a_84720_11701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4475 a_65414_8719# a_66035_8611# a_66243_8611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4476 vdd d0 a_52595_4670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4477 a_40543_4000# a_41636_4662# a_41591_4675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4478 a_9205_7148# a_9209_6203# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4479 a_76740_7011# a_76527_7011# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4480 a_64817_433# a_75531_444# a_75853_444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4481 a_33610_12251# a_33397_12251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4482 a_83670_7144# a_83927_6954# a_82227_6200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4483 a_4965_4733# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4484 gnd d1 a_8414_5515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4485 a_23737_12253# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4486 vdd a_84976_3983# a_84768_3983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4487 a_61998_4179# a_62255_3989# a_60555_3235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4488 a_61998_4179# a_63095_3985# a_63046_4175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4489 vdd d1 a_73222_10001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4490 a_72966_6973# a_74059_7635# a_74010_7825# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4491 a_44570_10739# a_44149_10739# a_43741_10423# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4492 a_2483_6247# a_2062_6247# a_1435_5572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4493 a_19914_2728# a_20171_2538# a_18866_2732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4494 a_72967_2559# a_73220_2546# a_71516_3416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4495 a_68679_5567# a_68315_4045# a_67289_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4496 a_60556_12210# a_60809_12197# a_60514_10688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4497 gnd a_81372_7638# a_81164_7638# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4498 a_52341_6203# a_52594_6190# a_51293_5528# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4499 a_66241_4050# a_65820_4050# a_65412_4158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4500 a_36257_11569# a_36148_11569# a_36356_11569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4501 gnd d0 a_20173_8546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4502 a_6674_10694# a_6761_12203# a_6716_12216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4503 a_33397_11572# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4504 vdd a_63305_10672# a_63097_10672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4505 a_44359_7019# a_44146_7019# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4506 a_67289_3278# a_66868_3278# a_66241_3282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4507 a_22900_5570# a_22687_5570# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4508 a_47013_11696# a_46899_11577# a_47107_11577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4509 a_84720_11701# a_84725_10683# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4510 a_22280_4413# a_22901_4729# a_23109_4729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4511 vdd a_6925_4673# a_6717_4673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4512 a_71522_9247# a_73014_10001# a_72965_10191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4513 a_12143_5566# a_11722_5566# a_11315_5060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4514 gnd a_30089_12968# a_29881_12968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4515 a_8164_8569# a_8417_8556# a_6713_9426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4516 a_84721_8734# a_84722_7642# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4517 vdd a_40795_5507# a_40587_5507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4518 a_34867_10727# a_34446_10727# a_33819_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4519 a_60553_9420# a_62049_8550# a_62004_8563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4520 a_66034_13025# a_65821_13025# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4521 a_22281_12592# a_22281_12336# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4522 a_23735_6245# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4523 vdd d2 a_28641_3226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4524 a_82225_12385# a_83721_11515# a_83676_11528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4525 a_9212_10691# a_9465_10678# a_8164_10016# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4526 a_45618_10735# a_45197_10735# a_44570_10060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4527 a_2065_9288# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4528 gnd a_63302_5505# a_63094_5505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4529 a_33818_11572# a_34658_12247# a_34866_12247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4530 a_11317_9621# a_11317_9365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4531 a_34656_6239# a_34443_6239# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4532 a_3723_4047# a_3510_4047# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4533 a_39051_10863# a_39143_9228# a_39098_9241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4534 a_55904_13696# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4535 a_11314_6324# a_11935_6245# a_12143_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4536 a_609_9627# a_609_9371# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4537 a_14584_11571# a_14475_11571# a_14683_11571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4538 vdd a_50099_6195# a_49891_6195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4539 a_66033_4729# a_65820_4729# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4540 gnd a_31137_12196# a_30929_12196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4541 a_16314_7653# a_16567_7640# a_15995_4727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4542 a_22282_9369# a_22903_9290# a_23111_9290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4543 a_609_2614# a_1228_2605# a_1436_2605# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4544 a_83672_11705# a_84769_11511# a_84724_11524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4545 a_45408_4727# a_45195_4727# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4546 a_30885_9242# a_30881_9419# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4547 a_82181_4855# a_82273_3220# a_82224_3410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4548 a_22280_2711# a_22282_2612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4549 a_11723_4725# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4550 a_43740_13785# a_44361_13706# a_44569_13706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4551 vdd d1 a_8414_5515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4552 vdd d2 a_50101_12203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4553 gnd d2 a_6968_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4554 vdd a_8415_3995# a_8207_3995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4555 a_18869_6969# a_19962_7631# a_19913_7821# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4556 a_72966_6973# a_74059_7635# a_74014_7648# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4557 a_55276_4046# a_54855_4046# a_54447_4154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4558 a_1228_4731# a_1015_4731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4559 gnd d0 a_41845_12190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4560 a_3876_11577# a_3767_11577# a_3975_11577# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4561 a_72963_2736# a_73220_2546# a_71516_3416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4562 a_76948_6243# a_76527_6243# a_76119_6322# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4563 a_68317_10053# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4564 a_11314_8027# a_11314_7771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4565 gnd d1 a_73221_12968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4566 a_43741_9627# a_44362_10060# a_44570_10060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4567 vdd d0 a_20173_8546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4568 a_19913_7142# a_19917_6197# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4569 a_43738_5935# a_44359_6251# a_44567_6251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4570 a_607_4415# a_607_4160# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4571 a_23949_3278# a_23736_3278# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4572 a_2486_10735# a_2065_10735# a_1438_10739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4573 a_66035_9290# a_65822_9290# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4574 a_11722_7013# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4575 gnd d1 a_30088_2546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4576 a_30879_4179# a_31136_3989# a_29831_4183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4577 a_8160_8746# a_8417_8556# a_6713_9426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4578 a_47107_11577# a_47965_8604# a_48173_8604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4579 a_30883_2555# a_30879_2732# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4580 a_22690_10737# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4581 gnd a_74270_9229# a_74062_9229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4582 vdd d2 a_17675_6189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4583 vdd a_52595_3991# a_52387_3991# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4584 gnd d1 a_19122_5509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4585 a_60554_6202# a_60807_6189# a_60512_4680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4586 a_6711_3418# a_6968_3228# a_6668_4863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4587 gnd a_19123_3989# a_18915_3989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4588 a_52340_9421# a_52344_8565# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4589 a_23108_7017# a_22687_7017# a_22279_6584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4590 a_9206_4860# a_9210_4004# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4591 a_41590_5516# a_41586_5693# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4592 a_33397_13019# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4593 a_76527_7690# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4594 a_49846_6208# a_51338_6962# a_51293_6975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4595 a_44148_13027# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4596 a_33611_10731# a_33398_10731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4597 a_14587_5682# a_14217_7008# a_13191_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4598 a_43738_7127# a_44359_7019# a_44567_7019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4599 a_49800_4863# a_49892_3228# a_49847_3241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
C0 d0 vdd 85.85fF
C1 d5 d4 60.70fF
C2 d6 d7 59.65fF
C3 vdd d2 42.21fF
C4 vdd d4 2.34fF
C5 d0 d1 56.56fF
C6 d3 d2 62.10fF
C7 d3 d4 68.59fF
C8 d1 d2 51.15fF
C9 d6 a_21784_433# 5.71fF
C10 d0 d2 3.70fF
C11 d6 d8 12.82fF
C12 d5 vdd 2.38fF
C13 d3 d5 16.52fF
C14 d3 vdd 46.01fF
C15 d1 vdd 76.21fF
C16 a_64817_433# gnd 12.30fF
C17 a_54279_446# gnd 12.71fF
C18 a_43118_401# gnd 27.41fF
C19 d8 gnd 47.51fF
C20 a_21685_433# gnd 12.30fF
C21 a_21784_433# gnd 24.05fF
C22 d7 gnd 56.60fF
C23 a_11147_446# gnd 12.71fF
C24 d6 gnd 123.66fF
C25 a_84719_2726# gnd 2.27fF
C26 a_83671_2730# gnd 2.80fF
C27 a_76122_2606# gnd 17.59fF
C28 a_74011_2732# gnd 2.27fF
C29 a_72963_2736# gnd 2.80fF
C30 a_76120_2705# gnd 2.28fF
C31 a_65414_2612# gnd 17.59fF
C32 a_63046_2728# gnd 2.27fF
C33 a_61998_2732# gnd 2.80fF
C34 a_65412_2711# gnd 2.28fF
C35 a_54449_2608# gnd 17.59fF
C36 a_52338_2734# gnd 2.27fF
C37 a_51290_2738# gnd 2.80fF
C38 a_54447_2707# gnd 2.28fF
C39 a_43741_2614# gnd 17.59fF
C40 a_41587_2726# gnd 2.27fF
C41 a_40539_2730# gnd 2.80fF
C42 a_32990_2606# gnd 17.59fF
C43 a_30879_2732# gnd 2.27fF
C44 a_29831_2736# gnd 2.80fF
C45 a_43739_2713# gnd 2.28fF
C46 a_32988_2705# gnd 2.28fF
C47 a_22282_2612# gnd 17.59fF
C48 a_19914_2728# gnd 2.27fF
C49 a_18866_2732# gnd 2.80fF
C50 a_22280_2711# gnd 2.28fF
C51 a_11317_2608# gnd 17.59fF
C52 a_9206_2734# gnd 2.27fF
C53 a_8158_2738# gnd 2.80fF
C54 a_11315_2707# gnd 2.28fF
C55 a_609_2614# gnd 17.59fF
C56 a_607_2713# gnd 2.28fF
C57 a_84723_2549# gnd 3.17fF
C58 a_74015_2555# gnd 3.17fF
C59 a_63050_2551# gnd 3.17fF
C60 a_52342_2557# gnd 3.17fF
C61 a_41591_2549# gnd 3.17fF
C62 a_30883_2555# gnd 3.17fF
C63 a_83675_2553# gnd 3.33fF
C64 a_84719_3405# gnd 2.33fF
C65 a_82224_3410# gnd 4.37fF
C66 a_76949_2597# gnd 3.33fF
C67 a_19918_2551# gnd 3.17fF
C68 a_9210_2557# gnd 3.17fF
C69 a_76120_2960# gnd 3.17fF
C70 a_76949_3276# gnd 2.80fF
C71 a_72967_2559# gnd 3.33fF
C72 a_74011_3411# gnd 2.33fF
C73 a_71516_3416# gnd 4.37fF
C74 a_66241_2603# gnd 3.33fF
C75 a_76120_3355# gnd 2.27fF
C76 a_65412_2966# gnd 3.17fF
C77 a_66241_3282# gnd 2.80fF
C78 a_62002_2555# gnd 3.33fF
C79 a_63046_3407# gnd 2.33fF
C80 a_60551_3412# gnd 4.37fF
C81 a_55276_2599# gnd 3.33fF
C82 a_65412_3361# gnd 2.27fF
C83 a_54447_2962# gnd 3.17fF
C84 a_55276_3278# gnd 2.80fF
C85 a_51294_2561# gnd 3.33fF
C86 a_52338_3413# gnd 2.33fF
C87 a_49843_3418# gnd 4.37fF
C88 a_44568_2605# gnd 3.33fF
C89 a_54447_3357# gnd 2.27fF
C90 a_43739_2968# gnd 3.17fF
C91 a_44568_3284# gnd 2.80fF
C92 a_40543_2553# gnd 3.33fF
C93 a_41587_3405# gnd 2.33fF
C94 a_39092_3410# gnd 4.37fF
C95 a_33817_2597# gnd 3.33fF
C96 a_43739_3363# gnd 2.27fF
C97 a_32988_2960# gnd 3.17fF
C98 a_33817_3276# gnd 2.80fF
C99 a_29835_2559# gnd 3.33fF
C100 a_30879_3411# gnd 2.33fF
C101 a_28384_3416# gnd 4.37fF
C102 a_23109_2603# gnd 3.33fF
C103 a_32988_3355# gnd 2.27fF
C104 a_22280_2966# gnd 3.17fF
C105 a_23109_3282# gnd 2.80fF
C106 a_18870_2555# gnd 3.33fF
C107 a_19914_3407# gnd 2.33fF
C108 a_17419_3412# gnd 4.37fF
C109 a_12144_2599# gnd 3.33fF
C110 a_22280_3361# gnd 2.27fF
C111 a_11315_2962# gnd 3.17fF
C112 a_12144_3278# gnd 2.80fF
C113 a_8162_2561# gnd 3.33fF
C114 a_9206_3413# gnd 2.33fF
C115 a_6711_3418# gnd 4.37fF
C116 a_1436_2605# gnd 3.33fF
C117 a_11315_3357# gnd 2.27fF
C118 a_607_2968# gnd 3.17fF
C119 a_1436_3284# gnd 2.80fF
C120 a_607_3363# gnd 2.27fF
C121 a_84723_3228# gnd 3.43fF
C122 a_74015_3234# gnd 3.43fF
C123 a_63050_3230# gnd 3.43fF
C124 a_52342_3236# gnd 3.43fF
C125 a_41591_3228# gnd 3.43fF
C126 a_30883_3234# gnd 3.43fF
C127 a_84719_4173# gnd 2.27fF
C128 a_82228_3233# gnd 3.43fF
C129 a_83671_4177# gnd 2.80fF
C130 a_77997_3272# gnd 3.16fF
C131 a_76120_3611# gnd 3.43fF
C132 a_74011_4179# gnd 2.27fF
C133 a_71520_3239# gnd 3.43fF
C134 a_72963_4183# gnd 2.80fF
C135 a_67289_3278# gnd 3.16fF
C136 a_19918_3230# gnd 3.43fF
C137 a_9210_3236# gnd 3.43fF
C138 a_76120_4152# gnd 2.33fF
C139 a_65412_3617# gnd 3.43fF
C140 a_63046_4175# gnd 2.27fF
C141 a_60555_3235# gnd 3.43fF
C142 a_61998_4179# gnd 2.80fF
C143 a_56324_3274# gnd 3.16fF
C144 a_65412_4158# gnd 2.33fF
C145 a_54447_3613# gnd 3.43fF
C146 a_52338_4181# gnd 2.27fF
C147 a_49847_3241# gnd 3.43fF
C148 a_51290_4185# gnd 2.80fF
C149 a_45616_3280# gnd 3.16fF
C150 a_54447_4154# gnd 2.33fF
C151 a_43739_3619# gnd 3.43fF
C152 a_41587_4173# gnd 2.27fF
C153 a_39096_3233# gnd 3.43fF
C154 a_40539_4177# gnd 2.80fF
C155 a_34865_3272# gnd 3.16fF
C156 a_32988_3611# gnd 3.43fF
C157 a_30879_4179# gnd 2.27fF
C158 a_28388_3239# gnd 3.43fF
C159 a_29831_4183# gnd 2.80fF
C160 a_24157_3278# gnd 3.16fF
C161 a_43739_4160# gnd 2.33fF
C162 a_32988_4152# gnd 2.33fF
C163 a_22280_3617# gnd 3.43fF
C164 a_19914_4175# gnd 2.27fF
C165 a_17423_3235# gnd 3.43fF
C166 a_18866_4179# gnd 2.80fF
C167 a_13192_3274# gnd 3.16fF
C168 a_22280_4158# gnd 2.33fF
C169 a_11315_3613# gnd 3.43fF
C170 a_9206_4181# gnd 2.27fF
C171 a_6715_3241# gnd 3.43fF
C172 a_8158_4185# gnd 2.80fF
C173 a_2484_3280# gnd 3.16fF
C174 a_11315_4154# gnd 2.33fF
C175 a_607_3619# gnd 3.43fF
C176 a_607_4160# gnd 2.33fF
C177 a_84723_3996# gnd 3.17fF
C178 a_74015_4002# gnd 3.17fF
C179 a_63050_3998# gnd 3.17fF
C180 a_52342_4004# gnd 3.17fF
C181 a_41591_3996# gnd 3.17fF
C182 a_30883_4002# gnd 3.17fF
C183 a_83675_4000# gnd 3.33fF
C184 a_84719_4852# gnd 2.33fF
C185 a_82181_4855# gnd 3.27fF
C186 a_75853_444# gnd 10.85fF
C187 a_76949_4044# gnd 3.33fF
C188 a_77997_4719# gnd 3.64fF
C189 a_76120_4407# gnd 3.17fF
C190 a_76949_4723# gnd 2.80fF
C191 a_19918_3998# gnd 3.17fF
C192 a_9210_4004# gnd 3.17fF
C193 a_72967_4006# gnd 3.33fF
C194 a_74011_4858# gnd 2.33fF
C195 a_71473_4861# gnd 3.27fF
C196 a_76120_4802# gnd 2.27fF
C197 a_70191_4731# gnd 11.63fF
C198 a_66241_4050# gnd 3.33fF
C199 a_67289_4725# gnd 3.64fF
C200 a_65412_4413# gnd 3.17fF
C201 a_66241_4729# gnd 2.80fF
C202 a_62002_4002# gnd 3.33fF
C203 a_63046_4854# gnd 2.33fF
C204 a_60508_4857# gnd 3.27fF
C205 a_65412_4808# gnd 2.27fF
C206 a_54180_446# gnd 10.85fF
C207 a_55276_4046# gnd 3.33fF
C208 a_56324_4721# gnd 3.64fF
C209 a_54447_4409# gnd 3.17fF
C210 a_55276_4725# gnd 2.80fF
C211 a_51294_4008# gnd 3.33fF
C212 a_52338_4860# gnd 2.33fF
C213 a_49800_4863# gnd 3.27fF
C214 a_54447_4804# gnd 2.27fF
C215 a_48518_4733# gnd 11.63fF
C216 a_44568_4052# gnd 3.33fF
C217 a_45616_4727# gnd 3.64fF
C218 a_43739_4415# gnd 3.17fF
C219 a_44568_4731# gnd 2.80fF
C220 a_40543_4000# gnd 3.33fF
C221 a_41587_4852# gnd 2.33fF
C222 a_39049_4855# gnd 3.27fF
C223 a_43739_4810# gnd 2.27fF
C224 a_32721_444# gnd 10.85fF
C225 a_33817_4044# gnd 3.33fF
C226 a_34865_4719# gnd 3.64fF
C227 a_32988_4407# gnd 3.17fF
C228 a_33817_4723# gnd 2.80fF
C229 a_29835_4006# gnd 3.33fF
C230 a_30879_4858# gnd 2.33fF
C231 a_28341_4861# gnd 3.27fF
C232 a_32988_4802# gnd 2.27fF
C233 a_27059_4731# gnd 11.63fF
C234 a_23109_4050# gnd 3.33fF
C235 a_24157_4725# gnd 3.64fF
C236 a_22280_4413# gnd 3.17fF
C237 a_23109_4729# gnd 2.80fF
C238 a_18870_4002# gnd 3.33fF
C239 a_19914_4854# gnd 2.33fF
C240 a_17376_4857# gnd 3.27fF
C241 a_22280_4808# gnd 2.27fF
C242 a_11048_446# gnd 10.85fF
C243 a_12144_4046# gnd 3.33fF
C244 a_13192_4721# gnd 3.64fF
C245 a_11315_4409# gnd 3.17fF
C246 a_12144_4725# gnd 2.80fF
C247 a_8162_4008# gnd 3.33fF
C248 a_9206_4860# gnd 2.33fF
C249 a_6668_4863# gnd 3.27fF
C250 a_11315_4804# gnd 2.27fF
C251 a_5386_4733# gnd 11.63fF
C252 a_1436_4052# gnd 3.33fF
C253 a_2484_4727# gnd 3.64fF
C254 d5 gnd 178.70fF
C255 a_607_4415# gnd 3.17fF
C256 a_1436_4731# gnd 2.80fF
C257 a_607_4810# gnd 2.27fF
C258 a_84723_4675# gnd 3.52fF
C259 a_74015_4681# gnd 3.52fF
C260 a_63050_4677# gnd 3.52fF
C261 a_52342_4683# gnd 3.52fF
C262 a_41591_4675# gnd 3.52fF
C263 a_30883_4681# gnd 3.52fF
C264 a_84718_5693# gnd 2.27fF
C265 a_83670_5697# gnd 2.80fF
C266 a_79387_5561# gnd 3.19fF
C267 a_76120_5058# gnd 3.52fF
C268 a_74010_5699# gnd 2.27fF
C269 a_72962_5703# gnd 2.80fF
C270 a_68679_5567# gnd 3.19fF
C271 a_19918_4677# gnd 3.52fF
C272 a_9210_4683# gnd 3.52fF
C273 a_76119_5672# gnd 2.33fF
C274 a_65412_5064# gnd 3.52fF
C275 a_63045_5695# gnd 2.27fF
C276 a_61997_5699# gnd 2.80fF
C277 a_57714_5563# gnd 3.19fF
C278 a_65411_5678# gnd 2.33fF
C279 a_54447_5060# gnd 3.52fF
C280 a_52337_5701# gnd 2.27fF
C281 a_51289_5705# gnd 2.80fF
C282 a_47006_5569# gnd 3.19fF
C283 a_54446_5674# gnd 2.33fF
C284 a_43739_5066# gnd 3.52fF
C285 a_41586_5693# gnd 2.27fF
C286 a_40538_5697# gnd 2.80fF
C287 a_36255_5561# gnd 3.19fF
C288 a_32988_5058# gnd 3.52fF
C289 a_30878_5699# gnd 2.27fF
C290 a_29830_5703# gnd 2.80fF
C291 a_25547_5567# gnd 3.19fF
C292 a_43738_5680# gnd 2.33fF
C293 a_32987_5672# gnd 2.33fF
C294 a_22280_5064# gnd 3.52fF
C295 a_19913_5695# gnd 2.27fF
C296 a_18865_5699# gnd 2.80fF
C297 a_14582_5563# gnd 3.19fF
C298 a_22279_5678# gnd 2.33fF
C299 a_11315_5060# gnd 3.52fF
C300 a_9205_5701# gnd 2.27fF
C301 a_8157_5705# gnd 2.80fF
C302 a_3874_5569# gnd 3.19fF
C303 a_11314_5674# gnd 2.33fF
C304 a_607_5066# gnd 3.52fF
C305 a_606_5680# gnd 2.33fF
C306 a_84722_5516# gnd 3.17fF
C307 a_74014_5522# gnd 3.17fF
C308 a_63049_5518# gnd 3.17fF
C309 a_52341_5524# gnd 3.17fF
C310 a_41590_5516# gnd 3.17fF
C311 a_30882_5522# gnd 3.17fF
C312 a_83674_5520# gnd 3.33fF
C313 a_84718_6372# gnd 2.33fF
C314 a_82185_4678# gnd 3.19fF
C315 a_82223_6377# gnd 3.65fF
C316 a_76948_5564# gnd 3.33fF
C317 a_19917_5518# gnd 3.17fF
C318 a_9209_5524# gnd 3.17fF
C319 a_76119_5927# gnd 3.17fF
C320 a_76948_6243# gnd 2.80fF
C321 a_72966_5526# gnd 3.33fF
C322 a_74010_6378# gnd 2.33fF
C323 a_71477_4684# gnd 3.19fF
C324 a_71515_6383# gnd 3.65fF
C325 a_66240_5570# gnd 3.33fF
C326 a_76119_6322# gnd 2.27fF
C327 a_65411_5933# gnd 3.17fF
C328 a_66240_6249# gnd 2.80fF
C329 a_62001_5522# gnd 3.33fF
C330 a_63045_6374# gnd 2.33fF
C331 a_60512_4680# gnd 3.19fF
C332 a_60550_6379# gnd 3.65fF
C333 a_55275_5566# gnd 3.33fF
C334 a_65411_6328# gnd 2.27fF
C335 a_54446_5929# gnd 3.17fF
C336 a_55275_6245# gnd 2.80fF
C337 a_51293_5528# gnd 3.33fF
C338 a_52337_6380# gnd 2.33fF
C339 a_49804_4686# gnd 3.19fF
C340 a_49842_6385# gnd 3.65fF
C341 a_44567_5572# gnd 3.33fF
C342 a_54446_6324# gnd 2.27fF
C343 a_43738_5935# gnd 3.17fF
C344 a_44567_6251# gnd 2.80fF
C345 a_40542_5520# gnd 3.33fF
C346 a_41586_6372# gnd 2.33fF
C347 a_39053_4678# gnd 3.19fF
C348 a_39091_6377# gnd 3.65fF
C349 a_33816_5564# gnd 3.33fF
C350 a_43738_6330# gnd 2.27fF
C351 a_32987_5927# gnd 3.17fF
C352 a_33816_6243# gnd 2.80fF
C353 a_29834_5526# gnd 3.33fF
C354 a_30878_6378# gnd 2.33fF
C355 a_28345_4684# gnd 3.19fF
C356 a_28383_6383# gnd 3.65fF
C357 a_23108_5570# gnd 3.33fF
C358 a_32987_6322# gnd 2.27fF
C359 a_22279_5933# gnd 3.17fF
C360 a_23108_6249# gnd 2.80fF
C361 a_18869_5522# gnd 3.33fF
C362 a_19913_6374# gnd 2.33fF
C363 a_17380_4680# gnd 3.19fF
C364 a_17418_6379# gnd 3.65fF
C365 a_12143_5566# gnd 3.33fF
C366 a_22279_6328# gnd 2.27fF
C367 a_11314_5929# gnd 3.17fF
C368 a_12143_6245# gnd 2.80fF
C369 a_8161_5528# gnd 3.33fF
C370 a_9205_6380# gnd 2.33fF
C371 a_6672_4686# gnd 3.19fF
C372 a_6710_6385# gnd 3.65fF
C373 a_1435_5572# gnd 3.33fF
C374 a_11314_6324# gnd 2.27fF
C375 a_606_5935# gnd 3.17fF
C376 a_1435_6251# gnd 2.80fF
C377 a_606_6330# gnd 2.27fF
C378 a_84722_6195# gnd 3.43fF
C379 a_74014_6201# gnd 3.43fF
C380 a_63049_6197# gnd 3.43fF
C381 a_52341_6203# gnd 3.43fF
C382 a_41590_6195# gnd 3.43fF
C383 a_30882_6201# gnd 3.43fF
C384 a_84718_7140# gnd 2.27fF
C385 a_82227_6200# gnd 3.20fF
C386 a_83670_7144# gnd 2.80fF
C387 a_77996_6239# gnd 3.43fF
C388 a_79392_5680# gnd 3.27fF
C389 a_76119_6578# gnd 3.43fF
C390 a_74010_7146# gnd 2.27fF
C391 a_71519_6206# gnd 3.20fF
C392 a_72962_7150# gnd 2.80fF
C393 a_67288_6245# gnd 3.43fF
C394 a_68684_5686# gnd 3.27fF
C395 a_19917_6197# gnd 3.43fF
C396 a_9209_6203# gnd 3.43fF
C397 a_76119_7119# gnd 2.33fF
C398 a_65411_6584# gnd 3.43fF
C399 a_63045_7142# gnd 2.27fF
C400 a_60554_6202# gnd 3.20fF
C401 a_61997_7146# gnd 2.80fF
C402 a_56323_6241# gnd 3.43fF
C403 a_57719_5682# gnd 3.27fF
C404 a_65411_7125# gnd 2.33fF
C405 a_54446_6580# gnd 3.43fF
C406 a_52337_7148# gnd 2.27fF
C407 a_49846_6208# gnd 3.20fF
C408 a_51289_7152# gnd 2.80fF
C409 a_45615_6247# gnd 3.43fF
C410 a_47011_5688# gnd 3.27fF
C411 a_54446_7121# gnd 2.33fF
C412 a_43738_6586# gnd 3.43fF
C413 a_41586_7140# gnd 2.27fF
C414 a_39095_6200# gnd 3.20fF
C415 a_40538_7144# gnd 2.80fF
C416 a_34864_6239# gnd 3.43fF
C417 a_36260_5680# gnd 3.27fF
C418 a_32987_6578# gnd 3.43fF
C419 a_30878_7146# gnd 2.27fF
C420 a_28387_6206# gnd 3.20fF
C421 a_29830_7150# gnd 2.80fF
C422 a_24156_6245# gnd 3.43fF
C423 a_25552_5686# gnd 3.27fF
C424 a_43738_7127# gnd 2.33fF
C425 a_32987_7119# gnd 2.33fF
C426 a_22279_6584# gnd 3.43fF
C427 a_19913_7142# gnd 2.27fF
C428 a_17422_6202# gnd 3.20fF
C429 a_18865_7146# gnd 2.80fF
C430 a_13191_6241# gnd 3.43fF
C431 a_14587_5682# gnd 3.27fF
C432 a_22279_7125# gnd 2.33fF
C433 a_11314_6580# gnd 3.43fF
C434 a_9205_7148# gnd 2.27fF
C435 a_6714_6208# gnd 3.20fF
C436 a_8157_7152# gnd 2.80fF
C437 a_2483_6247# gnd 3.43fF
C438 a_3879_5688# gnd 3.27fF
C439 a_11314_7121# gnd 2.33fF
C440 a_606_6586# gnd 3.43fF
C441 a_606_7127# gnd 2.33fF
C442 a_84722_6963# gnd 3.17fF
C443 a_74014_6969# gnd 3.17fF
C444 a_63049_6965# gnd 3.17fF
C445 a_52341_6971# gnd 3.17fF
C446 a_41590_6963# gnd 3.17fF
C447 a_30882_6969# gnd 3.17fF
C448 a_83674_6967# gnd 3.33fF
C449 a_84718_7819# gnd 2.33fF
C450 a_80800_4725# gnd 4.30fF
C451 a_81115_7828# gnd 7.03fF
C452 a_76948_7011# gnd 3.33fF
C453 a_77996_7686# gnd 4.35fF
C454 a_19917_6965# gnd 3.17fF
C455 a_9209_6971# gnd 3.17fF
C456 a_76119_7374# gnd 3.17fF
C457 a_76948_7690# gnd 2.80fF
C458 a_72966_6973# gnd 3.33fF
C459 a_74010_7825# gnd 2.33fF
C460 a_70092_4731# gnd 4.30fF
C461 a_70407_7834# gnd 7.03fF
C462 a_66240_7017# gnd 3.33fF
C463 a_67288_7692# gnd 4.35fF
C464 a_76119_7769# gnd 2.27fF
C465 a_65411_7380# gnd 3.17fF
C466 a_66240_7696# gnd 2.80fF
C467 a_62001_6969# gnd 3.33fF
C468 a_63045_7821# gnd 2.33fF
C469 a_59127_4727# gnd 4.30fF
C470 a_59442_7830# gnd 7.03fF
C471 a_55275_7013# gnd 3.33fF
C472 a_56323_7688# gnd 4.35fF
C473 a_65411_7775# gnd 2.27fF
C474 a_54446_7376# gnd 3.17fF
C475 a_55275_7692# gnd 2.80fF
C476 a_51293_6975# gnd 3.33fF
C477 a_52337_7827# gnd 2.33fF
C478 a_48419_4733# gnd 4.30fF
C479 a_48734_7836# gnd 7.03fF
C480 a_44567_7019# gnd 3.33fF
C481 a_45615_7694# gnd 4.35fF
C482 a_54446_7771# gnd 2.27fF
C483 a_43738_7382# gnd 3.17fF
C484 a_44567_7698# gnd 2.80fF
C485 a_40542_6967# gnd 3.33fF
C486 a_41586_7819# gnd 2.33fF
C487 a_37668_4725# gnd 4.30fF
C488 a_37983_7828# gnd 7.03fF
C489 a_33816_7011# gnd 3.33fF
C490 a_34864_7686# gnd 4.35fF
C491 a_43738_7777# gnd 2.27fF
C492 a_32987_7374# gnd 3.17fF
C493 a_33816_7690# gnd 2.80fF
C494 a_29834_6973# gnd 3.33fF
C495 a_30878_7825# gnd 2.33fF
C496 a_26960_4731# gnd 4.30fF
C497 a_27275_7834# gnd 7.03fF
C498 a_23108_7017# gnd 3.33fF
C499 a_24156_7692# gnd 4.35fF
C500 a_32987_7769# gnd 2.27fF
C501 a_22279_7380# gnd 3.17fF
C502 a_23108_7696# gnd 2.80fF
C503 a_18869_6969# gnd 3.33fF
C504 a_19913_7821# gnd 2.33fF
C505 a_15995_4727# gnd 4.30fF
C506 a_16310_7830# gnd 7.03fF
C507 a_12143_7013# gnd 3.33fF
C508 a_13191_7688# gnd 4.35fF
C509 a_22279_7775# gnd 2.27fF
C510 a_11314_7376# gnd 3.17fF
C511 a_12143_7692# gnd 2.80fF
C512 a_8161_6975# gnd 3.33fF
C513 a_9205_7827# gnd 2.33fF
C514 a_5287_4733# gnd 4.30fF
C515 a_5602_7836# gnd 7.03fF
C516 a_1435_7019# gnd 3.33fF
C517 a_2483_7694# gnd 4.35fF
C518 a_11314_7771# gnd 2.27fF
C519 a_606_7382# gnd 3.17fF
C520 a_1435_7698# gnd 2.80fF
C521 a_606_7777# gnd 2.27fF
C522 a_84722_7642# gnd 3.62fF
C523 a_74014_7648# gnd 3.62fF
C524 a_63049_7644# gnd 3.62fF
C525 a_52341_7650# gnd 3.62fF
C526 a_41590_7642# gnd 3.62fF
C527 a_30882_7648# gnd 3.62fF
C528 a_84721_8734# gnd 2.27fF
C529 a_83673_8738# gnd 2.80fF
C530 a_79486_5561# gnd 4.97fF
C531 a_80554_8596# gnd 4.72fF
C532 a_76119_8025# gnd 3.62fF
C533 a_74013_8740# gnd 2.27fF
C534 a_72965_8744# gnd 2.80fF
C535 a_68778_5567# gnd 4.97fF
C536 a_69846_8602# gnd 4.72fF
C537 a_19917_7644# gnd 3.62fF
C538 a_9209_7650# gnd 3.62fF
C539 a_76122_8713# gnd 2.33fF
C540 a_65411_8031# gnd 3.62fF
C541 a_63048_8736# gnd 2.27fF
C542 a_62000_8740# gnd 2.80fF
C543 a_57813_5563# gnd 4.97fF
C544 a_58881_8598# gnd 4.72fF
C545 a_65414_8719# gnd 2.33fF
C546 a_54446_8027# gnd 3.62fF
C547 a_52340_8742# gnd 2.27fF
C548 a_51292_8746# gnd 2.80fF
C549 a_47105_5569# gnd 4.97fF
C550 a_48173_8604# gnd 4.72fF
C551 a_54449_8715# gnd 2.33fF
C552 a_43738_8033# gnd 3.62fF
C553 a_41589_8734# gnd 2.27fF
C554 a_40541_8738# gnd 2.80fF
C555 a_36354_5561# gnd 4.97fF
C556 a_37422_8596# gnd 4.72fF
C557 a_32987_8025# gnd 3.62fF
C558 a_30881_8740# gnd 2.27fF
C559 a_29833_8744# gnd 2.80fF
C560 a_25646_5567# gnd 4.97fF
C561 a_26714_8602# gnd 4.72fF
C562 a_43741_8721# gnd 2.33fF
C563 a_32990_8713# gnd 2.33fF
C564 a_22279_8031# gnd 3.62fF
C565 a_19916_8736# gnd 2.27fF
C566 a_18868_8740# gnd 2.80fF
C567 a_14681_5563# gnd 4.97fF
C568 a_15749_8598# gnd 4.72fF
C569 a_22282_8719# gnd 2.33fF
C570 a_11314_8027# gnd 3.62fF
C571 a_9208_8742# gnd 2.27fF
C572 a_8160_8746# gnd 2.80fF
C573 a_3973_5569# gnd 4.97fF
C574 a_5041_8604# gnd 4.72fF
C575 a_11317_8715# gnd 2.33fF
C576 d4 gnd 224.03fF
C577 a_606_8033# gnd 3.62fF
C578 a_609_8721# gnd 2.33fF
C579 a_84725_8557# gnd 3.17fF
C580 a_74017_8563# gnd 3.17fF
C581 a_63052_8559# gnd 3.17fF
C582 a_52344_8565# gnd 3.17fF
C583 a_41593_8557# gnd 3.17fF
C584 a_30885_8563# gnd 3.17fF
C585 a_83677_8561# gnd 3.33fF
C586 a_84721_9413# gnd 2.33fF
C587 a_82226_9418# gnd 4.35fF
C588 a_76951_8605# gnd 3.33fF
C589 a_19920_8559# gnd 3.17fF
C590 a_9212_8565# gnd 3.17fF
C591 a_76122_8968# gnd 3.17fF
C592 a_76951_9284# gnd 2.80fF
C593 a_72969_8567# gnd 3.33fF
C594 a_74013_9419# gnd 2.33fF
C595 a_71518_9424# gnd 4.35fF
C596 a_66243_8611# gnd 3.33fF
C597 a_76122_9363# gnd 2.27fF
C598 a_65414_8974# gnd 3.17fF
C599 a_66243_9290# gnd 2.80fF
C600 a_62004_8563# gnd 3.33fF
C601 a_63048_9415# gnd 2.33fF
C602 a_60553_9420# gnd 4.35fF
C603 a_55278_8607# gnd 3.33fF
C604 a_65414_9369# gnd 2.27fF
C605 a_54449_8970# gnd 3.17fF
C606 a_55278_9286# gnd 2.80fF
C607 a_51296_8569# gnd 3.33fF
C608 a_52340_9421# gnd 2.33fF
C609 a_49845_9426# gnd 4.35fF
C610 a_44570_8613# gnd 3.33fF
C611 a_54449_9365# gnd 2.27fF
C612 a_43741_8976# gnd 3.17fF
C613 a_44570_9292# gnd 2.80fF
C614 a_40545_8561# gnd 3.33fF
C615 a_41589_9413# gnd 2.33fF
C616 a_39094_9418# gnd 4.35fF
C617 a_33819_8605# gnd 3.33fF
C618 a_43741_9371# gnd 2.27fF
C619 a_32990_8968# gnd 3.17fF
C620 a_33819_9284# gnd 2.80fF
C621 a_29837_8567# gnd 3.33fF
C622 a_30881_9419# gnd 2.33fF
C623 a_28386_9424# gnd 4.35fF
C624 a_23111_8611# gnd 3.33fF
C625 a_32990_9363# gnd 2.27fF
C626 a_22282_8974# gnd 3.17fF
C627 a_23111_9290# gnd 2.80fF
C628 a_18872_8563# gnd 3.33fF
C629 a_19916_9415# gnd 2.33fF
C630 a_17421_9420# gnd 4.35fF
C631 a_12146_8607# gnd 3.33fF
C632 a_22282_9369# gnd 2.27fF
C633 a_11317_8970# gnd 3.17fF
C634 a_12146_9286# gnd 2.80fF
C635 a_8164_8569# gnd 3.33fF
C636 a_9208_9421# gnd 2.33fF
C637 a_6713_9426# gnd 4.35fF
C638 a_1438_8613# gnd 3.33fF
C639 a_11317_9365# gnd 2.27fF
C640 a_609_8976# gnd 3.17fF
C641 a_1438_9292# gnd 2.80fF
C642 a_609_9371# gnd 2.27fF
C643 a_84725_9236# gnd 3.43fF
C644 a_74017_9242# gnd 3.43fF
C645 a_63052_9238# gnd 3.43fF
C646 a_52344_9244# gnd 3.43fF
C647 a_41593_9236# gnd 3.43fF
C648 a_30885_9242# gnd 3.43fF
C649 a_84721_10181# gnd 2.27fF
C650 a_82230_9241# gnd 3.43fF
C651 a_83673_10185# gnd 2.80fF
C652 a_77999_9280# gnd 3.20fF
C653 a_76122_9619# gnd 3.43fF
C654 a_74013_10187# gnd 2.27fF
C655 a_71522_9247# gnd 3.43fF
C656 a_72965_10191# gnd 2.80fF
C657 a_67291_9286# gnd 3.20fF
C658 a_19920_9238# gnd 3.43fF
C659 a_9212_9244# gnd 3.43fF
C660 a_76122_10160# gnd 2.33fF
C661 a_65414_9625# gnd 3.43fF
C662 a_63048_10183# gnd 2.27fF
C663 a_60557_9243# gnd 3.43fF
C664 a_62000_10187# gnd 2.80fF
C665 a_56326_9282# gnd 3.20fF
C666 a_65414_10166# gnd 2.33fF
C667 a_54449_9621# gnd 3.43fF
C668 a_52340_10189# gnd 2.27fF
C669 a_49849_9249# gnd 3.43fF
C670 a_51292_10193# gnd 2.80fF
C671 a_45618_9288# gnd 3.20fF
C672 a_54449_10162# gnd 2.33fF
C673 a_43741_9627# gnd 3.43fF
C674 a_41589_10181# gnd 2.27fF
C675 a_39098_9241# gnd 3.43fF
C676 a_40541_10185# gnd 2.80fF
C677 a_34867_9280# gnd 3.20fF
C678 a_32990_9619# gnd 3.43fF
C679 a_30881_10187# gnd 2.27fF
C680 a_28390_9247# gnd 3.43fF
C681 a_29833_10191# gnd 2.80fF
C682 a_24159_9286# gnd 3.20fF
C683 a_43741_10168# gnd 2.33fF
C684 a_32990_10160# gnd 2.33fF
C685 a_22282_9625# gnd 3.43fF
C686 a_19916_10183# gnd 2.27fF
C687 a_17425_9243# gnd 3.43fF
C688 a_18868_10187# gnd 2.80fF
C689 a_13194_9282# gnd 3.20fF
C690 a_22282_10166# gnd 2.33fF
C691 a_11317_9621# gnd 3.43fF
C692 a_9208_10189# gnd 2.27fF
C693 a_6717_9249# gnd 3.43fF
C694 a_8160_10193# gnd 2.80fF
C695 a_2486_9288# gnd 3.20fF
C696 a_11317_10162# gnd 2.33fF
C697 a_609_9627# gnd 3.43fF
C698 a_609_10168# gnd 2.33fF
C699 a_84725_10004# gnd 3.17fF
C700 a_74017_10010# gnd 3.17fF
C701 a_63052_10006# gnd 3.17fF
C702 a_52344_10012# gnd 3.17fF
C703 a_41593_10004# gnd 3.17fF
C704 a_30885_10010# gnd 3.17fF
C705 a_83677_10008# gnd 3.33fF
C706 a_84721_10860# gnd 2.33fF
C707 a_81119_7651# gnd 4.90fF
C708 a_82183_10863# gnd 3.27fF
C709 a_76951_10052# gnd 3.33fF
C710 a_77999_10727# gnd 3.65fF
C711 a_19920_10006# gnd 3.17fF
C712 a_9212_10012# gnd 3.17fF
C713 a_76122_10415# gnd 3.17fF
C714 a_76951_10731# gnd 2.80fF
C715 a_72969_10014# gnd 3.33fF
C716 a_74013_10866# gnd 2.33fF
C717 a_70411_7657# gnd 4.90fF
C718 a_71475_10869# gnd 3.27fF
C719 a_66243_10058# gnd 3.33fF
C720 a_67291_10733# gnd 3.65fF
C721 a_76122_10810# gnd 2.27fF
C722 a_65414_10421# gnd 3.17fF
C723 a_66243_10737# gnd 2.80fF
C724 a_62004_10010# gnd 3.33fF
C725 a_63048_10862# gnd 2.33fF
C726 a_59446_7653# gnd 4.90fF
C727 a_60510_10865# gnd 3.27fF
C728 a_55278_10054# gnd 3.33fF
C729 a_56326_10729# gnd 3.65fF
C730 a_65414_10816# gnd 2.27fF
C731 a_54449_10417# gnd 3.17fF
C732 a_55278_10733# gnd 2.80fF
C733 a_51296_10016# gnd 3.33fF
C734 a_52340_10868# gnd 2.33fF
C735 a_48738_7659# gnd 4.90fF
C736 a_49802_10871# gnd 3.27fF
C737 a_44570_10060# gnd 3.33fF
C738 a_45618_10735# gnd 3.65fF
C739 a_54449_10812# gnd 2.27fF
C740 a_43741_10423# gnd 3.17fF
C741 a_44570_10739# gnd 2.80fF
C742 a_40545_10008# gnd 3.33fF
C743 a_41589_10860# gnd 2.33fF
C744 a_37987_7651# gnd 4.90fF
C745 a_39051_10863# gnd 3.27fF
C746 a_33819_10052# gnd 3.33fF
C747 a_34867_10727# gnd 3.65fF
C748 a_43741_10818# gnd 2.27fF
C749 a_32990_10415# gnd 3.17fF
C750 a_33819_10731# gnd 2.80fF
C751 a_29837_10014# gnd 3.33fF
C752 a_30881_10866# gnd 2.33fF
C753 a_27279_7657# gnd 4.90fF
C754 a_28343_10869# gnd 3.27fF
C755 a_23111_10058# gnd 3.33fF
C756 a_24159_10733# gnd 3.65fF
C757 a_32990_10810# gnd 2.27fF
C758 a_22282_10421# gnd 3.17fF
C759 a_23111_10737# gnd 2.80fF
C760 a_18872_10010# gnd 3.33fF
C761 a_19916_10862# gnd 2.33fF
C762 a_16314_7653# gnd 4.90fF
C763 a_17378_10865# gnd 3.27fF
C764 a_12146_10054# gnd 3.33fF
C765 a_13194_10729# gnd 3.65fF
C766 a_22282_10816# gnd 2.27fF
C767 a_11317_10417# gnd 3.17fF
C768 a_12146_10733# gnd 2.80fF
C769 a_8164_10016# gnd 3.33fF
C770 a_9208_10868# gnd 2.33fF
C771 a_5606_7659# gnd 4.90fF
C772 a_6670_10871# gnd 3.27fF
C773 a_1438_10060# gnd 3.33fF
C774 a_2486_10735# gnd 3.65fF
C775 a_11317_10812# gnd 2.27fF
C776 a_609_10423# gnd 3.17fF
C777 a_1438_10739# gnd 2.80fF
C778 a_609_10818# gnd 2.27fF
C779 a_84725_10683# gnd 3.52fF
C780 a_74017_10689# gnd 3.52fF
C781 a_63052_10685# gnd 3.52fF
C782 a_52344_10691# gnd 3.52fF
C783 a_41593_10683# gnd 3.52fF
C784 a_30885_10689# gnd 3.52fF
C785 a_84720_11701# gnd 2.27fF
C786 a_83672_11705# gnd 2.80fF
C787 a_79389_11569# gnd 3.19fF
C788 a_79488_11569# gnd 7.02fF
C789 a_76122_11066# gnd 3.52fF
C790 a_74012_11707# gnd 2.27fF
C791 a_72964_11711# gnd 2.80fF
C792 a_68681_11575# gnd 3.19fF
C793 a_68780_11575# gnd 7.02fF
C794 a_19920_10685# gnd 3.52fF
C795 a_9212_10691# gnd 3.52fF
C796 a_76121_11680# gnd 2.33fF
C797 a_65414_11072# gnd 3.52fF
C798 a_63047_11703# gnd 2.27fF
C799 a_61999_11707# gnd 2.80fF
C800 a_57716_11571# gnd 3.19fF
C801 a_57815_11571# gnd 7.02fF
C802 a_65413_11686# gnd 2.33fF
C803 a_54449_11068# gnd 3.52fF
C804 a_52339_11709# gnd 2.27fF
C805 a_51291_11713# gnd 2.80fF
C806 a_47008_11577# gnd 3.19fF
C807 a_47107_11577# gnd 7.02fF
C808 a_54448_11682# gnd 2.33fF
C809 a_43741_11074# gnd 3.52fF
C810 a_41588_11701# gnd 2.27fF
C811 a_40540_11705# gnd 2.80fF
C812 a_36257_11569# gnd 3.19fF
C813 a_36356_11569# gnd 7.02fF
C814 a_32990_11066# gnd 3.52fF
C815 a_30880_11707# gnd 2.27fF
C816 a_29832_11711# gnd 2.80fF
C817 a_25549_11575# gnd 3.19fF
C818 a_25648_11575# gnd 7.02fF
C819 a_43740_11688# gnd 2.33fF
C820 a_32989_11680# gnd 2.33fF
C821 a_22282_11072# gnd 3.52fF
C822 a_19915_11703# gnd 2.27fF
C823 a_18867_11707# gnd 2.80fF
C824 a_14584_11571# gnd 3.19fF
C825 a_14683_11571# gnd 7.02fF
C826 a_22281_11686# gnd 2.33fF
C827 a_11317_11068# gnd 3.52fF
C828 a_9207_11709# gnd 2.27fF
C829 a_8159_11713# gnd 2.80fF
C830 a_3876_11577# gnd 3.19fF
C831 a_3975_11577# gnd 7.02fF
C832 a_11316_11682# gnd 2.33fF
C833 d3 gnd 423.95fF
C834 a_609_11074# gnd 3.52fF
C835 a_608_11688# gnd 2.33fF
C836 a_84724_11524# gnd 3.17fF
C837 a_74016_11530# gnd 3.17fF
C838 a_63051_11526# gnd 3.17fF
C839 a_52343_11532# gnd 3.17fF
C840 a_41592_11524# gnd 3.17fF
C841 a_30884_11530# gnd 3.17fF
C842 a_83676_11528# gnd 3.33fF
C843 a_84720_12380# gnd 2.33fF
C844 a_82187_10686# gnd 3.19fF
C845 a_82225_12385# gnd 3.73fF
C846 a_76950_11572# gnd 3.33fF
C847 a_19919_11526# gnd 3.17fF
C848 a_9211_11532# gnd 3.17fF
C849 a_76121_11935# gnd 3.17fF
C850 a_76950_12251# gnd 2.80fF
C851 a_72968_11534# gnd 3.33fF
C852 a_74012_12386# gnd 2.33fF
C853 a_71479_10692# gnd 3.19fF
C854 a_71517_12391# gnd 3.73fF
C855 a_66242_11578# gnd 3.33fF
C856 a_76121_12330# gnd 2.27fF
C857 a_65413_11941# gnd 3.17fF
C858 a_66242_12257# gnd 2.80fF
C859 a_62003_11530# gnd 3.33fF
C860 a_63047_12382# gnd 2.33fF
C861 a_60514_10688# gnd 3.19fF
C862 a_60552_12387# gnd 3.73fF
C863 a_55277_11574# gnd 3.33fF
C864 a_65413_12336# gnd 2.27fF
C865 a_54448_11937# gnd 3.17fF
C866 a_55277_12253# gnd 2.80fF
C867 a_51295_11536# gnd 3.33fF
C868 a_52339_12388# gnd 2.33fF
C869 a_49806_10694# gnd 3.19fF
C870 a_49844_12393# gnd 3.73fF
C871 a_44569_11580# gnd 3.33fF
C872 a_54448_12332# gnd 2.27fF
C873 a_43740_11943# gnd 3.17fF
C874 a_44569_12259# gnd 2.80fF
C875 a_40544_11528# gnd 3.33fF
C876 a_41588_12380# gnd 2.33fF
C877 a_39055_10686# gnd 3.19fF
C878 a_39093_12385# gnd 3.73fF
C879 a_33818_11572# gnd 3.33fF
C880 a_43740_12338# gnd 2.27fF
C881 a_32989_11935# gnd 3.17fF
C882 a_33818_12251# gnd 2.80fF
C883 a_29836_11534# gnd 3.33fF
C884 a_30880_12386# gnd 2.33fF
C885 a_28347_10692# gnd 3.19fF
C886 a_28385_12391# gnd 3.73fF
C887 a_23110_11578# gnd 3.33fF
C888 a_32989_12330# gnd 2.27fF
C889 a_22281_11941# gnd 3.17fF
C890 a_23110_12257# gnd 2.80fF
C891 a_18871_11530# gnd 3.33fF
C892 a_19915_12382# gnd 2.33fF
C893 a_17382_10688# gnd 3.19fF
C894 a_17420_12387# gnd 3.73fF
C895 a_12145_11574# gnd 3.33fF
C896 a_22281_12336# gnd 2.27fF
C897 a_11316_11937# gnd 3.17fF
C898 a_12145_12253# gnd 2.80fF
C899 a_8163_11536# gnd 3.33fF
C900 a_9207_12388# gnd 2.33fF
C901 a_6674_10694# gnd 3.19fF
C902 a_6712_12393# gnd 3.73fF
C903 a_1437_11580# gnd 3.33fF
C904 a_11316_12332# gnd 2.27fF
C905 a_608_11943# gnd 3.17fF
C906 a_1437_12259# gnd 2.80fF
C907 a_608_12338# gnd 2.27fF
C908 a_84724_12203# gnd 3.43fF
C909 a_74016_12209# gnd 3.43fF
C910 a_63051_12205# gnd 3.43fF
C911 a_52343_12211# gnd 3.43fF
C912 a_41592_12203# gnd 3.43fF
C913 a_30884_12209# gnd 3.43fF
C914 a_84720_13148# gnd 2.27fF
C915 a_82229_12208# gnd 3.35fF
C916 a_83672_13152# gnd 2.80fF
C917 a_77998_12247# gnd 3.43fF
C918 a_79394_11688# gnd 3.27fF
C919 a_76121_12586# gnd 3.43fF
C920 a_74012_13154# gnd 2.27fF
C921 a_71521_12214# gnd 3.35fF
C922 a_72964_13158# gnd 2.80fF
C923 a_67290_12253# gnd 3.43fF
C924 a_68686_11694# gnd 3.27fF
C925 a_19919_12205# gnd 3.43fF
C926 a_9211_12211# gnd 3.43fF
C927 a_76121_13127# gnd 2.33fF
C928 a_65413_12592# gnd 3.43fF
C929 a_63047_13150# gnd 2.27fF
C930 a_60556_12210# gnd 3.35fF
C931 a_61999_13154# gnd 2.80fF
C932 a_56325_12249# gnd 3.43fF
C933 a_57721_11690# gnd 3.27fF
C934 a_65413_13133# gnd 2.33fF
C935 a_54448_12588# gnd 3.43fF
C936 a_52339_13156# gnd 2.27fF
C937 a_49848_12216# gnd 3.35fF
C938 a_51291_13160# gnd 2.80fF
C939 a_45617_12255# gnd 3.43fF
C940 a_47013_11696# gnd 3.27fF
C941 a_54448_13129# gnd 2.33fF
C942 a_43740_12594# gnd 3.43fF
C943 a_41588_13148# gnd 2.27fF
C944 a_39097_12208# gnd 3.35fF
C945 a_40540_13152# gnd 2.80fF
C946 a_34866_12247# gnd 3.43fF
C947 a_36262_11688# gnd 3.27fF
C948 a_32989_12586# gnd 3.43fF
C949 a_30880_13154# gnd 2.27fF
C950 a_28389_12214# gnd 3.35fF
C951 a_29832_13158# gnd 2.80fF
C952 a_24158_12253# gnd 3.43fF
C953 a_25554_11694# gnd 3.27fF
C954 a_43740_13135# gnd 2.33fF
C955 a_32989_13127# gnd 2.33fF
C956 a_22281_12592# gnd 3.43fF
C957 a_19915_13150# gnd 2.27fF
C958 a_17424_12210# gnd 3.35fF
C959 a_18867_13154# gnd 2.80fF
C960 a_13193_12249# gnd 3.43fF
C961 a_14589_11690# gnd 3.27fF
C962 a_22281_13133# gnd 2.33fF
C963 a_11316_12588# gnd 3.43fF
C964 a_9207_13156# gnd 2.27fF
C965 a_6716_12216# gnd 3.35fF
C966 a_8159_13160# gnd 2.80fF
C967 a_2485_12255# gnd 3.43fF
C968 a_3881_11696# gnd 3.27fF
C969 a_11316_13129# gnd 2.33fF
C970 d2 gnd 428.42fF
C971 a_608_12594# gnd 3.43fF
C972 a_608_13135# gnd 2.33fF
C973 a_84724_12971# gnd 3.17fF
C974 a_74016_12977# gnd 3.17fF
C975 a_63051_12973# gnd 3.17fF
C976 a_52343_12979# gnd 3.17fF
C977 a_41592_12971# gnd 3.17fF
C978 a_30884_12977# gnd 3.17fF
C979 a_83676_12975# gnd 3.40fF
C980 a_84720_13827# gnd 2.73fF
C981 a_76950_13019# gnd 3.33fF
C982 a_77998_13694# gnd 4.35fF
C983 a_19919_12973# gnd 3.17fF
C984 a_9211_12979# gnd 3.17fF
C985 a_76121_13382# gnd 3.17fF
C986 a_76950_13698# gnd 2.80fF
C987 a_72968_12981# gnd 3.33fF
C988 a_74012_13833# gnd 2.33fF
C989 a_66242_13025# gnd 3.33fF
C990 a_67290_13700# gnd 4.35fF
C991 a_76121_13777# gnd 2.27fF
C992 a_65413_13388# gnd 3.17fF
C993 a_66242_13704# gnd 2.80fF
C994 a_62003_12977# gnd 3.33fF
C995 a_63047_13829# gnd 2.33fF
C996 a_55277_13021# gnd 3.33fF
C997 a_56325_13696# gnd 4.35fF
C998 a_65413_13783# gnd 2.27fF
C999 a_54448_13384# gnd 3.17fF
C1000 a_55277_13700# gnd 2.80fF
C1001 a_51295_12983# gnd 3.33fF
C1002 a_52339_13835# gnd 2.33fF
C1003 a_44569_13027# gnd 3.33fF
C1004 a_45617_13702# gnd 4.35fF
C1005 a_54448_13779# gnd 2.27fF
C1006 a_43740_13390# gnd 3.17fF
C1007 a_44569_13706# gnd 2.80fF
C1008 a_40544_12975# gnd 3.33fF
C1009 a_41588_13827# gnd 2.33fF
C1010 a_33818_13019# gnd 3.33fF
C1011 a_34866_13694# gnd 4.35fF
C1012 a_43740_13785# gnd 2.27fF
C1013 a_32989_13382# gnd 3.17fF
C1014 a_33818_13698# gnd 2.80fF
C1015 a_29836_12981# gnd 3.33fF
C1016 a_30880_13833# gnd 2.33fF
C1017 a_23110_13025# gnd 3.33fF
C1018 a_24158_13700# gnd 4.35fF
C1019 a_74016_13656# gnd 4.89fF
C1020 a_63051_13652# gnd 5.08fF
C1021 a_32989_13777# gnd 2.27fF
C1022 a_22281_13388# gnd 3.17fF
C1023 a_23110_13704# gnd 2.80fF
C1024 a_18871_12977# gnd 3.33fF
C1025 a_19915_13829# gnd 2.33fF
C1026 a_12145_13021# gnd 3.33fF
C1027 a_13193_13696# gnd 4.35fF
C1028 a_22281_13783# gnd 2.27fF
C1029 a_11316_13384# gnd 3.17fF
C1030 a_12145_13700# gnd 2.80fF
C1031 a_8163_12983# gnd 3.33fF
C1032 a_9207_13835# gnd 2.33fF
C1033 a_1437_13027# gnd 3.33fF
C1034 a_2485_13702# gnd 4.35fF
C1035 a_52343_13658# gnd 4.89fF
C1036 a_41592_13650# gnd 4.85fF
C1037 a_11316_13779# gnd 2.27fF
C1038 d1 gnd 498.39fF
C1039 a_608_13390# gnd 3.17fF
C1040 a_1437_13706# gnd 2.80fF
C1041 d0 gnd 616.94fF
C1042 a_608_13785# gnd 2.27fF
C1043 a_30884_13656# gnd 4.89fF
C1044 a_19919_13652# gnd 5.08fF
C1045 a_9211_13658# gnd 4.89fF
C1046 vdd gnd 2614.00fF
