* SPICE3 file created from 7bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 vdd d1 a_19017_11974# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1 a_502_10084# a_1122_10590# a_1330_10590# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X2 a_11831_9064# a_11618_9064# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X3 a_14574_4573# a_15434_7608# a_15642_7608# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X4 a_1120_4582# a_907_4582# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X5 a_6607_5218# a_6860_5205# a_6565_3696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X6 gnd d0 a_9356_1554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X7 a_6603_5395# a_8099_4525# a_8050_4715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X8 a_2170_12712# a_1957_12712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X9 a_18760_10717# a_19857_10523# a_19808_10713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X10 a_6561_3873# a_6818_3683# a_5495_6846# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X11 a_9104_11989# a_9357_11976# a_8052_12170# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X12 a_19813_8248# a_20066_8235# a_18765_7573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X13 a_11616_3056# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X14 gnd d0 a_20064_3674# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X15 a_11828_4576# a_11615_4576# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X16 a_11830_11263# a_11617_11263# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X17 a_17275_9698# a_17362_11207# a_17317_11220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X18 a_8054_5985# a_9147_6647# a_9102_6660# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X19 a_18758_6156# a_19855_5962# a_19806_6152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X20 a_11207_5334# a_11207_4939# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X21 a_8052_10723# a_9149_10529# a_9100_10719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X22 gnd d1 a_8310_7566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X23 a_12037_2288# a_12877_2284# a_13085_2284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X24 a_1122_11269# a_909_11269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X25 gnd a_9358_8241# a_9150_8241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X26 a_2379_8298# a_1958_8298# a_1331_8302# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X27 a_9102_6660# a_9098_6837# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X28 gnd d4 a_16460_6650# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X29 vdd d0 a_9356_1554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X30 a_14475_4573# a_14366_4573# a_14574_4573# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X31 a_6603_5395# a_8099_4525# a_8054_4538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X32 vdd d0 a_20063_5194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X33 a_2376_6704# a_1955_6704# a_1328_6029# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X34 a_18760_10717# a_19857_10523# a_19812_10536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X35 a_14111_3051# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X36 a_17317_11220# a_18809_11974# a_18764_11987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X37 a_1123_8302# a_910_8302# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X38 a_19809_8425# a_20066_8235# a_18765_7573# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X39 a_15434_7608# a_15221_7608# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X40 vdd d0 a_20064_3674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X41 a_14477_10581# a_14368_10581# a_14576_10581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X42 vdd d1 a_8310_7566# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X43 a_19811_1561# a_20064_1548# a_18759_1742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X44 vdd a_9358_8241# a_9150_8241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X45 a_3769_10587# a_3660_10587# a_3868_10587# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X46 vdd a_9357_10529# a_9149_10529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X47 a_11210_9427# a_11831_9743# a_12039_9743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X48 vdd d4 a_16460_6650# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X49 a_11208_3164# a_11208_2623# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X50 a_3774_10706# a_3404_12032# a_2378_11265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X51 vdd a_8309_11980# a_8101_11980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X52 gnd a_9356_1554# a_9148_1554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X53 a_499_6787# a_1120_6708# a_1328_6708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X54 a_907_5261# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X55 a_1955_5257# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X56 a_14477_10581# a_14113_9059# a_13087_8292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X57 a_13084_6698# a_12663_6698# a_12036_6023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X58 gnd a_20064_3674# a_19856_3674# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X59 a_11615_4576# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X60 a_14323_6018# a_14110_6018# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X61 a_1121_1615# a_908_1615# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X62 a_15779_3737# a_15566_3737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X63 gnd d0 a_9357_11208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X64 a_1329_3062# a_2169_3737# a_2377_3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X65 vdd a_9356_1554# a_9148_1554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X66 vdd a_20063_5194# a_19855_5194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X67 a_14325_12026# a_14112_12026# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X68 vdd d3 a_6820_9691# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X69 a_9098_5390# a_9102_4534# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X70 a_19809_9872# a_19813_9016# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X71 vdd d1 a_19015_5966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X72 vdd a_20064_3674# a_19856_3674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X73 a_15221_7608# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X74 a_9099_3191# a_9103_2246# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X75 gnd d0 a_20064_2995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X76 a_17311_5389# a_17568_5199# a_17273_3690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X77 a_8055_3018# a_8308_3005# a_6608_2251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X78 a_9103_2246# a_9356_2233# a_8055_1571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X79 gnd d1 a_8309_11980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X80 a_2169_2290# a_1956_2290# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X81 vdd d0 a_9358_9688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X82 a_11209_12394# a_11209_12139# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X83 gnd a_19017_11974# a_18809_11974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X84 a_9102_4534# a_9098_4711# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X85 a_18764_10540# a_19017_10527# a_17313_11397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X86 a_14110_6018# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X87 a_499_4945# a_1120_5261# a_1328_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X88 a_9099_2423# a_9356_2233# a_8055_1571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X89 a_15566_3737# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X90 a_9100_10719# a_9105_9701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X91 a_11210_8631# a_11831_9064# a_12039_9064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X92 a_3868_10587# a_4726_7614# a_4934_7614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X93 a_11208_3814# a_11208_3419# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X94 a_1123_9749# a_910_9749# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X95 a_10619_n544# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X96 a_499_6137# a_1120_6029# a_1328_6029# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X97 a_12037_3735# a_12877_3731# a_13085_3731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X98 a_3404_12032# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X99 vdd a_19015_5966# a_18807_5966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X100 a_1122_12716# a_909_12716# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X101 a_12039_9743# a_11618_9743# a_11210_9822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X102 a_9105_9022# a_9101_9199# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X103 gnd a_20064_2995# a_19856_2995# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X104 a_501_12400# a_501_12145# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X105 a_11208_1717# a_11829_1609# a_12037_1609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X106 a_8054_5985# a_9147_6647# a_9098_6837# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X107 a_13086_11259# a_12665_11259# a_12038_10584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X108 a_12876_6698# a_12663_6698# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X109 vdd a_9358_9688# a_9150_9688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X110 a_11207_6781# a_11207_6386# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X111 gnd a_6862_11213# a_6654_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X112 a_1958_8298# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X113 a_9101_7752# a_9102_6660# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X114 a_2377_2290# a_1956_2290# a_1329_1615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X115 a_1955_6704# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X116 a_17318_8253# a_17571_8240# a_17271_9875# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X117 a_11618_7617# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X118 a_13087_9739# a_12666_9739# a_12039_9743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X119 gnd a_9357_10529# a_9149_10529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X120 a_1122_10590# a_909_10590# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X121 gnd d0 a_9357_12655# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X122 vdd d0 a_9358_9009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X123 vdd d1 a_8308_1558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X124 vdd a_6862_11213# a_6654_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X125 a_9099_3870# a_9103_3014# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X126 a_19808_12160# a_19812_11215# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X127 gnd d0 a_9355_5200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X128 a_19807_2417# a_19811_1561# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X129 a_500_2373# a_1121_2294# a_1329_2294# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X130 a_9100_11398# a_9357_11208# a_8056_10546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X131 a_17314_8430# a_17571_8240# a_17271_9875# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X132 a_908_1615# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X133 a_3618_9065# a_3405_9065# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X134 a_11830_12031# a_11617_12031# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X135 gnd a_17570_11207# a_17362_11207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X136 a_1123_9070# a_910_9070# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X137 a_12663_6698# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X138 vdd d0 a_9357_12655# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X139 a_909_11269# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X140 a_502_7731# a_1123_7623# a_1331_7623# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X141 a_1122_12037# a_909_12037# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X142 a_11208_1717# a_11210_1618# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X143 a_500_2373# a_500_1978# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X144 a_12039_9064# a_11618_9064# a_11210_9172# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X145 a_4934_7614# a_4513_7614# a_3866_4579# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X146 a_12036_6023# a_12876_6698# a_13084_6698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X147 a_11829_3735# a_11616_3735# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X148 a_1328_4582# a_907_4582# a_499_4690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X149 a_6563_9881# a_6820_9691# a_5499_6669# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X150 a_2170_11265# a_1957_11265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X151 a_8050_6162# a_9147_5968# a_9098_6158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X152 vout a_10619_n544# a_10941_n544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X153 a_9100_11398# a_9104_10542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X154 a_19809_9193# a_20066_9003# a_18761_9197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X155 a_19811_1561# a_19807_1738# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X156 a_3767_4579# a_3658_4579# a_3866_4579# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X157 gnd d4 a_5752_6656# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X158 a_18762_5979# a_19015_5966# a_17315_5212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X159 a_19810_5207# a_20063_5194# a_18762_4532# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X160 vdd a_8308_1558# a_8100_1558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X161 a_12037_1609# a_11616_1609# a_11210_1618# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X162 a_19808_12160# a_20065_11970# a_18760_12164# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X163 vdd a_9358_9009# a_9150_9009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X164 vdd d0 a_20065_11202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X165 vdd d1 a_19017_10527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X166 a_1331_8302# a_2171_8298# a_2379_8298# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X167 a_13086_11259# a_14325_12026# a_14482_10700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X168 a_11209_11342# a_11209_10947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X169 a_18761_7750# a_19858_7556# a_19809_7746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X170 a_3772_4698# a_3402_6024# a_2376_5257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X171 gnd a_9355_5200# a_9147_5200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X172 a_2376_5257# a_1955_5257# a_1328_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X173 a_17269_3867# a_17361_2232# a_17312_2422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X174 a_8057_9026# a_9150_9688# a_9101_9878# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X175 a_8056_11993# a_8309_11980# a_6609_11226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X176 a_3405_9065# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X177 vdd d4 a_5752_6656# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X178 a_1120_5261# a_907_5261# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X179 a_501_11348# a_1122_11269# a_1330_11269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X180 a_9104_10542# a_9100_10719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X181 gnd d0 a_9357_11976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X182 a_12879_9739# a_12666_9739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X183 a_13086_12706# a_12665_12706# a_12038_12031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X184 a_18761_7750# a_19858_7556# a_19813_7569# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X185 a_11616_3735# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X186 a_17269_3867# a_17361_2232# a_17316_2245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X187 a_17313_11397# a_18809_10527# a_18764_10540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X188 a_11210_9172# a_11210_8631# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X189 vdd d0 a_20063_5962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X190 vdd d0 a_20064_2227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X191 vdd d1 a_19016_2999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X192 a_11209_10947# a_11209_10692# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X193 a_11830_12710# a_11617_12710# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X194 a_8050_6162# a_8307_5972# a_6607_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X195 a_1329_1615# a_908_1615# a_502_1624# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X196 a_2377_2290# a_3616_3057# a_3767_4579# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X197 a_11829_3056# a_11616_3056# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X198 a_11207_7037# a_11207_6781# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X199 a_19806_6152# a_19810_5207# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 a_8057_9026# a_8310_9013# a_6610_8259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X201 a_1956_2290# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X202 a_500_3820# a_1121_3741# a_1329_3741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X203 a_13084_5251# a_12663_5251# a_12036_4576# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X204 a_11831_8296# a_11618_8296# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X205 a_18765_7573# a_19018_7560# a_17314_8430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X206 a_9099_3191# a_9356_3001# a_8051_3195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X207 a_12666_9739# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X208 gnd d1 a_8308_1558# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X209 a_14324_3051# a_14111_3051# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X210 a_9103_2246# a_9099_2423# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X211 a_909_12716# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X212 a_1331_7623# a_910_7623# a_502_7731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X213 a_907_6708# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X214 a_3866_4579# a_3445_4579# a_3772_4698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X215 a_11830_10584# a_11617_10584# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X216 a_17315_5212# a_18807_5966# a_18758_6156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X217 vdd a_20063_5962# a_19855_5962# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X218 vdd a_20064_2227# a_19856_2227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X219 vdd a_19016_2999# a_18808_2999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X220 vdd d1 a_19015_4519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X221 a_8053_9203# a_9150_9009# a_9101_9199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X222 a_8053_9203# a_8310_9013# a_6610_8259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X223 vdd d0 a_9355_6647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X224 a_11207_5334# a_11828_5255# a_12036_5255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X225 a_2170_12712# a_1957_12712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X226 a_18761_7750# a_19018_7560# a_17314_8430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X227 a_3868_10587# a_3447_10587# a_3774_10706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X228 a_18763_3012# a_19856_3674# a_19807_3864# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X229 a_9102_4534# a_9355_4521# a_8050_4715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X230 a_11828_4576# a_11615_4576# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X231 a_501_12795# a_501_12400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X232 a_19810_6654# a_20063_6641# a_18762_5979# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X233 a_499_6137# a_499_5596# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X234 a_11616_3056# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X235 a_11210_9822# a_11210_9427# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X236 a_13085_3731# a_14324_3051# a_14475_4573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X237 a_1331_9749# a_2171_9745# a_2379_9745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X238 a_910_9070# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X239 a_18762_4532# a_19855_5194# a_19810_5207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X240 a_19813_9695# a_19809_9872# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X241 a_2376_6704# a_1955_6704# a_1328_6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X242 a_18763_3012# a_19856_3674# a_19811_3687# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X243 a_9098_4711# a_9355_4521# a_8050_4715# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X244 a_1123_8302# a_910_8302# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X245 gnd a_8308_1558# a_8100_1558# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X246 a_14111_3051# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X247 gnd d1 a_19017_10527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X248 a_19806_6831# a_20063_6641# a_18762_5979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X249 a_501_12795# a_1122_12716# a_1330_12716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X250 a_5499_6669# a_6612_9691# a_6563_9881# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X251 a_5499_6669# a_5752_6656# a_5180_3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X252 vdd a_19015_4519# a_18807_4519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X253 vdd a_9355_6647# a_9147_6647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X254 a_14574_4573# a_14153_4573# a_14475_4573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X255 a_1330_10590# a_909_10590# a_501_10698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X256 a_500_3170# a_1121_3062# a_1329_3062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X257 a_3774_10706# a_3404_12032# a_2378_12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X258 a_499_6392# a_1120_6708# a_1328_6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X259 a_499_5596# a_499_5340# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X260 a_14477_10581# a_14113_9059# a_13087_9739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X261 gnd a_17571_8240# a_17363_8240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X262 a_907_5261# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X263 a_1955_5257# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X264 a_3447_10587# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X265 vdd d2 a_6860_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X266 a_8055_3018# a_9148_3680# a_9099_3870# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X267 a_11615_4576# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X268 a_12876_5251# a_12663_5251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X269 a_909_12037# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X270 gnd d3 a_17528_9685# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X271 a_5495_6846# a_5752_6656# a_5180_3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X272 a_907_6029# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X273 a_1121_1615# a_908_1615# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X274 a_17269_3867# a_17526_3677# a_16203_6840# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X275 a_17313_11397# a_18809_10527# a_18760_10717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X276 gnd d0 a_20064_2227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X277 a_6608_2251# a_8100_3005# a_8055_3018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X278 a_15779_3737# a_15566_3737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X279 gnd a_20065_11202# a_19857_11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X280 a_8054_4538# a_9147_5200# a_9102_5213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X281 a_13087_8292# a_12666_8292# a_12039_8296# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X282 vdd a_17571_8240# a_17363_8240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X283 a_18759_3189# a_19856_2995# a_19807_3185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X284 a_8055_3018# a_9148_3680# a_9103_3693# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X285 gnd a_8309_10533# a_8101_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X286 vdd d3 a_17528_9685# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X287 a_19810_5975# a_20063_5962# a_18758_6156# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X288 a_12036_5255# a_11615_5255# a_11207_4939# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X289 a_910_9749# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X290 a_17318_8253# a_18810_9007# a_18761_9197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X291 a_2377_3737# a_1956_3737# a_1329_3062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X292 a_499_4690# a_1120_4582# a_1328_4582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X293 a_11618_8296# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X294 a_501_10698# a_502_10084# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X295 a_502_8381# a_502_7986# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X296 a_12878_11259# a_12665_11259# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X297 a_11210_7980# a_11831_8296# a_12039_8296# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X298 a_11207_6781# a_11828_6702# a_12036_6702# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X299 a_14112_12026# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X300 vdd a_8309_10533# a_8101_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X301 a_9099_2423# a_9103_1567# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X302 a_12663_5251# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X303 a_501_12145# a_1122_12037# a_1330_12037# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X304 a_6609_11226# a_6862_11213# a_6567_9704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X305 vdd d0 a_9357_11208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X306 a_19808_10713# a_19813_9695# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X307 gnd a_17528_9685# a_17320_9685# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X308 a_19813_7569# a_19809_7746# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X309 gnd a_20064_2227# a_19856_2227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X310 a_15566_3737# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X311 gnd d1 a_19015_4519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X312 a_1330_11269# a_2170_11265# a_2378_11265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X313 a_3866_4579# a_4726_7614# a_4934_7614# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X314 gnd d0 a_9355_6647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X315 a_908_2294# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X316 a_499_5596# a_1120_6029# a_1328_6029# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X317 a_12037_3056# a_12877_3731# a_13085_3731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X318 a_9105_9701# a_9358_9688# a_8057_9026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X319 a_6563_9881# a_6655_8246# a_6606_8436# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X320 a_17316_2245# a_17569_2232# a_17269_3867# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X321 a_1329_1615# a_2169_2290# a_2377_2290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X322 a_502_7986# a_502_7731# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X323 a_8051_3195# a_9148_3001# a_9099_3191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X324 a_6605_11403# a_6862_11213# a_6567_9704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X325 vdd a_17528_9685# a_17320_9685# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X326 a_1328_5261# a_907_5261# a_499_4945# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X327 a_11210_1618# a_11829_1609# a_12037_1609# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X328 a_13086_11259# a_12665_11259# a_12038_11263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X329 vdd d0 a_20065_11970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X330 a_8057_7579# a_9150_8241# a_9101_8431# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X331 a_11210_10078# a_11830_10584# a_12038_10584# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X332 a_6563_9881# a_6655_8246# a_6610_8259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X333 a_17312_2422# a_17569_2232# a_17269_3867# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X334 a_11208_1972# a_11208_1717# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X335 a_4934_7614# a_5071_3743# a_5279_3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X336 a_1957_11265# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X337 a_500_4076# a_500_3820# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X338 a_1955_6704# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X339 gnd a_6820_9691# a_6612_9691# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X340 a_12879_8292# a_12666_8292# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X341 gnd a_19015_4519# a_18807_4519# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X342 gnd d1 a_19018_9007# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X343 gnd a_9355_6647# a_9147_6647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X344 a_8057_7579# a_9150_8241# a_9105_8254# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X345 gnd a_8310_9013# a_8102_9013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X346 a_1120_6708# a_907_6708# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X347 a_11207_6131# a_11828_6023# a_12036_6023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X348 a_11617_10584# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X349 a_17273_3690# a_17526_3677# a_16203_6840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X350 a_12039_8296# a_11618_8296# a_11210_8375# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X351 a_6603_5395# a_6860_5205# a_6565_3696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X352 a_3618_9065# a_3405_9065# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X353 a_12036_6702# a_11615_6702# a_11207_6386# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X354 gnd d0 a_9355_5968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X355 a_10832_n544# a_10619_n544# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X356 a_909_11269# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X357 a_499_7043# a_1123_7623# a_1331_7623# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X358 vdd a_20065_12649# a_19857_12649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X359 a_11618_9743# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X360 a_9105_9022# a_9358_9009# a_8053_9203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X361 vdd a_8310_9013# a_8102_9013# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X362 a_4934_7614# a_4513_7614# a_3868_10587# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X363 a_12878_12706# a_12665_12706# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X364 a_19808_11392# a_19812_10536# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X365 a_12666_8292# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X366 a_9098_6158# a_9102_5213# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X367 a_19806_4705# a_19811_3687# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X368 gnd a_19018_9007# a_18810_9007# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X369 gnd d2 a_17569_2232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X370 a_12037_1609# a_11616_1609# a_11208_1717# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X371 a_19811_3008# a_19807_3185# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X372 a_2379_9745# a_3618_9065# a_3769_10587# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X373 a_1956_3737# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X374 a_1330_12716# a_2170_12712# a_2378_12712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X375 a_502_8637# a_502_8381# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X376 a_908_3741# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X377 a_14155_10581# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X378 a_3772_4698# a_3402_6024# a_2376_6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X379 vdd a_17570_11207# a_17362_11207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X380 a_500_3425# a_500_3170# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X381 a_3405_9065# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X382 gnd a_9355_5968# a_9147_5968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X383 vdd d2 a_17569_2232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X384 a_501_10953# a_1122_11269# a_1330_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X385 a_17317_11220# a_17570_11207# a_17275_9698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X386 a_1120_5261# a_907_5261# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X387 a_13086_12706# a_12665_12706# a_12038_12710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X388 a_9100_12166# a_9357_11976# a_8052_12170# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X389 gnd a_20065_11970# a_19857_11970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X390 a_18764_10540# a_19857_11202# a_19808_11392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X391 a_1120_6029# a_907_6029# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X392 a_18758_6156# a_19855_5962# a_19810_5975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X393 a_2168_5257# a_1955_5257# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X394 a_18763_1565# a_19856_2227# a_19811_2240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X395 a_1957_12712# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X396 a_19812_10536# a_20065_10523# a_18760_10717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X397 a_11210_8375# a_11210_7980# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X398 a_8056_10546# a_9149_11208# a_9100_11398# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X399 a_11829_2288# a_11616_2288# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X400 a_9105_9701# a_9101_9878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X401 gnd d0 a_9358_7562# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X402 a_12036_6023# a_11615_6023# a_11207_5590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X403 a_1329_1615# a_908_1615# a_500_1723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X404 vdd d0 a_20064_2995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X405 gnd d0 a_20066_9682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X406 a_499_6392# a_499_6137# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X407 a_11618_9064# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X408 a_11831_7617# a_11618_7617# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X409 a_8051_3195# a_8308_3005# a_6608_2251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X410 a_19808_10713# a_20065_10523# a_18760_10717# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X411 a_8057_9026# a_9150_9688# a_9105_9701# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X412 a_12039_8296# a_12879_8292# a_13087_8292# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X413 a_18763_3012# a_19016_2999# a_17316_2245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X414 a_500_3425# a_1121_3741# a_1329_3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X415 a_6609_11226# a_8101_11980# a_8052_12170# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X416 vdd d0 a_9358_7562# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X417 a_13084_5251# a_12663_5251# a_12036_5255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X418 vdd d2 a_6861_2238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X419 a_1330_11269# a_909_11269# a_501_10953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X420 vdd d0 a_20066_9682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X421 gnd d0 a_20063_4515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X422 a_3767_4579# a_3403_3057# a_2377_2290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X423 a_908_3062# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X424 a_8054_4538# a_8307_4525# a_6603_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X425 a_909_12716# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X426 a_19813_7569# a_20066_7556# a_18761_7750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X427 a_907_6708# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X428 a_8050_6162# a_9147_5968# a_9102_5981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X429 a_11616_2288# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X430 a_1121_2294# a_908_2294# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X431 a_19806_5384# a_19810_4528# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X432 gnd a_9358_7562# a_9150_7562# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X433 a_11207_4939# a_11828_5255# a_12036_5255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X434 a_19807_3185# a_19811_2240# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X435 a_910_8302# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X436 a_10941_n544# a_10832_n544# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X437 vdd a_20064_2995# a_19856_2995# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X438 vdd d0 a_20063_4515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X439 gnd a_20066_9682# a_19858_9682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X440 a_8050_4715# a_8307_4525# a_6603_5395# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X441 gnd a_20065_12649# a_19857_12649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X442 a_1123_7623# a_910_7623# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X443 a_19809_7746# a_20066_7556# a_18761_7750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X444 a_3658_4579# a_3445_4579# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X445 a_13085_2284# a_14324_3051# a_14475_4573# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X446 a_1331_9070# a_2171_9745# a_2379_9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X447 vdd d1 a_8309_11980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X448 vdd a_9358_7562# a_9150_7562# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X449 gnd d1 a_8307_5972# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X450 a_6565_3696# a_6652_5205# a_6603_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X451 vdd a_20066_9682# a_19858_9682# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X452 gnd a_20063_4515# a_19855_4515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X453 a_19808_12839# a_19812_11983# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X454 a_14482_10700# a_14112_12026# a_13086_11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X455 a_9100_12166# a_9104_11221# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X456 vdd a_19017_11974# a_18809_11974# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X457 a_909_10590# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X458 gnd d0 a_20066_9003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X459 a_907_4582# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X460 a_501_12400# a_1122_12716# a_1330_12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X461 a_8053_9203# a_9150_9009# a_9105_9022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X462 a_6604_2428# a_8100_1558# a_8055_1571# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X463 gnd d1 a_19016_1552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X464 a_9105_7575# a_9101_7752# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X465 a_13085_2284# a_12664_2284# a_12037_1609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X466 a_9105_8254# a_9358_8241# a_8057_7579# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X467 a_2171_8298# a_1958_8298# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X468 gnd d0 a_9356_3680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X469 a_500_2629# a_1121_3062# a_1329_3062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X470 a_14574_4573# a_14153_4573# a_14480_4692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X471 a_2168_6704# a_1955_6704# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X472 gnd d2 a_17568_5199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X473 vdd a_20063_4515# a_19855_4515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X474 a_8056_11993# a_9149_12655# a_9100_12845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X475 a_3660_10587# a_3447_10587# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X476 vdd d0 a_9355_5200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X477 a_12876_5251# a_12663_5251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X478 vdd d1 a_19016_1552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X479 a_17316_2245# a_18808_2999# a_18759_3189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X480 a_909_12037# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X481 a_9101_8431# a_9358_8241# a_8057_7579# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X482 a_907_6029# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X483 a_11208_2367# a_11829_2288# a_12037_2288# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X484 a_18763_1565# a_19856_2227# a_19807_2417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X485 vdd d0 a_9356_3680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X486 a_18764_11987# a_19857_12649# gnd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X487 a_11209_12139# a_11209_11598# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X488 a_19809_7746# a_19810_6654# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X489 a_1328_6708# a_907_6708# a_499_6392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X490 gnd a_8307_5972# a_8099_5972# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X491 a_9103_1567# a_9356_1554# a_8051_1748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X492 a_8056_11993# a_9149_12655# a_9104_12668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X493 a_14326_9059# a_14113_9059# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X494 a_11209_11342# a_11830_11263# a_12038_11263# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X495 a_501_10698# a_1122_10590# a_1330_10590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X496 gnd a_20066_9003# a_19858_9003# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X497 a_19811_3687# a_20064_3674# a_18763_3012# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X498 a_11210_7725# a_11831_7617# a_12039_7617# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X499 a_12036_5255# a_11615_5255# a_11207_5334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X500 gnd a_19016_1552# a_18808_1552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X501 a_1330_12716# a_909_12716# a_501_12400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X502 a_8057_7579# a_8310_7566# a_6606_8436# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X503 a_910_9749# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X504 a_15642_7608# a_15221_7608# a_14574_4573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X505 gnd a_9356_3680# a_9148_3680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X506 a_2377_3737# a_1956_3737# a_1329_3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X507 a_16207_6663# a_16460_6650# a_15888_3737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X508 gnd a_17568_5199# a_17360_5199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X509 a_9099_1744# a_9356_1554# a_8051_1748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X510 a_19806_5384# a_20063_5194# a_18762_4532# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X511 a_19807_3864# a_19811_3008# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X512 gnd a_9357_11208# a_9149_11208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X513 gnd d2 a_6861_2238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X514 a_1121_3741# a_908_3741# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X515 a_12878_11259# a_12665_11259# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X516 a_1331_9070# a_910_9070# a_502_8637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X517 vdd a_9355_5200# a_9147_5200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X518 a_19807_3864# a_20064_3674# a_18763_3012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X519 a_11207_6386# a_11828_6702# a_12036_6702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X520 a_12663_5251# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X521 vdd a_19016_1552# a_18808_1552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X522 a_501_11604# a_1122_12037# a_1330_12037# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X523 a_14112_12026# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X524 a_12038_10584# a_11617_10584# a_11209_10692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X525 a_14368_10581# a_14155_10581# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X526 a_8053_7756# a_8310_7566# a_6606_8436# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X527 a_6604_2428# a_6861_2238# a_6561_3873# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X528 a_11209_11598# a_11209_11342# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X529 a_6607_5218# a_8099_5972# a_8050_6162# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X530 vdd a_9356_3680# a_9148_3680# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X531 a_11617_11263# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X532 a_16203_6840# a_16460_6650# a_15888_3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X533 a_14480_4692# a_14110_6018# a_13084_5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X534 a_8055_1571# a_9148_2233# a_9099_2423# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X535 gnd d0 a_9356_3001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X536 a_18760_12164# a_19857_11970# a_19808_12160# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X537 a_1330_10590# a_2170_11265# a_2378_11265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X538 a_11207_6386# a_11207_6131# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X539 a_14113_9059# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X540 a_12877_2284# a_12664_2284# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X541 a_8052_12170# a_9149_11976# a_9100_12166# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X542 a_17318_8253# a_18810_9007# a_18765_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X543 a_1328_5261# a_907_5261# a_499_5340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X544 a_8055_1571# a_9148_2233# a_9103_2246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X545 gnd a_6860_5205# a_6652_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X546 a_13085_3731# a_12664_3731# a_12037_3056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X547 a_2171_9745# a_1958_9745# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X548 a_1328_6029# a_907_6029# a_499_5596# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X549 a_18758_6156# a_19015_5966# a_17315_5212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X550 a_9103_3014# a_9099_3191# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X551 a_1957_11265# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X552 a_499_6787# a_499_6392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X553 a_12037_2288# a_11616_2288# a_11208_1972# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X554 a_5180_3743# a_5071_3743# a_5279_3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X555 a_19812_11215# a_19808_11392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X556 a_19811_3008# a_20064_2995# a_18759_3189# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X557 a_14576_10581# a_14155_10581# a_14482_10700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X558 a_6604_2428# a_8100_1558# a_8051_1748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X559 a_1330_12037# a_909_12037# a_501_11604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X560 gnd a_9356_3001# a_9148_3001# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X561 a_9100_10719# a_9357_10529# a_8052_10723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X562 a_910_9070# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X563 a_3617_12032# a_3404_12032# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X564 a_8052_12170# a_8309_11980# a_6609_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X565 a_12039_7617# a_11618_7617# a_11207_7037# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X566 gnd d2 a_17570_11207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X567 a_9101_9878# a_9358_9688# a_8057_9026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X568 a_11208_3814# a_11829_3735# a_12037_3735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X569 a_1331_9749# a_910_9749# a_502_9433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X570 a_12664_2284# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X571 a_1121_3062# a_908_3062# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X572 vdd d0 a_9357_11976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X573 a_2169_2290# a_1956_2290# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X574 a_1120_6708# a_907_6708# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X575 a_11207_5590# a_11828_6023# a_12036_6023# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X576 gnd d0 a_20065_10523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X577 a_17271_9875# a_17363_8240# a_17314_8430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X578 a_12037_1609# a_12877_2284# a_13085_2284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X579 a_18764_11987# a_19857_12649# a_19808_12839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X580 a_11209_12789# a_11830_12710# a_12038_12710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X581 a_12036_6702# a_11615_6702# a_11207_6781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X582 a_11618_9743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X583 a_500_1723# a_502_1624# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X584 a_1329_2294# a_908_2294# a_500_1978# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X585 vdd d0 a_20065_10523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X586 a_17271_9875# a_17363_8240# a_17318_8253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X587 gnd a_9357_12655# a_9149_12655# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X588 a_12878_12706# a_12665_12706# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X589 vdd d1 a_19018_9007# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X590 a_11210_10078# a_11210_9822# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X591 a_12039_9743# a_12879_9739# a_13087_9739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X592 a_19811_2240# a_19807_2417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X593 a_11617_12710# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X594 a_18764_11987# a_19017_11974# a_17317_11220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X595 a_1120_4582# a_907_4582# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X596 a_1330_12037# a_2170_12712# a_2378_12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X597 a_2379_8298# a_3618_9065# a_3769_10587# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X598 a_4726_7614# a_4513_7614# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X599 a_13084_6698# a_12663_6698# a_12036_6702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X600 a_1956_3737# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X601 a_908_3741# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X602 a_5499_6669# a_6612_9691# a_6567_9704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X603 vdd a_9357_12655# a_9149_12655# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X604 a_10832_n544# a_10619_n544# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X605 a_12877_3731# a_12664_3731# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X606 a_17315_5212# a_18807_5966# a_18762_5979# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X607 a_6608_2251# a_6861_2238# a_6561_3873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X608 vdd d0 a_20064_1548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X609 a_499_4690# a_500_4076# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X610 a_16207_6663# a_17320_9685# a_17271_9875# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X611 a_11829_1609# a_11616_1609# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X612 a_9101_9199# a_9358_9009# a_8053_9203# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X613 a_8051_1748# a_8308_1558# a_6604_2428# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X614 a_11208_3164# a_11829_3056# a_12037_3056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X615 a_2379_8298# a_1958_8298# a_1331_7623# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X616 a_3615_6024# a_3402_6024# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X617 a_9102_5213# a_9355_5200# a_8054_4538# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X618 a_1120_6029# a_907_6029# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X619 a_2168_5257# a_1955_5257# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X620 a_19810_5207# a_19806_5384# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X621 vdd a_20065_11202# a_19857_11202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X622 a_502_9178# a_502_8637# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X623 vdd a_19018_9007# a_18810_9007# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X624 a_12037_3735# a_11616_3735# a_11208_3419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X625 a_1957_12712# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X626 a_11209_12139# a_11830_12031# a_12038_12031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X627 vdd a_19017_10527# a_18809_10527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X628 a_14482_10700# a_14368_10581# a_14576_10581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X629 a_16207_6663# a_17320_9685# a_17275_9698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X630 a_12036_6023# a_11615_6023# a_11207_6131# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X631 a_18759_3189# a_19856_2995# a_19811_3008# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X632 a_18765_9020# a_19858_9682# a_19809_9872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X633 a_3774_10706# a_3660_10587# a_3868_10587# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X634 a_11618_9064# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X635 a_4513_7614# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X636 a_11831_7617# a_11618_7617# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X637 a_11207_4939# a_11207_4684# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X638 a_499_7043# a_499_6787# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X639 a_12664_3731# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X640 a_5071_3743# a_4858_3743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X641 gnd a_9357_11976# a_9149_11976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X642 a_17313_11397# a_17570_11207# a_17275_9698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X643 a_9104_10542# a_9357_10529# a_8052_10723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X644 a_1328_5261# a_2168_5257# a_2376_5257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X645 vdd a_20064_1548# a_19856_1548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X646 vdd d0 a_9355_5968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X647 a_11616_1609# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X648 a_1330_11269# a_909_11269# a_501_11348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X649 a_18765_9020# a_19858_9682# a_19813_9695# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X650 gnd a_8310_7566# a_8102_7566# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X651 a_18758_4709# a_19855_4515# a_19806_4705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X652 a_11207_4684# a_11828_4576# a_12036_4576# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X653 a_11617_12031# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X654 a_11210_9427# a_11210_9172# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X655 a_3767_4579# a_3403_3057# a_2377_3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X656 a_3402_6024# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X657 a_908_3062# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X658 a_8056_10546# a_9149_11208# a_9104_11221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X659 gnd a_16460_6650# a_16252_6650# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X660 a_6610_8259# a_8102_9013# a_8053_9203# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X661 a_502_9178# a_1123_9070# a_1331_9070# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X662 a_12876_6698# a_12663_6698# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X663 a_1329_3741# a_908_3741# a_500_3425# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X664 a_18758_4709# a_19855_4515# a_19810_4528# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X665 vdd a_8310_7566# a_8102_7566# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X666 a_9104_11989# a_9100_12166# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X667 a_910_8302# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X668 a_8051_3195# a_9148_3001# a_9103_3014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X669 a_2378_12712# a_3617_12032# a_3774_10706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X670 a_13084_6698# a_14323_6018# a_14480_4692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X671 a_1123_7623# a_910_7623# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X672 vdd a_16460_6650# a_16252_6650# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X673 a_3658_4579# a_3445_4579# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X674 a_502_9828# a_502_9433# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X675 a_19806_6152# a_20063_5962# a_18758_6156# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X676 a_19807_2417# a_20064_2227# a_18763_1565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X677 a_18759_3189# a_19016_2999# a_17316_2245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X678 a_6610_8259# a_8102_9013# a_8057_9026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X679 gnd d0 a_20066_8235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X680 a_12037_3056# a_11616_3056# a_11208_2623# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X681 vdd a_9355_5968# a_9147_5968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X682 a_18761_9197# a_19858_9003# a_19809_9193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X683 a_8050_4715# a_9147_4521# a_9098_4711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X684 a_500_1978# a_1121_2294# a_1329_2294# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X685 a_14482_10700# a_14112_12026# a_13086_12706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X686 vdd a_6820_9691# a_6612_9691# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X687 a_14475_4573# a_14111_3051# a_13085_2284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X688 a_15642_7608# a_15779_3737# a_10941_n544# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X689 a_12038_11263# a_11617_11263# a_11209_10947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X690 a_2379_9745# a_1958_9745# a_1331_9070# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X691 vdd d0 a_20066_8235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X692 a_5279_3743# a_10832_n544# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X693 a_12663_6698# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X694 a_19811_3687# a_19807_3864# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X695 a_2168_6704# a_1955_6704# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X696 gnd d0 a_20064_1548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X697 a_8050_4715# a_9147_4521# a_9102_4534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X698 a_8055_1571# a_8308_1558# a_6604_2428# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X699 gnd d1 a_8309_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X700 a_9098_6837# a_9102_5981# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X701 a_5180_3743# a_5544_6656# a_5495_6846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X702 a_18758_4709# a_19015_4519# a_17311_5389# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X703 a_502_9828# a_1123_9749# a_1331_9749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X704 gnd a_20066_8235# a_19858_8235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X705 a_9098_6837# a_9355_6647# a_8054_5985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X706 a_14366_4573# a_14153_4573# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X707 a_12036_4576# a_11615_4576# a_11208_4070# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X708 gnd a_19017_10527# a_18809_10527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X709 a_1958_8298# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X710 a_1329_3062# a_908_3062# a_500_2629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X711 a_1328_6708# a_907_6708# a_499_6787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X712 a_9104_12668# a_9100_12845# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X713 a_14326_9059# a_14113_9059# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X714 a_1331_7623# a_2171_8298# a_2379_8298# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X715 a_1328_6708# a_2168_6704# a_2376_6704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X716 a_11209_10947# a_11830_11263# a_12038_11263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X717 vdd d1 a_8309_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X718 a_11207_7037# a_11831_7617# a_12039_7617# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X719 a_1330_12716# a_909_12716# a_501_12795# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X720 a_5180_3743# a_5544_6656# a_5499_6669# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X721 a_16203_6840# a_17318_3677# a_17273_3690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X722 a_11207_4684# a_11208_4070# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X723 a_1331_8302# a_910_8302# a_502_7986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X724 vdd a_20066_8235# a_19858_8235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X725 a_15642_7608# a_15221_7608# a_14576_10581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X726 vdd d2 a_17568_5199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X727 vdd d0 a_9357_10529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X728 gnd a_20064_1548# a_19856_1548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X729 gnd d1 a_8308_3005# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X730 gnd d0 a_9356_2233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X731 a_12038_11263# a_12878_11259# a_13086_11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X732 a_502_7731# a_499_7043# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X733 a_17316_2245# a_18808_2999# a_18763_3012# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X734 a_1121_3741# a_908_3741# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X735 a_501_11348# a_501_10953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X736 a_11828_5255# a_11615_5255# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X737 a_13087_9739# a_14326_9059# a_14477_10581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X738 a_11617_11263# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X739 a_12036_6702# a_12876_6698# a_13084_6698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X740 a_2169_3737# a_1956_3737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X741 a_14153_4573# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X742 a_19813_8248# a_19809_8425# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X743 a_14480_4692# a_14110_6018# a_13084_6698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X744 a_1328_4582# a_907_4582# a_500_4076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X745 vdd d0 a_9356_2233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X746 a_10941_n544# a_15566_3737# a_15888_3737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X747 a_14113_9059# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X748 a_18764_10540# a_19857_11202# a_19812_11215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X749 a_1330_10590# a_909_10590# a_502_10084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X750 a_8053_7756# a_9150_7562# a_9101_7752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X751 a_3445_4579# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X752 a_12665_11259# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X753 a_501_10953# a_501_10698# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X754 a_17275_9698# a_17528_9685# a_16207_6663# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X755 a_19811_2240# a_20064_2227# a_18763_1565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X756 vdd a_17568_5199# a_17360_5199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X757 a_9101_9199# a_9105_8254# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X758 vdd a_9357_11208# a_9149_11208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X759 gnd a_8308_3005# a_8100_3005# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X760 a_12038_12710# a_11617_12710# a_11209_12394# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X761 gnd d1 a_19017_11974# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X762 a_1328_6029# a_907_6029# a_499_6137# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X763 gnd a_9356_2233# a_9148_2233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X764 a_13085_3731# a_12664_3731# a_12037_3735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X765 a_2171_9745# a_1958_9745# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X766 a_500_1978# a_500_1723# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X767 a_2377_2290# a_1956_2290# a_1329_2294# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X768 a_17311_5389# a_18807_4519# a_18762_4532# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X769 a_8053_7756# a_9150_7562# a_9105_7575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X770 a_11615_5255# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X771 a_1330_12037# a_909_12037# a_501_12145# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X772 a_11830_10584# a_11617_10584# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X773 a_17271_9875# a_17528_9685# a_16207_6663# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X774 a_1122_10590# a_909_10590# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X775 a_3617_12032# a_3404_12032# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X776 gnd d2 a_17571_8240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X777 a_12039_7617# a_11618_7617# a_11210_7725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X778 vdd a_9356_2233# a_9148_2233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X779 a_11208_3419# a_11829_3735# a_12037_3735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X780 a_5279_3743# a_4858_3743# a_5180_3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X781 a_1331_9749# a_910_9749# a_502_9828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X782 a_1958_9745# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X783 a_1121_3062# a_908_3062# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X784 a_17317_11220# a_18809_11974# a_18760_12164# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X785 vdd a_20065_11970# a_19857_11970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X786 a_9102_5213# a_9098_5390# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X787 a_18762_4532# a_19015_4519# a_17311_5389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X788 a_19812_11215# a_20065_11202# a_18764_10540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X789 vdd d2 a_17571_8240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X790 a_9102_6660# a_9355_6647# a_8054_5985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X791 a_9100_12845# a_9104_11989# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X792 gnd a_8309_11980# a_8101_11980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X793 gnd d2 a_6862_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X794 a_8056_10546# a_8309_10533# a_6605_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X795 a_12038_12710# a_12878_12706# a_13086_12706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X796 a_11831_8296# a_11618_8296# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X797 a_1329_2294# a_2169_2290# a_2377_2290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X798 a_16203_6840# a_17318_3677# a_17269_3867# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X799 vdd d2 a_17570_11207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X800 a_6565_3696# a_6652_5205# a_6607_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X801 a_11209_12789# a_11209_12394# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X802 gnd d0 a_9357_10529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X803 a_11828_6702# a_11615_6702# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X804 a_6609_11226# a_8101_11980# a_8056_11993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X805 a_12039_9064# a_12879_9739# a_13087_9739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X806 a_12038_12031# a_11617_12031# a_11209_11598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X807 vdd d2 a_6862_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X808 a_3447_10587# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X809 vdd d0 a_20066_9003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X810 a_17273_3690# a_17360_5199# a_17311_5389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X811 a_8052_10723# a_8309_10533# a_6605_11403# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X812 a_4726_7614# a_4513_7614# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X813 a_17314_8430# a_18810_7560# a_18761_7750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X814 gnd d1 a_19015_5966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X815 gnd d0 a_20063_5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X816 a_6567_9704# a_6654_11213# a_6605_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X817 a_3868_10587# a_3447_10587# a_3769_10587# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X818 a_501_11604# a_501_11348# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X819 a_12877_3731# a_12664_3731# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X820 a_2378_11265# a_1957_11265# a_1330_10590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X821 a_9101_9878# a_9105_9022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X822 a_18765_9020# a_19018_9007# a_17318_8253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X823 a_18759_1742# a_19856_1548# a_19811_1561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X824 a_19809_8425# a_19813_7569# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X825 a_12665_12706# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X826 a_11829_1609# a_11616_1609# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X827 a_1331_9070# a_910_9070# a_502_9178# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X828 a_3769_10587# a_3405_9065# a_2379_8298# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X829 a_500_2629# a_500_2373# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X830 a_11208_2623# a_11829_3056# a_12037_3056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X831 a_17314_8430# a_18810_7560# a_18765_7573# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X832 a_6567_9704# a_6654_11213# a_6609_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X833 a_3615_6024# a_3402_6024# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X834 a_11618_8296# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X835 a_12037_3735# a_11616_3735# a_11208_3814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X836 a_500_4076# a_1120_4582# a_1328_4582# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X837 a_11209_11598# a_11830_12031# a_12038_12031# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X838 a_11210_7725# a_11207_7037# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X839 a_11615_6702# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X840 a_9102_5981# a_9355_5968# a_8050_6162# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X841 vdd a_20066_9003# a_19858_9003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X842 vdd d1 a_8307_5972# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X843 a_17311_5389# a_18807_4519# a_18758_4709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X844 a_4513_7614# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X845 gnd a_19015_5966# a_18807_5966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X846 gnd a_20063_5194# a_19855_5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X847 gnd d3 a_6820_9691# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X848 a_11208_2367# a_11208_1972# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X849 a_5071_3743# a_4858_3743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X850 a_12664_3731# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X851 a_2376_6704# a_3615_6024# a_3772_4698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X852 a_1956_2290# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X853 a_908_2294# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X854 a_9103_3693# a_9099_3870# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X855 a_11828_6023# a_11615_6023# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X856 a_1328_4582# a_2168_5257# a_2376_5257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X857 a_11616_1609# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X858 a_11617_12031# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X859 gnd d1 a_8310_9013# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X860 a_502_8381# a_1123_8302# a_1331_8302# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X861 a_11208_4070# a_11828_4576# a_12036_4576# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X862 a_11209_10692# a_11210_10078# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X863 a_910_7623# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X864 gnd d1 a_19018_7560# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X865 a_3402_6024# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X866 vdd d0 a_9356_3001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X867 a_13087_8292# a_12666_8292# a_12039_7617# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X868 a_4858_3743# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X869 a_1329_3741# a_908_3741# a_500_3820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X870 a_19812_11983# a_19808_12160# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X871 a_11831_9743# a_11618_9743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X872 vdd d1 a_8310_9013# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X873 a_19808_12839# a_20065_12649# a_18764_11987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X874 a_9104_11221# a_9100_11398# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X875 vdd a_8307_5972# a_8099_5972# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X876 a_3616_3057# a_3403_3057# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X877 a_2378_11265# a_3617_12032# a_3774_10706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X878 vdd d1 a_19018_7560# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X879 a_13084_5251# a_14323_6018# a_14480_4692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X880 a_18765_7573# a_19858_8235# a_19809_8425# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X881 a_500_1723# a_1121_1615# a_1329_1615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X882 gnd d0 a_9355_4521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X883 a_11210_8375# a_11831_8296# a_12039_8296# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X884 a_11209_12394# a_11830_12710# a_12038_12710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X885 gnd d0 a_20063_6641# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X886 vdd a_6860_5205# a_6652_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X887 a_12037_3056# a_11616_3056# a_11208_3164# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X888 a_9105_7575# a_9358_7562# a_8053_7756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X889 a_11615_6023# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X890 a_19807_3185# a_20064_2995# a_18759_3189# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X891 a_9104_12668# a_11209_12789# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X892 a_19813_9695# a_20066_9682# a_18765_9020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X893 a_12036_5255# a_12876_5251# a_13084_5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X894 a_2378_12712# a_1957_12712# a_1330_12037# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X895 a_18765_7573# a_19858_8235# a_19813_8248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X896 gnd a_19018_7560# a_18810_7560# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X897 vdd a_9356_3001# a_9148_3001# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X898 a_15888_3737# a_15779_3737# a_10941_n544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X899 vdd d0 a_9355_4521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X900 a_14475_4573# a_14111_3051# a_13085_3731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X901 a_12038_11263# a_11617_11263# a_11209_11342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X902 a_2379_9745# a_1958_9745# a_1331_9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X903 vdd d0 a_20063_6641# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X904 a_6607_5218# a_8099_5972# a_8054_5985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X905 a_9105_8254# a_9101_8431# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X906 a_9101_7752# a_9358_7562# a_8053_7756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X907 a_18759_1742# a_19856_1548# a_19807_1738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X908 a_18760_12164# a_19857_11970# a_19812_11983# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X909 a_17275_9698# a_17362_11207# a_17313_11397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X910 gnd d2 a_6863_8246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X911 a_19809_9872# a_20066_9682# a_18765_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X912 a_19810_4528# a_20063_4515# a_18758_4709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X913 a_11617_12710# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X914 a_3403_3057# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X915 vref a_501_12795# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X916 a_8052_12170# a_9149_11976# a_9104_11989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X917 a_19812_11983# a_20065_11970# a_18760_12164# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X918 vdd a_19018_7560# a_18810_7560# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X919 a_9103_1567# a_9099_1744# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X920 a_11209_10692# a_11830_10584# a_12038_10584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X921 gnd a_9355_4521# a_9147_4521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X922 a_12036_4576# a_11615_4576# a_11207_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X923 a_502_9433# a_1123_9749# a_1331_9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X924 gnd a_20063_6641# a_19855_6641# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X925 a_1329_3062# a_908_3062# a_500_3170# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X926 a_14366_4573# a_14153_4573# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X927 gnd a_19808_12839# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X928 vdd d2 a_6863_8246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X929 vdd d3 a_17526_3677# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X930 a_11831_9064# a_11618_9064# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X931 a_12879_8292# a_12666_8292# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X932 a_14576_10581# a_15434_7608# a_15642_7608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X933 a_19806_4705# a_20063_4515# a_18758_4709# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X934 a_1328_6029# a_2168_6704# a_2376_6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X935 vdd a_9355_4521# a_9147_4521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X936 a_1331_8302# a_910_8302# a_502_8381# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X937 a_11830_11263# a_11617_11263# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X938 vdd a_20063_6641# a_19855_6641# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X939 a_11207_6131# a_11207_5590# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X940 gnd d0 a_20063_5962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X941 a_19807_1738# a_11210_1618# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X942 a_11208_2623# a_11208_2367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X943 a_11617_10584# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X944 a_6567_9704# a_6820_9691# a_5499_6669# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X945 gnd a_6863_8246# a_6655_8246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X946 gnd a_5752_6656# a_5544_6656# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X947 a_8051_1748# a_9148_1554# a_9099_1744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X948 a_1122_11269# a_909_11269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X949 a_12039_8296# a_11618_8296# a_11210_7980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X950 a_8054_5985# a_8307_5972# a_6607_5218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X951 a_14480_4692# a_14366_4573# a_14574_4573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X952 a_12038_10584# a_12878_11259# a_13086_11259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X953 a_19813_9016# a_20066_9003# a_18761_9197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X954 a_19810_5975# a_19806_6152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X955 a_11828_5255# a_11615_5255# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X956 a_18763_1565# a_19016_1552# a_17312_2422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X957 a_13087_8292# a_14326_9059# a_14477_10581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X958 a_6606_8436# a_8102_7566# a_8053_7756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X959 a_15434_7608# a_15221_7608# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X960 a_9103_3693# a_9356_3680# a_8055_3018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X961 gnd d0 a_20065_11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X962 a_15888_3737# a_16252_6650# a_16203_6840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X963 a_2169_3737# a_1956_3737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X964 a_14153_4573# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X965 vdd a_6863_8246# a_6655_8246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X966 vdd a_5752_6656# a_5544_6656# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X967 a_17315_5212# a_17568_5199# a_17273_3690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X968 a_8051_1748# a_9148_1554# a_9103_1567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X969 vdd a_17526_3677# a_17318_3677# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X970 a_11210_9822# a_11831_9743# a_12039_9743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X971 a_12666_8292# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X972 a_10941_n544# a_15566_3737# a_15642_7608# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X973 a_1123_9070# a_910_9070# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X974 a_9098_5390# a_9355_5200# a_8054_4538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X975 gnd a_20065_12649# a_18764_11987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X976 a_11207_5590# a_11207_5334# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X977 a_18759_1742# a_19016_1552# a_17312_2422# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X978 a_3445_4579# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X979 a_12039_7617# a_12879_8292# a_13087_8292# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X980 a_6606_8436# a_8102_7566# a_8057_7579# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X981 a_12665_11259# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X982 gnd d0 a_9358_9688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X983 a_6561_3873# a_6653_2238# a_6608_2251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X984 a_9099_3870# a_9356_3680# a_8055_3018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X985 a_15888_3737# a_16252_6650# a_16207_6663# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X986 a_14323_6018# a_14110_6018# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X987 a_502_8637# a_1123_9070# a_1331_9070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X988 gnd a_20063_5962# a_19855_5962# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X989 a_14155_10581# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X990 a_1329_3741# a_2169_3737# a_2377_3737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X991 a_14325_12026# a_14112_12026# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X992 a_18760_12164# a_19017_11974# a_17317_11220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X993 a_11615_5255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X994 a_19812_10536# a_19808_10713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X995 a_10619_n544# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X996 a_15221_7608# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X997 a_1121_2294# a_908_2294# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X998 a_9101_8431# a_9105_7575# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X999 a_19810_6654# a_19806_6831# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1000 a_5495_6846# a_6610_3683# a_6561_3873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1001 a_11829_2288# a_11616_2288# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1002 a_5279_3743# a_4858_3743# a_4934_7614# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1003 a_1958_9745# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1004 gnd a_9358_9688# a_9150_9688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1005 a_6610_8259# a_6863_8246# a_6563_9881# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1006 gnd a_17569_2232# a_17361_2232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1007 a_14110_6018# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1008 a_9103_3014# a_9356_3001# a_8051_3195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1009 a_499_5340# a_1120_5261# a_1328_5261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1010 a_17312_2422# a_18808_1552# a_18759_1742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1011 gnd d3 a_17526_3677# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1012 a_5495_6846# a_6610_3683# a_6565_3696# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1013 a_11830_12710# a_11617_12710# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1014 a_1123_9749# a_910_9749# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1015 a_11210_9172# a_11831_9064# a_12039_9064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1016 a_907_4582# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1017 a_3404_12032# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1018 a_1122_12716# a_909_12716# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1019 a_2171_8298# a_1958_8298# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1020 a_6606_8436# a_6863_8246# a_6563_9881# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1021 a_13085_2284# a_12664_2284# a_12037_2288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1022 vdd a_17569_2232# a_17361_2232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1023 a_12038_12031# a_12878_12706# a_13086_12706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1024 a_12039_9743# a_11618_9743# a_11210_9427# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1025 gnd d0 a_9358_9009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1026 a_11210_7980# a_11210_7725# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1027 vdd a_9357_11976# a_9149_11976# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1028 a_502_10084# a_502_9828# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1029 gnd a_20065_10523# a_19857_10523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1030 a_18761_9197# a_19858_9003# a_19813_9016# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1031 a_11828_6702# a_11615_6702# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1032 a_17312_2422# a_18808_1552# a_18763_1565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1033 a_9104_11221# a_9357_11208# a_8056_10546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1034 a_12038_12031# a_11617_12031# a_11209_12139# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1035 a_11616_2288# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1036 a_18762_4532# a_19855_5194# a_19806_5384# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1037 a_11208_1972# a_11829_2288# a_12037_2288# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1038 a_11208_4070# a_11208_3814# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1039 a_2378_11265# a_1957_11265# a_1330_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1040 vdd a_20065_10523# a_19857_10523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1041 a_13087_9739# a_12666_9739# a_12039_9064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1042 a_11618_7617# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1043 gnd a_17526_3677# a_17318_3677# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1044 a_12665_12706# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1045 vdd d0 a_20065_12649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1046 a_499_5340# a_499_4945# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1047 gnd d3 a_6818_3683# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1048 a_3769_10587# a_3405_9065# a_2379_9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1049 vout a_10619_n544# a_5279_3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1050 a_6605_11403# a_8101_10533# a_8052_10723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1051 vdd a_6861_2238# a_6653_2238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1052 gnd a_9358_9009# a_9150_9009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1053 a_6561_3873# a_6653_2238# a_6604_2428# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1054 a_19810_4528# a_19806_4705# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1055 gnd d2 a_6860_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1056 a_501_12145# a_501_11604# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1057 a_11615_6702# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1058 a_908_1615# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1059 vdd d3 a_6818_3683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1060 a_17273_3690# a_17360_5199# a_17315_5212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1061 a_11830_12031# a_11617_12031# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1062 a_6608_2251# a_8100_3005# a_8051_3195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1063 a_8054_4538# a_9147_5200# a_9098_5390# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1064 a_6605_11403# a_8101_10533# a_8056_10546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1065 a_14368_10581# a_14155_10581# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1066 a_19813_9016# a_19809_9193# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1067 a_500_3170# a_500_2629# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1068 a_499_4945# a_499_4690# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1069 a_1122_12037# a_909_12037# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1070 a_3660_10587# a_3447_10587# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1071 a_18761_9197# a_19018_9007# a_17318_8253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1072 a_11829_3735# a_11616_3735# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1073 a_8052_10723# a_9149_10529# a_9104_10542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1074 a_12039_9064# a_11618_9064# a_11210_8631# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1075 vdd d1 a_8308_3005# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1076 a_2376_5257# a_3615_6024# a_3772_4698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1077 a_11828_6023# a_11615_6023# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1078 a_2170_11265# a_1957_11265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1079 a_12877_2284# a_12664_2284# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1080 a_12038_12710# a_11617_12710# a_11209_12789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1081 a_19806_6831# a_19810_5975# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1082 gnd d1 a_19016_2999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1083 gnd a_6818_3683# a_6610_3683# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1084 gnd d0 a_20065_11970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1085 a_502_9433# a_502_9178# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1086 a_502_7986# a_1123_8302# a_1331_8302# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1087 a_3772_4698# a_3658_4579# a_3866_4579# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1088 a_910_7623# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1089 a_11210_8631# a_11210_8375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1090 a_13086_12706# a_14325_12026# a_14482_10700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1091 a_4858_3743# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1092 gnd d1 a_8307_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1093 a_2376_5257# a_1955_5257# a_1328_4582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1094 a_19807_1738# a_20064_1548# a_18759_1742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1095 gnd d0 a_20066_7556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1096 a_11831_9743# a_11618_9743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1097 a_12037_2288# a_11616_2288# a_11208_2367# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1098 a_11208_3419# a_11208_3164# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1099 vdd a_6818_3683# a_6610_3683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1100 a_3616_3057# a_3403_3057# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1101 a_502_1624# a_1121_1615# a_1329_1615# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1102 a_9104_12668# a_9357_12655# a_8056_11993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1103 a_12879_9739# a_12666_9739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1104 vdd a_8308_3005# a_8100_3005# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1105 a_11616_3735# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1106 vdd d1 a_8307_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1107 a_18762_5979# a_19855_6641# a_19806_6831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1108 a_12038_10584# a_11617_10584# a_11210_10078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1109 vdd d0 a_20066_7556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1110 a_11615_6023# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1111 a_9099_1744# a_502_1624# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1112 a_12664_2284# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1113 a_12036_4576# a_12876_5251# a_13084_5251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1114 gnd a_19016_2999# a_18808_2999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1115 a_2378_12712# a_1957_12712# a_1330_12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1116 a_909_10590# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1117 a_9102_5981# a_9098_6158# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1118 a_500_3820# a_500_3425# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1119 a_9100_12845# a_9357_12655# a_8056_11993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1120 a_2377_3737# a_3616_3057# a_3767_4579# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1121 a_18762_5979# a_19855_6641# a_19810_6654# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1122 a_11829_3056# a_11616_3056# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1123 gnd a_8307_4525# a_8099_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1124 gnd a_20066_7556# a_19858_7556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1125 gnd d0 a_9358_8241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1126 a_9098_6158# a_9355_5968# a_8050_6162# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1127 gnd d0 a_20065_12649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1128 a_1329_2294# a_908_2294# a_500_2373# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1129 a_3403_3057# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1130 a_9098_4711# a_9103_3693# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1131 a_19809_9193# a_19813_8248# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1132 a_14324_3051# a_14111_3051# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1133 a_19808_11392# a_20065_11202# a_18764_10540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1134 a_12666_9739# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1135 a_6565_3696# a_6818_3683# a_5495_6846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1136 vdd a_8307_4525# a_8099_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1137 a_18760_10717# a_19017_10527# a_17313_11397# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1138 gnd a_6861_2238# a_6653_2238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1139 a_14576_10581# a_14155_10581# a_14477_10581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1140 a_1331_7623# a_910_7623# a_499_7043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1141 vdd a_20066_7556# a_19858_7556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
X1142 a_3866_4579# a_3445_4579# a_3767_4579# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1143 vdd d0 a_9358_8241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.50
C0 d3 d5 2.69fF
C1 d1 d0 11.64fF
C2 d3 vdd 10.84fF
C3 d1 d2 9.86fF
C4 d3 d2 15.70fF
C5 vdd d0 20.57fF
C6 vdd d2 9.78fF
C7 vdd d1 18.18fF
C8 d3 d4 8.57fF
C9 d4 d5 8.69fF
C10 d6 gnd 11.35fF
C11 a_19807_1738# gnd 2.27fF
C12 a_18759_1742# gnd 2.80fF
C13 a_11210_1618# gnd 17.59fF
C14 a_9099_1744# gnd 2.27fF
C15 a_8051_1748# gnd 2.80fF
C16 a_11208_1717# gnd 2.28fF
C17 a_502_1624# gnd 17.59fF
C18 a_500_1723# gnd 2.28fF
C19 a_19811_1561# gnd 3.17fF
C20 a_9103_1567# gnd 3.17fF
C21 a_18763_1565# gnd 3.33fF
C22 a_19807_2417# gnd 2.33fF
C23 a_17312_2422# gnd 4.37fF
C24 a_12037_1609# gnd 3.33fF
C25 a_11208_1972# gnd 3.17fF
C26 a_12037_2288# gnd 2.80fF
C27 a_8055_1571# gnd 3.33fF
C28 a_9099_2423# gnd 2.33fF
C29 a_6604_2428# gnd 4.37fF
C30 a_1329_1615# gnd 3.33fF
C31 a_11208_2367# gnd 2.27fF
C32 a_500_1978# gnd 3.17fF
C33 a_1329_2294# gnd 2.80fF
C34 a_500_2373# gnd 2.27fF
C35 a_19811_2240# gnd 3.43fF
C36 a_9103_2246# gnd 3.43fF
C37 a_19807_3185# gnd 2.27fF
C38 a_17316_2245# gnd 3.43fF
C39 a_18759_3189# gnd 2.80fF
C40 a_13085_2284# gnd 3.16fF
C41 a_11208_2623# gnd 3.43fF
C42 a_9099_3191# gnd 2.27fF
C43 a_6608_2251# gnd 3.43fF
C44 a_8051_3195# gnd 2.80fF
C45 a_2377_2290# gnd 3.16fF
C46 a_11208_3164# gnd 2.33fF
C47 a_500_2629# gnd 3.43fF
C48 a_500_3170# gnd 2.33fF
C49 a_19811_3008# gnd 3.17fF
C50 a_9103_3014# gnd 3.17fF
C51 a_18763_3012# gnd 3.33fF
C52 a_19807_3864# gnd 2.33fF
C53 a_17269_3867# gnd 3.27fF
C54 a_10941_n544# gnd 10.85fF
C55 a_12037_3056# gnd 3.33fF
C56 a_13085_3731# gnd 3.64fF
C57 a_11208_3419# gnd 3.17fF
C58 a_12037_3735# gnd 2.80fF
C59 a_8055_3018# gnd 3.33fF
C60 a_9099_3870# gnd 2.33fF
C61 a_6561_3873# gnd 3.27fF
C62 a_11208_3814# gnd 2.27fF
C63 a_5279_3743# gnd 11.63fF
C64 a_1329_3062# gnd 3.33fF
C65 a_2377_3737# gnd 3.64fF
C66 d5 gnd 37.29fF
C67 a_500_3425# gnd 3.17fF
C68 a_1329_3741# gnd 2.80fF
C69 a_500_3820# gnd 2.27fF
C70 a_19811_3687# gnd 3.52fF
C71 a_9103_3693# gnd 3.52fF
C72 a_19806_4705# gnd 2.27fF
C73 a_18758_4709# gnd 2.80fF
C74 a_14475_4573# gnd 3.19fF
C75 a_11208_4070# gnd 3.52fF
C76 a_9098_4711# gnd 2.27fF
C77 a_8050_4715# gnd 2.80fF
C78 a_3767_4579# gnd 3.19fF
C79 a_11207_4684# gnd 2.33fF
C80 a_500_4076# gnd 3.52fF
C81 a_499_4690# gnd 2.33fF
C82 a_19810_4528# gnd 3.17fF
C83 a_9102_4534# gnd 3.17fF
C84 a_18762_4532# gnd 3.33fF
C85 a_19806_5384# gnd 2.33fF
C86 a_17273_3690# gnd 3.19fF
C87 a_17311_5389# gnd 3.65fF
C88 a_12036_4576# gnd 3.33fF
C89 a_11207_4939# gnd 3.17fF
C90 a_12036_5255# gnd 2.80fF
C91 a_8054_4538# gnd 3.33fF
C92 a_9098_5390# gnd 2.33fF
C93 a_6565_3696# gnd 3.19fF
C94 a_6603_5395# gnd 3.65fF
C95 a_1328_4582# gnd 3.33fF
C96 a_11207_5334# gnd 2.27fF
C97 a_499_4945# gnd 3.17fF
C98 a_1328_5261# gnd 2.80fF
C99 a_499_5340# gnd 2.27fF
C100 a_19810_5207# gnd 3.43fF
C101 a_9102_5213# gnd 3.43fF
C102 a_19806_6152# gnd 2.27fF
C103 a_17315_5212# gnd 3.20fF
C104 a_18758_6156# gnd 2.80fF
C105 a_13084_5251# gnd 3.43fF
C106 a_14480_4692# gnd 3.27fF
C107 a_11207_5590# gnd 3.43fF
C108 a_9098_6158# gnd 2.27fF
C109 a_6607_5218# gnd 3.20fF
C110 a_8050_6162# gnd 2.80fF
C111 a_2376_5257# gnd 3.43fF
C112 a_3772_4698# gnd 3.27fF
C113 a_11207_6131# gnd 2.33fF
C114 a_499_5596# gnd 3.43fF
C115 a_499_6137# gnd 2.33fF
C116 a_19810_5975# gnd 3.17fF
C117 a_9102_5981# gnd 3.17fF
C118 a_18762_5979# gnd 3.33fF
C119 a_19806_6831# gnd 2.33fF
C120 a_15888_3737# gnd 4.30fF
C121 a_16203_6840# gnd 7.03fF
C122 a_12036_6023# gnd 3.33fF
C123 a_13084_6698# gnd 4.35fF
C124 a_11207_6386# gnd 3.17fF
C125 a_12036_6702# gnd 2.80fF
C126 a_8054_5985# gnd 3.33fF
C127 a_9098_6837# gnd 2.33fF
C128 a_5180_3743# gnd 4.30fF
C129 a_5495_6846# gnd 7.03fF
C130 a_1328_6029# gnd 3.33fF
C131 a_2376_6704# gnd 4.35fF
C132 a_11207_6781# gnd 2.27fF
C133 a_499_6392# gnd 3.17fF
C134 a_1328_6708# gnd 2.80fF
C135 a_499_6787# gnd 2.27fF
C136 a_19810_6654# gnd 3.62fF
C137 a_9102_6660# gnd 3.62fF
C138 a_19809_7746# gnd 2.27fF
C139 a_18761_7750# gnd 2.80fF
C140 a_14574_4573# gnd 4.97fF
C141 a_15642_7608# gnd 4.72fF
C142 a_11207_7037# gnd 3.62fF
C143 a_9101_7752# gnd 2.27fF
C144 a_8053_7756# gnd 2.80fF
C145 a_3866_4579# gnd 4.97fF
C146 a_4934_7614# gnd 4.72fF
C147 a_11210_7725# gnd 2.33fF
C148 d4 gnd 48.75fF
C149 a_499_7043# gnd 3.62fF
C150 a_502_7731# gnd 2.33fF
C151 a_19813_7569# gnd 3.17fF
C152 a_9105_7575# gnd 3.17fF
C153 a_18765_7573# gnd 3.33fF
C154 a_19809_8425# gnd 2.33fF
C155 a_17314_8430# gnd 4.35fF
C156 a_12039_7617# gnd 3.33fF
C157 a_11210_7980# gnd 3.17fF
C158 a_12039_8296# gnd 2.80fF
C159 a_8057_7579# gnd 3.33fF
C160 a_9101_8431# gnd 2.33fF
C161 a_6606_8436# gnd 4.35fF
C162 a_1331_7623# gnd 3.33fF
C163 a_11210_8375# gnd 2.27fF
C164 a_502_7986# gnd 3.17fF
C165 a_1331_8302# gnd 2.80fF
C166 a_502_8381# gnd 2.27fF
C167 a_19813_8248# gnd 3.43fF
C168 a_9105_8254# gnd 3.43fF
C169 a_19809_9193# gnd 2.27fF
C170 a_17318_8253# gnd 3.43fF
C171 a_18761_9197# gnd 2.80fF
C172 a_13087_8292# gnd 3.20fF
C173 a_11210_8631# gnd 3.43fF
C174 a_9101_9199# gnd 2.27fF
C175 a_6610_8259# gnd 3.43fF
C176 a_8053_9203# gnd 2.80fF
C177 a_2379_8298# gnd 3.20fF
C178 a_11210_9172# gnd 2.33fF
C179 a_502_8637# gnd 3.43fF
C180 a_502_9178# gnd 2.33fF
C181 a_19813_9016# gnd 3.17fF
C182 a_9105_9022# gnd 3.17fF
C183 a_18765_9020# gnd 3.33fF
C184 a_19809_9872# gnd 2.33fF
C185 a_16207_6663# gnd 4.90fF
C186 a_17271_9875# gnd 3.27fF
C187 a_12039_9064# gnd 3.33fF
C188 a_13087_9739# gnd 3.65fF
C189 a_11210_9427# gnd 3.17fF
C190 a_12039_9743# gnd 2.80fF
C191 a_8057_9026# gnd 3.33fF
C192 a_9101_9878# gnd 2.33fF
C193 a_5499_6669# gnd 4.90fF
C194 a_6563_9881# gnd 3.27fF
C195 a_1331_9070# gnd 3.33fF
C196 a_2379_9745# gnd 3.65fF
C197 a_11210_9822# gnd 2.27fF
C198 a_502_9433# gnd 3.17fF
C199 a_1331_9749# gnd 2.80fF
C200 a_502_9828# gnd 2.27fF
C201 a_19813_9695# gnd 3.52fF
C202 a_9105_9701# gnd 3.52fF
C203 a_19808_10713# gnd 2.27fF
C204 a_18760_10717# gnd 2.80fF
C205 a_14477_10581# gnd 3.19fF
C206 a_14576_10581# gnd 7.02fF
C207 a_11210_10078# gnd 3.52fF
C208 a_9100_10719# gnd 2.27fF
C209 a_8052_10723# gnd 2.80fF
C210 a_3769_10587# gnd 3.19fF
C211 a_3868_10587# gnd 7.02fF
C212 a_11209_10692# gnd 2.33fF
C213 d3 gnd 98.77fF
C214 a_502_10084# gnd 3.52fF
C215 a_501_10698# gnd 2.33fF
C216 a_19812_10536# gnd 3.17fF
C217 a_9104_10542# gnd 3.17fF
C218 a_18764_10540# gnd 3.33fF
C219 a_19808_11392# gnd 2.33fF
C220 a_17275_9698# gnd 3.19fF
C221 a_17313_11397# gnd 3.73fF
C222 a_12038_10584# gnd 3.33fF
C223 a_11209_10947# gnd 3.17fF
C224 a_12038_11263# gnd 2.80fF
C225 a_8056_10546# gnd 3.33fF
C226 a_9100_11398# gnd 2.33fF
C227 a_6567_9704# gnd 3.19fF
C228 a_6605_11403# gnd 3.73fF
C229 a_1330_10590# gnd 3.33fF
C230 a_11209_11342# gnd 2.27fF
C231 a_501_10953# gnd 3.17fF
C232 a_1330_11269# gnd 2.80fF
C233 a_501_11348# gnd 2.27fF
C234 a_19812_11215# gnd 3.43fF
C235 a_9104_11221# gnd 3.43fF
C236 a_19808_12160# gnd 2.27fF
C237 a_17317_11220# gnd 3.35fF
C238 a_18760_12164# gnd 2.80fF
C239 a_13086_11259# gnd 3.43fF
C240 a_14482_10700# gnd 3.27fF
C241 a_11209_11598# gnd 3.43fF
C242 a_9100_12166# gnd 2.27fF
C243 a_6609_11226# gnd 3.35fF
C244 a_8052_12170# gnd 2.80fF
C245 a_2378_11265# gnd 3.43fF
C246 a_3774_10706# gnd 3.27fF
C247 a_11209_12139# gnd 2.33fF
C248 d2 gnd 103.51fF
C249 a_501_11604# gnd 3.43fF
C250 a_501_12145# gnd 2.33fF
C251 a_19812_11983# gnd 3.17fF
C252 a_9104_11989# gnd 3.17fF
C253 a_18764_11987# gnd 3.40fF
C254 a_19808_12839# gnd 2.73fF
C255 a_12038_12031# gnd 3.33fF
C256 a_13086_12706# gnd 4.35fF
C257 a_11209_12394# gnd 3.17fF
C258 a_12038_12710# gnd 2.80fF
C259 a_8056_11993# gnd 3.33fF
C260 a_9100_12845# gnd 2.33fF
C261 a_1330_12037# gnd 3.33fF
C262 a_2378_12712# gnd 4.35fF
C263 a_11209_12789# gnd 2.27fF
C264 d1 gnd 121.94fF
C265 a_501_12400# gnd 3.17fF
C266 a_1330_12716# gnd 2.80fF
C267 d0 gnd 152.21fF
C268 a_501_12795# gnd 2.27fF
C269 a_9104_12668# gnd 4.89fF
C270 vdd gnd 655.73fF
