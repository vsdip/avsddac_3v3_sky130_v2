magic
tech sky130A
timestamp 1616446538
<< metal1 >>
rect -339 -218 2408 2552
<< metal3 >>
rect -339 -218 2408 2552
<< mimcap >>
rect -256 -57 2300 2433
<< end >>
