magic
tech sky130A
timestamp 1616156947
<< nwell >>
rect 41 156 852 306
rect 1053 -25 1864 125
rect 40 -259 851 -109
<< nmos >>
rect 105 55 155 97
rect 318 55 368 97
rect 526 55 576 97
rect 734 55 784 97
rect 1117 -126 1167 -84
rect 1330 -126 1380 -84
rect 1538 -126 1588 -84
rect 1746 -126 1796 -84
rect 104 -360 154 -318
rect 317 -360 367 -318
rect 525 -360 575 -318
rect 733 -360 783 -318
<< pmos >>
rect 105 174 155 274
rect 318 174 368 274
rect 526 174 576 274
rect 734 174 784 274
rect 1117 -7 1167 93
rect 1330 -7 1380 93
rect 1538 -7 1588 93
rect 1746 -7 1796 93
rect 104 -241 154 -141
rect 317 -241 367 -141
rect 525 -241 575 -141
rect 733 -241 783 -141
<< ndiff >>
rect 56 87 105 97
rect 56 67 67 87
rect 87 67 105 87
rect 56 55 105 67
rect 155 91 199 97
rect 155 71 170 91
rect 190 71 199 91
rect 155 55 199 71
rect 269 87 318 97
rect 269 67 280 87
rect 300 67 318 87
rect 269 55 318 67
rect 368 91 412 97
rect 368 71 383 91
rect 403 71 412 91
rect 368 55 412 71
rect 477 87 526 97
rect 477 67 488 87
rect 508 67 526 87
rect 477 55 526 67
rect 576 91 620 97
rect 576 71 591 91
rect 611 71 620 91
rect 576 55 620 71
rect 690 91 734 97
rect 690 71 699 91
rect 719 71 734 91
rect 690 55 734 71
rect 784 87 833 97
rect 784 67 802 87
rect 822 67 833 87
rect 784 55 833 67
rect 1068 -94 1117 -84
rect 1068 -114 1079 -94
rect 1099 -114 1117 -94
rect 1068 -126 1117 -114
rect 1167 -90 1211 -84
rect 1167 -110 1182 -90
rect 1202 -110 1211 -90
rect 1167 -126 1211 -110
rect 1281 -94 1330 -84
rect 1281 -114 1292 -94
rect 1312 -114 1330 -94
rect 1281 -126 1330 -114
rect 1380 -90 1424 -84
rect 1380 -110 1395 -90
rect 1415 -110 1424 -90
rect 1380 -126 1424 -110
rect 1489 -94 1538 -84
rect 1489 -114 1500 -94
rect 1520 -114 1538 -94
rect 1489 -126 1538 -114
rect 1588 -90 1632 -84
rect 1588 -110 1603 -90
rect 1623 -110 1632 -90
rect 1588 -126 1632 -110
rect 1702 -90 1746 -84
rect 1702 -110 1711 -90
rect 1731 -110 1746 -90
rect 1702 -126 1746 -110
rect 1796 -94 1845 -84
rect 1796 -114 1814 -94
rect 1834 -114 1845 -94
rect 1796 -126 1845 -114
rect 55 -328 104 -318
rect 55 -348 66 -328
rect 86 -348 104 -328
rect 55 -360 104 -348
rect 154 -324 198 -318
rect 154 -344 169 -324
rect 189 -344 198 -324
rect 154 -360 198 -344
rect 268 -328 317 -318
rect 268 -348 279 -328
rect 299 -348 317 -328
rect 268 -360 317 -348
rect 367 -324 411 -318
rect 367 -344 382 -324
rect 402 -344 411 -324
rect 367 -360 411 -344
rect 476 -328 525 -318
rect 476 -348 487 -328
rect 507 -348 525 -328
rect 476 -360 525 -348
rect 575 -324 619 -318
rect 575 -344 590 -324
rect 610 -344 619 -324
rect 575 -360 619 -344
rect 689 -324 733 -318
rect 689 -344 698 -324
rect 718 -344 733 -324
rect 689 -360 733 -344
rect 783 -328 832 -318
rect 783 -348 801 -328
rect 821 -348 832 -328
rect 783 -360 832 -348
<< pdiff >>
rect 61 236 105 274
rect 61 216 73 236
rect 93 216 105 236
rect 61 174 105 216
rect 155 236 197 274
rect 155 216 169 236
rect 189 216 197 236
rect 155 174 197 216
rect 274 236 318 274
rect 274 216 286 236
rect 306 216 318 236
rect 274 174 318 216
rect 368 236 410 274
rect 368 216 382 236
rect 402 216 410 236
rect 368 174 410 216
rect 482 236 526 274
rect 482 216 494 236
rect 514 216 526 236
rect 482 174 526 216
rect 576 236 618 274
rect 576 216 590 236
rect 610 216 618 236
rect 576 174 618 216
rect 692 236 734 274
rect 692 216 700 236
rect 720 216 734 236
rect 692 174 734 216
rect 784 243 829 274
rect 784 236 828 243
rect 784 216 796 236
rect 816 216 828 236
rect 784 174 828 216
rect 1073 55 1117 93
rect 1073 35 1085 55
rect 1105 35 1117 55
rect 1073 -7 1117 35
rect 1167 55 1209 93
rect 1167 35 1181 55
rect 1201 35 1209 55
rect 1167 -7 1209 35
rect 1286 55 1330 93
rect 1286 35 1298 55
rect 1318 35 1330 55
rect 1286 -7 1330 35
rect 1380 55 1422 93
rect 1380 35 1394 55
rect 1414 35 1422 55
rect 1380 -7 1422 35
rect 1494 55 1538 93
rect 1494 35 1506 55
rect 1526 35 1538 55
rect 1494 -7 1538 35
rect 1588 55 1630 93
rect 1588 35 1602 55
rect 1622 35 1630 55
rect 1588 -7 1630 35
rect 1704 55 1746 93
rect 1704 35 1712 55
rect 1732 35 1746 55
rect 1704 -7 1746 35
rect 1796 62 1841 93
rect 1796 55 1840 62
rect 1796 35 1808 55
rect 1828 35 1840 55
rect 1796 -7 1840 35
rect 60 -179 104 -141
rect 60 -199 72 -179
rect 92 -199 104 -179
rect 60 -241 104 -199
rect 154 -179 196 -141
rect 154 -199 168 -179
rect 188 -199 196 -179
rect 154 -241 196 -199
rect 273 -179 317 -141
rect 273 -199 285 -179
rect 305 -199 317 -179
rect 273 -241 317 -199
rect 367 -179 409 -141
rect 367 -199 381 -179
rect 401 -199 409 -179
rect 367 -241 409 -199
rect 481 -179 525 -141
rect 481 -199 493 -179
rect 513 -199 525 -179
rect 481 -241 525 -199
rect 575 -179 617 -141
rect 575 -199 589 -179
rect 609 -199 617 -179
rect 575 -241 617 -199
rect 691 -179 733 -141
rect 691 -199 699 -179
rect 719 -199 733 -179
rect 691 -241 733 -199
rect 783 -172 828 -141
rect 783 -179 827 -172
rect 783 -199 795 -179
rect 815 -199 827 -179
rect 783 -241 827 -199
<< ndiffc >>
rect -119 451 -101 469
rect -117 352 -99 370
rect -121 237 -103 255
rect -119 138 -101 156
rect 67 67 87 87
rect 170 71 190 91
rect 280 67 300 87
rect 383 71 403 91
rect 488 67 508 87
rect 591 71 611 91
rect 699 71 719 91
rect 802 67 822 87
rect -121 -45 -103 -27
rect 1079 -114 1099 -94
rect 1182 -110 1202 -90
rect 1292 -114 1312 -94
rect 1395 -110 1415 -90
rect 1500 -114 1520 -94
rect 1603 -110 1623 -90
rect 1711 -110 1731 -90
rect 1814 -114 1834 -94
rect -119 -144 -101 -126
rect -114 -246 -96 -228
rect -112 -345 -94 -327
rect 66 -348 86 -328
rect 169 -344 189 -324
rect 279 -348 299 -328
rect 382 -344 402 -324
rect 487 -348 507 -328
rect 590 -344 610 -324
rect 698 -344 718 -324
rect 801 -348 821 -328
<< pdiffc >>
rect 73 216 93 236
rect 169 216 189 236
rect 286 216 306 236
rect 382 216 402 236
rect 494 216 514 236
rect 590 216 610 236
rect 700 216 720 236
rect 796 216 816 236
rect 1085 35 1105 55
rect 1181 35 1201 55
rect 1298 35 1318 55
rect 1394 35 1414 55
rect 1506 35 1526 55
rect 1602 35 1622 55
rect 1712 35 1732 55
rect 1808 35 1828 55
rect 72 -199 92 -179
rect 168 -199 188 -179
rect 285 -199 305 -179
rect 381 -199 401 -179
rect 493 -199 513 -179
rect 589 -199 609 -179
rect 699 -199 719 -179
rect 795 -199 815 -179
<< poly >>
rect 105 274 155 287
rect 318 274 368 287
rect 526 274 576 287
rect 734 274 784 287
rect 105 146 155 174
rect 105 126 118 146
rect 138 126 155 146
rect 105 97 155 126
rect 318 145 368 174
rect 318 121 329 145
rect 353 121 368 145
rect 318 97 368 121
rect 526 150 576 174
rect 526 126 538 150
rect 562 126 576 150
rect 526 97 576 126
rect 734 148 784 174
rect 734 122 752 148
rect 778 122 784 148
rect 734 97 784 122
rect 1117 93 1167 106
rect 1330 93 1380 106
rect 1538 93 1588 106
rect 1746 93 1796 106
rect 105 39 155 55
rect 318 39 368 55
rect 526 39 576 55
rect 734 39 784 55
rect 1117 -35 1167 -7
rect 1117 -55 1130 -35
rect 1150 -55 1167 -35
rect 1117 -84 1167 -55
rect 1330 -36 1380 -7
rect 1330 -60 1341 -36
rect 1365 -60 1380 -36
rect 1330 -84 1380 -60
rect 1538 -31 1588 -7
rect 1538 -55 1550 -31
rect 1574 -55 1588 -31
rect 1538 -84 1588 -55
rect 1746 -33 1796 -7
rect 1746 -59 1764 -33
rect 1790 -59 1796 -33
rect 1746 -84 1796 -59
rect 104 -141 154 -128
rect 317 -141 367 -128
rect 525 -141 575 -128
rect 733 -141 783 -128
rect 1117 -142 1167 -126
rect 1330 -142 1380 -126
rect 1538 -142 1588 -126
rect 1746 -142 1796 -126
rect 104 -269 154 -241
rect 104 -289 117 -269
rect 137 -289 154 -269
rect 104 -318 154 -289
rect 317 -270 367 -241
rect 317 -294 328 -270
rect 352 -294 367 -270
rect 317 -318 367 -294
rect 525 -265 575 -241
rect 525 -289 537 -265
rect 561 -289 575 -265
rect 525 -318 575 -289
rect 733 -267 783 -241
rect 733 -293 751 -267
rect 777 -293 783 -267
rect 733 -318 783 -293
rect 104 -376 154 -360
rect 317 -376 367 -360
rect 525 -376 575 -360
rect 733 -376 783 -360
<< polycont >>
rect 118 126 138 146
rect 329 121 353 145
rect 538 126 562 150
rect 752 122 778 148
rect 1130 -55 1150 -35
rect 1341 -60 1365 -36
rect 1550 -55 1574 -31
rect 1764 -59 1790 -33
rect 117 -289 137 -269
rect 328 -294 352 -270
rect 537 -289 561 -265
rect 751 -293 777 -267
<< ndiffres >>
rect -140 469 -83 488
rect -140 466 -119 469
rect -234 451 -119 466
rect -101 451 -83 469
rect -234 428 -83 451
rect -234 392 -192 428
rect -235 391 -135 392
rect -235 370 -79 391
rect -235 352 -117 370
rect -99 352 -79 370
rect -235 348 -79 352
rect -140 332 -79 348
rect -142 255 -85 274
rect -142 252 -121 255
rect -236 237 -121 252
rect -103 237 -85 255
rect -236 214 -85 237
rect -236 178 -194 214
rect -237 177 -137 178
rect -237 156 -81 177
rect -237 138 -119 156
rect -101 138 -81 156
rect -237 134 -81 138
rect -142 118 -81 134
rect -142 -27 -85 -8
rect -142 -30 -121 -27
rect -236 -45 -121 -30
rect -103 -45 -85 -27
rect -236 -68 -85 -45
rect -236 -104 -194 -68
rect -237 -105 -137 -104
rect -237 -126 -81 -105
rect -237 -144 -119 -126
rect -101 -144 -81 -126
rect -237 -148 -81 -144
rect -142 -164 -81 -148
rect -135 -228 -78 -209
rect -135 -231 -114 -228
rect -229 -246 -114 -231
rect -96 -246 -78 -228
rect -229 -269 -78 -246
rect -229 -305 -187 -269
rect -230 -306 -130 -305
rect -230 -327 -74 -306
rect -230 -345 -112 -327
rect -94 -345 -74 -327
rect -230 -349 -74 -345
rect -135 -365 -74 -349
<< locali >>
rect -127 478 -92 526
rect -129 469 -92 478
rect -129 451 -119 469
rect -101 451 -92 469
rect -129 441 -92 451
rect -126 377 -89 379
rect -126 376 522 377
rect -127 370 522 376
rect -127 352 -117 370
rect -99 356 522 370
rect -99 352 -89 356
rect 352 355 522 356
rect -127 342 -89 352
rect -127 264 -92 342
rect 485 332 522 355
rect -131 255 -92 264
rect -131 237 -121 255
rect -103 237 -92 255
rect -131 231 -92 237
rect 64 307 314 331
rect 64 236 101 307
rect 216 246 247 247
rect -131 227 -94 231
rect 64 216 73 236
rect 93 216 101 236
rect 64 206 101 216
rect 160 236 247 246
rect 160 216 169 236
rect 189 216 247 236
rect 160 207 247 216
rect 160 206 197 207
rect -128 156 -91 165
rect -130 138 -119 156
rect -101 138 -91 156
rect 216 154 247 207
rect 277 236 314 307
rect 485 312 878 332
rect 898 312 901 332
rect 485 307 901 312
rect 485 306 826 307
rect 429 246 460 247
rect 277 216 286 236
rect 306 216 314 236
rect 277 206 314 216
rect 373 239 460 246
rect 373 236 434 239
rect 373 216 382 236
rect 402 219 434 236
rect 455 219 460 239
rect 402 216 460 219
rect 373 209 460 216
rect 485 236 522 306
rect 788 305 825 306
rect 637 246 673 247
rect 485 216 494 236
rect 514 216 522 236
rect 373 207 429 209
rect 373 206 410 207
rect 485 206 522 216
rect 581 236 729 246
rect 829 243 925 245
rect 581 216 590 236
rect 610 216 700 236
rect 720 216 729 236
rect 581 207 729 216
rect 787 236 925 243
rect 787 216 796 236
rect 816 216 925 236
rect 787 207 925 216
rect 581 206 618 207
rect 637 155 673 207
rect 692 206 729 207
rect 788 206 825 207
rect 108 153 149 154
rect -130 -11 -91 138
rect 0 146 149 153
rect 0 126 118 146
rect 138 126 149 146
rect 0 118 149 126
rect 216 150 575 154
rect 216 145 538 150
rect 216 121 329 145
rect 353 126 538 145
rect 562 126 575 150
rect 353 121 575 126
rect 216 118 575 121
rect 637 118 672 155
rect 740 152 840 155
rect 740 148 807 152
rect 740 122 752 148
rect 778 126 807 148
rect 833 126 840 152
rect 778 122 840 126
rect 740 118 840 122
rect 216 97 247 118
rect 637 97 673 118
rect 59 96 96 97
rect 58 87 96 96
rect 58 67 67 87
rect 87 67 96 87
rect 58 59 96 67
rect 162 91 247 97
rect 272 96 309 97
rect 162 71 170 91
rect 190 71 247 91
rect 162 63 247 71
rect 271 87 309 96
rect 271 67 280 87
rect 300 67 309 87
rect 162 62 198 63
rect 271 59 309 67
rect 375 91 460 97
rect 480 96 517 97
rect 375 71 383 91
rect 403 90 460 91
rect 403 71 432 90
rect 375 70 432 71
rect 453 70 460 90
rect 375 63 460 70
rect 479 87 517 96
rect 479 67 488 87
rect 508 67 517 87
rect 375 62 411 63
rect 479 59 517 67
rect 583 92 727 97
rect 583 91 648 92
rect 583 71 591 91
rect 611 71 648 91
rect 670 91 727 92
rect 670 71 699 91
rect 719 71 727 91
rect 583 63 727 71
rect 583 62 619 63
rect 691 62 727 63
rect 793 96 830 97
rect 793 95 831 96
rect 793 87 857 95
rect 793 67 802 87
rect 822 73 857 87
rect 877 73 880 93
rect 822 68 880 73
rect 822 67 857 68
rect 59 30 96 59
rect 60 28 96 30
rect 272 28 309 59
rect 60 6 309 28
rect 480 27 517 59
rect 793 55 857 67
rect 897 29 924 207
rect 756 27 924 29
rect 480 1 924 27
rect 1076 126 1326 150
rect 1076 55 1113 126
rect 1228 65 1259 66
rect 1076 35 1085 55
rect 1105 35 1113 55
rect 1076 25 1113 35
rect 1172 55 1259 65
rect 1172 35 1181 55
rect 1201 35 1259 55
rect 1172 26 1259 35
rect 1172 25 1209 26
rect 480 -9 502 1
rect 756 0 924 1
rect 440 -11 502 -9
rect -130 -18 502 -11
rect -131 -27 502 -18
rect 1228 -27 1259 26
rect 1289 55 1326 126
rect 1497 131 1890 151
rect 1910 131 1913 151
rect 1497 126 1913 131
rect 1497 125 1838 126
rect 1441 65 1472 66
rect 1289 35 1298 55
rect 1318 35 1326 55
rect 1289 25 1326 35
rect 1385 58 1472 65
rect 1385 55 1446 58
rect 1385 35 1394 55
rect 1414 38 1446 55
rect 1467 38 1472 58
rect 1414 35 1472 38
rect 1385 28 1472 35
rect 1497 55 1534 125
rect 1800 124 1837 125
rect 1649 65 1685 66
rect 1497 35 1506 55
rect 1526 35 1534 55
rect 1385 26 1441 28
rect 1385 25 1422 26
rect 1497 25 1534 35
rect 1593 55 1741 65
rect 1841 62 1937 64
rect 1593 35 1602 55
rect 1622 35 1712 55
rect 1732 35 1741 55
rect 1593 26 1741 35
rect 1799 55 1937 62
rect 1799 35 1808 55
rect 1828 35 1937 55
rect 1799 26 1937 35
rect 1593 25 1630 26
rect 1649 -26 1685 26
rect 1704 25 1741 26
rect 1800 25 1837 26
rect -131 -45 -121 -27
rect -103 -28 502 -27
rect 1120 -28 1161 -27
rect -103 -33 -82 -28
rect -103 -45 -91 -33
rect 1012 -35 1161 -28
rect -131 -53 -91 -45
rect -48 -46 -22 -45
rect -131 -55 -94 -53
rect -48 -64 506 -46
rect 1012 -55 1130 -35
rect 1150 -55 1161 -35
rect 1012 -63 1161 -55
rect 1228 -31 1587 -27
rect 1228 -36 1550 -31
rect 1228 -60 1341 -36
rect 1365 -55 1550 -36
rect 1574 -55 1587 -31
rect 1365 -60 1587 -55
rect 1228 -63 1587 -60
rect 1649 -63 1684 -26
rect 1752 -29 1852 -26
rect 1752 -33 1819 -29
rect 1752 -59 1764 -33
rect 1790 -55 1819 -33
rect 1845 -55 1852 -29
rect 1790 -59 1852 -55
rect 1752 -63 1852 -59
rect -128 -123 -91 -117
rect -48 -123 -22 -64
rect 485 -83 506 -64
rect -128 -126 -22 -123
rect -128 -144 -119 -126
rect -101 -140 -22 -126
rect 63 -108 313 -84
rect -101 -142 -25 -140
rect -101 -144 -91 -142
rect -128 -154 -91 -144
rect -123 -219 -92 -154
rect 63 -179 100 -108
rect 215 -169 246 -168
rect 63 -199 72 -179
rect 92 -199 100 -179
rect 63 -209 100 -199
rect 159 -179 246 -169
rect 159 -199 168 -179
rect 188 -199 246 -179
rect 159 -208 246 -199
rect 159 -209 196 -208
rect -124 -228 -87 -219
rect -124 -246 -114 -228
rect -96 -246 -87 -228
rect -124 -256 -87 -246
rect 215 -261 246 -208
rect 276 -179 313 -108
rect 484 -103 877 -83
rect 897 -103 900 -83
rect 1228 -84 1259 -63
rect 1649 -84 1685 -63
rect 1071 -85 1108 -84
rect 484 -108 900 -103
rect 1070 -94 1108 -85
rect 484 -109 825 -108
rect 428 -169 459 -168
rect 276 -199 285 -179
rect 305 -199 313 -179
rect 276 -209 313 -199
rect 372 -176 459 -169
rect 372 -179 433 -176
rect 372 -199 381 -179
rect 401 -196 433 -179
rect 454 -196 459 -176
rect 401 -199 459 -196
rect 372 -206 459 -199
rect 484 -179 521 -109
rect 787 -110 824 -109
rect 1070 -114 1079 -94
rect 1099 -114 1108 -94
rect 1070 -122 1108 -114
rect 1174 -90 1259 -84
rect 1284 -85 1321 -84
rect 1174 -110 1182 -90
rect 1202 -110 1259 -90
rect 1174 -118 1259 -110
rect 1283 -94 1321 -85
rect 1283 -114 1292 -94
rect 1312 -114 1321 -94
rect 1174 -119 1210 -118
rect 1283 -122 1321 -114
rect 1387 -90 1472 -84
rect 1492 -85 1529 -84
rect 1387 -110 1395 -90
rect 1415 -91 1472 -90
rect 1415 -110 1444 -91
rect 1387 -111 1444 -110
rect 1465 -111 1472 -91
rect 1387 -118 1472 -111
rect 1491 -94 1529 -85
rect 1491 -114 1500 -94
rect 1520 -114 1529 -94
rect 1387 -119 1423 -118
rect 1491 -122 1529 -114
rect 1595 -90 1739 -84
rect 1595 -110 1603 -90
rect 1623 -110 1711 -90
rect 1731 -110 1739 -90
rect 1595 -118 1739 -110
rect 1595 -119 1631 -118
rect 1703 -119 1739 -118
rect 1805 -85 1842 -84
rect 1805 -86 1843 -85
rect 1805 -94 1869 -86
rect 1805 -114 1814 -94
rect 1834 -108 1869 -94
rect 1889 -108 1892 -88
rect 1834 -113 1892 -108
rect 1834 -114 1869 -113
rect 1071 -151 1108 -122
rect 1072 -153 1108 -151
rect 1284 -153 1321 -122
rect 636 -169 672 -168
rect 484 -199 493 -179
rect 513 -199 521 -179
rect 372 -208 428 -206
rect 372 -209 409 -208
rect 484 -209 521 -199
rect 580 -179 728 -169
rect 828 -172 924 -170
rect 580 -199 589 -179
rect 609 -199 699 -179
rect 719 -199 728 -179
rect 580 -208 728 -199
rect 786 -179 924 -172
rect 1072 -175 1321 -153
rect 1492 -154 1529 -122
rect 1805 -126 1869 -114
rect 1909 -152 1936 26
rect 1768 -154 1936 -152
rect 1492 -158 1936 -154
rect 786 -199 795 -179
rect 815 -199 924 -179
rect 1492 -177 1541 -158
rect 1561 -177 1936 -158
rect 1492 -180 1936 -177
rect 1768 -181 1936 -180
rect 786 -208 924 -199
rect 580 -209 617 -208
rect 636 -260 672 -208
rect 691 -209 728 -208
rect 787 -209 824 -208
rect 107 -262 148 -261
rect -1 -269 148 -262
rect -1 -289 117 -269
rect 137 -289 148 -269
rect -1 -297 148 -289
rect 215 -265 574 -261
rect 215 -270 537 -265
rect 215 -294 328 -270
rect 352 -289 537 -270
rect 561 -289 574 -265
rect 352 -294 574 -289
rect 215 -297 574 -294
rect 636 -297 671 -260
rect 739 -263 839 -260
rect 739 -267 806 -263
rect 739 -293 751 -267
rect 777 -289 806 -267
rect 832 -289 839 -263
rect 777 -293 839 -289
rect 739 -297 839 -293
rect 215 -318 246 -297
rect 636 -318 672 -297
rect -121 -327 -84 -318
rect 58 -319 95 -318
rect -121 -345 -112 -327
rect -94 -345 -84 -327
rect -121 -355 -84 -345
rect -120 -390 -84 -355
rect 57 -328 95 -319
rect 57 -348 66 -328
rect 86 -348 95 -328
rect 57 -356 95 -348
rect 161 -324 246 -318
rect 271 -319 308 -318
rect 161 -344 169 -324
rect 189 -344 246 -324
rect 161 -352 246 -344
rect 270 -328 308 -319
rect 270 -348 279 -328
rect 299 -348 308 -328
rect 161 -353 197 -352
rect 270 -356 308 -348
rect 374 -324 459 -318
rect 479 -319 516 -318
rect 374 -344 382 -324
rect 402 -325 459 -324
rect 402 -344 431 -325
rect 374 -345 431 -344
rect 452 -345 459 -325
rect 374 -352 459 -345
rect 478 -328 516 -319
rect 478 -348 487 -328
rect 507 -348 516 -328
rect 374 -353 410 -352
rect 478 -356 516 -348
rect 582 -324 726 -318
rect 582 -344 590 -324
rect 610 -325 698 -324
rect 610 -344 638 -325
rect 582 -346 638 -344
rect 660 -344 698 -325
rect 718 -344 726 -324
rect 660 -346 726 -344
rect 582 -352 726 -346
rect 582 -353 618 -352
rect 690 -353 726 -352
rect 792 -319 829 -318
rect 792 -320 830 -319
rect 792 -328 856 -320
rect 792 -348 801 -328
rect 821 -342 856 -328
rect 876 -342 879 -322
rect 821 -347 879 -342
rect 821 -348 856 -347
rect 58 -385 95 -356
rect -122 -431 -84 -390
rect 59 -387 95 -385
rect 271 -387 308 -356
rect 59 -409 308 -387
rect 479 -388 516 -356
rect 792 -360 856 -348
rect 896 -386 923 -208
rect 755 -388 923 -386
rect 479 -414 923 -388
rect 480 -431 504 -414
rect 755 -415 923 -414
rect -122 -449 505 -431
rect -122 -455 -84 -449
<< viali >>
rect 878 312 898 332
rect 434 219 455 239
rect 807 126 833 152
rect 432 70 453 90
rect 648 71 670 92
rect 857 73 877 93
rect 1890 131 1910 151
rect 1446 38 1467 58
rect 1819 -55 1845 -29
rect 877 -103 897 -83
rect 433 -196 454 -176
rect 1444 -111 1465 -91
rect 1869 -108 1889 -88
rect 1541 -177 1561 -158
rect 806 -289 832 -263
rect 431 -345 452 -325
rect 638 -346 660 -325
rect 856 -342 876 -322
<< metal1 >>
rect 874 337 906 338
rect 871 332 906 337
rect 871 312 878 332
rect 898 312 906 332
rect 871 304 906 312
rect 427 239 459 246
rect 427 219 434 239
rect 455 219 459 239
rect 427 154 459 219
rect 797 154 837 155
rect 427 152 839 154
rect 427 126 807 152
rect 833 126 839 152
rect 427 118 839 126
rect 427 90 459 118
rect 872 98 906 304
rect 427 70 432 90
rect 453 70 459 90
rect 427 63 459 70
rect 636 92 676 97
rect 636 71 648 92
rect 670 71 676 92
rect 636 59 676 71
rect 850 93 906 98
rect 850 73 857 93
rect 877 73 906 93
rect 850 66 906 73
rect 963 167 1920 186
rect 850 65 885 66
rect 642 27 670 59
rect 963 27 994 167
rect 1883 151 1918 167
rect 1883 131 1890 151
rect 1910 131 1918 151
rect 1883 123 1918 131
rect 642 -4 994 27
rect 1439 58 1471 65
rect 1439 38 1446 58
rect 1467 38 1471 58
rect 1439 -27 1471 38
rect 1809 -27 1849 -26
rect 1439 -29 1851 -27
rect 1439 -55 1819 -29
rect 1845 -55 1851 -29
rect 1439 -63 1851 -55
rect 873 -78 905 -77
rect 870 -83 905 -78
rect 870 -103 877 -83
rect 897 -103 905 -83
rect 870 -111 905 -103
rect 426 -176 458 -169
rect 426 -196 433 -176
rect 454 -196 458 -176
rect 426 -261 458 -196
rect 796 -261 836 -260
rect 426 -263 838 -261
rect 426 -289 806 -263
rect 832 -289 838 -263
rect 426 -297 838 -289
rect 426 -325 458 -297
rect 426 -345 431 -325
rect 452 -345 458 -325
rect 426 -352 458 -345
rect 626 -325 676 -316
rect 871 -317 905 -111
rect 1439 -91 1471 -63
rect 1884 -83 1918 123
rect 1439 -111 1444 -91
rect 1465 -111 1471 -91
rect 1439 -118 1471 -111
rect 1862 -88 1918 -83
rect 1862 -108 1869 -88
rect 1889 -108 1918 -88
rect 1862 -115 1918 -108
rect 1862 -116 1897 -115
rect 1533 -158 1569 -154
rect 1533 -177 1541 -158
rect 1561 -177 1569 -158
rect 1533 -180 1569 -177
rect 1534 -208 1568 -180
rect 626 -346 638 -325
rect 660 -346 676 -325
rect 626 -354 676 -346
rect 849 -322 905 -317
rect 849 -342 856 -322
rect 876 -342 905 -322
rect 849 -349 905 -342
rect 1006 -236 1569 -208
rect 849 -350 884 -349
rect 631 -387 672 -354
rect 1006 -387 1046 -236
rect 631 -416 1046 -387
rect 631 -417 1040 -416
<< labels >>
rlabel locali 67 316 96 322 1 vdd
rlabel locali 280 313 309 319 1 vdd
rlabel locali 13 128 35 143 1 d0
rlabel nwell 434 283 457 286 1 vdd
rlabel locali 64 17 93 23 1 gnd
rlabel locali 277 17 306 23 1 gnd
rlabel space 374 12 403 21 1 gnd
rlabel locali 66 -99 95 -93 1 vdd
rlabel locali 279 -102 308 -96 1 vdd
rlabel locali 12 -287 34 -272 1 d0
rlabel nwell 433 -132 456 -129 1 vdd
rlabel locali 63 -398 92 -392 1 gnd
rlabel locali 276 -398 305 -392 1 gnd
rlabel space 373 -403 402 -394 1 gnd
rlabel locali 1079 135 1108 141 1 vdd
rlabel locali 1292 132 1321 138 1 vdd
rlabel locali 1655 -18 1677 -3 1 vout
rlabel nwell 1446 102 1469 105 1 vdd
rlabel locali 1076 -164 1105 -158 1 gnd
rlabel locali 1289 -164 1318 -158 1 gnd
rlabel space 1386 -169 1415 -160 1 gnd
rlabel locali 1017 -54 1064 -33 1 d1
rlabel locali -121 508 -96 517 1 vref
rlabel locali -116 -447 -89 -434 1 gnd
<< end >>
