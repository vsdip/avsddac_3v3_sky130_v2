magic
tech sky130A
timestamp 1633161908
<< nwell >>
rect 795 12817 1606 13041
rect 1843 12813 2654 13037
rect 11503 12811 12314 13035
rect 12551 12807 13362 13031
rect 9081 12562 9892 12786
rect 19789 12556 20600 12780
rect 795 12138 1606 12362
rect 3290 12133 4101 12357
rect 11503 12132 12314 12356
rect 13998 12127 14809 12351
rect 8033 11887 8844 12111
rect 9081 11883 9892 12107
rect 18741 11881 19552 12105
rect 19789 11877 20600 12101
rect 795 11370 1606 11594
rect 1843 11366 2654 11590
rect 11503 11364 12314 11588
rect 12551 11360 13362 11584
rect 6586 11120 7397 11344
rect 9081 11115 9892 11339
rect 17294 11114 18105 11338
rect 19789 11109 20600 11333
rect 795 10691 1606 10915
rect 3333 10688 4144 10912
rect 11503 10685 12314 10909
rect 14041 10682 14852 10906
rect 8033 10440 8844 10664
rect 9081 10436 9892 10660
rect 18741 10434 19552 10658
rect 19789 10430 20600 10654
rect 796 9850 1607 10074
rect 1844 9846 2655 10070
rect 11504 9844 12315 10068
rect 12552 9840 13363 10064
rect 6544 9598 7355 9822
rect 9082 9595 9893 9819
rect 17252 9592 18063 9816
rect 19790 9589 20601 9813
rect 796 9171 1607 9395
rect 3291 9166 4102 9390
rect 11504 9165 12315 9389
rect 13999 9160 14810 9384
rect 8034 8920 8845 9144
rect 9082 8916 9893 9140
rect 18742 8914 19553 9138
rect 19790 8910 20601 9134
rect 796 8403 1607 8627
rect 1844 8399 2655 8623
rect 11504 8397 12315 8621
rect 12552 8393 13363 8617
rect 6587 8153 7398 8377
rect 9082 8148 9893 8372
rect 17295 8147 18106 8371
rect 19790 8142 20601 8366
rect 796 7724 1607 7948
rect 4399 7715 5210 7939
rect 11504 7718 12315 7942
rect 15107 7709 15918 7933
rect 8034 7473 8845 7697
rect 9082 7469 9893 7693
rect 18742 7467 19553 7691
rect 19790 7463 20601 7687
rect 793 6809 1604 7033
rect 1841 6805 2652 7029
rect 11501 6803 12312 7027
rect 12549 6799 13360 7023
rect 5476 6563 6287 6787
rect 9079 6554 9890 6778
rect 16184 6557 16995 6781
rect 19787 6548 20598 6772
rect 793 6130 1604 6354
rect 3288 6125 4099 6349
rect 11501 6124 12312 6348
rect 13996 6119 14807 6343
rect 8031 5879 8842 6103
rect 9079 5875 9890 6099
rect 18739 5873 19550 6097
rect 19787 5869 20598 6093
rect 793 5362 1604 5586
rect 1841 5358 2652 5582
rect 11501 5356 12312 5580
rect 12549 5352 13360 5576
rect 6584 5112 7395 5336
rect 9079 5107 9890 5331
rect 17292 5106 18103 5330
rect 19787 5101 20598 5325
rect 793 4683 1604 4907
rect 3331 4680 4142 4904
rect 11501 4677 12312 4901
rect 14039 4674 14850 4898
rect 8031 4432 8842 4656
rect 9079 4428 9890 4652
rect 18739 4426 19550 4650
rect 19787 4422 20598 4646
rect 794 3842 1605 4066
rect 1842 3838 2653 4062
rect 4744 3844 5555 4068
rect 11502 3836 12313 4060
rect 12550 3832 13361 4056
rect 15452 3838 16263 4062
rect 6542 3590 7353 3814
rect 9080 3587 9891 3811
rect 17250 3584 18061 3808
rect 19788 3581 20599 3805
rect 794 3163 1605 3387
rect 3289 3158 4100 3382
rect 11502 3157 12313 3381
rect 13997 3152 14808 3376
rect 8032 2912 8843 3136
rect 9080 2908 9891 3132
rect 18740 2906 19551 3130
rect 19788 2902 20599 3126
rect 794 2395 1605 2619
rect 1842 2391 2653 2615
rect 11502 2389 12313 2613
rect 12550 2385 13361 2609
rect 6585 2145 7396 2369
rect 9080 2140 9891 2364
rect 17293 2139 18104 2363
rect 19788 2134 20599 2358
rect 794 1716 1605 1940
rect 11502 1710 12313 1934
rect 8032 1465 8843 1689
rect 9080 1461 9891 1685
rect 18740 1459 19551 1683
rect 19788 1455 20599 1679
rect 10505 -443 11316 -219
<< nmos >>
rect 9149 12845 9199 12887
rect 9357 12845 9407 12887
rect 9565 12845 9615 12887
rect 9778 12845 9828 12887
rect 859 12716 909 12758
rect 1072 12716 1122 12758
rect 1280 12716 1330 12758
rect 1488 12716 1538 12758
rect 1907 12712 1957 12754
rect 2120 12712 2170 12754
rect 2328 12712 2378 12754
rect 2536 12712 2586 12754
rect 19857 12839 19907 12881
rect 20065 12839 20115 12881
rect 20273 12839 20323 12881
rect 20486 12839 20536 12881
rect 11567 12710 11617 12752
rect 11780 12710 11830 12752
rect 11988 12710 12038 12752
rect 12196 12710 12246 12752
rect 12615 12706 12665 12748
rect 12828 12706 12878 12748
rect 13036 12706 13086 12748
rect 13244 12706 13294 12748
rect 8101 12170 8151 12212
rect 8309 12170 8359 12212
rect 8517 12170 8567 12212
rect 8730 12170 8780 12212
rect 859 12037 909 12079
rect 1072 12037 1122 12079
rect 1280 12037 1330 12079
rect 1488 12037 1538 12079
rect 9149 12166 9199 12208
rect 9357 12166 9407 12208
rect 9565 12166 9615 12208
rect 9778 12166 9828 12208
rect 3354 12032 3404 12074
rect 3567 12032 3617 12074
rect 3775 12032 3825 12074
rect 3983 12032 4033 12074
rect 18809 12164 18859 12206
rect 19017 12164 19067 12206
rect 19225 12164 19275 12206
rect 19438 12164 19488 12206
rect 11567 12031 11617 12073
rect 11780 12031 11830 12073
rect 11988 12031 12038 12073
rect 12196 12031 12246 12073
rect 19857 12160 19907 12202
rect 20065 12160 20115 12202
rect 20273 12160 20323 12202
rect 20486 12160 20536 12202
rect 14062 12026 14112 12068
rect 14275 12026 14325 12068
rect 14483 12026 14533 12068
rect 14691 12026 14741 12068
rect 6654 11403 6704 11445
rect 6862 11403 6912 11445
rect 7070 11403 7120 11445
rect 7283 11403 7333 11445
rect 859 11269 909 11311
rect 1072 11269 1122 11311
rect 1280 11269 1330 11311
rect 1488 11269 1538 11311
rect 9149 11398 9199 11440
rect 9357 11398 9407 11440
rect 9565 11398 9615 11440
rect 9778 11398 9828 11440
rect 1907 11265 1957 11307
rect 2120 11265 2170 11307
rect 2328 11265 2378 11307
rect 2536 11265 2586 11307
rect 17362 11397 17412 11439
rect 17570 11397 17620 11439
rect 17778 11397 17828 11439
rect 17991 11397 18041 11439
rect 11567 11263 11617 11305
rect 11780 11263 11830 11305
rect 11988 11263 12038 11305
rect 12196 11263 12246 11305
rect 19857 11392 19907 11434
rect 20065 11392 20115 11434
rect 20273 11392 20323 11434
rect 20486 11392 20536 11434
rect 12615 11259 12665 11301
rect 12828 11259 12878 11301
rect 13036 11259 13086 11301
rect 13244 11259 13294 11301
rect 8101 10723 8151 10765
rect 8309 10723 8359 10765
rect 8517 10723 8567 10765
rect 8730 10723 8780 10765
rect 859 10590 909 10632
rect 1072 10590 1122 10632
rect 1280 10590 1330 10632
rect 1488 10590 1538 10632
rect 9149 10719 9199 10761
rect 9357 10719 9407 10761
rect 9565 10719 9615 10761
rect 9778 10719 9828 10761
rect 3397 10587 3447 10629
rect 3610 10587 3660 10629
rect 3818 10587 3868 10629
rect 4026 10587 4076 10629
rect 18809 10717 18859 10759
rect 19017 10717 19067 10759
rect 19225 10717 19275 10759
rect 19438 10717 19488 10759
rect 11567 10584 11617 10626
rect 11780 10584 11830 10626
rect 11988 10584 12038 10626
rect 12196 10584 12246 10626
rect 19857 10713 19907 10755
rect 20065 10713 20115 10755
rect 20273 10713 20323 10755
rect 20486 10713 20536 10755
rect 14105 10581 14155 10623
rect 14318 10581 14368 10623
rect 14526 10581 14576 10623
rect 14734 10581 14784 10623
rect 6612 9881 6662 9923
rect 6820 9881 6870 9923
rect 7028 9881 7078 9923
rect 7241 9881 7291 9923
rect 860 9749 910 9791
rect 1073 9749 1123 9791
rect 1281 9749 1331 9791
rect 1489 9749 1539 9791
rect 9150 9878 9200 9920
rect 9358 9878 9408 9920
rect 9566 9878 9616 9920
rect 9779 9878 9829 9920
rect 1908 9745 1958 9787
rect 2121 9745 2171 9787
rect 2329 9745 2379 9787
rect 2537 9745 2587 9787
rect 17320 9875 17370 9917
rect 17528 9875 17578 9917
rect 17736 9875 17786 9917
rect 17949 9875 17999 9917
rect 11568 9743 11618 9785
rect 11781 9743 11831 9785
rect 11989 9743 12039 9785
rect 12197 9743 12247 9785
rect 19858 9872 19908 9914
rect 20066 9872 20116 9914
rect 20274 9872 20324 9914
rect 20487 9872 20537 9914
rect 12616 9739 12666 9781
rect 12829 9739 12879 9781
rect 13037 9739 13087 9781
rect 13245 9739 13295 9781
rect 8102 9203 8152 9245
rect 8310 9203 8360 9245
rect 8518 9203 8568 9245
rect 8731 9203 8781 9245
rect 860 9070 910 9112
rect 1073 9070 1123 9112
rect 1281 9070 1331 9112
rect 1489 9070 1539 9112
rect 9150 9199 9200 9241
rect 9358 9199 9408 9241
rect 9566 9199 9616 9241
rect 9779 9199 9829 9241
rect 3355 9065 3405 9107
rect 3568 9065 3618 9107
rect 3776 9065 3826 9107
rect 3984 9065 4034 9107
rect 18810 9197 18860 9239
rect 19018 9197 19068 9239
rect 19226 9197 19276 9239
rect 19439 9197 19489 9239
rect 11568 9064 11618 9106
rect 11781 9064 11831 9106
rect 11989 9064 12039 9106
rect 12197 9064 12247 9106
rect 19858 9193 19908 9235
rect 20066 9193 20116 9235
rect 20274 9193 20324 9235
rect 20487 9193 20537 9235
rect 14063 9059 14113 9101
rect 14276 9059 14326 9101
rect 14484 9059 14534 9101
rect 14692 9059 14742 9101
rect 6655 8436 6705 8478
rect 6863 8436 6913 8478
rect 7071 8436 7121 8478
rect 7284 8436 7334 8478
rect 860 8302 910 8344
rect 1073 8302 1123 8344
rect 1281 8302 1331 8344
rect 1489 8302 1539 8344
rect 9150 8431 9200 8473
rect 9358 8431 9408 8473
rect 9566 8431 9616 8473
rect 9779 8431 9829 8473
rect 1908 8298 1958 8340
rect 2121 8298 2171 8340
rect 2329 8298 2379 8340
rect 2537 8298 2587 8340
rect 17363 8430 17413 8472
rect 17571 8430 17621 8472
rect 17779 8430 17829 8472
rect 17992 8430 18042 8472
rect 11568 8296 11618 8338
rect 11781 8296 11831 8338
rect 11989 8296 12039 8338
rect 12197 8296 12247 8338
rect 19858 8425 19908 8467
rect 20066 8425 20116 8467
rect 20274 8425 20324 8467
rect 20487 8425 20537 8467
rect 12616 8292 12666 8334
rect 12829 8292 12879 8334
rect 13037 8292 13087 8334
rect 13245 8292 13295 8334
rect 8102 7756 8152 7798
rect 8310 7756 8360 7798
rect 8518 7756 8568 7798
rect 8731 7756 8781 7798
rect 860 7623 910 7665
rect 1073 7623 1123 7665
rect 1281 7623 1331 7665
rect 1489 7623 1539 7665
rect 9150 7752 9200 7794
rect 9358 7752 9408 7794
rect 9566 7752 9616 7794
rect 9779 7752 9829 7794
rect 4463 7614 4513 7656
rect 4676 7614 4726 7656
rect 4884 7614 4934 7656
rect 5092 7614 5142 7656
rect 18810 7750 18860 7792
rect 19018 7750 19068 7792
rect 19226 7750 19276 7792
rect 19439 7750 19489 7792
rect 11568 7617 11618 7659
rect 11781 7617 11831 7659
rect 11989 7617 12039 7659
rect 12197 7617 12247 7659
rect 19858 7746 19908 7788
rect 20066 7746 20116 7788
rect 20274 7746 20324 7788
rect 20487 7746 20537 7788
rect 15171 7608 15221 7650
rect 15384 7608 15434 7650
rect 15592 7608 15642 7650
rect 15800 7608 15850 7650
rect 5544 6846 5594 6888
rect 5752 6846 5802 6888
rect 5960 6846 6010 6888
rect 6173 6846 6223 6888
rect 857 6708 907 6750
rect 1070 6708 1120 6750
rect 1278 6708 1328 6750
rect 1486 6708 1536 6750
rect 9147 6837 9197 6879
rect 9355 6837 9405 6879
rect 9563 6837 9613 6879
rect 9776 6837 9826 6879
rect 1905 6704 1955 6746
rect 2118 6704 2168 6746
rect 2326 6704 2376 6746
rect 2534 6704 2584 6746
rect 16252 6840 16302 6882
rect 16460 6840 16510 6882
rect 16668 6840 16718 6882
rect 16881 6840 16931 6882
rect 11565 6702 11615 6744
rect 11778 6702 11828 6744
rect 11986 6702 12036 6744
rect 12194 6702 12244 6744
rect 19855 6831 19905 6873
rect 20063 6831 20113 6873
rect 20271 6831 20321 6873
rect 20484 6831 20534 6873
rect 12613 6698 12663 6740
rect 12826 6698 12876 6740
rect 13034 6698 13084 6740
rect 13242 6698 13292 6740
rect 8099 6162 8149 6204
rect 8307 6162 8357 6204
rect 8515 6162 8565 6204
rect 8728 6162 8778 6204
rect 857 6029 907 6071
rect 1070 6029 1120 6071
rect 1278 6029 1328 6071
rect 1486 6029 1536 6071
rect 9147 6158 9197 6200
rect 9355 6158 9405 6200
rect 9563 6158 9613 6200
rect 9776 6158 9826 6200
rect 3352 6024 3402 6066
rect 3565 6024 3615 6066
rect 3773 6024 3823 6066
rect 3981 6024 4031 6066
rect 18807 6156 18857 6198
rect 19015 6156 19065 6198
rect 19223 6156 19273 6198
rect 19436 6156 19486 6198
rect 11565 6023 11615 6065
rect 11778 6023 11828 6065
rect 11986 6023 12036 6065
rect 12194 6023 12244 6065
rect 19855 6152 19905 6194
rect 20063 6152 20113 6194
rect 20271 6152 20321 6194
rect 20484 6152 20534 6194
rect 14060 6018 14110 6060
rect 14273 6018 14323 6060
rect 14481 6018 14531 6060
rect 14689 6018 14739 6060
rect 6652 5395 6702 5437
rect 6860 5395 6910 5437
rect 7068 5395 7118 5437
rect 7281 5395 7331 5437
rect 857 5261 907 5303
rect 1070 5261 1120 5303
rect 1278 5261 1328 5303
rect 1486 5261 1536 5303
rect 9147 5390 9197 5432
rect 9355 5390 9405 5432
rect 9563 5390 9613 5432
rect 9776 5390 9826 5432
rect 1905 5257 1955 5299
rect 2118 5257 2168 5299
rect 2326 5257 2376 5299
rect 2534 5257 2584 5299
rect 17360 5389 17410 5431
rect 17568 5389 17618 5431
rect 17776 5389 17826 5431
rect 17989 5389 18039 5431
rect 11565 5255 11615 5297
rect 11778 5255 11828 5297
rect 11986 5255 12036 5297
rect 12194 5255 12244 5297
rect 19855 5384 19905 5426
rect 20063 5384 20113 5426
rect 20271 5384 20321 5426
rect 20484 5384 20534 5426
rect 12613 5251 12663 5293
rect 12826 5251 12876 5293
rect 13034 5251 13084 5293
rect 13242 5251 13292 5293
rect 8099 4715 8149 4757
rect 8307 4715 8357 4757
rect 8515 4715 8565 4757
rect 8728 4715 8778 4757
rect 857 4582 907 4624
rect 1070 4582 1120 4624
rect 1278 4582 1328 4624
rect 1486 4582 1536 4624
rect 9147 4711 9197 4753
rect 9355 4711 9405 4753
rect 9563 4711 9613 4753
rect 9776 4711 9826 4753
rect 3395 4579 3445 4621
rect 3608 4579 3658 4621
rect 3816 4579 3866 4621
rect 4024 4579 4074 4621
rect 18807 4709 18857 4751
rect 19015 4709 19065 4751
rect 19223 4709 19273 4751
rect 19436 4709 19486 4751
rect 11565 4576 11615 4618
rect 11778 4576 11828 4618
rect 11986 4576 12036 4618
rect 12194 4576 12244 4618
rect 19855 4705 19905 4747
rect 20063 4705 20113 4747
rect 20271 4705 20321 4747
rect 20484 4705 20534 4747
rect 14103 4573 14153 4615
rect 14316 4573 14366 4615
rect 14524 4573 14574 4615
rect 14732 4573 14782 4615
rect 6610 3873 6660 3915
rect 6818 3873 6868 3915
rect 7026 3873 7076 3915
rect 7239 3873 7289 3915
rect 858 3741 908 3783
rect 1071 3741 1121 3783
rect 1279 3741 1329 3783
rect 1487 3741 1537 3783
rect 9148 3870 9198 3912
rect 9356 3870 9406 3912
rect 9564 3870 9614 3912
rect 9777 3870 9827 3912
rect 1906 3737 1956 3779
rect 2119 3737 2169 3779
rect 2327 3737 2377 3779
rect 2535 3737 2585 3779
rect 4808 3743 4858 3785
rect 5021 3743 5071 3785
rect 5229 3743 5279 3785
rect 5437 3743 5487 3785
rect 17318 3867 17368 3909
rect 17526 3867 17576 3909
rect 17734 3867 17784 3909
rect 17947 3867 17997 3909
rect 11566 3735 11616 3777
rect 11779 3735 11829 3777
rect 11987 3735 12037 3777
rect 12195 3735 12245 3777
rect 19856 3864 19906 3906
rect 20064 3864 20114 3906
rect 20272 3864 20322 3906
rect 20485 3864 20535 3906
rect 12614 3731 12664 3773
rect 12827 3731 12877 3773
rect 13035 3731 13085 3773
rect 13243 3731 13293 3773
rect 15516 3737 15566 3779
rect 15729 3737 15779 3779
rect 15937 3737 15987 3779
rect 16145 3737 16195 3779
rect 8100 3195 8150 3237
rect 8308 3195 8358 3237
rect 8516 3195 8566 3237
rect 8729 3195 8779 3237
rect 858 3062 908 3104
rect 1071 3062 1121 3104
rect 1279 3062 1329 3104
rect 1487 3062 1537 3104
rect 9148 3191 9198 3233
rect 9356 3191 9406 3233
rect 9564 3191 9614 3233
rect 9777 3191 9827 3233
rect 3353 3057 3403 3099
rect 3566 3057 3616 3099
rect 3774 3057 3824 3099
rect 3982 3057 4032 3099
rect 18808 3189 18858 3231
rect 19016 3189 19066 3231
rect 19224 3189 19274 3231
rect 19437 3189 19487 3231
rect 11566 3056 11616 3098
rect 11779 3056 11829 3098
rect 11987 3056 12037 3098
rect 12195 3056 12245 3098
rect 19856 3185 19906 3227
rect 20064 3185 20114 3227
rect 20272 3185 20322 3227
rect 20485 3185 20535 3227
rect 14061 3051 14111 3093
rect 14274 3051 14324 3093
rect 14482 3051 14532 3093
rect 14690 3051 14740 3093
rect 6653 2428 6703 2470
rect 6861 2428 6911 2470
rect 7069 2428 7119 2470
rect 7282 2428 7332 2470
rect 858 2294 908 2336
rect 1071 2294 1121 2336
rect 1279 2294 1329 2336
rect 1487 2294 1537 2336
rect 9148 2423 9198 2465
rect 9356 2423 9406 2465
rect 9564 2423 9614 2465
rect 9777 2423 9827 2465
rect 1906 2290 1956 2332
rect 2119 2290 2169 2332
rect 2327 2290 2377 2332
rect 2535 2290 2585 2332
rect 17361 2422 17411 2464
rect 17569 2422 17619 2464
rect 17777 2422 17827 2464
rect 17990 2422 18040 2464
rect 11566 2288 11616 2330
rect 11779 2288 11829 2330
rect 11987 2288 12037 2330
rect 12195 2288 12245 2330
rect 19856 2417 19906 2459
rect 20064 2417 20114 2459
rect 20272 2417 20322 2459
rect 20485 2417 20535 2459
rect 12614 2284 12664 2326
rect 12827 2284 12877 2326
rect 13035 2284 13085 2326
rect 13243 2284 13293 2326
rect 8100 1748 8150 1790
rect 8308 1748 8358 1790
rect 8516 1748 8566 1790
rect 8729 1748 8779 1790
rect 9148 1744 9198 1786
rect 9356 1744 9406 1786
rect 9564 1744 9614 1786
rect 9777 1744 9827 1786
rect 858 1615 908 1657
rect 1071 1615 1121 1657
rect 1279 1615 1329 1657
rect 1487 1615 1537 1657
rect 18808 1742 18858 1784
rect 19016 1742 19066 1784
rect 19224 1742 19274 1784
rect 19437 1742 19487 1784
rect 19856 1738 19906 1780
rect 20064 1738 20114 1780
rect 20272 1738 20322 1780
rect 20485 1738 20535 1780
rect 11566 1609 11616 1651
rect 11779 1609 11829 1651
rect 11987 1609 12037 1651
rect 12195 1609 12245 1651
rect 10569 -544 10619 -502
rect 10782 -544 10832 -502
rect 10990 -544 11040 -502
rect 11198 -544 11248 -502
<< pmos >>
rect 859 12835 909 12935
rect 1072 12835 1122 12935
rect 1280 12835 1330 12935
rect 1488 12835 1538 12935
rect 1907 12831 1957 12931
rect 2120 12831 2170 12931
rect 2328 12831 2378 12931
rect 2536 12831 2586 12931
rect 11567 12829 11617 12929
rect 11780 12829 11830 12929
rect 11988 12829 12038 12929
rect 12196 12829 12246 12929
rect 9149 12668 9199 12768
rect 9357 12668 9407 12768
rect 9565 12668 9615 12768
rect 9778 12668 9828 12768
rect 12615 12825 12665 12925
rect 12828 12825 12878 12925
rect 13036 12825 13086 12925
rect 13244 12825 13294 12925
rect 19857 12662 19907 12762
rect 20065 12662 20115 12762
rect 20273 12662 20323 12762
rect 20486 12662 20536 12762
rect 859 12156 909 12256
rect 1072 12156 1122 12256
rect 1280 12156 1330 12256
rect 1488 12156 1538 12256
rect 3354 12151 3404 12251
rect 3567 12151 3617 12251
rect 3775 12151 3825 12251
rect 3983 12151 4033 12251
rect 8101 11993 8151 12093
rect 8309 11993 8359 12093
rect 8517 11993 8567 12093
rect 8730 11993 8780 12093
rect 11567 12150 11617 12250
rect 11780 12150 11830 12250
rect 11988 12150 12038 12250
rect 12196 12150 12246 12250
rect 9149 11989 9199 12089
rect 9357 11989 9407 12089
rect 9565 11989 9615 12089
rect 9778 11989 9828 12089
rect 14062 12145 14112 12245
rect 14275 12145 14325 12245
rect 14483 12145 14533 12245
rect 14691 12145 14741 12245
rect 18809 11987 18859 12087
rect 19017 11987 19067 12087
rect 19225 11987 19275 12087
rect 19438 11987 19488 12087
rect 19857 11983 19907 12083
rect 20065 11983 20115 12083
rect 20273 11983 20323 12083
rect 20486 11983 20536 12083
rect 859 11388 909 11488
rect 1072 11388 1122 11488
rect 1280 11388 1330 11488
rect 1488 11388 1538 11488
rect 1907 11384 1957 11484
rect 2120 11384 2170 11484
rect 2328 11384 2378 11484
rect 2536 11384 2586 11484
rect 6654 11226 6704 11326
rect 6862 11226 6912 11326
rect 7070 11226 7120 11326
rect 7283 11226 7333 11326
rect 11567 11382 11617 11482
rect 11780 11382 11830 11482
rect 11988 11382 12038 11482
rect 12196 11382 12246 11482
rect 9149 11221 9199 11321
rect 9357 11221 9407 11321
rect 9565 11221 9615 11321
rect 9778 11221 9828 11321
rect 12615 11378 12665 11478
rect 12828 11378 12878 11478
rect 13036 11378 13086 11478
rect 13244 11378 13294 11478
rect 17362 11220 17412 11320
rect 17570 11220 17620 11320
rect 17778 11220 17828 11320
rect 17991 11220 18041 11320
rect 19857 11215 19907 11315
rect 20065 11215 20115 11315
rect 20273 11215 20323 11315
rect 20486 11215 20536 11315
rect 859 10709 909 10809
rect 1072 10709 1122 10809
rect 1280 10709 1330 10809
rect 1488 10709 1538 10809
rect 3397 10706 3447 10806
rect 3610 10706 3660 10806
rect 3818 10706 3868 10806
rect 4026 10706 4076 10806
rect 8101 10546 8151 10646
rect 8309 10546 8359 10646
rect 8517 10546 8567 10646
rect 8730 10546 8780 10646
rect 11567 10703 11617 10803
rect 11780 10703 11830 10803
rect 11988 10703 12038 10803
rect 12196 10703 12246 10803
rect 9149 10542 9199 10642
rect 9357 10542 9407 10642
rect 9565 10542 9615 10642
rect 9778 10542 9828 10642
rect 14105 10700 14155 10800
rect 14318 10700 14368 10800
rect 14526 10700 14576 10800
rect 14734 10700 14784 10800
rect 18809 10540 18859 10640
rect 19017 10540 19067 10640
rect 19225 10540 19275 10640
rect 19438 10540 19488 10640
rect 19857 10536 19907 10636
rect 20065 10536 20115 10636
rect 20273 10536 20323 10636
rect 20486 10536 20536 10636
rect 860 9868 910 9968
rect 1073 9868 1123 9968
rect 1281 9868 1331 9968
rect 1489 9868 1539 9968
rect 1908 9864 1958 9964
rect 2121 9864 2171 9964
rect 2329 9864 2379 9964
rect 2537 9864 2587 9964
rect 6612 9704 6662 9804
rect 6820 9704 6870 9804
rect 7028 9704 7078 9804
rect 7241 9704 7291 9804
rect 11568 9862 11618 9962
rect 11781 9862 11831 9962
rect 11989 9862 12039 9962
rect 12197 9862 12247 9962
rect 9150 9701 9200 9801
rect 9358 9701 9408 9801
rect 9566 9701 9616 9801
rect 9779 9701 9829 9801
rect 12616 9858 12666 9958
rect 12829 9858 12879 9958
rect 13037 9858 13087 9958
rect 13245 9858 13295 9958
rect 17320 9698 17370 9798
rect 17528 9698 17578 9798
rect 17736 9698 17786 9798
rect 17949 9698 17999 9798
rect 19858 9695 19908 9795
rect 20066 9695 20116 9795
rect 20274 9695 20324 9795
rect 20487 9695 20537 9795
rect 860 9189 910 9289
rect 1073 9189 1123 9289
rect 1281 9189 1331 9289
rect 1489 9189 1539 9289
rect 3355 9184 3405 9284
rect 3568 9184 3618 9284
rect 3776 9184 3826 9284
rect 3984 9184 4034 9284
rect 8102 9026 8152 9126
rect 8310 9026 8360 9126
rect 8518 9026 8568 9126
rect 8731 9026 8781 9126
rect 11568 9183 11618 9283
rect 11781 9183 11831 9283
rect 11989 9183 12039 9283
rect 12197 9183 12247 9283
rect 9150 9022 9200 9122
rect 9358 9022 9408 9122
rect 9566 9022 9616 9122
rect 9779 9022 9829 9122
rect 14063 9178 14113 9278
rect 14276 9178 14326 9278
rect 14484 9178 14534 9278
rect 14692 9178 14742 9278
rect 18810 9020 18860 9120
rect 19018 9020 19068 9120
rect 19226 9020 19276 9120
rect 19439 9020 19489 9120
rect 19858 9016 19908 9116
rect 20066 9016 20116 9116
rect 20274 9016 20324 9116
rect 20487 9016 20537 9116
rect 860 8421 910 8521
rect 1073 8421 1123 8521
rect 1281 8421 1331 8521
rect 1489 8421 1539 8521
rect 1908 8417 1958 8517
rect 2121 8417 2171 8517
rect 2329 8417 2379 8517
rect 2537 8417 2587 8517
rect 6655 8259 6705 8359
rect 6863 8259 6913 8359
rect 7071 8259 7121 8359
rect 7284 8259 7334 8359
rect 11568 8415 11618 8515
rect 11781 8415 11831 8515
rect 11989 8415 12039 8515
rect 12197 8415 12247 8515
rect 9150 8254 9200 8354
rect 9358 8254 9408 8354
rect 9566 8254 9616 8354
rect 9779 8254 9829 8354
rect 12616 8411 12666 8511
rect 12829 8411 12879 8511
rect 13037 8411 13087 8511
rect 13245 8411 13295 8511
rect 17363 8253 17413 8353
rect 17571 8253 17621 8353
rect 17779 8253 17829 8353
rect 17992 8253 18042 8353
rect 19858 8248 19908 8348
rect 20066 8248 20116 8348
rect 20274 8248 20324 8348
rect 20487 8248 20537 8348
rect 860 7742 910 7842
rect 1073 7742 1123 7842
rect 1281 7742 1331 7842
rect 1489 7742 1539 7842
rect 4463 7733 4513 7833
rect 4676 7733 4726 7833
rect 4884 7733 4934 7833
rect 5092 7733 5142 7833
rect 8102 7579 8152 7679
rect 8310 7579 8360 7679
rect 8518 7579 8568 7679
rect 8731 7579 8781 7679
rect 11568 7736 11618 7836
rect 11781 7736 11831 7836
rect 11989 7736 12039 7836
rect 12197 7736 12247 7836
rect 9150 7575 9200 7675
rect 9358 7575 9408 7675
rect 9566 7575 9616 7675
rect 9779 7575 9829 7675
rect 15171 7727 15221 7827
rect 15384 7727 15434 7827
rect 15592 7727 15642 7827
rect 15800 7727 15850 7827
rect 18810 7573 18860 7673
rect 19018 7573 19068 7673
rect 19226 7573 19276 7673
rect 19439 7573 19489 7673
rect 19858 7569 19908 7669
rect 20066 7569 20116 7669
rect 20274 7569 20324 7669
rect 20487 7569 20537 7669
rect 857 6827 907 6927
rect 1070 6827 1120 6927
rect 1278 6827 1328 6927
rect 1486 6827 1536 6927
rect 1905 6823 1955 6923
rect 2118 6823 2168 6923
rect 2326 6823 2376 6923
rect 2534 6823 2584 6923
rect 5544 6669 5594 6769
rect 5752 6669 5802 6769
rect 5960 6669 6010 6769
rect 6173 6669 6223 6769
rect 11565 6821 11615 6921
rect 11778 6821 11828 6921
rect 11986 6821 12036 6921
rect 12194 6821 12244 6921
rect 9147 6660 9197 6760
rect 9355 6660 9405 6760
rect 9563 6660 9613 6760
rect 9776 6660 9826 6760
rect 12613 6817 12663 6917
rect 12826 6817 12876 6917
rect 13034 6817 13084 6917
rect 13242 6817 13292 6917
rect 16252 6663 16302 6763
rect 16460 6663 16510 6763
rect 16668 6663 16718 6763
rect 16881 6663 16931 6763
rect 19855 6654 19905 6754
rect 20063 6654 20113 6754
rect 20271 6654 20321 6754
rect 20484 6654 20534 6754
rect 857 6148 907 6248
rect 1070 6148 1120 6248
rect 1278 6148 1328 6248
rect 1486 6148 1536 6248
rect 3352 6143 3402 6243
rect 3565 6143 3615 6243
rect 3773 6143 3823 6243
rect 3981 6143 4031 6243
rect 8099 5985 8149 6085
rect 8307 5985 8357 6085
rect 8515 5985 8565 6085
rect 8728 5985 8778 6085
rect 11565 6142 11615 6242
rect 11778 6142 11828 6242
rect 11986 6142 12036 6242
rect 12194 6142 12244 6242
rect 9147 5981 9197 6081
rect 9355 5981 9405 6081
rect 9563 5981 9613 6081
rect 9776 5981 9826 6081
rect 14060 6137 14110 6237
rect 14273 6137 14323 6237
rect 14481 6137 14531 6237
rect 14689 6137 14739 6237
rect 18807 5979 18857 6079
rect 19015 5979 19065 6079
rect 19223 5979 19273 6079
rect 19436 5979 19486 6079
rect 19855 5975 19905 6075
rect 20063 5975 20113 6075
rect 20271 5975 20321 6075
rect 20484 5975 20534 6075
rect 857 5380 907 5480
rect 1070 5380 1120 5480
rect 1278 5380 1328 5480
rect 1486 5380 1536 5480
rect 1905 5376 1955 5476
rect 2118 5376 2168 5476
rect 2326 5376 2376 5476
rect 2534 5376 2584 5476
rect 6652 5218 6702 5318
rect 6860 5218 6910 5318
rect 7068 5218 7118 5318
rect 7281 5218 7331 5318
rect 11565 5374 11615 5474
rect 11778 5374 11828 5474
rect 11986 5374 12036 5474
rect 12194 5374 12244 5474
rect 9147 5213 9197 5313
rect 9355 5213 9405 5313
rect 9563 5213 9613 5313
rect 9776 5213 9826 5313
rect 12613 5370 12663 5470
rect 12826 5370 12876 5470
rect 13034 5370 13084 5470
rect 13242 5370 13292 5470
rect 17360 5212 17410 5312
rect 17568 5212 17618 5312
rect 17776 5212 17826 5312
rect 17989 5212 18039 5312
rect 19855 5207 19905 5307
rect 20063 5207 20113 5307
rect 20271 5207 20321 5307
rect 20484 5207 20534 5307
rect 857 4701 907 4801
rect 1070 4701 1120 4801
rect 1278 4701 1328 4801
rect 1486 4701 1536 4801
rect 3395 4698 3445 4798
rect 3608 4698 3658 4798
rect 3816 4698 3866 4798
rect 4024 4698 4074 4798
rect 8099 4538 8149 4638
rect 8307 4538 8357 4638
rect 8515 4538 8565 4638
rect 8728 4538 8778 4638
rect 11565 4695 11615 4795
rect 11778 4695 11828 4795
rect 11986 4695 12036 4795
rect 12194 4695 12244 4795
rect 9147 4534 9197 4634
rect 9355 4534 9405 4634
rect 9563 4534 9613 4634
rect 9776 4534 9826 4634
rect 14103 4692 14153 4792
rect 14316 4692 14366 4792
rect 14524 4692 14574 4792
rect 14732 4692 14782 4792
rect 18807 4532 18857 4632
rect 19015 4532 19065 4632
rect 19223 4532 19273 4632
rect 19436 4532 19486 4632
rect 19855 4528 19905 4628
rect 20063 4528 20113 4628
rect 20271 4528 20321 4628
rect 20484 4528 20534 4628
rect 858 3860 908 3960
rect 1071 3860 1121 3960
rect 1279 3860 1329 3960
rect 1487 3860 1537 3960
rect 1906 3856 1956 3956
rect 2119 3856 2169 3956
rect 2327 3856 2377 3956
rect 2535 3856 2585 3956
rect 4808 3862 4858 3962
rect 5021 3862 5071 3962
rect 5229 3862 5279 3962
rect 5437 3862 5487 3962
rect 6610 3696 6660 3796
rect 6818 3696 6868 3796
rect 7026 3696 7076 3796
rect 7239 3696 7289 3796
rect 11566 3854 11616 3954
rect 11779 3854 11829 3954
rect 11987 3854 12037 3954
rect 12195 3854 12245 3954
rect 9148 3693 9198 3793
rect 9356 3693 9406 3793
rect 9564 3693 9614 3793
rect 9777 3693 9827 3793
rect 12614 3850 12664 3950
rect 12827 3850 12877 3950
rect 13035 3850 13085 3950
rect 13243 3850 13293 3950
rect 15516 3856 15566 3956
rect 15729 3856 15779 3956
rect 15937 3856 15987 3956
rect 16145 3856 16195 3956
rect 17318 3690 17368 3790
rect 17526 3690 17576 3790
rect 17734 3690 17784 3790
rect 17947 3690 17997 3790
rect 19856 3687 19906 3787
rect 20064 3687 20114 3787
rect 20272 3687 20322 3787
rect 20485 3687 20535 3787
rect 858 3181 908 3281
rect 1071 3181 1121 3281
rect 1279 3181 1329 3281
rect 1487 3181 1537 3281
rect 3353 3176 3403 3276
rect 3566 3176 3616 3276
rect 3774 3176 3824 3276
rect 3982 3176 4032 3276
rect 8100 3018 8150 3118
rect 8308 3018 8358 3118
rect 8516 3018 8566 3118
rect 8729 3018 8779 3118
rect 11566 3175 11616 3275
rect 11779 3175 11829 3275
rect 11987 3175 12037 3275
rect 12195 3175 12245 3275
rect 9148 3014 9198 3114
rect 9356 3014 9406 3114
rect 9564 3014 9614 3114
rect 9777 3014 9827 3114
rect 14061 3170 14111 3270
rect 14274 3170 14324 3270
rect 14482 3170 14532 3270
rect 14690 3170 14740 3270
rect 18808 3012 18858 3112
rect 19016 3012 19066 3112
rect 19224 3012 19274 3112
rect 19437 3012 19487 3112
rect 19856 3008 19906 3108
rect 20064 3008 20114 3108
rect 20272 3008 20322 3108
rect 20485 3008 20535 3108
rect 858 2413 908 2513
rect 1071 2413 1121 2513
rect 1279 2413 1329 2513
rect 1487 2413 1537 2513
rect 1906 2409 1956 2509
rect 2119 2409 2169 2509
rect 2327 2409 2377 2509
rect 2535 2409 2585 2509
rect 6653 2251 6703 2351
rect 6861 2251 6911 2351
rect 7069 2251 7119 2351
rect 7282 2251 7332 2351
rect 11566 2407 11616 2507
rect 11779 2407 11829 2507
rect 11987 2407 12037 2507
rect 12195 2407 12245 2507
rect 9148 2246 9198 2346
rect 9356 2246 9406 2346
rect 9564 2246 9614 2346
rect 9777 2246 9827 2346
rect 12614 2403 12664 2503
rect 12827 2403 12877 2503
rect 13035 2403 13085 2503
rect 13243 2403 13293 2503
rect 17361 2245 17411 2345
rect 17569 2245 17619 2345
rect 17777 2245 17827 2345
rect 17990 2245 18040 2345
rect 19856 2240 19906 2340
rect 20064 2240 20114 2340
rect 20272 2240 20322 2340
rect 20485 2240 20535 2340
rect 858 1734 908 1834
rect 1071 1734 1121 1834
rect 1279 1734 1329 1834
rect 1487 1734 1537 1834
rect 8100 1571 8150 1671
rect 8308 1571 8358 1671
rect 8516 1571 8566 1671
rect 8729 1571 8779 1671
rect 11566 1728 11616 1828
rect 11779 1728 11829 1828
rect 11987 1728 12037 1828
rect 12195 1728 12245 1828
rect 9148 1567 9198 1667
rect 9356 1567 9406 1667
rect 9564 1567 9614 1667
rect 9777 1567 9827 1667
rect 18808 1565 18858 1665
rect 19016 1565 19066 1665
rect 19224 1565 19274 1665
rect 19437 1565 19487 1665
rect 19856 1561 19906 1661
rect 20064 1561 20114 1661
rect 20272 1561 20322 1661
rect 20485 1561 20535 1661
rect 10569 -425 10619 -325
rect 10782 -425 10832 -325
rect 10990 -425 11040 -325
rect 11198 -425 11248 -325
<< ndiff >>
rect 9100 12875 9149 12887
rect 9100 12855 9111 12875
rect 9131 12855 9149 12875
rect 9100 12845 9149 12855
rect 9199 12871 9243 12887
rect 9199 12851 9214 12871
rect 9234 12851 9243 12871
rect 9199 12845 9243 12851
rect 9313 12871 9357 12887
rect 9313 12851 9322 12871
rect 9342 12851 9357 12871
rect 9313 12845 9357 12851
rect 9407 12875 9456 12887
rect 9407 12855 9425 12875
rect 9445 12855 9456 12875
rect 9407 12845 9456 12855
rect 9521 12871 9565 12887
rect 9521 12851 9530 12871
rect 9550 12851 9565 12871
rect 9521 12845 9565 12851
rect 9615 12875 9664 12887
rect 9615 12855 9633 12875
rect 9653 12855 9664 12875
rect 9615 12845 9664 12855
rect 9734 12871 9778 12887
rect 9734 12851 9743 12871
rect 9763 12851 9778 12871
rect 9734 12845 9778 12851
rect 9828 12875 9877 12887
rect 9828 12855 9846 12875
rect 9866 12855 9877 12875
rect 9828 12845 9877 12855
rect 810 12748 859 12758
rect 810 12728 821 12748
rect 841 12728 859 12748
rect 810 12716 859 12728
rect 909 12752 953 12758
rect 909 12732 924 12752
rect 944 12732 953 12752
rect 909 12716 953 12732
rect 1023 12748 1072 12758
rect 1023 12728 1034 12748
rect 1054 12728 1072 12748
rect 1023 12716 1072 12728
rect 1122 12752 1166 12758
rect 1122 12732 1137 12752
rect 1157 12732 1166 12752
rect 1122 12716 1166 12732
rect 1231 12748 1280 12758
rect 1231 12728 1242 12748
rect 1262 12728 1280 12748
rect 1231 12716 1280 12728
rect 1330 12752 1374 12758
rect 1330 12732 1345 12752
rect 1365 12732 1374 12752
rect 1330 12716 1374 12732
rect 1444 12752 1488 12758
rect 1444 12732 1453 12752
rect 1473 12732 1488 12752
rect 1444 12716 1488 12732
rect 1538 12748 1587 12758
rect 1538 12728 1556 12748
rect 1576 12728 1587 12748
rect 1538 12716 1587 12728
rect 1858 12744 1907 12754
rect 1858 12724 1869 12744
rect 1889 12724 1907 12744
rect 1858 12712 1907 12724
rect 1957 12748 2001 12754
rect 1957 12728 1972 12748
rect 1992 12728 2001 12748
rect 1957 12712 2001 12728
rect 2071 12744 2120 12754
rect 2071 12724 2082 12744
rect 2102 12724 2120 12744
rect 2071 12712 2120 12724
rect 2170 12748 2214 12754
rect 2170 12728 2185 12748
rect 2205 12728 2214 12748
rect 2170 12712 2214 12728
rect 2279 12744 2328 12754
rect 2279 12724 2290 12744
rect 2310 12724 2328 12744
rect 2279 12712 2328 12724
rect 2378 12748 2422 12754
rect 2378 12728 2393 12748
rect 2413 12728 2422 12748
rect 2378 12712 2422 12728
rect 2492 12748 2536 12754
rect 2492 12728 2501 12748
rect 2521 12728 2536 12748
rect 2492 12712 2536 12728
rect 2586 12744 2635 12754
rect 2586 12724 2604 12744
rect 2624 12724 2635 12744
rect 2586 12712 2635 12724
rect 19808 12869 19857 12881
rect 19808 12849 19819 12869
rect 19839 12849 19857 12869
rect 19808 12839 19857 12849
rect 19907 12865 19951 12881
rect 19907 12845 19922 12865
rect 19942 12845 19951 12865
rect 19907 12839 19951 12845
rect 20021 12865 20065 12881
rect 20021 12845 20030 12865
rect 20050 12845 20065 12865
rect 20021 12839 20065 12845
rect 20115 12869 20164 12881
rect 20115 12849 20133 12869
rect 20153 12849 20164 12869
rect 20115 12839 20164 12849
rect 20229 12865 20273 12881
rect 20229 12845 20238 12865
rect 20258 12845 20273 12865
rect 20229 12839 20273 12845
rect 20323 12869 20372 12881
rect 20323 12849 20341 12869
rect 20361 12849 20372 12869
rect 20323 12839 20372 12849
rect 20442 12865 20486 12881
rect 20442 12845 20451 12865
rect 20471 12845 20486 12865
rect 20442 12839 20486 12845
rect 20536 12869 20585 12881
rect 20536 12849 20554 12869
rect 20574 12849 20585 12869
rect 20536 12839 20585 12849
rect 11518 12742 11567 12752
rect 11518 12722 11529 12742
rect 11549 12722 11567 12742
rect 11518 12710 11567 12722
rect 11617 12746 11661 12752
rect 11617 12726 11632 12746
rect 11652 12726 11661 12746
rect 11617 12710 11661 12726
rect 11731 12742 11780 12752
rect 11731 12722 11742 12742
rect 11762 12722 11780 12742
rect 11731 12710 11780 12722
rect 11830 12746 11874 12752
rect 11830 12726 11845 12746
rect 11865 12726 11874 12746
rect 11830 12710 11874 12726
rect 11939 12742 11988 12752
rect 11939 12722 11950 12742
rect 11970 12722 11988 12742
rect 11939 12710 11988 12722
rect 12038 12746 12082 12752
rect 12038 12726 12053 12746
rect 12073 12726 12082 12746
rect 12038 12710 12082 12726
rect 12152 12746 12196 12752
rect 12152 12726 12161 12746
rect 12181 12726 12196 12746
rect 12152 12710 12196 12726
rect 12246 12742 12295 12752
rect 12246 12722 12264 12742
rect 12284 12722 12295 12742
rect 12246 12710 12295 12722
rect 12566 12738 12615 12748
rect 12566 12718 12577 12738
rect 12597 12718 12615 12738
rect 12566 12706 12615 12718
rect 12665 12742 12709 12748
rect 12665 12722 12680 12742
rect 12700 12722 12709 12742
rect 12665 12706 12709 12722
rect 12779 12738 12828 12748
rect 12779 12718 12790 12738
rect 12810 12718 12828 12738
rect 12779 12706 12828 12718
rect 12878 12742 12922 12748
rect 12878 12722 12893 12742
rect 12913 12722 12922 12742
rect 12878 12706 12922 12722
rect 12987 12738 13036 12748
rect 12987 12718 12998 12738
rect 13018 12718 13036 12738
rect 12987 12706 13036 12718
rect 13086 12742 13130 12748
rect 13086 12722 13101 12742
rect 13121 12722 13130 12742
rect 13086 12706 13130 12722
rect 13200 12742 13244 12748
rect 13200 12722 13209 12742
rect 13229 12722 13244 12742
rect 13200 12706 13244 12722
rect 13294 12738 13343 12748
rect 13294 12718 13312 12738
rect 13332 12718 13343 12738
rect 13294 12706 13343 12718
rect 8052 12200 8101 12212
rect 8052 12180 8063 12200
rect 8083 12180 8101 12200
rect 8052 12170 8101 12180
rect 8151 12196 8195 12212
rect 8151 12176 8166 12196
rect 8186 12176 8195 12196
rect 8151 12170 8195 12176
rect 8265 12196 8309 12212
rect 8265 12176 8274 12196
rect 8294 12176 8309 12196
rect 8265 12170 8309 12176
rect 8359 12200 8408 12212
rect 8359 12180 8377 12200
rect 8397 12180 8408 12200
rect 8359 12170 8408 12180
rect 8473 12196 8517 12212
rect 8473 12176 8482 12196
rect 8502 12176 8517 12196
rect 8473 12170 8517 12176
rect 8567 12200 8616 12212
rect 8567 12180 8585 12200
rect 8605 12180 8616 12200
rect 8567 12170 8616 12180
rect 8686 12196 8730 12212
rect 8686 12176 8695 12196
rect 8715 12176 8730 12196
rect 8686 12170 8730 12176
rect 8780 12200 8829 12212
rect 8780 12180 8798 12200
rect 8818 12180 8829 12200
rect 8780 12170 8829 12180
rect 9100 12196 9149 12208
rect 9100 12176 9111 12196
rect 9131 12176 9149 12196
rect 810 12069 859 12079
rect 810 12049 821 12069
rect 841 12049 859 12069
rect 810 12037 859 12049
rect 909 12073 953 12079
rect 909 12053 924 12073
rect 944 12053 953 12073
rect 909 12037 953 12053
rect 1023 12069 1072 12079
rect 1023 12049 1034 12069
rect 1054 12049 1072 12069
rect 1023 12037 1072 12049
rect 1122 12073 1166 12079
rect 1122 12053 1137 12073
rect 1157 12053 1166 12073
rect 1122 12037 1166 12053
rect 1231 12069 1280 12079
rect 1231 12049 1242 12069
rect 1262 12049 1280 12069
rect 1231 12037 1280 12049
rect 1330 12073 1374 12079
rect 1330 12053 1345 12073
rect 1365 12053 1374 12073
rect 1330 12037 1374 12053
rect 1444 12073 1488 12079
rect 1444 12053 1453 12073
rect 1473 12053 1488 12073
rect 1444 12037 1488 12053
rect 1538 12069 1587 12079
rect 9100 12166 9149 12176
rect 9199 12192 9243 12208
rect 9199 12172 9214 12192
rect 9234 12172 9243 12192
rect 9199 12166 9243 12172
rect 9313 12192 9357 12208
rect 9313 12172 9322 12192
rect 9342 12172 9357 12192
rect 9313 12166 9357 12172
rect 9407 12196 9456 12208
rect 9407 12176 9425 12196
rect 9445 12176 9456 12196
rect 9407 12166 9456 12176
rect 9521 12192 9565 12208
rect 9521 12172 9530 12192
rect 9550 12172 9565 12192
rect 9521 12166 9565 12172
rect 9615 12196 9664 12208
rect 9615 12176 9633 12196
rect 9653 12176 9664 12196
rect 9615 12166 9664 12176
rect 9734 12192 9778 12208
rect 9734 12172 9743 12192
rect 9763 12172 9778 12192
rect 9734 12166 9778 12172
rect 9828 12196 9877 12208
rect 9828 12176 9846 12196
rect 9866 12176 9877 12196
rect 9828 12166 9877 12176
rect 1538 12049 1556 12069
rect 1576 12049 1587 12069
rect 1538 12037 1587 12049
rect 3305 12064 3354 12074
rect 3305 12044 3316 12064
rect 3336 12044 3354 12064
rect 3305 12032 3354 12044
rect 3404 12068 3448 12074
rect 3404 12048 3419 12068
rect 3439 12048 3448 12068
rect 3404 12032 3448 12048
rect 3518 12064 3567 12074
rect 3518 12044 3529 12064
rect 3549 12044 3567 12064
rect 3518 12032 3567 12044
rect 3617 12068 3661 12074
rect 3617 12048 3632 12068
rect 3652 12048 3661 12068
rect 3617 12032 3661 12048
rect 3726 12064 3775 12074
rect 3726 12044 3737 12064
rect 3757 12044 3775 12064
rect 3726 12032 3775 12044
rect 3825 12068 3869 12074
rect 3825 12048 3840 12068
rect 3860 12048 3869 12068
rect 3825 12032 3869 12048
rect 3939 12068 3983 12074
rect 3939 12048 3948 12068
rect 3968 12048 3983 12068
rect 3939 12032 3983 12048
rect 4033 12064 4082 12074
rect 4033 12044 4051 12064
rect 4071 12044 4082 12064
rect 4033 12032 4082 12044
rect 18760 12194 18809 12206
rect 18760 12174 18771 12194
rect 18791 12174 18809 12194
rect 18760 12164 18809 12174
rect 18859 12190 18903 12206
rect 18859 12170 18874 12190
rect 18894 12170 18903 12190
rect 18859 12164 18903 12170
rect 18973 12190 19017 12206
rect 18973 12170 18982 12190
rect 19002 12170 19017 12190
rect 18973 12164 19017 12170
rect 19067 12194 19116 12206
rect 19067 12174 19085 12194
rect 19105 12174 19116 12194
rect 19067 12164 19116 12174
rect 19181 12190 19225 12206
rect 19181 12170 19190 12190
rect 19210 12170 19225 12190
rect 19181 12164 19225 12170
rect 19275 12194 19324 12206
rect 19275 12174 19293 12194
rect 19313 12174 19324 12194
rect 19275 12164 19324 12174
rect 19394 12190 19438 12206
rect 19394 12170 19403 12190
rect 19423 12170 19438 12190
rect 19394 12164 19438 12170
rect 19488 12194 19537 12206
rect 19488 12174 19506 12194
rect 19526 12174 19537 12194
rect 19488 12164 19537 12174
rect 19808 12190 19857 12202
rect 19808 12170 19819 12190
rect 19839 12170 19857 12190
rect 11518 12063 11567 12073
rect 11518 12043 11529 12063
rect 11549 12043 11567 12063
rect 11518 12031 11567 12043
rect 11617 12067 11661 12073
rect 11617 12047 11632 12067
rect 11652 12047 11661 12067
rect 11617 12031 11661 12047
rect 11731 12063 11780 12073
rect 11731 12043 11742 12063
rect 11762 12043 11780 12063
rect 11731 12031 11780 12043
rect 11830 12067 11874 12073
rect 11830 12047 11845 12067
rect 11865 12047 11874 12067
rect 11830 12031 11874 12047
rect 11939 12063 11988 12073
rect 11939 12043 11950 12063
rect 11970 12043 11988 12063
rect 11939 12031 11988 12043
rect 12038 12067 12082 12073
rect 12038 12047 12053 12067
rect 12073 12047 12082 12067
rect 12038 12031 12082 12047
rect 12152 12067 12196 12073
rect 12152 12047 12161 12067
rect 12181 12047 12196 12067
rect 12152 12031 12196 12047
rect 12246 12063 12295 12073
rect 19808 12160 19857 12170
rect 19907 12186 19951 12202
rect 19907 12166 19922 12186
rect 19942 12166 19951 12186
rect 19907 12160 19951 12166
rect 20021 12186 20065 12202
rect 20021 12166 20030 12186
rect 20050 12166 20065 12186
rect 20021 12160 20065 12166
rect 20115 12190 20164 12202
rect 20115 12170 20133 12190
rect 20153 12170 20164 12190
rect 20115 12160 20164 12170
rect 20229 12186 20273 12202
rect 20229 12166 20238 12186
rect 20258 12166 20273 12186
rect 20229 12160 20273 12166
rect 20323 12190 20372 12202
rect 20323 12170 20341 12190
rect 20361 12170 20372 12190
rect 20323 12160 20372 12170
rect 20442 12186 20486 12202
rect 20442 12166 20451 12186
rect 20471 12166 20486 12186
rect 20442 12160 20486 12166
rect 20536 12190 20585 12202
rect 20536 12170 20554 12190
rect 20574 12170 20585 12190
rect 20536 12160 20585 12170
rect 12246 12043 12264 12063
rect 12284 12043 12295 12063
rect 12246 12031 12295 12043
rect 14013 12058 14062 12068
rect 14013 12038 14024 12058
rect 14044 12038 14062 12058
rect 14013 12026 14062 12038
rect 14112 12062 14156 12068
rect 14112 12042 14127 12062
rect 14147 12042 14156 12062
rect 14112 12026 14156 12042
rect 14226 12058 14275 12068
rect 14226 12038 14237 12058
rect 14257 12038 14275 12058
rect 14226 12026 14275 12038
rect 14325 12062 14369 12068
rect 14325 12042 14340 12062
rect 14360 12042 14369 12062
rect 14325 12026 14369 12042
rect 14434 12058 14483 12068
rect 14434 12038 14445 12058
rect 14465 12038 14483 12058
rect 14434 12026 14483 12038
rect 14533 12062 14577 12068
rect 14533 12042 14548 12062
rect 14568 12042 14577 12062
rect 14533 12026 14577 12042
rect 14647 12062 14691 12068
rect 14647 12042 14656 12062
rect 14676 12042 14691 12062
rect 14647 12026 14691 12042
rect 14741 12058 14790 12068
rect 14741 12038 14759 12058
rect 14779 12038 14790 12058
rect 14741 12026 14790 12038
rect 6605 11433 6654 11445
rect 6605 11413 6616 11433
rect 6636 11413 6654 11433
rect 6605 11403 6654 11413
rect 6704 11429 6748 11445
rect 6704 11409 6719 11429
rect 6739 11409 6748 11429
rect 6704 11403 6748 11409
rect 6818 11429 6862 11445
rect 6818 11409 6827 11429
rect 6847 11409 6862 11429
rect 6818 11403 6862 11409
rect 6912 11433 6961 11445
rect 6912 11413 6930 11433
rect 6950 11413 6961 11433
rect 6912 11403 6961 11413
rect 7026 11429 7070 11445
rect 7026 11409 7035 11429
rect 7055 11409 7070 11429
rect 7026 11403 7070 11409
rect 7120 11433 7169 11445
rect 7120 11413 7138 11433
rect 7158 11413 7169 11433
rect 7120 11403 7169 11413
rect 7239 11429 7283 11445
rect 7239 11409 7248 11429
rect 7268 11409 7283 11429
rect 7239 11403 7283 11409
rect 7333 11433 7382 11445
rect 7333 11413 7351 11433
rect 7371 11413 7382 11433
rect 7333 11403 7382 11413
rect 9100 11428 9149 11440
rect 9100 11408 9111 11428
rect 9131 11408 9149 11428
rect 810 11301 859 11311
rect 810 11281 821 11301
rect 841 11281 859 11301
rect 810 11269 859 11281
rect 909 11305 953 11311
rect 909 11285 924 11305
rect 944 11285 953 11305
rect 909 11269 953 11285
rect 1023 11301 1072 11311
rect 1023 11281 1034 11301
rect 1054 11281 1072 11301
rect 1023 11269 1072 11281
rect 1122 11305 1166 11311
rect 1122 11285 1137 11305
rect 1157 11285 1166 11305
rect 1122 11269 1166 11285
rect 1231 11301 1280 11311
rect 1231 11281 1242 11301
rect 1262 11281 1280 11301
rect 1231 11269 1280 11281
rect 1330 11305 1374 11311
rect 1330 11285 1345 11305
rect 1365 11285 1374 11305
rect 1330 11269 1374 11285
rect 1444 11305 1488 11311
rect 1444 11285 1453 11305
rect 1473 11285 1488 11305
rect 1444 11269 1488 11285
rect 1538 11301 1587 11311
rect 9100 11398 9149 11408
rect 9199 11424 9243 11440
rect 9199 11404 9214 11424
rect 9234 11404 9243 11424
rect 9199 11398 9243 11404
rect 9313 11424 9357 11440
rect 9313 11404 9322 11424
rect 9342 11404 9357 11424
rect 9313 11398 9357 11404
rect 9407 11428 9456 11440
rect 9407 11408 9425 11428
rect 9445 11408 9456 11428
rect 9407 11398 9456 11408
rect 9521 11424 9565 11440
rect 9521 11404 9530 11424
rect 9550 11404 9565 11424
rect 9521 11398 9565 11404
rect 9615 11428 9664 11440
rect 9615 11408 9633 11428
rect 9653 11408 9664 11428
rect 9615 11398 9664 11408
rect 9734 11424 9778 11440
rect 9734 11404 9743 11424
rect 9763 11404 9778 11424
rect 9734 11398 9778 11404
rect 9828 11428 9877 11440
rect 9828 11408 9846 11428
rect 9866 11408 9877 11428
rect 9828 11398 9877 11408
rect 1538 11281 1556 11301
rect 1576 11281 1587 11301
rect 1538 11269 1587 11281
rect 1858 11297 1907 11307
rect 1858 11277 1869 11297
rect 1889 11277 1907 11297
rect 1858 11265 1907 11277
rect 1957 11301 2001 11307
rect 1957 11281 1972 11301
rect 1992 11281 2001 11301
rect 1957 11265 2001 11281
rect 2071 11297 2120 11307
rect 2071 11277 2082 11297
rect 2102 11277 2120 11297
rect 2071 11265 2120 11277
rect 2170 11301 2214 11307
rect 2170 11281 2185 11301
rect 2205 11281 2214 11301
rect 2170 11265 2214 11281
rect 2279 11297 2328 11307
rect 2279 11277 2290 11297
rect 2310 11277 2328 11297
rect 2279 11265 2328 11277
rect 2378 11301 2422 11307
rect 2378 11281 2393 11301
rect 2413 11281 2422 11301
rect 2378 11265 2422 11281
rect 2492 11301 2536 11307
rect 2492 11281 2501 11301
rect 2521 11281 2536 11301
rect 2492 11265 2536 11281
rect 2586 11297 2635 11307
rect 2586 11277 2604 11297
rect 2624 11277 2635 11297
rect 2586 11265 2635 11277
rect 17313 11427 17362 11439
rect 17313 11407 17324 11427
rect 17344 11407 17362 11427
rect 17313 11397 17362 11407
rect 17412 11423 17456 11439
rect 17412 11403 17427 11423
rect 17447 11403 17456 11423
rect 17412 11397 17456 11403
rect 17526 11423 17570 11439
rect 17526 11403 17535 11423
rect 17555 11403 17570 11423
rect 17526 11397 17570 11403
rect 17620 11427 17669 11439
rect 17620 11407 17638 11427
rect 17658 11407 17669 11427
rect 17620 11397 17669 11407
rect 17734 11423 17778 11439
rect 17734 11403 17743 11423
rect 17763 11403 17778 11423
rect 17734 11397 17778 11403
rect 17828 11427 17877 11439
rect 17828 11407 17846 11427
rect 17866 11407 17877 11427
rect 17828 11397 17877 11407
rect 17947 11423 17991 11439
rect 17947 11403 17956 11423
rect 17976 11403 17991 11423
rect 17947 11397 17991 11403
rect 18041 11427 18090 11439
rect 18041 11407 18059 11427
rect 18079 11407 18090 11427
rect 18041 11397 18090 11407
rect 19808 11422 19857 11434
rect 19808 11402 19819 11422
rect 19839 11402 19857 11422
rect 11518 11295 11567 11305
rect 11518 11275 11529 11295
rect 11549 11275 11567 11295
rect 11518 11263 11567 11275
rect 11617 11299 11661 11305
rect 11617 11279 11632 11299
rect 11652 11279 11661 11299
rect 11617 11263 11661 11279
rect 11731 11295 11780 11305
rect 11731 11275 11742 11295
rect 11762 11275 11780 11295
rect 11731 11263 11780 11275
rect 11830 11299 11874 11305
rect 11830 11279 11845 11299
rect 11865 11279 11874 11299
rect 11830 11263 11874 11279
rect 11939 11295 11988 11305
rect 11939 11275 11950 11295
rect 11970 11275 11988 11295
rect 11939 11263 11988 11275
rect 12038 11299 12082 11305
rect 12038 11279 12053 11299
rect 12073 11279 12082 11299
rect 12038 11263 12082 11279
rect 12152 11299 12196 11305
rect 12152 11279 12161 11299
rect 12181 11279 12196 11299
rect 12152 11263 12196 11279
rect 12246 11295 12295 11305
rect 19808 11392 19857 11402
rect 19907 11418 19951 11434
rect 19907 11398 19922 11418
rect 19942 11398 19951 11418
rect 19907 11392 19951 11398
rect 20021 11418 20065 11434
rect 20021 11398 20030 11418
rect 20050 11398 20065 11418
rect 20021 11392 20065 11398
rect 20115 11422 20164 11434
rect 20115 11402 20133 11422
rect 20153 11402 20164 11422
rect 20115 11392 20164 11402
rect 20229 11418 20273 11434
rect 20229 11398 20238 11418
rect 20258 11398 20273 11418
rect 20229 11392 20273 11398
rect 20323 11422 20372 11434
rect 20323 11402 20341 11422
rect 20361 11402 20372 11422
rect 20323 11392 20372 11402
rect 20442 11418 20486 11434
rect 20442 11398 20451 11418
rect 20471 11398 20486 11418
rect 20442 11392 20486 11398
rect 20536 11422 20585 11434
rect 20536 11402 20554 11422
rect 20574 11402 20585 11422
rect 20536 11392 20585 11402
rect 12246 11275 12264 11295
rect 12284 11275 12295 11295
rect 12246 11263 12295 11275
rect 12566 11291 12615 11301
rect 12566 11271 12577 11291
rect 12597 11271 12615 11291
rect 12566 11259 12615 11271
rect 12665 11295 12709 11301
rect 12665 11275 12680 11295
rect 12700 11275 12709 11295
rect 12665 11259 12709 11275
rect 12779 11291 12828 11301
rect 12779 11271 12790 11291
rect 12810 11271 12828 11291
rect 12779 11259 12828 11271
rect 12878 11295 12922 11301
rect 12878 11275 12893 11295
rect 12913 11275 12922 11295
rect 12878 11259 12922 11275
rect 12987 11291 13036 11301
rect 12987 11271 12998 11291
rect 13018 11271 13036 11291
rect 12987 11259 13036 11271
rect 13086 11295 13130 11301
rect 13086 11275 13101 11295
rect 13121 11275 13130 11295
rect 13086 11259 13130 11275
rect 13200 11295 13244 11301
rect 13200 11275 13209 11295
rect 13229 11275 13244 11295
rect 13200 11259 13244 11275
rect 13294 11291 13343 11301
rect 13294 11271 13312 11291
rect 13332 11271 13343 11291
rect 13294 11259 13343 11271
rect 8052 10753 8101 10765
rect 8052 10733 8063 10753
rect 8083 10733 8101 10753
rect 8052 10723 8101 10733
rect 8151 10749 8195 10765
rect 8151 10729 8166 10749
rect 8186 10729 8195 10749
rect 8151 10723 8195 10729
rect 8265 10749 8309 10765
rect 8265 10729 8274 10749
rect 8294 10729 8309 10749
rect 8265 10723 8309 10729
rect 8359 10753 8408 10765
rect 8359 10733 8377 10753
rect 8397 10733 8408 10753
rect 8359 10723 8408 10733
rect 8473 10749 8517 10765
rect 8473 10729 8482 10749
rect 8502 10729 8517 10749
rect 8473 10723 8517 10729
rect 8567 10753 8616 10765
rect 8567 10733 8585 10753
rect 8605 10733 8616 10753
rect 8567 10723 8616 10733
rect 8686 10749 8730 10765
rect 8686 10729 8695 10749
rect 8715 10729 8730 10749
rect 8686 10723 8730 10729
rect 8780 10753 8829 10765
rect 8780 10733 8798 10753
rect 8818 10733 8829 10753
rect 8780 10723 8829 10733
rect 9100 10749 9149 10761
rect 9100 10729 9111 10749
rect 9131 10729 9149 10749
rect 810 10622 859 10632
rect 810 10602 821 10622
rect 841 10602 859 10622
rect 810 10590 859 10602
rect 909 10626 953 10632
rect 909 10606 924 10626
rect 944 10606 953 10626
rect 909 10590 953 10606
rect 1023 10622 1072 10632
rect 1023 10602 1034 10622
rect 1054 10602 1072 10622
rect 1023 10590 1072 10602
rect 1122 10626 1166 10632
rect 1122 10606 1137 10626
rect 1157 10606 1166 10626
rect 1122 10590 1166 10606
rect 1231 10622 1280 10632
rect 1231 10602 1242 10622
rect 1262 10602 1280 10622
rect 1231 10590 1280 10602
rect 1330 10626 1374 10632
rect 1330 10606 1345 10626
rect 1365 10606 1374 10626
rect 1330 10590 1374 10606
rect 1444 10626 1488 10632
rect 1444 10606 1453 10626
rect 1473 10606 1488 10626
rect 1444 10590 1488 10606
rect 1538 10622 1587 10632
rect 9100 10719 9149 10729
rect 9199 10745 9243 10761
rect 9199 10725 9214 10745
rect 9234 10725 9243 10745
rect 9199 10719 9243 10725
rect 9313 10745 9357 10761
rect 9313 10725 9322 10745
rect 9342 10725 9357 10745
rect 9313 10719 9357 10725
rect 9407 10749 9456 10761
rect 9407 10729 9425 10749
rect 9445 10729 9456 10749
rect 9407 10719 9456 10729
rect 9521 10745 9565 10761
rect 9521 10725 9530 10745
rect 9550 10725 9565 10745
rect 9521 10719 9565 10725
rect 9615 10749 9664 10761
rect 9615 10729 9633 10749
rect 9653 10729 9664 10749
rect 9615 10719 9664 10729
rect 9734 10745 9778 10761
rect 9734 10725 9743 10745
rect 9763 10725 9778 10745
rect 9734 10719 9778 10725
rect 9828 10749 9877 10761
rect 9828 10729 9846 10749
rect 9866 10729 9877 10749
rect 9828 10719 9877 10729
rect 1538 10602 1556 10622
rect 1576 10602 1587 10622
rect 1538 10590 1587 10602
rect 3348 10619 3397 10629
rect 3348 10599 3359 10619
rect 3379 10599 3397 10619
rect 3348 10587 3397 10599
rect 3447 10623 3491 10629
rect 3447 10603 3462 10623
rect 3482 10603 3491 10623
rect 3447 10587 3491 10603
rect 3561 10619 3610 10629
rect 3561 10599 3572 10619
rect 3592 10599 3610 10619
rect 3561 10587 3610 10599
rect 3660 10623 3704 10629
rect 3660 10603 3675 10623
rect 3695 10603 3704 10623
rect 3660 10587 3704 10603
rect 3769 10619 3818 10629
rect 3769 10599 3780 10619
rect 3800 10599 3818 10619
rect 3769 10587 3818 10599
rect 3868 10623 3912 10629
rect 3868 10603 3883 10623
rect 3903 10603 3912 10623
rect 3868 10587 3912 10603
rect 3982 10623 4026 10629
rect 3982 10603 3991 10623
rect 4011 10603 4026 10623
rect 3982 10587 4026 10603
rect 4076 10619 4125 10629
rect 4076 10599 4094 10619
rect 4114 10599 4125 10619
rect 4076 10587 4125 10599
rect 18760 10747 18809 10759
rect 18760 10727 18771 10747
rect 18791 10727 18809 10747
rect 18760 10717 18809 10727
rect 18859 10743 18903 10759
rect 18859 10723 18874 10743
rect 18894 10723 18903 10743
rect 18859 10717 18903 10723
rect 18973 10743 19017 10759
rect 18973 10723 18982 10743
rect 19002 10723 19017 10743
rect 18973 10717 19017 10723
rect 19067 10747 19116 10759
rect 19067 10727 19085 10747
rect 19105 10727 19116 10747
rect 19067 10717 19116 10727
rect 19181 10743 19225 10759
rect 19181 10723 19190 10743
rect 19210 10723 19225 10743
rect 19181 10717 19225 10723
rect 19275 10747 19324 10759
rect 19275 10727 19293 10747
rect 19313 10727 19324 10747
rect 19275 10717 19324 10727
rect 19394 10743 19438 10759
rect 19394 10723 19403 10743
rect 19423 10723 19438 10743
rect 19394 10717 19438 10723
rect 19488 10747 19537 10759
rect 19488 10727 19506 10747
rect 19526 10727 19537 10747
rect 19488 10717 19537 10727
rect 19808 10743 19857 10755
rect 19808 10723 19819 10743
rect 19839 10723 19857 10743
rect 11518 10616 11567 10626
rect 11518 10596 11529 10616
rect 11549 10596 11567 10616
rect 11518 10584 11567 10596
rect 11617 10620 11661 10626
rect 11617 10600 11632 10620
rect 11652 10600 11661 10620
rect 11617 10584 11661 10600
rect 11731 10616 11780 10626
rect 11731 10596 11742 10616
rect 11762 10596 11780 10616
rect 11731 10584 11780 10596
rect 11830 10620 11874 10626
rect 11830 10600 11845 10620
rect 11865 10600 11874 10620
rect 11830 10584 11874 10600
rect 11939 10616 11988 10626
rect 11939 10596 11950 10616
rect 11970 10596 11988 10616
rect 11939 10584 11988 10596
rect 12038 10620 12082 10626
rect 12038 10600 12053 10620
rect 12073 10600 12082 10620
rect 12038 10584 12082 10600
rect 12152 10620 12196 10626
rect 12152 10600 12161 10620
rect 12181 10600 12196 10620
rect 12152 10584 12196 10600
rect 12246 10616 12295 10626
rect 19808 10713 19857 10723
rect 19907 10739 19951 10755
rect 19907 10719 19922 10739
rect 19942 10719 19951 10739
rect 19907 10713 19951 10719
rect 20021 10739 20065 10755
rect 20021 10719 20030 10739
rect 20050 10719 20065 10739
rect 20021 10713 20065 10719
rect 20115 10743 20164 10755
rect 20115 10723 20133 10743
rect 20153 10723 20164 10743
rect 20115 10713 20164 10723
rect 20229 10739 20273 10755
rect 20229 10719 20238 10739
rect 20258 10719 20273 10739
rect 20229 10713 20273 10719
rect 20323 10743 20372 10755
rect 20323 10723 20341 10743
rect 20361 10723 20372 10743
rect 20323 10713 20372 10723
rect 20442 10739 20486 10755
rect 20442 10719 20451 10739
rect 20471 10719 20486 10739
rect 20442 10713 20486 10719
rect 20536 10743 20585 10755
rect 20536 10723 20554 10743
rect 20574 10723 20585 10743
rect 20536 10713 20585 10723
rect 12246 10596 12264 10616
rect 12284 10596 12295 10616
rect 12246 10584 12295 10596
rect 14056 10613 14105 10623
rect 14056 10593 14067 10613
rect 14087 10593 14105 10613
rect 14056 10581 14105 10593
rect 14155 10617 14199 10623
rect 14155 10597 14170 10617
rect 14190 10597 14199 10617
rect 14155 10581 14199 10597
rect 14269 10613 14318 10623
rect 14269 10593 14280 10613
rect 14300 10593 14318 10613
rect 14269 10581 14318 10593
rect 14368 10617 14412 10623
rect 14368 10597 14383 10617
rect 14403 10597 14412 10617
rect 14368 10581 14412 10597
rect 14477 10613 14526 10623
rect 14477 10593 14488 10613
rect 14508 10593 14526 10613
rect 14477 10581 14526 10593
rect 14576 10617 14620 10623
rect 14576 10597 14591 10617
rect 14611 10597 14620 10617
rect 14576 10581 14620 10597
rect 14690 10617 14734 10623
rect 14690 10597 14699 10617
rect 14719 10597 14734 10617
rect 14690 10581 14734 10597
rect 14784 10613 14833 10623
rect 14784 10593 14802 10613
rect 14822 10593 14833 10613
rect 14784 10581 14833 10593
rect 6563 9911 6612 9923
rect 6563 9891 6574 9911
rect 6594 9891 6612 9911
rect 6563 9881 6612 9891
rect 6662 9907 6706 9923
rect 6662 9887 6677 9907
rect 6697 9887 6706 9907
rect 6662 9881 6706 9887
rect 6776 9907 6820 9923
rect 6776 9887 6785 9907
rect 6805 9887 6820 9907
rect 6776 9881 6820 9887
rect 6870 9911 6919 9923
rect 6870 9891 6888 9911
rect 6908 9891 6919 9911
rect 6870 9881 6919 9891
rect 6984 9907 7028 9923
rect 6984 9887 6993 9907
rect 7013 9887 7028 9907
rect 6984 9881 7028 9887
rect 7078 9911 7127 9923
rect 7078 9891 7096 9911
rect 7116 9891 7127 9911
rect 7078 9881 7127 9891
rect 7197 9907 7241 9923
rect 7197 9887 7206 9907
rect 7226 9887 7241 9907
rect 7197 9881 7241 9887
rect 7291 9911 7340 9923
rect 7291 9891 7309 9911
rect 7329 9891 7340 9911
rect 7291 9881 7340 9891
rect 9101 9908 9150 9920
rect 9101 9888 9112 9908
rect 9132 9888 9150 9908
rect 811 9781 860 9791
rect 811 9761 822 9781
rect 842 9761 860 9781
rect 811 9749 860 9761
rect 910 9785 954 9791
rect 910 9765 925 9785
rect 945 9765 954 9785
rect 910 9749 954 9765
rect 1024 9781 1073 9791
rect 1024 9761 1035 9781
rect 1055 9761 1073 9781
rect 1024 9749 1073 9761
rect 1123 9785 1167 9791
rect 1123 9765 1138 9785
rect 1158 9765 1167 9785
rect 1123 9749 1167 9765
rect 1232 9781 1281 9791
rect 1232 9761 1243 9781
rect 1263 9761 1281 9781
rect 1232 9749 1281 9761
rect 1331 9785 1375 9791
rect 1331 9765 1346 9785
rect 1366 9765 1375 9785
rect 1331 9749 1375 9765
rect 1445 9785 1489 9791
rect 1445 9765 1454 9785
rect 1474 9765 1489 9785
rect 1445 9749 1489 9765
rect 1539 9781 1588 9791
rect 9101 9878 9150 9888
rect 9200 9904 9244 9920
rect 9200 9884 9215 9904
rect 9235 9884 9244 9904
rect 9200 9878 9244 9884
rect 9314 9904 9358 9920
rect 9314 9884 9323 9904
rect 9343 9884 9358 9904
rect 9314 9878 9358 9884
rect 9408 9908 9457 9920
rect 9408 9888 9426 9908
rect 9446 9888 9457 9908
rect 9408 9878 9457 9888
rect 9522 9904 9566 9920
rect 9522 9884 9531 9904
rect 9551 9884 9566 9904
rect 9522 9878 9566 9884
rect 9616 9908 9665 9920
rect 9616 9888 9634 9908
rect 9654 9888 9665 9908
rect 9616 9878 9665 9888
rect 9735 9904 9779 9920
rect 9735 9884 9744 9904
rect 9764 9884 9779 9904
rect 9735 9878 9779 9884
rect 9829 9908 9878 9920
rect 9829 9888 9847 9908
rect 9867 9888 9878 9908
rect 9829 9878 9878 9888
rect 1539 9761 1557 9781
rect 1577 9761 1588 9781
rect 1539 9749 1588 9761
rect 1859 9777 1908 9787
rect 1859 9757 1870 9777
rect 1890 9757 1908 9777
rect 1859 9745 1908 9757
rect 1958 9781 2002 9787
rect 1958 9761 1973 9781
rect 1993 9761 2002 9781
rect 1958 9745 2002 9761
rect 2072 9777 2121 9787
rect 2072 9757 2083 9777
rect 2103 9757 2121 9777
rect 2072 9745 2121 9757
rect 2171 9781 2215 9787
rect 2171 9761 2186 9781
rect 2206 9761 2215 9781
rect 2171 9745 2215 9761
rect 2280 9777 2329 9787
rect 2280 9757 2291 9777
rect 2311 9757 2329 9777
rect 2280 9745 2329 9757
rect 2379 9781 2423 9787
rect 2379 9761 2394 9781
rect 2414 9761 2423 9781
rect 2379 9745 2423 9761
rect 2493 9781 2537 9787
rect 2493 9761 2502 9781
rect 2522 9761 2537 9781
rect 2493 9745 2537 9761
rect 2587 9777 2636 9787
rect 2587 9757 2605 9777
rect 2625 9757 2636 9777
rect 2587 9745 2636 9757
rect 17271 9905 17320 9917
rect 17271 9885 17282 9905
rect 17302 9885 17320 9905
rect 17271 9875 17320 9885
rect 17370 9901 17414 9917
rect 17370 9881 17385 9901
rect 17405 9881 17414 9901
rect 17370 9875 17414 9881
rect 17484 9901 17528 9917
rect 17484 9881 17493 9901
rect 17513 9881 17528 9901
rect 17484 9875 17528 9881
rect 17578 9905 17627 9917
rect 17578 9885 17596 9905
rect 17616 9885 17627 9905
rect 17578 9875 17627 9885
rect 17692 9901 17736 9917
rect 17692 9881 17701 9901
rect 17721 9881 17736 9901
rect 17692 9875 17736 9881
rect 17786 9905 17835 9917
rect 17786 9885 17804 9905
rect 17824 9885 17835 9905
rect 17786 9875 17835 9885
rect 17905 9901 17949 9917
rect 17905 9881 17914 9901
rect 17934 9881 17949 9901
rect 17905 9875 17949 9881
rect 17999 9905 18048 9917
rect 17999 9885 18017 9905
rect 18037 9885 18048 9905
rect 17999 9875 18048 9885
rect 19809 9902 19858 9914
rect 19809 9882 19820 9902
rect 19840 9882 19858 9902
rect 11519 9775 11568 9785
rect 11519 9755 11530 9775
rect 11550 9755 11568 9775
rect 11519 9743 11568 9755
rect 11618 9779 11662 9785
rect 11618 9759 11633 9779
rect 11653 9759 11662 9779
rect 11618 9743 11662 9759
rect 11732 9775 11781 9785
rect 11732 9755 11743 9775
rect 11763 9755 11781 9775
rect 11732 9743 11781 9755
rect 11831 9779 11875 9785
rect 11831 9759 11846 9779
rect 11866 9759 11875 9779
rect 11831 9743 11875 9759
rect 11940 9775 11989 9785
rect 11940 9755 11951 9775
rect 11971 9755 11989 9775
rect 11940 9743 11989 9755
rect 12039 9779 12083 9785
rect 12039 9759 12054 9779
rect 12074 9759 12083 9779
rect 12039 9743 12083 9759
rect 12153 9779 12197 9785
rect 12153 9759 12162 9779
rect 12182 9759 12197 9779
rect 12153 9743 12197 9759
rect 12247 9775 12296 9785
rect 19809 9872 19858 9882
rect 19908 9898 19952 9914
rect 19908 9878 19923 9898
rect 19943 9878 19952 9898
rect 19908 9872 19952 9878
rect 20022 9898 20066 9914
rect 20022 9878 20031 9898
rect 20051 9878 20066 9898
rect 20022 9872 20066 9878
rect 20116 9902 20165 9914
rect 20116 9882 20134 9902
rect 20154 9882 20165 9902
rect 20116 9872 20165 9882
rect 20230 9898 20274 9914
rect 20230 9878 20239 9898
rect 20259 9878 20274 9898
rect 20230 9872 20274 9878
rect 20324 9902 20373 9914
rect 20324 9882 20342 9902
rect 20362 9882 20373 9902
rect 20324 9872 20373 9882
rect 20443 9898 20487 9914
rect 20443 9878 20452 9898
rect 20472 9878 20487 9898
rect 20443 9872 20487 9878
rect 20537 9902 20586 9914
rect 20537 9882 20555 9902
rect 20575 9882 20586 9902
rect 20537 9872 20586 9882
rect 12247 9755 12265 9775
rect 12285 9755 12296 9775
rect 12247 9743 12296 9755
rect 12567 9771 12616 9781
rect 12567 9751 12578 9771
rect 12598 9751 12616 9771
rect 12567 9739 12616 9751
rect 12666 9775 12710 9781
rect 12666 9755 12681 9775
rect 12701 9755 12710 9775
rect 12666 9739 12710 9755
rect 12780 9771 12829 9781
rect 12780 9751 12791 9771
rect 12811 9751 12829 9771
rect 12780 9739 12829 9751
rect 12879 9775 12923 9781
rect 12879 9755 12894 9775
rect 12914 9755 12923 9775
rect 12879 9739 12923 9755
rect 12988 9771 13037 9781
rect 12988 9751 12999 9771
rect 13019 9751 13037 9771
rect 12988 9739 13037 9751
rect 13087 9775 13131 9781
rect 13087 9755 13102 9775
rect 13122 9755 13131 9775
rect 13087 9739 13131 9755
rect 13201 9775 13245 9781
rect 13201 9755 13210 9775
rect 13230 9755 13245 9775
rect 13201 9739 13245 9755
rect 13295 9771 13344 9781
rect 13295 9751 13313 9771
rect 13333 9751 13344 9771
rect 13295 9739 13344 9751
rect 8053 9233 8102 9245
rect 8053 9213 8064 9233
rect 8084 9213 8102 9233
rect 8053 9203 8102 9213
rect 8152 9229 8196 9245
rect 8152 9209 8167 9229
rect 8187 9209 8196 9229
rect 8152 9203 8196 9209
rect 8266 9229 8310 9245
rect 8266 9209 8275 9229
rect 8295 9209 8310 9229
rect 8266 9203 8310 9209
rect 8360 9233 8409 9245
rect 8360 9213 8378 9233
rect 8398 9213 8409 9233
rect 8360 9203 8409 9213
rect 8474 9229 8518 9245
rect 8474 9209 8483 9229
rect 8503 9209 8518 9229
rect 8474 9203 8518 9209
rect 8568 9233 8617 9245
rect 8568 9213 8586 9233
rect 8606 9213 8617 9233
rect 8568 9203 8617 9213
rect 8687 9229 8731 9245
rect 8687 9209 8696 9229
rect 8716 9209 8731 9229
rect 8687 9203 8731 9209
rect 8781 9233 8830 9245
rect 8781 9213 8799 9233
rect 8819 9213 8830 9233
rect 8781 9203 8830 9213
rect 9101 9229 9150 9241
rect 9101 9209 9112 9229
rect 9132 9209 9150 9229
rect 811 9102 860 9112
rect 811 9082 822 9102
rect 842 9082 860 9102
rect 811 9070 860 9082
rect 910 9106 954 9112
rect 910 9086 925 9106
rect 945 9086 954 9106
rect 910 9070 954 9086
rect 1024 9102 1073 9112
rect 1024 9082 1035 9102
rect 1055 9082 1073 9102
rect 1024 9070 1073 9082
rect 1123 9106 1167 9112
rect 1123 9086 1138 9106
rect 1158 9086 1167 9106
rect 1123 9070 1167 9086
rect 1232 9102 1281 9112
rect 1232 9082 1243 9102
rect 1263 9082 1281 9102
rect 1232 9070 1281 9082
rect 1331 9106 1375 9112
rect 1331 9086 1346 9106
rect 1366 9086 1375 9106
rect 1331 9070 1375 9086
rect 1445 9106 1489 9112
rect 1445 9086 1454 9106
rect 1474 9086 1489 9106
rect 1445 9070 1489 9086
rect 1539 9102 1588 9112
rect 9101 9199 9150 9209
rect 9200 9225 9244 9241
rect 9200 9205 9215 9225
rect 9235 9205 9244 9225
rect 9200 9199 9244 9205
rect 9314 9225 9358 9241
rect 9314 9205 9323 9225
rect 9343 9205 9358 9225
rect 9314 9199 9358 9205
rect 9408 9229 9457 9241
rect 9408 9209 9426 9229
rect 9446 9209 9457 9229
rect 9408 9199 9457 9209
rect 9522 9225 9566 9241
rect 9522 9205 9531 9225
rect 9551 9205 9566 9225
rect 9522 9199 9566 9205
rect 9616 9229 9665 9241
rect 9616 9209 9634 9229
rect 9654 9209 9665 9229
rect 9616 9199 9665 9209
rect 9735 9225 9779 9241
rect 9735 9205 9744 9225
rect 9764 9205 9779 9225
rect 9735 9199 9779 9205
rect 9829 9229 9878 9241
rect 9829 9209 9847 9229
rect 9867 9209 9878 9229
rect 9829 9199 9878 9209
rect 1539 9082 1557 9102
rect 1577 9082 1588 9102
rect 1539 9070 1588 9082
rect 3306 9097 3355 9107
rect 3306 9077 3317 9097
rect 3337 9077 3355 9097
rect 3306 9065 3355 9077
rect 3405 9101 3449 9107
rect 3405 9081 3420 9101
rect 3440 9081 3449 9101
rect 3405 9065 3449 9081
rect 3519 9097 3568 9107
rect 3519 9077 3530 9097
rect 3550 9077 3568 9097
rect 3519 9065 3568 9077
rect 3618 9101 3662 9107
rect 3618 9081 3633 9101
rect 3653 9081 3662 9101
rect 3618 9065 3662 9081
rect 3727 9097 3776 9107
rect 3727 9077 3738 9097
rect 3758 9077 3776 9097
rect 3727 9065 3776 9077
rect 3826 9101 3870 9107
rect 3826 9081 3841 9101
rect 3861 9081 3870 9101
rect 3826 9065 3870 9081
rect 3940 9101 3984 9107
rect 3940 9081 3949 9101
rect 3969 9081 3984 9101
rect 3940 9065 3984 9081
rect 4034 9097 4083 9107
rect 4034 9077 4052 9097
rect 4072 9077 4083 9097
rect 4034 9065 4083 9077
rect 18761 9227 18810 9239
rect 18761 9207 18772 9227
rect 18792 9207 18810 9227
rect 18761 9197 18810 9207
rect 18860 9223 18904 9239
rect 18860 9203 18875 9223
rect 18895 9203 18904 9223
rect 18860 9197 18904 9203
rect 18974 9223 19018 9239
rect 18974 9203 18983 9223
rect 19003 9203 19018 9223
rect 18974 9197 19018 9203
rect 19068 9227 19117 9239
rect 19068 9207 19086 9227
rect 19106 9207 19117 9227
rect 19068 9197 19117 9207
rect 19182 9223 19226 9239
rect 19182 9203 19191 9223
rect 19211 9203 19226 9223
rect 19182 9197 19226 9203
rect 19276 9227 19325 9239
rect 19276 9207 19294 9227
rect 19314 9207 19325 9227
rect 19276 9197 19325 9207
rect 19395 9223 19439 9239
rect 19395 9203 19404 9223
rect 19424 9203 19439 9223
rect 19395 9197 19439 9203
rect 19489 9227 19538 9239
rect 19489 9207 19507 9227
rect 19527 9207 19538 9227
rect 19489 9197 19538 9207
rect 19809 9223 19858 9235
rect 19809 9203 19820 9223
rect 19840 9203 19858 9223
rect 11519 9096 11568 9106
rect 11519 9076 11530 9096
rect 11550 9076 11568 9096
rect 11519 9064 11568 9076
rect 11618 9100 11662 9106
rect 11618 9080 11633 9100
rect 11653 9080 11662 9100
rect 11618 9064 11662 9080
rect 11732 9096 11781 9106
rect 11732 9076 11743 9096
rect 11763 9076 11781 9096
rect 11732 9064 11781 9076
rect 11831 9100 11875 9106
rect 11831 9080 11846 9100
rect 11866 9080 11875 9100
rect 11831 9064 11875 9080
rect 11940 9096 11989 9106
rect 11940 9076 11951 9096
rect 11971 9076 11989 9096
rect 11940 9064 11989 9076
rect 12039 9100 12083 9106
rect 12039 9080 12054 9100
rect 12074 9080 12083 9100
rect 12039 9064 12083 9080
rect 12153 9100 12197 9106
rect 12153 9080 12162 9100
rect 12182 9080 12197 9100
rect 12153 9064 12197 9080
rect 12247 9096 12296 9106
rect 19809 9193 19858 9203
rect 19908 9219 19952 9235
rect 19908 9199 19923 9219
rect 19943 9199 19952 9219
rect 19908 9193 19952 9199
rect 20022 9219 20066 9235
rect 20022 9199 20031 9219
rect 20051 9199 20066 9219
rect 20022 9193 20066 9199
rect 20116 9223 20165 9235
rect 20116 9203 20134 9223
rect 20154 9203 20165 9223
rect 20116 9193 20165 9203
rect 20230 9219 20274 9235
rect 20230 9199 20239 9219
rect 20259 9199 20274 9219
rect 20230 9193 20274 9199
rect 20324 9223 20373 9235
rect 20324 9203 20342 9223
rect 20362 9203 20373 9223
rect 20324 9193 20373 9203
rect 20443 9219 20487 9235
rect 20443 9199 20452 9219
rect 20472 9199 20487 9219
rect 20443 9193 20487 9199
rect 20537 9223 20586 9235
rect 20537 9203 20555 9223
rect 20575 9203 20586 9223
rect 20537 9193 20586 9203
rect 12247 9076 12265 9096
rect 12285 9076 12296 9096
rect 12247 9064 12296 9076
rect 14014 9091 14063 9101
rect 14014 9071 14025 9091
rect 14045 9071 14063 9091
rect 14014 9059 14063 9071
rect 14113 9095 14157 9101
rect 14113 9075 14128 9095
rect 14148 9075 14157 9095
rect 14113 9059 14157 9075
rect 14227 9091 14276 9101
rect 14227 9071 14238 9091
rect 14258 9071 14276 9091
rect 14227 9059 14276 9071
rect 14326 9095 14370 9101
rect 14326 9075 14341 9095
rect 14361 9075 14370 9095
rect 14326 9059 14370 9075
rect 14435 9091 14484 9101
rect 14435 9071 14446 9091
rect 14466 9071 14484 9091
rect 14435 9059 14484 9071
rect 14534 9095 14578 9101
rect 14534 9075 14549 9095
rect 14569 9075 14578 9095
rect 14534 9059 14578 9075
rect 14648 9095 14692 9101
rect 14648 9075 14657 9095
rect 14677 9075 14692 9095
rect 14648 9059 14692 9075
rect 14742 9091 14791 9101
rect 14742 9071 14760 9091
rect 14780 9071 14791 9091
rect 14742 9059 14791 9071
rect 6606 8466 6655 8478
rect 6606 8446 6617 8466
rect 6637 8446 6655 8466
rect 6606 8436 6655 8446
rect 6705 8462 6749 8478
rect 6705 8442 6720 8462
rect 6740 8442 6749 8462
rect 6705 8436 6749 8442
rect 6819 8462 6863 8478
rect 6819 8442 6828 8462
rect 6848 8442 6863 8462
rect 6819 8436 6863 8442
rect 6913 8466 6962 8478
rect 6913 8446 6931 8466
rect 6951 8446 6962 8466
rect 6913 8436 6962 8446
rect 7027 8462 7071 8478
rect 7027 8442 7036 8462
rect 7056 8442 7071 8462
rect 7027 8436 7071 8442
rect 7121 8466 7170 8478
rect 7121 8446 7139 8466
rect 7159 8446 7170 8466
rect 7121 8436 7170 8446
rect 7240 8462 7284 8478
rect 7240 8442 7249 8462
rect 7269 8442 7284 8462
rect 7240 8436 7284 8442
rect 7334 8466 7383 8478
rect 7334 8446 7352 8466
rect 7372 8446 7383 8466
rect 7334 8436 7383 8446
rect 9101 8461 9150 8473
rect 9101 8441 9112 8461
rect 9132 8441 9150 8461
rect 811 8334 860 8344
rect 811 8314 822 8334
rect 842 8314 860 8334
rect 811 8302 860 8314
rect 910 8338 954 8344
rect 910 8318 925 8338
rect 945 8318 954 8338
rect 910 8302 954 8318
rect 1024 8334 1073 8344
rect 1024 8314 1035 8334
rect 1055 8314 1073 8334
rect 1024 8302 1073 8314
rect 1123 8338 1167 8344
rect 1123 8318 1138 8338
rect 1158 8318 1167 8338
rect 1123 8302 1167 8318
rect 1232 8334 1281 8344
rect 1232 8314 1243 8334
rect 1263 8314 1281 8334
rect 1232 8302 1281 8314
rect 1331 8338 1375 8344
rect 1331 8318 1346 8338
rect 1366 8318 1375 8338
rect 1331 8302 1375 8318
rect 1445 8338 1489 8344
rect 1445 8318 1454 8338
rect 1474 8318 1489 8338
rect 1445 8302 1489 8318
rect 1539 8334 1588 8344
rect 9101 8431 9150 8441
rect 9200 8457 9244 8473
rect 9200 8437 9215 8457
rect 9235 8437 9244 8457
rect 9200 8431 9244 8437
rect 9314 8457 9358 8473
rect 9314 8437 9323 8457
rect 9343 8437 9358 8457
rect 9314 8431 9358 8437
rect 9408 8461 9457 8473
rect 9408 8441 9426 8461
rect 9446 8441 9457 8461
rect 9408 8431 9457 8441
rect 9522 8457 9566 8473
rect 9522 8437 9531 8457
rect 9551 8437 9566 8457
rect 9522 8431 9566 8437
rect 9616 8461 9665 8473
rect 9616 8441 9634 8461
rect 9654 8441 9665 8461
rect 9616 8431 9665 8441
rect 9735 8457 9779 8473
rect 9735 8437 9744 8457
rect 9764 8437 9779 8457
rect 9735 8431 9779 8437
rect 9829 8461 9878 8473
rect 9829 8441 9847 8461
rect 9867 8441 9878 8461
rect 9829 8431 9878 8441
rect 1539 8314 1557 8334
rect 1577 8314 1588 8334
rect 1539 8302 1588 8314
rect 1859 8330 1908 8340
rect 1859 8310 1870 8330
rect 1890 8310 1908 8330
rect 1859 8298 1908 8310
rect 1958 8334 2002 8340
rect 1958 8314 1973 8334
rect 1993 8314 2002 8334
rect 1958 8298 2002 8314
rect 2072 8330 2121 8340
rect 2072 8310 2083 8330
rect 2103 8310 2121 8330
rect 2072 8298 2121 8310
rect 2171 8334 2215 8340
rect 2171 8314 2186 8334
rect 2206 8314 2215 8334
rect 2171 8298 2215 8314
rect 2280 8330 2329 8340
rect 2280 8310 2291 8330
rect 2311 8310 2329 8330
rect 2280 8298 2329 8310
rect 2379 8334 2423 8340
rect 2379 8314 2394 8334
rect 2414 8314 2423 8334
rect 2379 8298 2423 8314
rect 2493 8334 2537 8340
rect 2493 8314 2502 8334
rect 2522 8314 2537 8334
rect 2493 8298 2537 8314
rect 2587 8330 2636 8340
rect 2587 8310 2605 8330
rect 2625 8310 2636 8330
rect 2587 8298 2636 8310
rect 17314 8460 17363 8472
rect 17314 8440 17325 8460
rect 17345 8440 17363 8460
rect 17314 8430 17363 8440
rect 17413 8456 17457 8472
rect 17413 8436 17428 8456
rect 17448 8436 17457 8456
rect 17413 8430 17457 8436
rect 17527 8456 17571 8472
rect 17527 8436 17536 8456
rect 17556 8436 17571 8456
rect 17527 8430 17571 8436
rect 17621 8460 17670 8472
rect 17621 8440 17639 8460
rect 17659 8440 17670 8460
rect 17621 8430 17670 8440
rect 17735 8456 17779 8472
rect 17735 8436 17744 8456
rect 17764 8436 17779 8456
rect 17735 8430 17779 8436
rect 17829 8460 17878 8472
rect 17829 8440 17847 8460
rect 17867 8440 17878 8460
rect 17829 8430 17878 8440
rect 17948 8456 17992 8472
rect 17948 8436 17957 8456
rect 17977 8436 17992 8456
rect 17948 8430 17992 8436
rect 18042 8460 18091 8472
rect 18042 8440 18060 8460
rect 18080 8440 18091 8460
rect 18042 8430 18091 8440
rect 19809 8455 19858 8467
rect 19809 8435 19820 8455
rect 19840 8435 19858 8455
rect 11519 8328 11568 8338
rect 11519 8308 11530 8328
rect 11550 8308 11568 8328
rect 11519 8296 11568 8308
rect 11618 8332 11662 8338
rect 11618 8312 11633 8332
rect 11653 8312 11662 8332
rect 11618 8296 11662 8312
rect 11732 8328 11781 8338
rect 11732 8308 11743 8328
rect 11763 8308 11781 8328
rect 11732 8296 11781 8308
rect 11831 8332 11875 8338
rect 11831 8312 11846 8332
rect 11866 8312 11875 8332
rect 11831 8296 11875 8312
rect 11940 8328 11989 8338
rect 11940 8308 11951 8328
rect 11971 8308 11989 8328
rect 11940 8296 11989 8308
rect 12039 8332 12083 8338
rect 12039 8312 12054 8332
rect 12074 8312 12083 8332
rect 12039 8296 12083 8312
rect 12153 8332 12197 8338
rect 12153 8312 12162 8332
rect 12182 8312 12197 8332
rect 12153 8296 12197 8312
rect 12247 8328 12296 8338
rect 19809 8425 19858 8435
rect 19908 8451 19952 8467
rect 19908 8431 19923 8451
rect 19943 8431 19952 8451
rect 19908 8425 19952 8431
rect 20022 8451 20066 8467
rect 20022 8431 20031 8451
rect 20051 8431 20066 8451
rect 20022 8425 20066 8431
rect 20116 8455 20165 8467
rect 20116 8435 20134 8455
rect 20154 8435 20165 8455
rect 20116 8425 20165 8435
rect 20230 8451 20274 8467
rect 20230 8431 20239 8451
rect 20259 8431 20274 8451
rect 20230 8425 20274 8431
rect 20324 8455 20373 8467
rect 20324 8435 20342 8455
rect 20362 8435 20373 8455
rect 20324 8425 20373 8435
rect 20443 8451 20487 8467
rect 20443 8431 20452 8451
rect 20472 8431 20487 8451
rect 20443 8425 20487 8431
rect 20537 8455 20586 8467
rect 20537 8435 20555 8455
rect 20575 8435 20586 8455
rect 20537 8425 20586 8435
rect 12247 8308 12265 8328
rect 12285 8308 12296 8328
rect 12247 8296 12296 8308
rect 12567 8324 12616 8334
rect 12567 8304 12578 8324
rect 12598 8304 12616 8324
rect 12567 8292 12616 8304
rect 12666 8328 12710 8334
rect 12666 8308 12681 8328
rect 12701 8308 12710 8328
rect 12666 8292 12710 8308
rect 12780 8324 12829 8334
rect 12780 8304 12791 8324
rect 12811 8304 12829 8324
rect 12780 8292 12829 8304
rect 12879 8328 12923 8334
rect 12879 8308 12894 8328
rect 12914 8308 12923 8328
rect 12879 8292 12923 8308
rect 12988 8324 13037 8334
rect 12988 8304 12999 8324
rect 13019 8304 13037 8324
rect 12988 8292 13037 8304
rect 13087 8328 13131 8334
rect 13087 8308 13102 8328
rect 13122 8308 13131 8328
rect 13087 8292 13131 8308
rect 13201 8328 13245 8334
rect 13201 8308 13210 8328
rect 13230 8308 13245 8328
rect 13201 8292 13245 8308
rect 13295 8324 13344 8334
rect 13295 8304 13313 8324
rect 13333 8304 13344 8324
rect 13295 8292 13344 8304
rect 8053 7786 8102 7798
rect 8053 7766 8064 7786
rect 8084 7766 8102 7786
rect 8053 7756 8102 7766
rect 8152 7782 8196 7798
rect 8152 7762 8167 7782
rect 8187 7762 8196 7782
rect 8152 7756 8196 7762
rect 8266 7782 8310 7798
rect 8266 7762 8275 7782
rect 8295 7762 8310 7782
rect 8266 7756 8310 7762
rect 8360 7786 8409 7798
rect 8360 7766 8378 7786
rect 8398 7766 8409 7786
rect 8360 7756 8409 7766
rect 8474 7782 8518 7798
rect 8474 7762 8483 7782
rect 8503 7762 8518 7782
rect 8474 7756 8518 7762
rect 8568 7786 8617 7798
rect 8568 7766 8586 7786
rect 8606 7766 8617 7786
rect 8568 7756 8617 7766
rect 8687 7782 8731 7798
rect 8687 7762 8696 7782
rect 8716 7762 8731 7782
rect 8687 7756 8731 7762
rect 8781 7786 8830 7798
rect 8781 7766 8799 7786
rect 8819 7766 8830 7786
rect 8781 7756 8830 7766
rect 9101 7782 9150 7794
rect 9101 7762 9112 7782
rect 9132 7762 9150 7782
rect 811 7655 860 7665
rect 811 7635 822 7655
rect 842 7635 860 7655
rect 811 7623 860 7635
rect 910 7659 954 7665
rect 910 7639 925 7659
rect 945 7639 954 7659
rect 910 7623 954 7639
rect 1024 7655 1073 7665
rect 1024 7635 1035 7655
rect 1055 7635 1073 7655
rect 1024 7623 1073 7635
rect 1123 7659 1167 7665
rect 1123 7639 1138 7659
rect 1158 7639 1167 7659
rect 1123 7623 1167 7639
rect 1232 7655 1281 7665
rect 1232 7635 1243 7655
rect 1263 7635 1281 7655
rect 1232 7623 1281 7635
rect 1331 7659 1375 7665
rect 1331 7639 1346 7659
rect 1366 7639 1375 7659
rect 1331 7623 1375 7639
rect 1445 7659 1489 7665
rect 1445 7639 1454 7659
rect 1474 7639 1489 7659
rect 1445 7623 1489 7639
rect 1539 7655 1588 7665
rect 9101 7752 9150 7762
rect 9200 7778 9244 7794
rect 9200 7758 9215 7778
rect 9235 7758 9244 7778
rect 9200 7752 9244 7758
rect 9314 7778 9358 7794
rect 9314 7758 9323 7778
rect 9343 7758 9358 7778
rect 9314 7752 9358 7758
rect 9408 7782 9457 7794
rect 9408 7762 9426 7782
rect 9446 7762 9457 7782
rect 9408 7752 9457 7762
rect 9522 7778 9566 7794
rect 9522 7758 9531 7778
rect 9551 7758 9566 7778
rect 9522 7752 9566 7758
rect 9616 7782 9665 7794
rect 9616 7762 9634 7782
rect 9654 7762 9665 7782
rect 9616 7752 9665 7762
rect 9735 7778 9779 7794
rect 9735 7758 9744 7778
rect 9764 7758 9779 7778
rect 9735 7752 9779 7758
rect 9829 7782 9878 7794
rect 9829 7762 9847 7782
rect 9867 7762 9878 7782
rect 9829 7752 9878 7762
rect 1539 7635 1557 7655
rect 1577 7635 1588 7655
rect 1539 7623 1588 7635
rect 4414 7646 4463 7656
rect 4414 7626 4425 7646
rect 4445 7626 4463 7646
rect 4414 7614 4463 7626
rect 4513 7650 4557 7656
rect 4513 7630 4528 7650
rect 4548 7630 4557 7650
rect 4513 7614 4557 7630
rect 4627 7646 4676 7656
rect 4627 7626 4638 7646
rect 4658 7626 4676 7646
rect 4627 7614 4676 7626
rect 4726 7650 4770 7656
rect 4726 7630 4741 7650
rect 4761 7630 4770 7650
rect 4726 7614 4770 7630
rect 4835 7646 4884 7656
rect 4835 7626 4846 7646
rect 4866 7626 4884 7646
rect 4835 7614 4884 7626
rect 4934 7650 4978 7656
rect 4934 7630 4949 7650
rect 4969 7630 4978 7650
rect 4934 7614 4978 7630
rect 5048 7650 5092 7656
rect 5048 7630 5057 7650
rect 5077 7630 5092 7650
rect 5048 7614 5092 7630
rect 5142 7646 5191 7656
rect 5142 7626 5160 7646
rect 5180 7626 5191 7646
rect 5142 7614 5191 7626
rect 18761 7780 18810 7792
rect 18761 7760 18772 7780
rect 18792 7760 18810 7780
rect 18761 7750 18810 7760
rect 18860 7776 18904 7792
rect 18860 7756 18875 7776
rect 18895 7756 18904 7776
rect 18860 7750 18904 7756
rect 18974 7776 19018 7792
rect 18974 7756 18983 7776
rect 19003 7756 19018 7776
rect 18974 7750 19018 7756
rect 19068 7780 19117 7792
rect 19068 7760 19086 7780
rect 19106 7760 19117 7780
rect 19068 7750 19117 7760
rect 19182 7776 19226 7792
rect 19182 7756 19191 7776
rect 19211 7756 19226 7776
rect 19182 7750 19226 7756
rect 19276 7780 19325 7792
rect 19276 7760 19294 7780
rect 19314 7760 19325 7780
rect 19276 7750 19325 7760
rect 19395 7776 19439 7792
rect 19395 7756 19404 7776
rect 19424 7756 19439 7776
rect 19395 7750 19439 7756
rect 19489 7780 19538 7792
rect 19489 7760 19507 7780
rect 19527 7760 19538 7780
rect 19489 7750 19538 7760
rect 19809 7776 19858 7788
rect 19809 7756 19820 7776
rect 19840 7756 19858 7776
rect 11519 7649 11568 7659
rect 11519 7629 11530 7649
rect 11550 7629 11568 7649
rect 11519 7617 11568 7629
rect 11618 7653 11662 7659
rect 11618 7633 11633 7653
rect 11653 7633 11662 7653
rect 11618 7617 11662 7633
rect 11732 7649 11781 7659
rect 11732 7629 11743 7649
rect 11763 7629 11781 7649
rect 11732 7617 11781 7629
rect 11831 7653 11875 7659
rect 11831 7633 11846 7653
rect 11866 7633 11875 7653
rect 11831 7617 11875 7633
rect 11940 7649 11989 7659
rect 11940 7629 11951 7649
rect 11971 7629 11989 7649
rect 11940 7617 11989 7629
rect 12039 7653 12083 7659
rect 12039 7633 12054 7653
rect 12074 7633 12083 7653
rect 12039 7617 12083 7633
rect 12153 7653 12197 7659
rect 12153 7633 12162 7653
rect 12182 7633 12197 7653
rect 12153 7617 12197 7633
rect 12247 7649 12296 7659
rect 19809 7746 19858 7756
rect 19908 7772 19952 7788
rect 19908 7752 19923 7772
rect 19943 7752 19952 7772
rect 19908 7746 19952 7752
rect 20022 7772 20066 7788
rect 20022 7752 20031 7772
rect 20051 7752 20066 7772
rect 20022 7746 20066 7752
rect 20116 7776 20165 7788
rect 20116 7756 20134 7776
rect 20154 7756 20165 7776
rect 20116 7746 20165 7756
rect 20230 7772 20274 7788
rect 20230 7752 20239 7772
rect 20259 7752 20274 7772
rect 20230 7746 20274 7752
rect 20324 7776 20373 7788
rect 20324 7756 20342 7776
rect 20362 7756 20373 7776
rect 20324 7746 20373 7756
rect 20443 7772 20487 7788
rect 20443 7752 20452 7772
rect 20472 7752 20487 7772
rect 20443 7746 20487 7752
rect 20537 7776 20586 7788
rect 20537 7756 20555 7776
rect 20575 7756 20586 7776
rect 20537 7746 20586 7756
rect 12247 7629 12265 7649
rect 12285 7629 12296 7649
rect 12247 7617 12296 7629
rect 15122 7640 15171 7650
rect 15122 7620 15133 7640
rect 15153 7620 15171 7640
rect 15122 7608 15171 7620
rect 15221 7644 15265 7650
rect 15221 7624 15236 7644
rect 15256 7624 15265 7644
rect 15221 7608 15265 7624
rect 15335 7640 15384 7650
rect 15335 7620 15346 7640
rect 15366 7620 15384 7640
rect 15335 7608 15384 7620
rect 15434 7644 15478 7650
rect 15434 7624 15449 7644
rect 15469 7624 15478 7644
rect 15434 7608 15478 7624
rect 15543 7640 15592 7650
rect 15543 7620 15554 7640
rect 15574 7620 15592 7640
rect 15543 7608 15592 7620
rect 15642 7644 15686 7650
rect 15642 7624 15657 7644
rect 15677 7624 15686 7644
rect 15642 7608 15686 7624
rect 15756 7644 15800 7650
rect 15756 7624 15765 7644
rect 15785 7624 15800 7644
rect 15756 7608 15800 7624
rect 15850 7640 15899 7650
rect 15850 7620 15868 7640
rect 15888 7620 15899 7640
rect 15850 7608 15899 7620
rect 5495 6876 5544 6888
rect 5495 6856 5506 6876
rect 5526 6856 5544 6876
rect 5495 6846 5544 6856
rect 5594 6872 5638 6888
rect 5594 6852 5609 6872
rect 5629 6852 5638 6872
rect 5594 6846 5638 6852
rect 5708 6872 5752 6888
rect 5708 6852 5717 6872
rect 5737 6852 5752 6872
rect 5708 6846 5752 6852
rect 5802 6876 5851 6888
rect 5802 6856 5820 6876
rect 5840 6856 5851 6876
rect 5802 6846 5851 6856
rect 5916 6872 5960 6888
rect 5916 6852 5925 6872
rect 5945 6852 5960 6872
rect 5916 6846 5960 6852
rect 6010 6876 6059 6888
rect 6010 6856 6028 6876
rect 6048 6856 6059 6876
rect 6010 6846 6059 6856
rect 6129 6872 6173 6888
rect 6129 6852 6138 6872
rect 6158 6852 6173 6872
rect 6129 6846 6173 6852
rect 6223 6876 6272 6888
rect 6223 6856 6241 6876
rect 6261 6856 6272 6876
rect 6223 6846 6272 6856
rect 9098 6867 9147 6879
rect 9098 6847 9109 6867
rect 9129 6847 9147 6867
rect 808 6740 857 6750
rect 808 6720 819 6740
rect 839 6720 857 6740
rect 808 6708 857 6720
rect 907 6744 951 6750
rect 907 6724 922 6744
rect 942 6724 951 6744
rect 907 6708 951 6724
rect 1021 6740 1070 6750
rect 1021 6720 1032 6740
rect 1052 6720 1070 6740
rect 1021 6708 1070 6720
rect 1120 6744 1164 6750
rect 1120 6724 1135 6744
rect 1155 6724 1164 6744
rect 1120 6708 1164 6724
rect 1229 6740 1278 6750
rect 1229 6720 1240 6740
rect 1260 6720 1278 6740
rect 1229 6708 1278 6720
rect 1328 6744 1372 6750
rect 1328 6724 1343 6744
rect 1363 6724 1372 6744
rect 1328 6708 1372 6724
rect 1442 6744 1486 6750
rect 1442 6724 1451 6744
rect 1471 6724 1486 6744
rect 1442 6708 1486 6724
rect 1536 6740 1585 6750
rect 9098 6837 9147 6847
rect 9197 6863 9241 6879
rect 9197 6843 9212 6863
rect 9232 6843 9241 6863
rect 9197 6837 9241 6843
rect 9311 6863 9355 6879
rect 9311 6843 9320 6863
rect 9340 6843 9355 6863
rect 9311 6837 9355 6843
rect 9405 6867 9454 6879
rect 9405 6847 9423 6867
rect 9443 6847 9454 6867
rect 9405 6837 9454 6847
rect 9519 6863 9563 6879
rect 9519 6843 9528 6863
rect 9548 6843 9563 6863
rect 9519 6837 9563 6843
rect 9613 6867 9662 6879
rect 9613 6847 9631 6867
rect 9651 6847 9662 6867
rect 9613 6837 9662 6847
rect 9732 6863 9776 6879
rect 9732 6843 9741 6863
rect 9761 6843 9776 6863
rect 9732 6837 9776 6843
rect 9826 6867 9875 6879
rect 9826 6847 9844 6867
rect 9864 6847 9875 6867
rect 9826 6837 9875 6847
rect 1536 6720 1554 6740
rect 1574 6720 1585 6740
rect 1536 6708 1585 6720
rect 1856 6736 1905 6746
rect 1856 6716 1867 6736
rect 1887 6716 1905 6736
rect 1856 6704 1905 6716
rect 1955 6740 1999 6746
rect 1955 6720 1970 6740
rect 1990 6720 1999 6740
rect 1955 6704 1999 6720
rect 2069 6736 2118 6746
rect 2069 6716 2080 6736
rect 2100 6716 2118 6736
rect 2069 6704 2118 6716
rect 2168 6740 2212 6746
rect 2168 6720 2183 6740
rect 2203 6720 2212 6740
rect 2168 6704 2212 6720
rect 2277 6736 2326 6746
rect 2277 6716 2288 6736
rect 2308 6716 2326 6736
rect 2277 6704 2326 6716
rect 2376 6740 2420 6746
rect 2376 6720 2391 6740
rect 2411 6720 2420 6740
rect 2376 6704 2420 6720
rect 2490 6740 2534 6746
rect 2490 6720 2499 6740
rect 2519 6720 2534 6740
rect 2490 6704 2534 6720
rect 2584 6736 2633 6746
rect 2584 6716 2602 6736
rect 2622 6716 2633 6736
rect 2584 6704 2633 6716
rect 16203 6870 16252 6882
rect 16203 6850 16214 6870
rect 16234 6850 16252 6870
rect 16203 6840 16252 6850
rect 16302 6866 16346 6882
rect 16302 6846 16317 6866
rect 16337 6846 16346 6866
rect 16302 6840 16346 6846
rect 16416 6866 16460 6882
rect 16416 6846 16425 6866
rect 16445 6846 16460 6866
rect 16416 6840 16460 6846
rect 16510 6870 16559 6882
rect 16510 6850 16528 6870
rect 16548 6850 16559 6870
rect 16510 6840 16559 6850
rect 16624 6866 16668 6882
rect 16624 6846 16633 6866
rect 16653 6846 16668 6866
rect 16624 6840 16668 6846
rect 16718 6870 16767 6882
rect 16718 6850 16736 6870
rect 16756 6850 16767 6870
rect 16718 6840 16767 6850
rect 16837 6866 16881 6882
rect 16837 6846 16846 6866
rect 16866 6846 16881 6866
rect 16837 6840 16881 6846
rect 16931 6870 16980 6882
rect 16931 6850 16949 6870
rect 16969 6850 16980 6870
rect 16931 6840 16980 6850
rect 19806 6861 19855 6873
rect 19806 6841 19817 6861
rect 19837 6841 19855 6861
rect 11516 6734 11565 6744
rect 11516 6714 11527 6734
rect 11547 6714 11565 6734
rect 11516 6702 11565 6714
rect 11615 6738 11659 6744
rect 11615 6718 11630 6738
rect 11650 6718 11659 6738
rect 11615 6702 11659 6718
rect 11729 6734 11778 6744
rect 11729 6714 11740 6734
rect 11760 6714 11778 6734
rect 11729 6702 11778 6714
rect 11828 6738 11872 6744
rect 11828 6718 11843 6738
rect 11863 6718 11872 6738
rect 11828 6702 11872 6718
rect 11937 6734 11986 6744
rect 11937 6714 11948 6734
rect 11968 6714 11986 6734
rect 11937 6702 11986 6714
rect 12036 6738 12080 6744
rect 12036 6718 12051 6738
rect 12071 6718 12080 6738
rect 12036 6702 12080 6718
rect 12150 6738 12194 6744
rect 12150 6718 12159 6738
rect 12179 6718 12194 6738
rect 12150 6702 12194 6718
rect 12244 6734 12293 6744
rect 19806 6831 19855 6841
rect 19905 6857 19949 6873
rect 19905 6837 19920 6857
rect 19940 6837 19949 6857
rect 19905 6831 19949 6837
rect 20019 6857 20063 6873
rect 20019 6837 20028 6857
rect 20048 6837 20063 6857
rect 20019 6831 20063 6837
rect 20113 6861 20162 6873
rect 20113 6841 20131 6861
rect 20151 6841 20162 6861
rect 20113 6831 20162 6841
rect 20227 6857 20271 6873
rect 20227 6837 20236 6857
rect 20256 6837 20271 6857
rect 20227 6831 20271 6837
rect 20321 6861 20370 6873
rect 20321 6841 20339 6861
rect 20359 6841 20370 6861
rect 20321 6831 20370 6841
rect 20440 6857 20484 6873
rect 20440 6837 20449 6857
rect 20469 6837 20484 6857
rect 20440 6831 20484 6837
rect 20534 6861 20583 6873
rect 20534 6841 20552 6861
rect 20572 6841 20583 6861
rect 20534 6831 20583 6841
rect 12244 6714 12262 6734
rect 12282 6714 12293 6734
rect 12244 6702 12293 6714
rect 12564 6730 12613 6740
rect 12564 6710 12575 6730
rect 12595 6710 12613 6730
rect 12564 6698 12613 6710
rect 12663 6734 12707 6740
rect 12663 6714 12678 6734
rect 12698 6714 12707 6734
rect 12663 6698 12707 6714
rect 12777 6730 12826 6740
rect 12777 6710 12788 6730
rect 12808 6710 12826 6730
rect 12777 6698 12826 6710
rect 12876 6734 12920 6740
rect 12876 6714 12891 6734
rect 12911 6714 12920 6734
rect 12876 6698 12920 6714
rect 12985 6730 13034 6740
rect 12985 6710 12996 6730
rect 13016 6710 13034 6730
rect 12985 6698 13034 6710
rect 13084 6734 13128 6740
rect 13084 6714 13099 6734
rect 13119 6714 13128 6734
rect 13084 6698 13128 6714
rect 13198 6734 13242 6740
rect 13198 6714 13207 6734
rect 13227 6714 13242 6734
rect 13198 6698 13242 6714
rect 13292 6730 13341 6740
rect 13292 6710 13310 6730
rect 13330 6710 13341 6730
rect 13292 6698 13341 6710
rect 8050 6192 8099 6204
rect 8050 6172 8061 6192
rect 8081 6172 8099 6192
rect 8050 6162 8099 6172
rect 8149 6188 8193 6204
rect 8149 6168 8164 6188
rect 8184 6168 8193 6188
rect 8149 6162 8193 6168
rect 8263 6188 8307 6204
rect 8263 6168 8272 6188
rect 8292 6168 8307 6188
rect 8263 6162 8307 6168
rect 8357 6192 8406 6204
rect 8357 6172 8375 6192
rect 8395 6172 8406 6192
rect 8357 6162 8406 6172
rect 8471 6188 8515 6204
rect 8471 6168 8480 6188
rect 8500 6168 8515 6188
rect 8471 6162 8515 6168
rect 8565 6192 8614 6204
rect 8565 6172 8583 6192
rect 8603 6172 8614 6192
rect 8565 6162 8614 6172
rect 8684 6188 8728 6204
rect 8684 6168 8693 6188
rect 8713 6168 8728 6188
rect 8684 6162 8728 6168
rect 8778 6192 8827 6204
rect 8778 6172 8796 6192
rect 8816 6172 8827 6192
rect 8778 6162 8827 6172
rect 9098 6188 9147 6200
rect 9098 6168 9109 6188
rect 9129 6168 9147 6188
rect 808 6061 857 6071
rect 808 6041 819 6061
rect 839 6041 857 6061
rect 808 6029 857 6041
rect 907 6065 951 6071
rect 907 6045 922 6065
rect 942 6045 951 6065
rect 907 6029 951 6045
rect 1021 6061 1070 6071
rect 1021 6041 1032 6061
rect 1052 6041 1070 6061
rect 1021 6029 1070 6041
rect 1120 6065 1164 6071
rect 1120 6045 1135 6065
rect 1155 6045 1164 6065
rect 1120 6029 1164 6045
rect 1229 6061 1278 6071
rect 1229 6041 1240 6061
rect 1260 6041 1278 6061
rect 1229 6029 1278 6041
rect 1328 6065 1372 6071
rect 1328 6045 1343 6065
rect 1363 6045 1372 6065
rect 1328 6029 1372 6045
rect 1442 6065 1486 6071
rect 1442 6045 1451 6065
rect 1471 6045 1486 6065
rect 1442 6029 1486 6045
rect 1536 6061 1585 6071
rect 9098 6158 9147 6168
rect 9197 6184 9241 6200
rect 9197 6164 9212 6184
rect 9232 6164 9241 6184
rect 9197 6158 9241 6164
rect 9311 6184 9355 6200
rect 9311 6164 9320 6184
rect 9340 6164 9355 6184
rect 9311 6158 9355 6164
rect 9405 6188 9454 6200
rect 9405 6168 9423 6188
rect 9443 6168 9454 6188
rect 9405 6158 9454 6168
rect 9519 6184 9563 6200
rect 9519 6164 9528 6184
rect 9548 6164 9563 6184
rect 9519 6158 9563 6164
rect 9613 6188 9662 6200
rect 9613 6168 9631 6188
rect 9651 6168 9662 6188
rect 9613 6158 9662 6168
rect 9732 6184 9776 6200
rect 9732 6164 9741 6184
rect 9761 6164 9776 6184
rect 9732 6158 9776 6164
rect 9826 6188 9875 6200
rect 9826 6168 9844 6188
rect 9864 6168 9875 6188
rect 9826 6158 9875 6168
rect 1536 6041 1554 6061
rect 1574 6041 1585 6061
rect 1536 6029 1585 6041
rect 3303 6056 3352 6066
rect 3303 6036 3314 6056
rect 3334 6036 3352 6056
rect 3303 6024 3352 6036
rect 3402 6060 3446 6066
rect 3402 6040 3417 6060
rect 3437 6040 3446 6060
rect 3402 6024 3446 6040
rect 3516 6056 3565 6066
rect 3516 6036 3527 6056
rect 3547 6036 3565 6056
rect 3516 6024 3565 6036
rect 3615 6060 3659 6066
rect 3615 6040 3630 6060
rect 3650 6040 3659 6060
rect 3615 6024 3659 6040
rect 3724 6056 3773 6066
rect 3724 6036 3735 6056
rect 3755 6036 3773 6056
rect 3724 6024 3773 6036
rect 3823 6060 3867 6066
rect 3823 6040 3838 6060
rect 3858 6040 3867 6060
rect 3823 6024 3867 6040
rect 3937 6060 3981 6066
rect 3937 6040 3946 6060
rect 3966 6040 3981 6060
rect 3937 6024 3981 6040
rect 4031 6056 4080 6066
rect 4031 6036 4049 6056
rect 4069 6036 4080 6056
rect 4031 6024 4080 6036
rect 18758 6186 18807 6198
rect 18758 6166 18769 6186
rect 18789 6166 18807 6186
rect 18758 6156 18807 6166
rect 18857 6182 18901 6198
rect 18857 6162 18872 6182
rect 18892 6162 18901 6182
rect 18857 6156 18901 6162
rect 18971 6182 19015 6198
rect 18971 6162 18980 6182
rect 19000 6162 19015 6182
rect 18971 6156 19015 6162
rect 19065 6186 19114 6198
rect 19065 6166 19083 6186
rect 19103 6166 19114 6186
rect 19065 6156 19114 6166
rect 19179 6182 19223 6198
rect 19179 6162 19188 6182
rect 19208 6162 19223 6182
rect 19179 6156 19223 6162
rect 19273 6186 19322 6198
rect 19273 6166 19291 6186
rect 19311 6166 19322 6186
rect 19273 6156 19322 6166
rect 19392 6182 19436 6198
rect 19392 6162 19401 6182
rect 19421 6162 19436 6182
rect 19392 6156 19436 6162
rect 19486 6186 19535 6198
rect 19486 6166 19504 6186
rect 19524 6166 19535 6186
rect 19486 6156 19535 6166
rect 19806 6182 19855 6194
rect 19806 6162 19817 6182
rect 19837 6162 19855 6182
rect 11516 6055 11565 6065
rect 11516 6035 11527 6055
rect 11547 6035 11565 6055
rect 11516 6023 11565 6035
rect 11615 6059 11659 6065
rect 11615 6039 11630 6059
rect 11650 6039 11659 6059
rect 11615 6023 11659 6039
rect 11729 6055 11778 6065
rect 11729 6035 11740 6055
rect 11760 6035 11778 6055
rect 11729 6023 11778 6035
rect 11828 6059 11872 6065
rect 11828 6039 11843 6059
rect 11863 6039 11872 6059
rect 11828 6023 11872 6039
rect 11937 6055 11986 6065
rect 11937 6035 11948 6055
rect 11968 6035 11986 6055
rect 11937 6023 11986 6035
rect 12036 6059 12080 6065
rect 12036 6039 12051 6059
rect 12071 6039 12080 6059
rect 12036 6023 12080 6039
rect 12150 6059 12194 6065
rect 12150 6039 12159 6059
rect 12179 6039 12194 6059
rect 12150 6023 12194 6039
rect 12244 6055 12293 6065
rect 19806 6152 19855 6162
rect 19905 6178 19949 6194
rect 19905 6158 19920 6178
rect 19940 6158 19949 6178
rect 19905 6152 19949 6158
rect 20019 6178 20063 6194
rect 20019 6158 20028 6178
rect 20048 6158 20063 6178
rect 20019 6152 20063 6158
rect 20113 6182 20162 6194
rect 20113 6162 20131 6182
rect 20151 6162 20162 6182
rect 20113 6152 20162 6162
rect 20227 6178 20271 6194
rect 20227 6158 20236 6178
rect 20256 6158 20271 6178
rect 20227 6152 20271 6158
rect 20321 6182 20370 6194
rect 20321 6162 20339 6182
rect 20359 6162 20370 6182
rect 20321 6152 20370 6162
rect 20440 6178 20484 6194
rect 20440 6158 20449 6178
rect 20469 6158 20484 6178
rect 20440 6152 20484 6158
rect 20534 6182 20583 6194
rect 20534 6162 20552 6182
rect 20572 6162 20583 6182
rect 20534 6152 20583 6162
rect 12244 6035 12262 6055
rect 12282 6035 12293 6055
rect 12244 6023 12293 6035
rect 14011 6050 14060 6060
rect 14011 6030 14022 6050
rect 14042 6030 14060 6050
rect 14011 6018 14060 6030
rect 14110 6054 14154 6060
rect 14110 6034 14125 6054
rect 14145 6034 14154 6054
rect 14110 6018 14154 6034
rect 14224 6050 14273 6060
rect 14224 6030 14235 6050
rect 14255 6030 14273 6050
rect 14224 6018 14273 6030
rect 14323 6054 14367 6060
rect 14323 6034 14338 6054
rect 14358 6034 14367 6054
rect 14323 6018 14367 6034
rect 14432 6050 14481 6060
rect 14432 6030 14443 6050
rect 14463 6030 14481 6050
rect 14432 6018 14481 6030
rect 14531 6054 14575 6060
rect 14531 6034 14546 6054
rect 14566 6034 14575 6054
rect 14531 6018 14575 6034
rect 14645 6054 14689 6060
rect 14645 6034 14654 6054
rect 14674 6034 14689 6054
rect 14645 6018 14689 6034
rect 14739 6050 14788 6060
rect 14739 6030 14757 6050
rect 14777 6030 14788 6050
rect 14739 6018 14788 6030
rect 6603 5425 6652 5437
rect 6603 5405 6614 5425
rect 6634 5405 6652 5425
rect 6603 5395 6652 5405
rect 6702 5421 6746 5437
rect 6702 5401 6717 5421
rect 6737 5401 6746 5421
rect 6702 5395 6746 5401
rect 6816 5421 6860 5437
rect 6816 5401 6825 5421
rect 6845 5401 6860 5421
rect 6816 5395 6860 5401
rect 6910 5425 6959 5437
rect 6910 5405 6928 5425
rect 6948 5405 6959 5425
rect 6910 5395 6959 5405
rect 7024 5421 7068 5437
rect 7024 5401 7033 5421
rect 7053 5401 7068 5421
rect 7024 5395 7068 5401
rect 7118 5425 7167 5437
rect 7118 5405 7136 5425
rect 7156 5405 7167 5425
rect 7118 5395 7167 5405
rect 7237 5421 7281 5437
rect 7237 5401 7246 5421
rect 7266 5401 7281 5421
rect 7237 5395 7281 5401
rect 7331 5425 7380 5437
rect 7331 5405 7349 5425
rect 7369 5405 7380 5425
rect 7331 5395 7380 5405
rect 9098 5420 9147 5432
rect 9098 5400 9109 5420
rect 9129 5400 9147 5420
rect 808 5293 857 5303
rect 808 5273 819 5293
rect 839 5273 857 5293
rect 808 5261 857 5273
rect 907 5297 951 5303
rect 907 5277 922 5297
rect 942 5277 951 5297
rect 907 5261 951 5277
rect 1021 5293 1070 5303
rect 1021 5273 1032 5293
rect 1052 5273 1070 5293
rect 1021 5261 1070 5273
rect 1120 5297 1164 5303
rect 1120 5277 1135 5297
rect 1155 5277 1164 5297
rect 1120 5261 1164 5277
rect 1229 5293 1278 5303
rect 1229 5273 1240 5293
rect 1260 5273 1278 5293
rect 1229 5261 1278 5273
rect 1328 5297 1372 5303
rect 1328 5277 1343 5297
rect 1363 5277 1372 5297
rect 1328 5261 1372 5277
rect 1442 5297 1486 5303
rect 1442 5277 1451 5297
rect 1471 5277 1486 5297
rect 1442 5261 1486 5277
rect 1536 5293 1585 5303
rect 9098 5390 9147 5400
rect 9197 5416 9241 5432
rect 9197 5396 9212 5416
rect 9232 5396 9241 5416
rect 9197 5390 9241 5396
rect 9311 5416 9355 5432
rect 9311 5396 9320 5416
rect 9340 5396 9355 5416
rect 9311 5390 9355 5396
rect 9405 5420 9454 5432
rect 9405 5400 9423 5420
rect 9443 5400 9454 5420
rect 9405 5390 9454 5400
rect 9519 5416 9563 5432
rect 9519 5396 9528 5416
rect 9548 5396 9563 5416
rect 9519 5390 9563 5396
rect 9613 5420 9662 5432
rect 9613 5400 9631 5420
rect 9651 5400 9662 5420
rect 9613 5390 9662 5400
rect 9732 5416 9776 5432
rect 9732 5396 9741 5416
rect 9761 5396 9776 5416
rect 9732 5390 9776 5396
rect 9826 5420 9875 5432
rect 9826 5400 9844 5420
rect 9864 5400 9875 5420
rect 9826 5390 9875 5400
rect 1536 5273 1554 5293
rect 1574 5273 1585 5293
rect 1536 5261 1585 5273
rect 1856 5289 1905 5299
rect 1856 5269 1867 5289
rect 1887 5269 1905 5289
rect 1856 5257 1905 5269
rect 1955 5293 1999 5299
rect 1955 5273 1970 5293
rect 1990 5273 1999 5293
rect 1955 5257 1999 5273
rect 2069 5289 2118 5299
rect 2069 5269 2080 5289
rect 2100 5269 2118 5289
rect 2069 5257 2118 5269
rect 2168 5293 2212 5299
rect 2168 5273 2183 5293
rect 2203 5273 2212 5293
rect 2168 5257 2212 5273
rect 2277 5289 2326 5299
rect 2277 5269 2288 5289
rect 2308 5269 2326 5289
rect 2277 5257 2326 5269
rect 2376 5293 2420 5299
rect 2376 5273 2391 5293
rect 2411 5273 2420 5293
rect 2376 5257 2420 5273
rect 2490 5293 2534 5299
rect 2490 5273 2499 5293
rect 2519 5273 2534 5293
rect 2490 5257 2534 5273
rect 2584 5289 2633 5299
rect 2584 5269 2602 5289
rect 2622 5269 2633 5289
rect 2584 5257 2633 5269
rect 17311 5419 17360 5431
rect 17311 5399 17322 5419
rect 17342 5399 17360 5419
rect 17311 5389 17360 5399
rect 17410 5415 17454 5431
rect 17410 5395 17425 5415
rect 17445 5395 17454 5415
rect 17410 5389 17454 5395
rect 17524 5415 17568 5431
rect 17524 5395 17533 5415
rect 17553 5395 17568 5415
rect 17524 5389 17568 5395
rect 17618 5419 17667 5431
rect 17618 5399 17636 5419
rect 17656 5399 17667 5419
rect 17618 5389 17667 5399
rect 17732 5415 17776 5431
rect 17732 5395 17741 5415
rect 17761 5395 17776 5415
rect 17732 5389 17776 5395
rect 17826 5419 17875 5431
rect 17826 5399 17844 5419
rect 17864 5399 17875 5419
rect 17826 5389 17875 5399
rect 17945 5415 17989 5431
rect 17945 5395 17954 5415
rect 17974 5395 17989 5415
rect 17945 5389 17989 5395
rect 18039 5419 18088 5431
rect 18039 5399 18057 5419
rect 18077 5399 18088 5419
rect 18039 5389 18088 5399
rect 19806 5414 19855 5426
rect 19806 5394 19817 5414
rect 19837 5394 19855 5414
rect 11516 5287 11565 5297
rect 11516 5267 11527 5287
rect 11547 5267 11565 5287
rect 11516 5255 11565 5267
rect 11615 5291 11659 5297
rect 11615 5271 11630 5291
rect 11650 5271 11659 5291
rect 11615 5255 11659 5271
rect 11729 5287 11778 5297
rect 11729 5267 11740 5287
rect 11760 5267 11778 5287
rect 11729 5255 11778 5267
rect 11828 5291 11872 5297
rect 11828 5271 11843 5291
rect 11863 5271 11872 5291
rect 11828 5255 11872 5271
rect 11937 5287 11986 5297
rect 11937 5267 11948 5287
rect 11968 5267 11986 5287
rect 11937 5255 11986 5267
rect 12036 5291 12080 5297
rect 12036 5271 12051 5291
rect 12071 5271 12080 5291
rect 12036 5255 12080 5271
rect 12150 5291 12194 5297
rect 12150 5271 12159 5291
rect 12179 5271 12194 5291
rect 12150 5255 12194 5271
rect 12244 5287 12293 5297
rect 19806 5384 19855 5394
rect 19905 5410 19949 5426
rect 19905 5390 19920 5410
rect 19940 5390 19949 5410
rect 19905 5384 19949 5390
rect 20019 5410 20063 5426
rect 20019 5390 20028 5410
rect 20048 5390 20063 5410
rect 20019 5384 20063 5390
rect 20113 5414 20162 5426
rect 20113 5394 20131 5414
rect 20151 5394 20162 5414
rect 20113 5384 20162 5394
rect 20227 5410 20271 5426
rect 20227 5390 20236 5410
rect 20256 5390 20271 5410
rect 20227 5384 20271 5390
rect 20321 5414 20370 5426
rect 20321 5394 20339 5414
rect 20359 5394 20370 5414
rect 20321 5384 20370 5394
rect 20440 5410 20484 5426
rect 20440 5390 20449 5410
rect 20469 5390 20484 5410
rect 20440 5384 20484 5390
rect 20534 5414 20583 5426
rect 20534 5394 20552 5414
rect 20572 5394 20583 5414
rect 20534 5384 20583 5394
rect 12244 5267 12262 5287
rect 12282 5267 12293 5287
rect 12244 5255 12293 5267
rect 12564 5283 12613 5293
rect 12564 5263 12575 5283
rect 12595 5263 12613 5283
rect 12564 5251 12613 5263
rect 12663 5287 12707 5293
rect 12663 5267 12678 5287
rect 12698 5267 12707 5287
rect 12663 5251 12707 5267
rect 12777 5283 12826 5293
rect 12777 5263 12788 5283
rect 12808 5263 12826 5283
rect 12777 5251 12826 5263
rect 12876 5287 12920 5293
rect 12876 5267 12891 5287
rect 12911 5267 12920 5287
rect 12876 5251 12920 5267
rect 12985 5283 13034 5293
rect 12985 5263 12996 5283
rect 13016 5263 13034 5283
rect 12985 5251 13034 5263
rect 13084 5287 13128 5293
rect 13084 5267 13099 5287
rect 13119 5267 13128 5287
rect 13084 5251 13128 5267
rect 13198 5287 13242 5293
rect 13198 5267 13207 5287
rect 13227 5267 13242 5287
rect 13198 5251 13242 5267
rect 13292 5283 13341 5293
rect 13292 5263 13310 5283
rect 13330 5263 13341 5283
rect 13292 5251 13341 5263
rect 8050 4745 8099 4757
rect 8050 4725 8061 4745
rect 8081 4725 8099 4745
rect 8050 4715 8099 4725
rect 8149 4741 8193 4757
rect 8149 4721 8164 4741
rect 8184 4721 8193 4741
rect 8149 4715 8193 4721
rect 8263 4741 8307 4757
rect 8263 4721 8272 4741
rect 8292 4721 8307 4741
rect 8263 4715 8307 4721
rect 8357 4745 8406 4757
rect 8357 4725 8375 4745
rect 8395 4725 8406 4745
rect 8357 4715 8406 4725
rect 8471 4741 8515 4757
rect 8471 4721 8480 4741
rect 8500 4721 8515 4741
rect 8471 4715 8515 4721
rect 8565 4745 8614 4757
rect 8565 4725 8583 4745
rect 8603 4725 8614 4745
rect 8565 4715 8614 4725
rect 8684 4741 8728 4757
rect 8684 4721 8693 4741
rect 8713 4721 8728 4741
rect 8684 4715 8728 4721
rect 8778 4745 8827 4757
rect 8778 4725 8796 4745
rect 8816 4725 8827 4745
rect 8778 4715 8827 4725
rect 9098 4741 9147 4753
rect 9098 4721 9109 4741
rect 9129 4721 9147 4741
rect 808 4614 857 4624
rect 808 4594 819 4614
rect 839 4594 857 4614
rect 808 4582 857 4594
rect 907 4618 951 4624
rect 907 4598 922 4618
rect 942 4598 951 4618
rect 907 4582 951 4598
rect 1021 4614 1070 4624
rect 1021 4594 1032 4614
rect 1052 4594 1070 4614
rect 1021 4582 1070 4594
rect 1120 4618 1164 4624
rect 1120 4598 1135 4618
rect 1155 4598 1164 4618
rect 1120 4582 1164 4598
rect 1229 4614 1278 4624
rect 1229 4594 1240 4614
rect 1260 4594 1278 4614
rect 1229 4582 1278 4594
rect 1328 4618 1372 4624
rect 1328 4598 1343 4618
rect 1363 4598 1372 4618
rect 1328 4582 1372 4598
rect 1442 4618 1486 4624
rect 1442 4598 1451 4618
rect 1471 4598 1486 4618
rect 1442 4582 1486 4598
rect 1536 4614 1585 4624
rect 9098 4711 9147 4721
rect 9197 4737 9241 4753
rect 9197 4717 9212 4737
rect 9232 4717 9241 4737
rect 9197 4711 9241 4717
rect 9311 4737 9355 4753
rect 9311 4717 9320 4737
rect 9340 4717 9355 4737
rect 9311 4711 9355 4717
rect 9405 4741 9454 4753
rect 9405 4721 9423 4741
rect 9443 4721 9454 4741
rect 9405 4711 9454 4721
rect 9519 4737 9563 4753
rect 9519 4717 9528 4737
rect 9548 4717 9563 4737
rect 9519 4711 9563 4717
rect 9613 4741 9662 4753
rect 9613 4721 9631 4741
rect 9651 4721 9662 4741
rect 9613 4711 9662 4721
rect 9732 4737 9776 4753
rect 9732 4717 9741 4737
rect 9761 4717 9776 4737
rect 9732 4711 9776 4717
rect 9826 4741 9875 4753
rect 9826 4721 9844 4741
rect 9864 4721 9875 4741
rect 9826 4711 9875 4721
rect 1536 4594 1554 4614
rect 1574 4594 1585 4614
rect 1536 4582 1585 4594
rect 3346 4611 3395 4621
rect 3346 4591 3357 4611
rect 3377 4591 3395 4611
rect 3346 4579 3395 4591
rect 3445 4615 3489 4621
rect 3445 4595 3460 4615
rect 3480 4595 3489 4615
rect 3445 4579 3489 4595
rect 3559 4611 3608 4621
rect 3559 4591 3570 4611
rect 3590 4591 3608 4611
rect 3559 4579 3608 4591
rect 3658 4615 3702 4621
rect 3658 4595 3673 4615
rect 3693 4595 3702 4615
rect 3658 4579 3702 4595
rect 3767 4611 3816 4621
rect 3767 4591 3778 4611
rect 3798 4591 3816 4611
rect 3767 4579 3816 4591
rect 3866 4615 3910 4621
rect 3866 4595 3881 4615
rect 3901 4595 3910 4615
rect 3866 4579 3910 4595
rect 3980 4615 4024 4621
rect 3980 4595 3989 4615
rect 4009 4595 4024 4615
rect 3980 4579 4024 4595
rect 4074 4611 4123 4621
rect 4074 4591 4092 4611
rect 4112 4591 4123 4611
rect 4074 4579 4123 4591
rect 18758 4739 18807 4751
rect 18758 4719 18769 4739
rect 18789 4719 18807 4739
rect 18758 4709 18807 4719
rect 18857 4735 18901 4751
rect 18857 4715 18872 4735
rect 18892 4715 18901 4735
rect 18857 4709 18901 4715
rect 18971 4735 19015 4751
rect 18971 4715 18980 4735
rect 19000 4715 19015 4735
rect 18971 4709 19015 4715
rect 19065 4739 19114 4751
rect 19065 4719 19083 4739
rect 19103 4719 19114 4739
rect 19065 4709 19114 4719
rect 19179 4735 19223 4751
rect 19179 4715 19188 4735
rect 19208 4715 19223 4735
rect 19179 4709 19223 4715
rect 19273 4739 19322 4751
rect 19273 4719 19291 4739
rect 19311 4719 19322 4739
rect 19273 4709 19322 4719
rect 19392 4735 19436 4751
rect 19392 4715 19401 4735
rect 19421 4715 19436 4735
rect 19392 4709 19436 4715
rect 19486 4739 19535 4751
rect 19486 4719 19504 4739
rect 19524 4719 19535 4739
rect 19486 4709 19535 4719
rect 19806 4735 19855 4747
rect 19806 4715 19817 4735
rect 19837 4715 19855 4735
rect 11516 4608 11565 4618
rect 11516 4588 11527 4608
rect 11547 4588 11565 4608
rect 11516 4576 11565 4588
rect 11615 4612 11659 4618
rect 11615 4592 11630 4612
rect 11650 4592 11659 4612
rect 11615 4576 11659 4592
rect 11729 4608 11778 4618
rect 11729 4588 11740 4608
rect 11760 4588 11778 4608
rect 11729 4576 11778 4588
rect 11828 4612 11872 4618
rect 11828 4592 11843 4612
rect 11863 4592 11872 4612
rect 11828 4576 11872 4592
rect 11937 4608 11986 4618
rect 11937 4588 11948 4608
rect 11968 4588 11986 4608
rect 11937 4576 11986 4588
rect 12036 4612 12080 4618
rect 12036 4592 12051 4612
rect 12071 4592 12080 4612
rect 12036 4576 12080 4592
rect 12150 4612 12194 4618
rect 12150 4592 12159 4612
rect 12179 4592 12194 4612
rect 12150 4576 12194 4592
rect 12244 4608 12293 4618
rect 19806 4705 19855 4715
rect 19905 4731 19949 4747
rect 19905 4711 19920 4731
rect 19940 4711 19949 4731
rect 19905 4705 19949 4711
rect 20019 4731 20063 4747
rect 20019 4711 20028 4731
rect 20048 4711 20063 4731
rect 20019 4705 20063 4711
rect 20113 4735 20162 4747
rect 20113 4715 20131 4735
rect 20151 4715 20162 4735
rect 20113 4705 20162 4715
rect 20227 4731 20271 4747
rect 20227 4711 20236 4731
rect 20256 4711 20271 4731
rect 20227 4705 20271 4711
rect 20321 4735 20370 4747
rect 20321 4715 20339 4735
rect 20359 4715 20370 4735
rect 20321 4705 20370 4715
rect 20440 4731 20484 4747
rect 20440 4711 20449 4731
rect 20469 4711 20484 4731
rect 20440 4705 20484 4711
rect 20534 4735 20583 4747
rect 20534 4715 20552 4735
rect 20572 4715 20583 4735
rect 20534 4705 20583 4715
rect 12244 4588 12262 4608
rect 12282 4588 12293 4608
rect 12244 4576 12293 4588
rect 14054 4605 14103 4615
rect 14054 4585 14065 4605
rect 14085 4585 14103 4605
rect 14054 4573 14103 4585
rect 14153 4609 14197 4615
rect 14153 4589 14168 4609
rect 14188 4589 14197 4609
rect 14153 4573 14197 4589
rect 14267 4605 14316 4615
rect 14267 4585 14278 4605
rect 14298 4585 14316 4605
rect 14267 4573 14316 4585
rect 14366 4609 14410 4615
rect 14366 4589 14381 4609
rect 14401 4589 14410 4609
rect 14366 4573 14410 4589
rect 14475 4605 14524 4615
rect 14475 4585 14486 4605
rect 14506 4585 14524 4605
rect 14475 4573 14524 4585
rect 14574 4609 14618 4615
rect 14574 4589 14589 4609
rect 14609 4589 14618 4609
rect 14574 4573 14618 4589
rect 14688 4609 14732 4615
rect 14688 4589 14697 4609
rect 14717 4589 14732 4609
rect 14688 4573 14732 4589
rect 14782 4605 14831 4615
rect 14782 4585 14800 4605
rect 14820 4585 14831 4605
rect 14782 4573 14831 4585
rect 6561 3903 6610 3915
rect 6561 3883 6572 3903
rect 6592 3883 6610 3903
rect 6561 3873 6610 3883
rect 6660 3899 6704 3915
rect 6660 3879 6675 3899
rect 6695 3879 6704 3899
rect 6660 3873 6704 3879
rect 6774 3899 6818 3915
rect 6774 3879 6783 3899
rect 6803 3879 6818 3899
rect 6774 3873 6818 3879
rect 6868 3903 6917 3915
rect 6868 3883 6886 3903
rect 6906 3883 6917 3903
rect 6868 3873 6917 3883
rect 6982 3899 7026 3915
rect 6982 3879 6991 3899
rect 7011 3879 7026 3899
rect 6982 3873 7026 3879
rect 7076 3903 7125 3915
rect 7076 3883 7094 3903
rect 7114 3883 7125 3903
rect 7076 3873 7125 3883
rect 7195 3899 7239 3915
rect 7195 3879 7204 3899
rect 7224 3879 7239 3899
rect 7195 3873 7239 3879
rect 7289 3903 7338 3915
rect 7289 3883 7307 3903
rect 7327 3883 7338 3903
rect 7289 3873 7338 3883
rect 9099 3900 9148 3912
rect 9099 3880 9110 3900
rect 9130 3880 9148 3900
rect 809 3773 858 3783
rect 809 3753 820 3773
rect 840 3753 858 3773
rect 809 3741 858 3753
rect 908 3777 952 3783
rect 908 3757 923 3777
rect 943 3757 952 3777
rect 908 3741 952 3757
rect 1022 3773 1071 3783
rect 1022 3753 1033 3773
rect 1053 3753 1071 3773
rect 1022 3741 1071 3753
rect 1121 3777 1165 3783
rect 1121 3757 1136 3777
rect 1156 3757 1165 3777
rect 1121 3741 1165 3757
rect 1230 3773 1279 3783
rect 1230 3753 1241 3773
rect 1261 3753 1279 3773
rect 1230 3741 1279 3753
rect 1329 3777 1373 3783
rect 1329 3757 1344 3777
rect 1364 3757 1373 3777
rect 1329 3741 1373 3757
rect 1443 3777 1487 3783
rect 1443 3757 1452 3777
rect 1472 3757 1487 3777
rect 1443 3741 1487 3757
rect 1537 3773 1586 3783
rect 9099 3870 9148 3880
rect 9198 3896 9242 3912
rect 9198 3876 9213 3896
rect 9233 3876 9242 3896
rect 9198 3870 9242 3876
rect 9312 3896 9356 3912
rect 9312 3876 9321 3896
rect 9341 3876 9356 3896
rect 9312 3870 9356 3876
rect 9406 3900 9455 3912
rect 9406 3880 9424 3900
rect 9444 3880 9455 3900
rect 9406 3870 9455 3880
rect 9520 3896 9564 3912
rect 9520 3876 9529 3896
rect 9549 3876 9564 3896
rect 9520 3870 9564 3876
rect 9614 3900 9663 3912
rect 9614 3880 9632 3900
rect 9652 3880 9663 3900
rect 9614 3870 9663 3880
rect 9733 3896 9777 3912
rect 9733 3876 9742 3896
rect 9762 3876 9777 3896
rect 9733 3870 9777 3876
rect 9827 3900 9876 3912
rect 9827 3880 9845 3900
rect 9865 3880 9876 3900
rect 9827 3870 9876 3880
rect 1537 3753 1555 3773
rect 1575 3753 1586 3773
rect 1537 3741 1586 3753
rect 1857 3769 1906 3779
rect 1857 3749 1868 3769
rect 1888 3749 1906 3769
rect 1857 3737 1906 3749
rect 1956 3773 2000 3779
rect 1956 3753 1971 3773
rect 1991 3753 2000 3773
rect 1956 3737 2000 3753
rect 2070 3769 2119 3779
rect 2070 3749 2081 3769
rect 2101 3749 2119 3769
rect 2070 3737 2119 3749
rect 2169 3773 2213 3779
rect 2169 3753 2184 3773
rect 2204 3753 2213 3773
rect 2169 3737 2213 3753
rect 2278 3769 2327 3779
rect 2278 3749 2289 3769
rect 2309 3749 2327 3769
rect 2278 3737 2327 3749
rect 2377 3773 2421 3779
rect 2377 3753 2392 3773
rect 2412 3753 2421 3773
rect 2377 3737 2421 3753
rect 2491 3773 2535 3779
rect 2491 3753 2500 3773
rect 2520 3753 2535 3773
rect 2491 3737 2535 3753
rect 2585 3769 2634 3779
rect 2585 3749 2603 3769
rect 2623 3749 2634 3769
rect 2585 3737 2634 3749
rect 4759 3775 4808 3785
rect 4759 3755 4770 3775
rect 4790 3755 4808 3775
rect 4759 3743 4808 3755
rect 4858 3779 4902 3785
rect 4858 3759 4873 3779
rect 4893 3759 4902 3779
rect 4858 3743 4902 3759
rect 4972 3775 5021 3785
rect 4972 3755 4983 3775
rect 5003 3755 5021 3775
rect 4972 3743 5021 3755
rect 5071 3779 5115 3785
rect 5071 3759 5086 3779
rect 5106 3759 5115 3779
rect 5071 3743 5115 3759
rect 5180 3775 5229 3785
rect 5180 3755 5191 3775
rect 5211 3755 5229 3775
rect 5180 3743 5229 3755
rect 5279 3779 5323 3785
rect 5279 3759 5294 3779
rect 5314 3759 5323 3779
rect 5279 3743 5323 3759
rect 5393 3779 5437 3785
rect 5393 3759 5402 3779
rect 5422 3759 5437 3779
rect 5393 3743 5437 3759
rect 5487 3775 5536 3785
rect 5487 3755 5505 3775
rect 5525 3755 5536 3775
rect 5487 3743 5536 3755
rect 17269 3897 17318 3909
rect 17269 3877 17280 3897
rect 17300 3877 17318 3897
rect 17269 3867 17318 3877
rect 17368 3893 17412 3909
rect 17368 3873 17383 3893
rect 17403 3873 17412 3893
rect 17368 3867 17412 3873
rect 17482 3893 17526 3909
rect 17482 3873 17491 3893
rect 17511 3873 17526 3893
rect 17482 3867 17526 3873
rect 17576 3897 17625 3909
rect 17576 3877 17594 3897
rect 17614 3877 17625 3897
rect 17576 3867 17625 3877
rect 17690 3893 17734 3909
rect 17690 3873 17699 3893
rect 17719 3873 17734 3893
rect 17690 3867 17734 3873
rect 17784 3897 17833 3909
rect 17784 3877 17802 3897
rect 17822 3877 17833 3897
rect 17784 3867 17833 3877
rect 17903 3893 17947 3909
rect 17903 3873 17912 3893
rect 17932 3873 17947 3893
rect 17903 3867 17947 3873
rect 17997 3897 18046 3909
rect 17997 3877 18015 3897
rect 18035 3877 18046 3897
rect 17997 3867 18046 3877
rect 19807 3894 19856 3906
rect 19807 3874 19818 3894
rect 19838 3874 19856 3894
rect 11517 3767 11566 3777
rect 11517 3747 11528 3767
rect 11548 3747 11566 3767
rect 11517 3735 11566 3747
rect 11616 3771 11660 3777
rect 11616 3751 11631 3771
rect 11651 3751 11660 3771
rect 11616 3735 11660 3751
rect 11730 3767 11779 3777
rect 11730 3747 11741 3767
rect 11761 3747 11779 3767
rect 11730 3735 11779 3747
rect 11829 3771 11873 3777
rect 11829 3751 11844 3771
rect 11864 3751 11873 3771
rect 11829 3735 11873 3751
rect 11938 3767 11987 3777
rect 11938 3747 11949 3767
rect 11969 3747 11987 3767
rect 11938 3735 11987 3747
rect 12037 3771 12081 3777
rect 12037 3751 12052 3771
rect 12072 3751 12081 3771
rect 12037 3735 12081 3751
rect 12151 3771 12195 3777
rect 12151 3751 12160 3771
rect 12180 3751 12195 3771
rect 12151 3735 12195 3751
rect 12245 3767 12294 3777
rect 19807 3864 19856 3874
rect 19906 3890 19950 3906
rect 19906 3870 19921 3890
rect 19941 3870 19950 3890
rect 19906 3864 19950 3870
rect 20020 3890 20064 3906
rect 20020 3870 20029 3890
rect 20049 3870 20064 3890
rect 20020 3864 20064 3870
rect 20114 3894 20163 3906
rect 20114 3874 20132 3894
rect 20152 3874 20163 3894
rect 20114 3864 20163 3874
rect 20228 3890 20272 3906
rect 20228 3870 20237 3890
rect 20257 3870 20272 3890
rect 20228 3864 20272 3870
rect 20322 3894 20371 3906
rect 20322 3874 20340 3894
rect 20360 3874 20371 3894
rect 20322 3864 20371 3874
rect 20441 3890 20485 3906
rect 20441 3870 20450 3890
rect 20470 3870 20485 3890
rect 20441 3864 20485 3870
rect 20535 3894 20584 3906
rect 20535 3874 20553 3894
rect 20573 3874 20584 3894
rect 20535 3864 20584 3874
rect 12245 3747 12263 3767
rect 12283 3747 12294 3767
rect 12245 3735 12294 3747
rect 12565 3763 12614 3773
rect 12565 3743 12576 3763
rect 12596 3743 12614 3763
rect 12565 3731 12614 3743
rect 12664 3767 12708 3773
rect 12664 3747 12679 3767
rect 12699 3747 12708 3767
rect 12664 3731 12708 3747
rect 12778 3763 12827 3773
rect 12778 3743 12789 3763
rect 12809 3743 12827 3763
rect 12778 3731 12827 3743
rect 12877 3767 12921 3773
rect 12877 3747 12892 3767
rect 12912 3747 12921 3767
rect 12877 3731 12921 3747
rect 12986 3763 13035 3773
rect 12986 3743 12997 3763
rect 13017 3743 13035 3763
rect 12986 3731 13035 3743
rect 13085 3767 13129 3773
rect 13085 3747 13100 3767
rect 13120 3747 13129 3767
rect 13085 3731 13129 3747
rect 13199 3767 13243 3773
rect 13199 3747 13208 3767
rect 13228 3747 13243 3767
rect 13199 3731 13243 3747
rect 13293 3763 13342 3773
rect 13293 3743 13311 3763
rect 13331 3743 13342 3763
rect 13293 3731 13342 3743
rect 15467 3769 15516 3779
rect 15467 3749 15478 3769
rect 15498 3749 15516 3769
rect 15467 3737 15516 3749
rect 15566 3773 15610 3779
rect 15566 3753 15581 3773
rect 15601 3753 15610 3773
rect 15566 3737 15610 3753
rect 15680 3769 15729 3779
rect 15680 3749 15691 3769
rect 15711 3749 15729 3769
rect 15680 3737 15729 3749
rect 15779 3773 15823 3779
rect 15779 3753 15794 3773
rect 15814 3753 15823 3773
rect 15779 3737 15823 3753
rect 15888 3769 15937 3779
rect 15888 3749 15899 3769
rect 15919 3749 15937 3769
rect 15888 3737 15937 3749
rect 15987 3773 16031 3779
rect 15987 3753 16002 3773
rect 16022 3753 16031 3773
rect 15987 3737 16031 3753
rect 16101 3773 16145 3779
rect 16101 3753 16110 3773
rect 16130 3753 16145 3773
rect 16101 3737 16145 3753
rect 16195 3769 16244 3779
rect 16195 3749 16213 3769
rect 16233 3749 16244 3769
rect 16195 3737 16244 3749
rect 8051 3225 8100 3237
rect 8051 3205 8062 3225
rect 8082 3205 8100 3225
rect 8051 3195 8100 3205
rect 8150 3221 8194 3237
rect 8150 3201 8165 3221
rect 8185 3201 8194 3221
rect 8150 3195 8194 3201
rect 8264 3221 8308 3237
rect 8264 3201 8273 3221
rect 8293 3201 8308 3221
rect 8264 3195 8308 3201
rect 8358 3225 8407 3237
rect 8358 3205 8376 3225
rect 8396 3205 8407 3225
rect 8358 3195 8407 3205
rect 8472 3221 8516 3237
rect 8472 3201 8481 3221
rect 8501 3201 8516 3221
rect 8472 3195 8516 3201
rect 8566 3225 8615 3237
rect 8566 3205 8584 3225
rect 8604 3205 8615 3225
rect 8566 3195 8615 3205
rect 8685 3221 8729 3237
rect 8685 3201 8694 3221
rect 8714 3201 8729 3221
rect 8685 3195 8729 3201
rect 8779 3225 8828 3237
rect 8779 3205 8797 3225
rect 8817 3205 8828 3225
rect 8779 3195 8828 3205
rect 9099 3221 9148 3233
rect 9099 3201 9110 3221
rect 9130 3201 9148 3221
rect 809 3094 858 3104
rect 809 3074 820 3094
rect 840 3074 858 3094
rect 809 3062 858 3074
rect 908 3098 952 3104
rect 908 3078 923 3098
rect 943 3078 952 3098
rect 908 3062 952 3078
rect 1022 3094 1071 3104
rect 1022 3074 1033 3094
rect 1053 3074 1071 3094
rect 1022 3062 1071 3074
rect 1121 3098 1165 3104
rect 1121 3078 1136 3098
rect 1156 3078 1165 3098
rect 1121 3062 1165 3078
rect 1230 3094 1279 3104
rect 1230 3074 1241 3094
rect 1261 3074 1279 3094
rect 1230 3062 1279 3074
rect 1329 3098 1373 3104
rect 1329 3078 1344 3098
rect 1364 3078 1373 3098
rect 1329 3062 1373 3078
rect 1443 3098 1487 3104
rect 1443 3078 1452 3098
rect 1472 3078 1487 3098
rect 1443 3062 1487 3078
rect 1537 3094 1586 3104
rect 9099 3191 9148 3201
rect 9198 3217 9242 3233
rect 9198 3197 9213 3217
rect 9233 3197 9242 3217
rect 9198 3191 9242 3197
rect 9312 3217 9356 3233
rect 9312 3197 9321 3217
rect 9341 3197 9356 3217
rect 9312 3191 9356 3197
rect 9406 3221 9455 3233
rect 9406 3201 9424 3221
rect 9444 3201 9455 3221
rect 9406 3191 9455 3201
rect 9520 3217 9564 3233
rect 9520 3197 9529 3217
rect 9549 3197 9564 3217
rect 9520 3191 9564 3197
rect 9614 3221 9663 3233
rect 9614 3201 9632 3221
rect 9652 3201 9663 3221
rect 9614 3191 9663 3201
rect 9733 3217 9777 3233
rect 9733 3197 9742 3217
rect 9762 3197 9777 3217
rect 9733 3191 9777 3197
rect 9827 3221 9876 3233
rect 9827 3201 9845 3221
rect 9865 3201 9876 3221
rect 9827 3191 9876 3201
rect 1537 3074 1555 3094
rect 1575 3074 1586 3094
rect 1537 3062 1586 3074
rect 3304 3089 3353 3099
rect 3304 3069 3315 3089
rect 3335 3069 3353 3089
rect 3304 3057 3353 3069
rect 3403 3093 3447 3099
rect 3403 3073 3418 3093
rect 3438 3073 3447 3093
rect 3403 3057 3447 3073
rect 3517 3089 3566 3099
rect 3517 3069 3528 3089
rect 3548 3069 3566 3089
rect 3517 3057 3566 3069
rect 3616 3093 3660 3099
rect 3616 3073 3631 3093
rect 3651 3073 3660 3093
rect 3616 3057 3660 3073
rect 3725 3089 3774 3099
rect 3725 3069 3736 3089
rect 3756 3069 3774 3089
rect 3725 3057 3774 3069
rect 3824 3093 3868 3099
rect 3824 3073 3839 3093
rect 3859 3073 3868 3093
rect 3824 3057 3868 3073
rect 3938 3093 3982 3099
rect 3938 3073 3947 3093
rect 3967 3073 3982 3093
rect 3938 3057 3982 3073
rect 4032 3089 4081 3099
rect 4032 3069 4050 3089
rect 4070 3069 4081 3089
rect 4032 3057 4081 3069
rect 18759 3219 18808 3231
rect 18759 3199 18770 3219
rect 18790 3199 18808 3219
rect 18759 3189 18808 3199
rect 18858 3215 18902 3231
rect 18858 3195 18873 3215
rect 18893 3195 18902 3215
rect 18858 3189 18902 3195
rect 18972 3215 19016 3231
rect 18972 3195 18981 3215
rect 19001 3195 19016 3215
rect 18972 3189 19016 3195
rect 19066 3219 19115 3231
rect 19066 3199 19084 3219
rect 19104 3199 19115 3219
rect 19066 3189 19115 3199
rect 19180 3215 19224 3231
rect 19180 3195 19189 3215
rect 19209 3195 19224 3215
rect 19180 3189 19224 3195
rect 19274 3219 19323 3231
rect 19274 3199 19292 3219
rect 19312 3199 19323 3219
rect 19274 3189 19323 3199
rect 19393 3215 19437 3231
rect 19393 3195 19402 3215
rect 19422 3195 19437 3215
rect 19393 3189 19437 3195
rect 19487 3219 19536 3231
rect 19487 3199 19505 3219
rect 19525 3199 19536 3219
rect 19487 3189 19536 3199
rect 19807 3215 19856 3227
rect 19807 3195 19818 3215
rect 19838 3195 19856 3215
rect 11517 3088 11566 3098
rect 11517 3068 11528 3088
rect 11548 3068 11566 3088
rect 11517 3056 11566 3068
rect 11616 3092 11660 3098
rect 11616 3072 11631 3092
rect 11651 3072 11660 3092
rect 11616 3056 11660 3072
rect 11730 3088 11779 3098
rect 11730 3068 11741 3088
rect 11761 3068 11779 3088
rect 11730 3056 11779 3068
rect 11829 3092 11873 3098
rect 11829 3072 11844 3092
rect 11864 3072 11873 3092
rect 11829 3056 11873 3072
rect 11938 3088 11987 3098
rect 11938 3068 11949 3088
rect 11969 3068 11987 3088
rect 11938 3056 11987 3068
rect 12037 3092 12081 3098
rect 12037 3072 12052 3092
rect 12072 3072 12081 3092
rect 12037 3056 12081 3072
rect 12151 3092 12195 3098
rect 12151 3072 12160 3092
rect 12180 3072 12195 3092
rect 12151 3056 12195 3072
rect 12245 3088 12294 3098
rect 19807 3185 19856 3195
rect 19906 3211 19950 3227
rect 19906 3191 19921 3211
rect 19941 3191 19950 3211
rect 19906 3185 19950 3191
rect 20020 3211 20064 3227
rect 20020 3191 20029 3211
rect 20049 3191 20064 3211
rect 20020 3185 20064 3191
rect 20114 3215 20163 3227
rect 20114 3195 20132 3215
rect 20152 3195 20163 3215
rect 20114 3185 20163 3195
rect 20228 3211 20272 3227
rect 20228 3191 20237 3211
rect 20257 3191 20272 3211
rect 20228 3185 20272 3191
rect 20322 3215 20371 3227
rect 20322 3195 20340 3215
rect 20360 3195 20371 3215
rect 20322 3185 20371 3195
rect 20441 3211 20485 3227
rect 20441 3191 20450 3211
rect 20470 3191 20485 3211
rect 20441 3185 20485 3191
rect 20535 3215 20584 3227
rect 20535 3195 20553 3215
rect 20573 3195 20584 3215
rect 20535 3185 20584 3195
rect 12245 3068 12263 3088
rect 12283 3068 12294 3088
rect 12245 3056 12294 3068
rect 14012 3083 14061 3093
rect 14012 3063 14023 3083
rect 14043 3063 14061 3083
rect 14012 3051 14061 3063
rect 14111 3087 14155 3093
rect 14111 3067 14126 3087
rect 14146 3067 14155 3087
rect 14111 3051 14155 3067
rect 14225 3083 14274 3093
rect 14225 3063 14236 3083
rect 14256 3063 14274 3083
rect 14225 3051 14274 3063
rect 14324 3087 14368 3093
rect 14324 3067 14339 3087
rect 14359 3067 14368 3087
rect 14324 3051 14368 3067
rect 14433 3083 14482 3093
rect 14433 3063 14444 3083
rect 14464 3063 14482 3083
rect 14433 3051 14482 3063
rect 14532 3087 14576 3093
rect 14532 3067 14547 3087
rect 14567 3067 14576 3087
rect 14532 3051 14576 3067
rect 14646 3087 14690 3093
rect 14646 3067 14655 3087
rect 14675 3067 14690 3087
rect 14646 3051 14690 3067
rect 14740 3083 14789 3093
rect 14740 3063 14758 3083
rect 14778 3063 14789 3083
rect 14740 3051 14789 3063
rect 6604 2458 6653 2470
rect 6604 2438 6615 2458
rect 6635 2438 6653 2458
rect 6604 2428 6653 2438
rect 6703 2454 6747 2470
rect 6703 2434 6718 2454
rect 6738 2434 6747 2454
rect 6703 2428 6747 2434
rect 6817 2454 6861 2470
rect 6817 2434 6826 2454
rect 6846 2434 6861 2454
rect 6817 2428 6861 2434
rect 6911 2458 6960 2470
rect 6911 2438 6929 2458
rect 6949 2438 6960 2458
rect 6911 2428 6960 2438
rect 7025 2454 7069 2470
rect 7025 2434 7034 2454
rect 7054 2434 7069 2454
rect 7025 2428 7069 2434
rect 7119 2458 7168 2470
rect 7119 2438 7137 2458
rect 7157 2438 7168 2458
rect 7119 2428 7168 2438
rect 7238 2454 7282 2470
rect 7238 2434 7247 2454
rect 7267 2434 7282 2454
rect 7238 2428 7282 2434
rect 7332 2458 7381 2470
rect 7332 2438 7350 2458
rect 7370 2438 7381 2458
rect 7332 2428 7381 2438
rect 9099 2453 9148 2465
rect 9099 2433 9110 2453
rect 9130 2433 9148 2453
rect 809 2326 858 2336
rect 809 2306 820 2326
rect 840 2306 858 2326
rect 809 2294 858 2306
rect 908 2330 952 2336
rect 908 2310 923 2330
rect 943 2310 952 2330
rect 908 2294 952 2310
rect 1022 2326 1071 2336
rect 1022 2306 1033 2326
rect 1053 2306 1071 2326
rect 1022 2294 1071 2306
rect 1121 2330 1165 2336
rect 1121 2310 1136 2330
rect 1156 2310 1165 2330
rect 1121 2294 1165 2310
rect 1230 2326 1279 2336
rect 1230 2306 1241 2326
rect 1261 2306 1279 2326
rect 1230 2294 1279 2306
rect 1329 2330 1373 2336
rect 1329 2310 1344 2330
rect 1364 2310 1373 2330
rect 1329 2294 1373 2310
rect 1443 2330 1487 2336
rect 1443 2310 1452 2330
rect 1472 2310 1487 2330
rect 1443 2294 1487 2310
rect 1537 2326 1586 2336
rect 9099 2423 9148 2433
rect 9198 2449 9242 2465
rect 9198 2429 9213 2449
rect 9233 2429 9242 2449
rect 9198 2423 9242 2429
rect 9312 2449 9356 2465
rect 9312 2429 9321 2449
rect 9341 2429 9356 2449
rect 9312 2423 9356 2429
rect 9406 2453 9455 2465
rect 9406 2433 9424 2453
rect 9444 2433 9455 2453
rect 9406 2423 9455 2433
rect 9520 2449 9564 2465
rect 9520 2429 9529 2449
rect 9549 2429 9564 2449
rect 9520 2423 9564 2429
rect 9614 2453 9663 2465
rect 9614 2433 9632 2453
rect 9652 2433 9663 2453
rect 9614 2423 9663 2433
rect 9733 2449 9777 2465
rect 9733 2429 9742 2449
rect 9762 2429 9777 2449
rect 9733 2423 9777 2429
rect 9827 2453 9876 2465
rect 9827 2433 9845 2453
rect 9865 2433 9876 2453
rect 9827 2423 9876 2433
rect 1537 2306 1555 2326
rect 1575 2306 1586 2326
rect 1537 2294 1586 2306
rect 1857 2322 1906 2332
rect 1857 2302 1868 2322
rect 1888 2302 1906 2322
rect 1857 2290 1906 2302
rect 1956 2326 2000 2332
rect 1956 2306 1971 2326
rect 1991 2306 2000 2326
rect 1956 2290 2000 2306
rect 2070 2322 2119 2332
rect 2070 2302 2081 2322
rect 2101 2302 2119 2322
rect 2070 2290 2119 2302
rect 2169 2326 2213 2332
rect 2169 2306 2184 2326
rect 2204 2306 2213 2326
rect 2169 2290 2213 2306
rect 2278 2322 2327 2332
rect 2278 2302 2289 2322
rect 2309 2302 2327 2322
rect 2278 2290 2327 2302
rect 2377 2326 2421 2332
rect 2377 2306 2392 2326
rect 2412 2306 2421 2326
rect 2377 2290 2421 2306
rect 2491 2326 2535 2332
rect 2491 2306 2500 2326
rect 2520 2306 2535 2326
rect 2491 2290 2535 2306
rect 2585 2322 2634 2332
rect 2585 2302 2603 2322
rect 2623 2302 2634 2322
rect 2585 2290 2634 2302
rect 17312 2452 17361 2464
rect 17312 2432 17323 2452
rect 17343 2432 17361 2452
rect 17312 2422 17361 2432
rect 17411 2448 17455 2464
rect 17411 2428 17426 2448
rect 17446 2428 17455 2448
rect 17411 2422 17455 2428
rect 17525 2448 17569 2464
rect 17525 2428 17534 2448
rect 17554 2428 17569 2448
rect 17525 2422 17569 2428
rect 17619 2452 17668 2464
rect 17619 2432 17637 2452
rect 17657 2432 17668 2452
rect 17619 2422 17668 2432
rect 17733 2448 17777 2464
rect 17733 2428 17742 2448
rect 17762 2428 17777 2448
rect 17733 2422 17777 2428
rect 17827 2452 17876 2464
rect 17827 2432 17845 2452
rect 17865 2432 17876 2452
rect 17827 2422 17876 2432
rect 17946 2448 17990 2464
rect 17946 2428 17955 2448
rect 17975 2428 17990 2448
rect 17946 2422 17990 2428
rect 18040 2452 18089 2464
rect 18040 2432 18058 2452
rect 18078 2432 18089 2452
rect 18040 2422 18089 2432
rect 19807 2447 19856 2459
rect 19807 2427 19818 2447
rect 19838 2427 19856 2447
rect 11517 2320 11566 2330
rect 11517 2300 11528 2320
rect 11548 2300 11566 2320
rect 11517 2288 11566 2300
rect 11616 2324 11660 2330
rect 11616 2304 11631 2324
rect 11651 2304 11660 2324
rect 11616 2288 11660 2304
rect 11730 2320 11779 2330
rect 11730 2300 11741 2320
rect 11761 2300 11779 2320
rect 11730 2288 11779 2300
rect 11829 2324 11873 2330
rect 11829 2304 11844 2324
rect 11864 2304 11873 2324
rect 11829 2288 11873 2304
rect 11938 2320 11987 2330
rect 11938 2300 11949 2320
rect 11969 2300 11987 2320
rect 11938 2288 11987 2300
rect 12037 2324 12081 2330
rect 12037 2304 12052 2324
rect 12072 2304 12081 2324
rect 12037 2288 12081 2304
rect 12151 2324 12195 2330
rect 12151 2304 12160 2324
rect 12180 2304 12195 2324
rect 12151 2288 12195 2304
rect 12245 2320 12294 2330
rect 19807 2417 19856 2427
rect 19906 2443 19950 2459
rect 19906 2423 19921 2443
rect 19941 2423 19950 2443
rect 19906 2417 19950 2423
rect 20020 2443 20064 2459
rect 20020 2423 20029 2443
rect 20049 2423 20064 2443
rect 20020 2417 20064 2423
rect 20114 2447 20163 2459
rect 20114 2427 20132 2447
rect 20152 2427 20163 2447
rect 20114 2417 20163 2427
rect 20228 2443 20272 2459
rect 20228 2423 20237 2443
rect 20257 2423 20272 2443
rect 20228 2417 20272 2423
rect 20322 2447 20371 2459
rect 20322 2427 20340 2447
rect 20360 2427 20371 2447
rect 20322 2417 20371 2427
rect 20441 2443 20485 2459
rect 20441 2423 20450 2443
rect 20470 2423 20485 2443
rect 20441 2417 20485 2423
rect 20535 2447 20584 2459
rect 20535 2427 20553 2447
rect 20573 2427 20584 2447
rect 20535 2417 20584 2427
rect 12245 2300 12263 2320
rect 12283 2300 12294 2320
rect 12245 2288 12294 2300
rect 12565 2316 12614 2326
rect 12565 2296 12576 2316
rect 12596 2296 12614 2316
rect 12565 2284 12614 2296
rect 12664 2320 12708 2326
rect 12664 2300 12679 2320
rect 12699 2300 12708 2320
rect 12664 2284 12708 2300
rect 12778 2316 12827 2326
rect 12778 2296 12789 2316
rect 12809 2296 12827 2316
rect 12778 2284 12827 2296
rect 12877 2320 12921 2326
rect 12877 2300 12892 2320
rect 12912 2300 12921 2320
rect 12877 2284 12921 2300
rect 12986 2316 13035 2326
rect 12986 2296 12997 2316
rect 13017 2296 13035 2316
rect 12986 2284 13035 2296
rect 13085 2320 13129 2326
rect 13085 2300 13100 2320
rect 13120 2300 13129 2320
rect 13085 2284 13129 2300
rect 13199 2320 13243 2326
rect 13199 2300 13208 2320
rect 13228 2300 13243 2320
rect 13199 2284 13243 2300
rect 13293 2316 13342 2326
rect 13293 2296 13311 2316
rect 13331 2296 13342 2316
rect 13293 2284 13342 2296
rect 8051 1778 8100 1790
rect 8051 1758 8062 1778
rect 8082 1758 8100 1778
rect 8051 1748 8100 1758
rect 8150 1774 8194 1790
rect 8150 1754 8165 1774
rect 8185 1754 8194 1774
rect 8150 1748 8194 1754
rect 8264 1774 8308 1790
rect 8264 1754 8273 1774
rect 8293 1754 8308 1774
rect 8264 1748 8308 1754
rect 8358 1778 8407 1790
rect 8358 1758 8376 1778
rect 8396 1758 8407 1778
rect 8358 1748 8407 1758
rect 8472 1774 8516 1790
rect 8472 1754 8481 1774
rect 8501 1754 8516 1774
rect 8472 1748 8516 1754
rect 8566 1778 8615 1790
rect 8566 1758 8584 1778
rect 8604 1758 8615 1778
rect 8566 1748 8615 1758
rect 8685 1774 8729 1790
rect 8685 1754 8694 1774
rect 8714 1754 8729 1774
rect 8685 1748 8729 1754
rect 8779 1778 8828 1790
rect 8779 1758 8797 1778
rect 8817 1758 8828 1778
rect 8779 1748 8828 1758
rect 9099 1774 9148 1786
rect 9099 1754 9110 1774
rect 9130 1754 9148 1774
rect 9099 1744 9148 1754
rect 9198 1770 9242 1786
rect 9198 1750 9213 1770
rect 9233 1750 9242 1770
rect 9198 1744 9242 1750
rect 9312 1770 9356 1786
rect 9312 1750 9321 1770
rect 9341 1750 9356 1770
rect 9312 1744 9356 1750
rect 9406 1774 9455 1786
rect 9406 1754 9424 1774
rect 9444 1754 9455 1774
rect 9406 1744 9455 1754
rect 9520 1770 9564 1786
rect 9520 1750 9529 1770
rect 9549 1750 9564 1770
rect 9520 1744 9564 1750
rect 9614 1774 9663 1786
rect 9614 1754 9632 1774
rect 9652 1754 9663 1774
rect 9614 1744 9663 1754
rect 9733 1770 9777 1786
rect 9733 1750 9742 1770
rect 9762 1750 9777 1770
rect 9733 1744 9777 1750
rect 9827 1774 9876 1786
rect 9827 1754 9845 1774
rect 9865 1754 9876 1774
rect 9827 1744 9876 1754
rect 809 1647 858 1657
rect 809 1627 820 1647
rect 840 1627 858 1647
rect 809 1615 858 1627
rect 908 1651 952 1657
rect 908 1631 923 1651
rect 943 1631 952 1651
rect 908 1615 952 1631
rect 1022 1647 1071 1657
rect 1022 1627 1033 1647
rect 1053 1627 1071 1647
rect 1022 1615 1071 1627
rect 1121 1651 1165 1657
rect 1121 1631 1136 1651
rect 1156 1631 1165 1651
rect 1121 1615 1165 1631
rect 1230 1647 1279 1657
rect 1230 1627 1241 1647
rect 1261 1627 1279 1647
rect 1230 1615 1279 1627
rect 1329 1651 1373 1657
rect 1329 1631 1344 1651
rect 1364 1631 1373 1651
rect 1329 1615 1373 1631
rect 1443 1651 1487 1657
rect 1443 1631 1452 1651
rect 1472 1631 1487 1651
rect 1443 1615 1487 1631
rect 1537 1647 1586 1657
rect 1537 1627 1555 1647
rect 1575 1627 1586 1647
rect 1537 1615 1586 1627
rect 18759 1772 18808 1784
rect 18759 1752 18770 1772
rect 18790 1752 18808 1772
rect 18759 1742 18808 1752
rect 18858 1768 18902 1784
rect 18858 1748 18873 1768
rect 18893 1748 18902 1768
rect 18858 1742 18902 1748
rect 18972 1768 19016 1784
rect 18972 1748 18981 1768
rect 19001 1748 19016 1768
rect 18972 1742 19016 1748
rect 19066 1772 19115 1784
rect 19066 1752 19084 1772
rect 19104 1752 19115 1772
rect 19066 1742 19115 1752
rect 19180 1768 19224 1784
rect 19180 1748 19189 1768
rect 19209 1748 19224 1768
rect 19180 1742 19224 1748
rect 19274 1772 19323 1784
rect 19274 1752 19292 1772
rect 19312 1752 19323 1772
rect 19274 1742 19323 1752
rect 19393 1768 19437 1784
rect 19393 1748 19402 1768
rect 19422 1748 19437 1768
rect 19393 1742 19437 1748
rect 19487 1772 19536 1784
rect 19487 1752 19505 1772
rect 19525 1752 19536 1772
rect 19487 1742 19536 1752
rect 19807 1768 19856 1780
rect 19807 1748 19818 1768
rect 19838 1748 19856 1768
rect 19807 1738 19856 1748
rect 19906 1764 19950 1780
rect 19906 1744 19921 1764
rect 19941 1744 19950 1764
rect 19906 1738 19950 1744
rect 20020 1764 20064 1780
rect 20020 1744 20029 1764
rect 20049 1744 20064 1764
rect 20020 1738 20064 1744
rect 20114 1768 20163 1780
rect 20114 1748 20132 1768
rect 20152 1748 20163 1768
rect 20114 1738 20163 1748
rect 20228 1764 20272 1780
rect 20228 1744 20237 1764
rect 20257 1744 20272 1764
rect 20228 1738 20272 1744
rect 20322 1768 20371 1780
rect 20322 1748 20340 1768
rect 20360 1748 20371 1768
rect 20322 1738 20371 1748
rect 20441 1764 20485 1780
rect 20441 1744 20450 1764
rect 20470 1744 20485 1764
rect 20441 1738 20485 1744
rect 20535 1768 20584 1780
rect 20535 1748 20553 1768
rect 20573 1748 20584 1768
rect 20535 1738 20584 1748
rect 11517 1641 11566 1651
rect 11517 1621 11528 1641
rect 11548 1621 11566 1641
rect 11517 1609 11566 1621
rect 11616 1645 11660 1651
rect 11616 1625 11631 1645
rect 11651 1625 11660 1645
rect 11616 1609 11660 1625
rect 11730 1641 11779 1651
rect 11730 1621 11741 1641
rect 11761 1621 11779 1641
rect 11730 1609 11779 1621
rect 11829 1645 11873 1651
rect 11829 1625 11844 1645
rect 11864 1625 11873 1645
rect 11829 1609 11873 1625
rect 11938 1641 11987 1651
rect 11938 1621 11949 1641
rect 11969 1621 11987 1641
rect 11938 1609 11987 1621
rect 12037 1645 12081 1651
rect 12037 1625 12052 1645
rect 12072 1625 12081 1645
rect 12037 1609 12081 1625
rect 12151 1645 12195 1651
rect 12151 1625 12160 1645
rect 12180 1625 12195 1645
rect 12151 1609 12195 1625
rect 12245 1641 12294 1651
rect 12245 1621 12263 1641
rect 12283 1621 12294 1641
rect 12245 1609 12294 1621
rect 10520 -512 10569 -502
rect 10520 -532 10531 -512
rect 10551 -532 10569 -512
rect 10520 -544 10569 -532
rect 10619 -508 10663 -502
rect 10619 -528 10634 -508
rect 10654 -528 10663 -508
rect 10619 -544 10663 -528
rect 10733 -512 10782 -502
rect 10733 -532 10744 -512
rect 10764 -532 10782 -512
rect 10733 -544 10782 -532
rect 10832 -508 10876 -502
rect 10832 -528 10847 -508
rect 10867 -528 10876 -508
rect 10832 -544 10876 -528
rect 10941 -512 10990 -502
rect 10941 -532 10952 -512
rect 10972 -532 10990 -512
rect 10941 -544 10990 -532
rect 11040 -508 11084 -502
rect 11040 -528 11055 -508
rect 11075 -528 11084 -508
rect 11040 -544 11084 -528
rect 11154 -508 11198 -502
rect 11154 -528 11163 -508
rect 11183 -528 11198 -508
rect 11154 -544 11198 -528
rect 11248 -512 11297 -502
rect 11248 -532 11266 -512
rect 11286 -532 11297 -512
rect 11248 -544 11297 -532
<< pdiff >>
rect 815 12897 859 12935
rect 815 12877 827 12897
rect 847 12877 859 12897
rect 815 12835 859 12877
rect 909 12897 951 12935
rect 909 12877 923 12897
rect 943 12877 951 12897
rect 909 12835 951 12877
rect 1028 12897 1072 12935
rect 1028 12877 1040 12897
rect 1060 12877 1072 12897
rect 1028 12835 1072 12877
rect 1122 12897 1164 12935
rect 1122 12877 1136 12897
rect 1156 12877 1164 12897
rect 1122 12835 1164 12877
rect 1236 12897 1280 12935
rect 1236 12877 1248 12897
rect 1268 12877 1280 12897
rect 1236 12835 1280 12877
rect 1330 12897 1372 12935
rect 1330 12877 1344 12897
rect 1364 12877 1372 12897
rect 1330 12835 1372 12877
rect 1446 12897 1488 12935
rect 1446 12877 1454 12897
rect 1474 12877 1488 12897
rect 1446 12835 1488 12877
rect 1538 12904 1583 12935
rect 1538 12897 1582 12904
rect 1538 12877 1550 12897
rect 1570 12877 1582 12897
rect 1538 12835 1582 12877
rect 1863 12893 1907 12931
rect 1863 12873 1875 12893
rect 1895 12873 1907 12893
rect 1863 12831 1907 12873
rect 1957 12893 1999 12931
rect 1957 12873 1971 12893
rect 1991 12873 1999 12893
rect 1957 12831 1999 12873
rect 2076 12893 2120 12931
rect 2076 12873 2088 12893
rect 2108 12873 2120 12893
rect 2076 12831 2120 12873
rect 2170 12893 2212 12931
rect 2170 12873 2184 12893
rect 2204 12873 2212 12893
rect 2170 12831 2212 12873
rect 2284 12893 2328 12931
rect 2284 12873 2296 12893
rect 2316 12873 2328 12893
rect 2284 12831 2328 12873
rect 2378 12893 2420 12931
rect 2378 12873 2392 12893
rect 2412 12873 2420 12893
rect 2378 12831 2420 12873
rect 2494 12893 2536 12931
rect 2494 12873 2502 12893
rect 2522 12873 2536 12893
rect 2494 12831 2536 12873
rect 2586 12900 2631 12931
rect 2586 12893 2630 12900
rect 2586 12873 2598 12893
rect 2618 12873 2630 12893
rect 2586 12831 2630 12873
rect 11523 12891 11567 12929
rect 11523 12871 11535 12891
rect 11555 12871 11567 12891
rect 11523 12829 11567 12871
rect 11617 12891 11659 12929
rect 11617 12871 11631 12891
rect 11651 12871 11659 12891
rect 11617 12829 11659 12871
rect 11736 12891 11780 12929
rect 11736 12871 11748 12891
rect 11768 12871 11780 12891
rect 11736 12829 11780 12871
rect 11830 12891 11872 12929
rect 11830 12871 11844 12891
rect 11864 12871 11872 12891
rect 11830 12829 11872 12871
rect 11944 12891 11988 12929
rect 11944 12871 11956 12891
rect 11976 12871 11988 12891
rect 11944 12829 11988 12871
rect 12038 12891 12080 12929
rect 12038 12871 12052 12891
rect 12072 12871 12080 12891
rect 12038 12829 12080 12871
rect 12154 12891 12196 12929
rect 12154 12871 12162 12891
rect 12182 12871 12196 12891
rect 12154 12829 12196 12871
rect 12246 12898 12291 12929
rect 12246 12891 12290 12898
rect 12246 12871 12258 12891
rect 12278 12871 12290 12891
rect 12246 12829 12290 12871
rect 12571 12887 12615 12925
rect 12571 12867 12583 12887
rect 12603 12867 12615 12887
rect 9105 12726 9149 12768
rect 9105 12706 9117 12726
rect 9137 12706 9149 12726
rect 9105 12699 9149 12706
rect 9104 12668 9149 12699
rect 9199 12726 9241 12768
rect 9199 12706 9213 12726
rect 9233 12706 9241 12726
rect 9199 12668 9241 12706
rect 9315 12726 9357 12768
rect 9315 12706 9323 12726
rect 9343 12706 9357 12726
rect 9315 12668 9357 12706
rect 9407 12726 9451 12768
rect 9407 12706 9419 12726
rect 9439 12706 9451 12726
rect 9407 12668 9451 12706
rect 9523 12726 9565 12768
rect 9523 12706 9531 12726
rect 9551 12706 9565 12726
rect 9523 12668 9565 12706
rect 9615 12726 9659 12768
rect 9615 12706 9627 12726
rect 9647 12706 9659 12726
rect 9615 12668 9659 12706
rect 9736 12726 9778 12768
rect 9736 12706 9744 12726
rect 9764 12706 9778 12726
rect 9736 12668 9778 12706
rect 9828 12726 9872 12768
rect 12571 12825 12615 12867
rect 12665 12887 12707 12925
rect 12665 12867 12679 12887
rect 12699 12867 12707 12887
rect 12665 12825 12707 12867
rect 12784 12887 12828 12925
rect 12784 12867 12796 12887
rect 12816 12867 12828 12887
rect 12784 12825 12828 12867
rect 12878 12887 12920 12925
rect 12878 12867 12892 12887
rect 12912 12867 12920 12887
rect 12878 12825 12920 12867
rect 12992 12887 13036 12925
rect 12992 12867 13004 12887
rect 13024 12867 13036 12887
rect 12992 12825 13036 12867
rect 13086 12887 13128 12925
rect 13086 12867 13100 12887
rect 13120 12867 13128 12887
rect 13086 12825 13128 12867
rect 13202 12887 13244 12925
rect 13202 12867 13210 12887
rect 13230 12867 13244 12887
rect 13202 12825 13244 12867
rect 13294 12894 13339 12925
rect 13294 12887 13338 12894
rect 13294 12867 13306 12887
rect 13326 12867 13338 12887
rect 13294 12825 13338 12867
rect 9828 12706 9840 12726
rect 9860 12706 9872 12726
rect 9828 12668 9872 12706
rect 19813 12720 19857 12762
rect 19813 12700 19825 12720
rect 19845 12700 19857 12720
rect 19813 12693 19857 12700
rect 19812 12662 19857 12693
rect 19907 12720 19949 12762
rect 19907 12700 19921 12720
rect 19941 12700 19949 12720
rect 19907 12662 19949 12700
rect 20023 12720 20065 12762
rect 20023 12700 20031 12720
rect 20051 12700 20065 12720
rect 20023 12662 20065 12700
rect 20115 12720 20159 12762
rect 20115 12700 20127 12720
rect 20147 12700 20159 12720
rect 20115 12662 20159 12700
rect 20231 12720 20273 12762
rect 20231 12700 20239 12720
rect 20259 12700 20273 12720
rect 20231 12662 20273 12700
rect 20323 12720 20367 12762
rect 20323 12700 20335 12720
rect 20355 12700 20367 12720
rect 20323 12662 20367 12700
rect 20444 12720 20486 12762
rect 20444 12700 20452 12720
rect 20472 12700 20486 12720
rect 20444 12662 20486 12700
rect 20536 12720 20580 12762
rect 20536 12700 20548 12720
rect 20568 12700 20580 12720
rect 20536 12662 20580 12700
rect 815 12218 859 12256
rect 815 12198 827 12218
rect 847 12198 859 12218
rect 815 12156 859 12198
rect 909 12218 951 12256
rect 909 12198 923 12218
rect 943 12198 951 12218
rect 909 12156 951 12198
rect 1028 12218 1072 12256
rect 1028 12198 1040 12218
rect 1060 12198 1072 12218
rect 1028 12156 1072 12198
rect 1122 12218 1164 12256
rect 1122 12198 1136 12218
rect 1156 12198 1164 12218
rect 1122 12156 1164 12198
rect 1236 12218 1280 12256
rect 1236 12198 1248 12218
rect 1268 12198 1280 12218
rect 1236 12156 1280 12198
rect 1330 12218 1372 12256
rect 1330 12198 1344 12218
rect 1364 12198 1372 12218
rect 1330 12156 1372 12198
rect 1446 12218 1488 12256
rect 1446 12198 1454 12218
rect 1474 12198 1488 12218
rect 1446 12156 1488 12198
rect 1538 12225 1583 12256
rect 1538 12218 1582 12225
rect 1538 12198 1550 12218
rect 1570 12198 1582 12218
rect 1538 12156 1582 12198
rect 3310 12213 3354 12251
rect 3310 12193 3322 12213
rect 3342 12193 3354 12213
rect 3310 12151 3354 12193
rect 3404 12213 3446 12251
rect 3404 12193 3418 12213
rect 3438 12193 3446 12213
rect 3404 12151 3446 12193
rect 3523 12213 3567 12251
rect 3523 12193 3535 12213
rect 3555 12193 3567 12213
rect 3523 12151 3567 12193
rect 3617 12213 3659 12251
rect 3617 12193 3631 12213
rect 3651 12193 3659 12213
rect 3617 12151 3659 12193
rect 3731 12213 3775 12251
rect 3731 12193 3743 12213
rect 3763 12193 3775 12213
rect 3731 12151 3775 12193
rect 3825 12213 3867 12251
rect 3825 12193 3839 12213
rect 3859 12193 3867 12213
rect 3825 12151 3867 12193
rect 3941 12213 3983 12251
rect 3941 12193 3949 12213
rect 3969 12193 3983 12213
rect 3941 12151 3983 12193
rect 4033 12220 4078 12251
rect 4033 12213 4077 12220
rect 4033 12193 4045 12213
rect 4065 12193 4077 12213
rect 4033 12151 4077 12193
rect 11523 12212 11567 12250
rect 11523 12192 11535 12212
rect 11555 12192 11567 12212
rect 8057 12051 8101 12093
rect 8057 12031 8069 12051
rect 8089 12031 8101 12051
rect 8057 12024 8101 12031
rect 8056 11993 8101 12024
rect 8151 12051 8193 12093
rect 8151 12031 8165 12051
rect 8185 12031 8193 12051
rect 8151 11993 8193 12031
rect 8267 12051 8309 12093
rect 8267 12031 8275 12051
rect 8295 12031 8309 12051
rect 8267 11993 8309 12031
rect 8359 12051 8403 12093
rect 8359 12031 8371 12051
rect 8391 12031 8403 12051
rect 8359 11993 8403 12031
rect 8475 12051 8517 12093
rect 8475 12031 8483 12051
rect 8503 12031 8517 12051
rect 8475 11993 8517 12031
rect 8567 12051 8611 12093
rect 8567 12031 8579 12051
rect 8599 12031 8611 12051
rect 8567 11993 8611 12031
rect 8688 12051 8730 12093
rect 8688 12031 8696 12051
rect 8716 12031 8730 12051
rect 8688 11993 8730 12031
rect 8780 12051 8824 12093
rect 11523 12150 11567 12192
rect 11617 12212 11659 12250
rect 11617 12192 11631 12212
rect 11651 12192 11659 12212
rect 11617 12150 11659 12192
rect 11736 12212 11780 12250
rect 11736 12192 11748 12212
rect 11768 12192 11780 12212
rect 11736 12150 11780 12192
rect 11830 12212 11872 12250
rect 11830 12192 11844 12212
rect 11864 12192 11872 12212
rect 11830 12150 11872 12192
rect 11944 12212 11988 12250
rect 11944 12192 11956 12212
rect 11976 12192 11988 12212
rect 11944 12150 11988 12192
rect 12038 12212 12080 12250
rect 12038 12192 12052 12212
rect 12072 12192 12080 12212
rect 12038 12150 12080 12192
rect 12154 12212 12196 12250
rect 12154 12192 12162 12212
rect 12182 12192 12196 12212
rect 12154 12150 12196 12192
rect 12246 12219 12291 12250
rect 12246 12212 12290 12219
rect 12246 12192 12258 12212
rect 12278 12192 12290 12212
rect 12246 12150 12290 12192
rect 14018 12207 14062 12245
rect 14018 12187 14030 12207
rect 14050 12187 14062 12207
rect 8780 12031 8792 12051
rect 8812 12031 8824 12051
rect 8780 11993 8824 12031
rect 9105 12047 9149 12089
rect 9105 12027 9117 12047
rect 9137 12027 9149 12047
rect 9105 12020 9149 12027
rect 9104 11989 9149 12020
rect 9199 12047 9241 12089
rect 9199 12027 9213 12047
rect 9233 12027 9241 12047
rect 9199 11989 9241 12027
rect 9315 12047 9357 12089
rect 9315 12027 9323 12047
rect 9343 12027 9357 12047
rect 9315 11989 9357 12027
rect 9407 12047 9451 12089
rect 9407 12027 9419 12047
rect 9439 12027 9451 12047
rect 9407 11989 9451 12027
rect 9523 12047 9565 12089
rect 9523 12027 9531 12047
rect 9551 12027 9565 12047
rect 9523 11989 9565 12027
rect 9615 12047 9659 12089
rect 9615 12027 9627 12047
rect 9647 12027 9659 12047
rect 9615 11989 9659 12027
rect 9736 12047 9778 12089
rect 9736 12027 9744 12047
rect 9764 12027 9778 12047
rect 9736 11989 9778 12027
rect 9828 12047 9872 12089
rect 9828 12027 9840 12047
rect 9860 12027 9872 12047
rect 14018 12145 14062 12187
rect 14112 12207 14154 12245
rect 14112 12187 14126 12207
rect 14146 12187 14154 12207
rect 14112 12145 14154 12187
rect 14231 12207 14275 12245
rect 14231 12187 14243 12207
rect 14263 12187 14275 12207
rect 14231 12145 14275 12187
rect 14325 12207 14367 12245
rect 14325 12187 14339 12207
rect 14359 12187 14367 12207
rect 14325 12145 14367 12187
rect 14439 12207 14483 12245
rect 14439 12187 14451 12207
rect 14471 12187 14483 12207
rect 14439 12145 14483 12187
rect 14533 12207 14575 12245
rect 14533 12187 14547 12207
rect 14567 12187 14575 12207
rect 14533 12145 14575 12187
rect 14649 12207 14691 12245
rect 14649 12187 14657 12207
rect 14677 12187 14691 12207
rect 14649 12145 14691 12187
rect 14741 12214 14786 12245
rect 14741 12207 14785 12214
rect 14741 12187 14753 12207
rect 14773 12187 14785 12207
rect 14741 12145 14785 12187
rect 9828 11989 9872 12027
rect 18765 12045 18809 12087
rect 18765 12025 18777 12045
rect 18797 12025 18809 12045
rect 18765 12018 18809 12025
rect 18764 11987 18809 12018
rect 18859 12045 18901 12087
rect 18859 12025 18873 12045
rect 18893 12025 18901 12045
rect 18859 11987 18901 12025
rect 18975 12045 19017 12087
rect 18975 12025 18983 12045
rect 19003 12025 19017 12045
rect 18975 11987 19017 12025
rect 19067 12045 19111 12087
rect 19067 12025 19079 12045
rect 19099 12025 19111 12045
rect 19067 11987 19111 12025
rect 19183 12045 19225 12087
rect 19183 12025 19191 12045
rect 19211 12025 19225 12045
rect 19183 11987 19225 12025
rect 19275 12045 19319 12087
rect 19275 12025 19287 12045
rect 19307 12025 19319 12045
rect 19275 11987 19319 12025
rect 19396 12045 19438 12087
rect 19396 12025 19404 12045
rect 19424 12025 19438 12045
rect 19396 11987 19438 12025
rect 19488 12045 19532 12087
rect 19488 12025 19500 12045
rect 19520 12025 19532 12045
rect 19488 11987 19532 12025
rect 19813 12041 19857 12083
rect 19813 12021 19825 12041
rect 19845 12021 19857 12041
rect 19813 12014 19857 12021
rect 19812 11983 19857 12014
rect 19907 12041 19949 12083
rect 19907 12021 19921 12041
rect 19941 12021 19949 12041
rect 19907 11983 19949 12021
rect 20023 12041 20065 12083
rect 20023 12021 20031 12041
rect 20051 12021 20065 12041
rect 20023 11983 20065 12021
rect 20115 12041 20159 12083
rect 20115 12021 20127 12041
rect 20147 12021 20159 12041
rect 20115 11983 20159 12021
rect 20231 12041 20273 12083
rect 20231 12021 20239 12041
rect 20259 12021 20273 12041
rect 20231 11983 20273 12021
rect 20323 12041 20367 12083
rect 20323 12021 20335 12041
rect 20355 12021 20367 12041
rect 20323 11983 20367 12021
rect 20444 12041 20486 12083
rect 20444 12021 20452 12041
rect 20472 12021 20486 12041
rect 20444 11983 20486 12021
rect 20536 12041 20580 12083
rect 20536 12021 20548 12041
rect 20568 12021 20580 12041
rect 20536 11983 20580 12021
rect 815 11450 859 11488
rect 815 11430 827 11450
rect 847 11430 859 11450
rect 815 11388 859 11430
rect 909 11450 951 11488
rect 909 11430 923 11450
rect 943 11430 951 11450
rect 909 11388 951 11430
rect 1028 11450 1072 11488
rect 1028 11430 1040 11450
rect 1060 11430 1072 11450
rect 1028 11388 1072 11430
rect 1122 11450 1164 11488
rect 1122 11430 1136 11450
rect 1156 11430 1164 11450
rect 1122 11388 1164 11430
rect 1236 11450 1280 11488
rect 1236 11430 1248 11450
rect 1268 11430 1280 11450
rect 1236 11388 1280 11430
rect 1330 11450 1372 11488
rect 1330 11430 1344 11450
rect 1364 11430 1372 11450
rect 1330 11388 1372 11430
rect 1446 11450 1488 11488
rect 1446 11430 1454 11450
rect 1474 11430 1488 11450
rect 1446 11388 1488 11430
rect 1538 11457 1583 11488
rect 1538 11450 1582 11457
rect 1538 11430 1550 11450
rect 1570 11430 1582 11450
rect 1538 11388 1582 11430
rect 1863 11446 1907 11484
rect 1863 11426 1875 11446
rect 1895 11426 1907 11446
rect 1863 11384 1907 11426
rect 1957 11446 1999 11484
rect 1957 11426 1971 11446
rect 1991 11426 1999 11446
rect 1957 11384 1999 11426
rect 2076 11446 2120 11484
rect 2076 11426 2088 11446
rect 2108 11426 2120 11446
rect 2076 11384 2120 11426
rect 2170 11446 2212 11484
rect 2170 11426 2184 11446
rect 2204 11426 2212 11446
rect 2170 11384 2212 11426
rect 2284 11446 2328 11484
rect 2284 11426 2296 11446
rect 2316 11426 2328 11446
rect 2284 11384 2328 11426
rect 2378 11446 2420 11484
rect 2378 11426 2392 11446
rect 2412 11426 2420 11446
rect 2378 11384 2420 11426
rect 2494 11446 2536 11484
rect 2494 11426 2502 11446
rect 2522 11426 2536 11446
rect 2494 11384 2536 11426
rect 2586 11453 2631 11484
rect 2586 11446 2630 11453
rect 2586 11426 2598 11446
rect 2618 11426 2630 11446
rect 2586 11384 2630 11426
rect 11523 11444 11567 11482
rect 6610 11284 6654 11326
rect 6610 11264 6622 11284
rect 6642 11264 6654 11284
rect 6610 11257 6654 11264
rect 6609 11226 6654 11257
rect 6704 11284 6746 11326
rect 6704 11264 6718 11284
rect 6738 11264 6746 11284
rect 6704 11226 6746 11264
rect 6820 11284 6862 11326
rect 6820 11264 6828 11284
rect 6848 11264 6862 11284
rect 6820 11226 6862 11264
rect 6912 11284 6956 11326
rect 6912 11264 6924 11284
rect 6944 11264 6956 11284
rect 6912 11226 6956 11264
rect 7028 11284 7070 11326
rect 7028 11264 7036 11284
rect 7056 11264 7070 11284
rect 7028 11226 7070 11264
rect 7120 11284 7164 11326
rect 7120 11264 7132 11284
rect 7152 11264 7164 11284
rect 7120 11226 7164 11264
rect 7241 11284 7283 11326
rect 7241 11264 7249 11284
rect 7269 11264 7283 11284
rect 7241 11226 7283 11264
rect 7333 11284 7377 11326
rect 11523 11424 11535 11444
rect 11555 11424 11567 11444
rect 11523 11382 11567 11424
rect 11617 11444 11659 11482
rect 11617 11424 11631 11444
rect 11651 11424 11659 11444
rect 11617 11382 11659 11424
rect 11736 11444 11780 11482
rect 11736 11424 11748 11444
rect 11768 11424 11780 11444
rect 11736 11382 11780 11424
rect 11830 11444 11872 11482
rect 11830 11424 11844 11444
rect 11864 11424 11872 11444
rect 11830 11382 11872 11424
rect 11944 11444 11988 11482
rect 11944 11424 11956 11444
rect 11976 11424 11988 11444
rect 11944 11382 11988 11424
rect 12038 11444 12080 11482
rect 12038 11424 12052 11444
rect 12072 11424 12080 11444
rect 12038 11382 12080 11424
rect 12154 11444 12196 11482
rect 12154 11424 12162 11444
rect 12182 11424 12196 11444
rect 12154 11382 12196 11424
rect 12246 11451 12291 11482
rect 12246 11444 12290 11451
rect 12246 11424 12258 11444
rect 12278 11424 12290 11444
rect 12246 11382 12290 11424
rect 12571 11440 12615 11478
rect 12571 11420 12583 11440
rect 12603 11420 12615 11440
rect 7333 11264 7345 11284
rect 7365 11264 7377 11284
rect 7333 11226 7377 11264
rect 9105 11279 9149 11321
rect 9105 11259 9117 11279
rect 9137 11259 9149 11279
rect 9105 11252 9149 11259
rect 9104 11221 9149 11252
rect 9199 11279 9241 11321
rect 9199 11259 9213 11279
rect 9233 11259 9241 11279
rect 9199 11221 9241 11259
rect 9315 11279 9357 11321
rect 9315 11259 9323 11279
rect 9343 11259 9357 11279
rect 9315 11221 9357 11259
rect 9407 11279 9451 11321
rect 9407 11259 9419 11279
rect 9439 11259 9451 11279
rect 9407 11221 9451 11259
rect 9523 11279 9565 11321
rect 9523 11259 9531 11279
rect 9551 11259 9565 11279
rect 9523 11221 9565 11259
rect 9615 11279 9659 11321
rect 9615 11259 9627 11279
rect 9647 11259 9659 11279
rect 9615 11221 9659 11259
rect 9736 11279 9778 11321
rect 9736 11259 9744 11279
rect 9764 11259 9778 11279
rect 9736 11221 9778 11259
rect 9828 11279 9872 11321
rect 12571 11378 12615 11420
rect 12665 11440 12707 11478
rect 12665 11420 12679 11440
rect 12699 11420 12707 11440
rect 12665 11378 12707 11420
rect 12784 11440 12828 11478
rect 12784 11420 12796 11440
rect 12816 11420 12828 11440
rect 12784 11378 12828 11420
rect 12878 11440 12920 11478
rect 12878 11420 12892 11440
rect 12912 11420 12920 11440
rect 12878 11378 12920 11420
rect 12992 11440 13036 11478
rect 12992 11420 13004 11440
rect 13024 11420 13036 11440
rect 12992 11378 13036 11420
rect 13086 11440 13128 11478
rect 13086 11420 13100 11440
rect 13120 11420 13128 11440
rect 13086 11378 13128 11420
rect 13202 11440 13244 11478
rect 13202 11420 13210 11440
rect 13230 11420 13244 11440
rect 13202 11378 13244 11420
rect 13294 11447 13339 11478
rect 13294 11440 13338 11447
rect 13294 11420 13306 11440
rect 13326 11420 13338 11440
rect 13294 11378 13338 11420
rect 9828 11259 9840 11279
rect 9860 11259 9872 11279
rect 9828 11221 9872 11259
rect 17318 11278 17362 11320
rect 17318 11258 17330 11278
rect 17350 11258 17362 11278
rect 17318 11251 17362 11258
rect 17317 11220 17362 11251
rect 17412 11278 17454 11320
rect 17412 11258 17426 11278
rect 17446 11258 17454 11278
rect 17412 11220 17454 11258
rect 17528 11278 17570 11320
rect 17528 11258 17536 11278
rect 17556 11258 17570 11278
rect 17528 11220 17570 11258
rect 17620 11278 17664 11320
rect 17620 11258 17632 11278
rect 17652 11258 17664 11278
rect 17620 11220 17664 11258
rect 17736 11278 17778 11320
rect 17736 11258 17744 11278
rect 17764 11258 17778 11278
rect 17736 11220 17778 11258
rect 17828 11278 17872 11320
rect 17828 11258 17840 11278
rect 17860 11258 17872 11278
rect 17828 11220 17872 11258
rect 17949 11278 17991 11320
rect 17949 11258 17957 11278
rect 17977 11258 17991 11278
rect 17949 11220 17991 11258
rect 18041 11278 18085 11320
rect 18041 11258 18053 11278
rect 18073 11258 18085 11278
rect 18041 11220 18085 11258
rect 19813 11273 19857 11315
rect 19813 11253 19825 11273
rect 19845 11253 19857 11273
rect 19813 11246 19857 11253
rect 19812 11215 19857 11246
rect 19907 11273 19949 11315
rect 19907 11253 19921 11273
rect 19941 11253 19949 11273
rect 19907 11215 19949 11253
rect 20023 11273 20065 11315
rect 20023 11253 20031 11273
rect 20051 11253 20065 11273
rect 20023 11215 20065 11253
rect 20115 11273 20159 11315
rect 20115 11253 20127 11273
rect 20147 11253 20159 11273
rect 20115 11215 20159 11253
rect 20231 11273 20273 11315
rect 20231 11253 20239 11273
rect 20259 11253 20273 11273
rect 20231 11215 20273 11253
rect 20323 11273 20367 11315
rect 20323 11253 20335 11273
rect 20355 11253 20367 11273
rect 20323 11215 20367 11253
rect 20444 11273 20486 11315
rect 20444 11253 20452 11273
rect 20472 11253 20486 11273
rect 20444 11215 20486 11253
rect 20536 11273 20580 11315
rect 20536 11253 20548 11273
rect 20568 11253 20580 11273
rect 20536 11215 20580 11253
rect 815 10771 859 10809
rect 815 10751 827 10771
rect 847 10751 859 10771
rect 815 10709 859 10751
rect 909 10771 951 10809
rect 909 10751 923 10771
rect 943 10751 951 10771
rect 909 10709 951 10751
rect 1028 10771 1072 10809
rect 1028 10751 1040 10771
rect 1060 10751 1072 10771
rect 1028 10709 1072 10751
rect 1122 10771 1164 10809
rect 1122 10751 1136 10771
rect 1156 10751 1164 10771
rect 1122 10709 1164 10751
rect 1236 10771 1280 10809
rect 1236 10751 1248 10771
rect 1268 10751 1280 10771
rect 1236 10709 1280 10751
rect 1330 10771 1372 10809
rect 1330 10751 1344 10771
rect 1364 10751 1372 10771
rect 1330 10709 1372 10751
rect 1446 10771 1488 10809
rect 1446 10751 1454 10771
rect 1474 10751 1488 10771
rect 1446 10709 1488 10751
rect 1538 10778 1583 10809
rect 1538 10771 1582 10778
rect 1538 10751 1550 10771
rect 1570 10751 1582 10771
rect 1538 10709 1582 10751
rect 3353 10768 3397 10806
rect 3353 10748 3365 10768
rect 3385 10748 3397 10768
rect 3353 10706 3397 10748
rect 3447 10768 3489 10806
rect 3447 10748 3461 10768
rect 3481 10748 3489 10768
rect 3447 10706 3489 10748
rect 3566 10768 3610 10806
rect 3566 10748 3578 10768
rect 3598 10748 3610 10768
rect 3566 10706 3610 10748
rect 3660 10768 3702 10806
rect 3660 10748 3674 10768
rect 3694 10748 3702 10768
rect 3660 10706 3702 10748
rect 3774 10768 3818 10806
rect 3774 10748 3786 10768
rect 3806 10748 3818 10768
rect 3774 10706 3818 10748
rect 3868 10768 3910 10806
rect 3868 10748 3882 10768
rect 3902 10748 3910 10768
rect 3868 10706 3910 10748
rect 3984 10768 4026 10806
rect 3984 10748 3992 10768
rect 4012 10748 4026 10768
rect 3984 10706 4026 10748
rect 4076 10775 4121 10806
rect 4076 10768 4120 10775
rect 4076 10748 4088 10768
rect 4108 10748 4120 10768
rect 4076 10706 4120 10748
rect 11523 10765 11567 10803
rect 11523 10745 11535 10765
rect 11555 10745 11567 10765
rect 8057 10604 8101 10646
rect 8057 10584 8069 10604
rect 8089 10584 8101 10604
rect 8057 10577 8101 10584
rect 8056 10546 8101 10577
rect 8151 10604 8193 10646
rect 8151 10584 8165 10604
rect 8185 10584 8193 10604
rect 8151 10546 8193 10584
rect 8267 10604 8309 10646
rect 8267 10584 8275 10604
rect 8295 10584 8309 10604
rect 8267 10546 8309 10584
rect 8359 10604 8403 10646
rect 8359 10584 8371 10604
rect 8391 10584 8403 10604
rect 8359 10546 8403 10584
rect 8475 10604 8517 10646
rect 8475 10584 8483 10604
rect 8503 10584 8517 10604
rect 8475 10546 8517 10584
rect 8567 10604 8611 10646
rect 8567 10584 8579 10604
rect 8599 10584 8611 10604
rect 8567 10546 8611 10584
rect 8688 10604 8730 10646
rect 8688 10584 8696 10604
rect 8716 10584 8730 10604
rect 8688 10546 8730 10584
rect 8780 10604 8824 10646
rect 11523 10703 11567 10745
rect 11617 10765 11659 10803
rect 11617 10745 11631 10765
rect 11651 10745 11659 10765
rect 11617 10703 11659 10745
rect 11736 10765 11780 10803
rect 11736 10745 11748 10765
rect 11768 10745 11780 10765
rect 11736 10703 11780 10745
rect 11830 10765 11872 10803
rect 11830 10745 11844 10765
rect 11864 10745 11872 10765
rect 11830 10703 11872 10745
rect 11944 10765 11988 10803
rect 11944 10745 11956 10765
rect 11976 10745 11988 10765
rect 11944 10703 11988 10745
rect 12038 10765 12080 10803
rect 12038 10745 12052 10765
rect 12072 10745 12080 10765
rect 12038 10703 12080 10745
rect 12154 10765 12196 10803
rect 12154 10745 12162 10765
rect 12182 10745 12196 10765
rect 12154 10703 12196 10745
rect 12246 10772 12291 10803
rect 12246 10765 12290 10772
rect 12246 10745 12258 10765
rect 12278 10745 12290 10765
rect 12246 10703 12290 10745
rect 14061 10762 14105 10800
rect 14061 10742 14073 10762
rect 14093 10742 14105 10762
rect 8780 10584 8792 10604
rect 8812 10584 8824 10604
rect 8780 10546 8824 10584
rect 9105 10600 9149 10642
rect 9105 10580 9117 10600
rect 9137 10580 9149 10600
rect 9105 10573 9149 10580
rect 9104 10542 9149 10573
rect 9199 10600 9241 10642
rect 9199 10580 9213 10600
rect 9233 10580 9241 10600
rect 9199 10542 9241 10580
rect 9315 10600 9357 10642
rect 9315 10580 9323 10600
rect 9343 10580 9357 10600
rect 9315 10542 9357 10580
rect 9407 10600 9451 10642
rect 9407 10580 9419 10600
rect 9439 10580 9451 10600
rect 9407 10542 9451 10580
rect 9523 10600 9565 10642
rect 9523 10580 9531 10600
rect 9551 10580 9565 10600
rect 9523 10542 9565 10580
rect 9615 10600 9659 10642
rect 9615 10580 9627 10600
rect 9647 10580 9659 10600
rect 9615 10542 9659 10580
rect 9736 10600 9778 10642
rect 9736 10580 9744 10600
rect 9764 10580 9778 10600
rect 9736 10542 9778 10580
rect 9828 10600 9872 10642
rect 9828 10580 9840 10600
rect 9860 10580 9872 10600
rect 14061 10700 14105 10742
rect 14155 10762 14197 10800
rect 14155 10742 14169 10762
rect 14189 10742 14197 10762
rect 14155 10700 14197 10742
rect 14274 10762 14318 10800
rect 14274 10742 14286 10762
rect 14306 10742 14318 10762
rect 14274 10700 14318 10742
rect 14368 10762 14410 10800
rect 14368 10742 14382 10762
rect 14402 10742 14410 10762
rect 14368 10700 14410 10742
rect 14482 10762 14526 10800
rect 14482 10742 14494 10762
rect 14514 10742 14526 10762
rect 14482 10700 14526 10742
rect 14576 10762 14618 10800
rect 14576 10742 14590 10762
rect 14610 10742 14618 10762
rect 14576 10700 14618 10742
rect 14692 10762 14734 10800
rect 14692 10742 14700 10762
rect 14720 10742 14734 10762
rect 14692 10700 14734 10742
rect 14784 10769 14829 10800
rect 14784 10762 14828 10769
rect 14784 10742 14796 10762
rect 14816 10742 14828 10762
rect 14784 10700 14828 10742
rect 9828 10542 9872 10580
rect 18765 10598 18809 10640
rect 18765 10578 18777 10598
rect 18797 10578 18809 10598
rect 18765 10571 18809 10578
rect 18764 10540 18809 10571
rect 18859 10598 18901 10640
rect 18859 10578 18873 10598
rect 18893 10578 18901 10598
rect 18859 10540 18901 10578
rect 18975 10598 19017 10640
rect 18975 10578 18983 10598
rect 19003 10578 19017 10598
rect 18975 10540 19017 10578
rect 19067 10598 19111 10640
rect 19067 10578 19079 10598
rect 19099 10578 19111 10598
rect 19067 10540 19111 10578
rect 19183 10598 19225 10640
rect 19183 10578 19191 10598
rect 19211 10578 19225 10598
rect 19183 10540 19225 10578
rect 19275 10598 19319 10640
rect 19275 10578 19287 10598
rect 19307 10578 19319 10598
rect 19275 10540 19319 10578
rect 19396 10598 19438 10640
rect 19396 10578 19404 10598
rect 19424 10578 19438 10598
rect 19396 10540 19438 10578
rect 19488 10598 19532 10640
rect 19488 10578 19500 10598
rect 19520 10578 19532 10598
rect 19488 10540 19532 10578
rect 19813 10594 19857 10636
rect 19813 10574 19825 10594
rect 19845 10574 19857 10594
rect 19813 10567 19857 10574
rect 19812 10536 19857 10567
rect 19907 10594 19949 10636
rect 19907 10574 19921 10594
rect 19941 10574 19949 10594
rect 19907 10536 19949 10574
rect 20023 10594 20065 10636
rect 20023 10574 20031 10594
rect 20051 10574 20065 10594
rect 20023 10536 20065 10574
rect 20115 10594 20159 10636
rect 20115 10574 20127 10594
rect 20147 10574 20159 10594
rect 20115 10536 20159 10574
rect 20231 10594 20273 10636
rect 20231 10574 20239 10594
rect 20259 10574 20273 10594
rect 20231 10536 20273 10574
rect 20323 10594 20367 10636
rect 20323 10574 20335 10594
rect 20355 10574 20367 10594
rect 20323 10536 20367 10574
rect 20444 10594 20486 10636
rect 20444 10574 20452 10594
rect 20472 10574 20486 10594
rect 20444 10536 20486 10574
rect 20536 10594 20580 10636
rect 20536 10574 20548 10594
rect 20568 10574 20580 10594
rect 20536 10536 20580 10574
rect 816 9930 860 9968
rect 816 9910 828 9930
rect 848 9910 860 9930
rect 816 9868 860 9910
rect 910 9930 952 9968
rect 910 9910 924 9930
rect 944 9910 952 9930
rect 910 9868 952 9910
rect 1029 9930 1073 9968
rect 1029 9910 1041 9930
rect 1061 9910 1073 9930
rect 1029 9868 1073 9910
rect 1123 9930 1165 9968
rect 1123 9910 1137 9930
rect 1157 9910 1165 9930
rect 1123 9868 1165 9910
rect 1237 9930 1281 9968
rect 1237 9910 1249 9930
rect 1269 9910 1281 9930
rect 1237 9868 1281 9910
rect 1331 9930 1373 9968
rect 1331 9910 1345 9930
rect 1365 9910 1373 9930
rect 1331 9868 1373 9910
rect 1447 9930 1489 9968
rect 1447 9910 1455 9930
rect 1475 9910 1489 9930
rect 1447 9868 1489 9910
rect 1539 9937 1584 9968
rect 1539 9930 1583 9937
rect 1539 9910 1551 9930
rect 1571 9910 1583 9930
rect 1539 9868 1583 9910
rect 1864 9926 1908 9964
rect 1864 9906 1876 9926
rect 1896 9906 1908 9926
rect 1864 9864 1908 9906
rect 1958 9926 2000 9964
rect 1958 9906 1972 9926
rect 1992 9906 2000 9926
rect 1958 9864 2000 9906
rect 2077 9926 2121 9964
rect 2077 9906 2089 9926
rect 2109 9906 2121 9926
rect 2077 9864 2121 9906
rect 2171 9926 2213 9964
rect 2171 9906 2185 9926
rect 2205 9906 2213 9926
rect 2171 9864 2213 9906
rect 2285 9926 2329 9964
rect 2285 9906 2297 9926
rect 2317 9906 2329 9926
rect 2285 9864 2329 9906
rect 2379 9926 2421 9964
rect 2379 9906 2393 9926
rect 2413 9906 2421 9926
rect 2379 9864 2421 9906
rect 2495 9926 2537 9964
rect 2495 9906 2503 9926
rect 2523 9906 2537 9926
rect 2495 9864 2537 9906
rect 2587 9933 2632 9964
rect 2587 9926 2631 9933
rect 2587 9906 2599 9926
rect 2619 9906 2631 9926
rect 2587 9864 2631 9906
rect 11524 9924 11568 9962
rect 6568 9762 6612 9804
rect 6568 9742 6580 9762
rect 6600 9742 6612 9762
rect 6568 9735 6612 9742
rect 6567 9704 6612 9735
rect 6662 9762 6704 9804
rect 6662 9742 6676 9762
rect 6696 9742 6704 9762
rect 6662 9704 6704 9742
rect 6778 9762 6820 9804
rect 6778 9742 6786 9762
rect 6806 9742 6820 9762
rect 6778 9704 6820 9742
rect 6870 9762 6914 9804
rect 6870 9742 6882 9762
rect 6902 9742 6914 9762
rect 6870 9704 6914 9742
rect 6986 9762 7028 9804
rect 6986 9742 6994 9762
rect 7014 9742 7028 9762
rect 6986 9704 7028 9742
rect 7078 9762 7122 9804
rect 7078 9742 7090 9762
rect 7110 9742 7122 9762
rect 7078 9704 7122 9742
rect 7199 9762 7241 9804
rect 7199 9742 7207 9762
rect 7227 9742 7241 9762
rect 7199 9704 7241 9742
rect 7291 9762 7335 9804
rect 11524 9904 11536 9924
rect 11556 9904 11568 9924
rect 11524 9862 11568 9904
rect 11618 9924 11660 9962
rect 11618 9904 11632 9924
rect 11652 9904 11660 9924
rect 11618 9862 11660 9904
rect 11737 9924 11781 9962
rect 11737 9904 11749 9924
rect 11769 9904 11781 9924
rect 11737 9862 11781 9904
rect 11831 9924 11873 9962
rect 11831 9904 11845 9924
rect 11865 9904 11873 9924
rect 11831 9862 11873 9904
rect 11945 9924 11989 9962
rect 11945 9904 11957 9924
rect 11977 9904 11989 9924
rect 11945 9862 11989 9904
rect 12039 9924 12081 9962
rect 12039 9904 12053 9924
rect 12073 9904 12081 9924
rect 12039 9862 12081 9904
rect 12155 9924 12197 9962
rect 12155 9904 12163 9924
rect 12183 9904 12197 9924
rect 12155 9862 12197 9904
rect 12247 9931 12292 9962
rect 12247 9924 12291 9931
rect 12247 9904 12259 9924
rect 12279 9904 12291 9924
rect 12247 9862 12291 9904
rect 12572 9920 12616 9958
rect 12572 9900 12584 9920
rect 12604 9900 12616 9920
rect 7291 9742 7303 9762
rect 7323 9742 7335 9762
rect 7291 9704 7335 9742
rect 9106 9759 9150 9801
rect 9106 9739 9118 9759
rect 9138 9739 9150 9759
rect 9106 9732 9150 9739
rect 9105 9701 9150 9732
rect 9200 9759 9242 9801
rect 9200 9739 9214 9759
rect 9234 9739 9242 9759
rect 9200 9701 9242 9739
rect 9316 9759 9358 9801
rect 9316 9739 9324 9759
rect 9344 9739 9358 9759
rect 9316 9701 9358 9739
rect 9408 9759 9452 9801
rect 9408 9739 9420 9759
rect 9440 9739 9452 9759
rect 9408 9701 9452 9739
rect 9524 9759 9566 9801
rect 9524 9739 9532 9759
rect 9552 9739 9566 9759
rect 9524 9701 9566 9739
rect 9616 9759 9660 9801
rect 9616 9739 9628 9759
rect 9648 9739 9660 9759
rect 9616 9701 9660 9739
rect 9737 9759 9779 9801
rect 9737 9739 9745 9759
rect 9765 9739 9779 9759
rect 9737 9701 9779 9739
rect 9829 9759 9873 9801
rect 12572 9858 12616 9900
rect 12666 9920 12708 9958
rect 12666 9900 12680 9920
rect 12700 9900 12708 9920
rect 12666 9858 12708 9900
rect 12785 9920 12829 9958
rect 12785 9900 12797 9920
rect 12817 9900 12829 9920
rect 12785 9858 12829 9900
rect 12879 9920 12921 9958
rect 12879 9900 12893 9920
rect 12913 9900 12921 9920
rect 12879 9858 12921 9900
rect 12993 9920 13037 9958
rect 12993 9900 13005 9920
rect 13025 9900 13037 9920
rect 12993 9858 13037 9900
rect 13087 9920 13129 9958
rect 13087 9900 13101 9920
rect 13121 9900 13129 9920
rect 13087 9858 13129 9900
rect 13203 9920 13245 9958
rect 13203 9900 13211 9920
rect 13231 9900 13245 9920
rect 13203 9858 13245 9900
rect 13295 9927 13340 9958
rect 13295 9920 13339 9927
rect 13295 9900 13307 9920
rect 13327 9900 13339 9920
rect 13295 9858 13339 9900
rect 9829 9739 9841 9759
rect 9861 9739 9873 9759
rect 9829 9701 9873 9739
rect 17276 9756 17320 9798
rect 17276 9736 17288 9756
rect 17308 9736 17320 9756
rect 17276 9729 17320 9736
rect 17275 9698 17320 9729
rect 17370 9756 17412 9798
rect 17370 9736 17384 9756
rect 17404 9736 17412 9756
rect 17370 9698 17412 9736
rect 17486 9756 17528 9798
rect 17486 9736 17494 9756
rect 17514 9736 17528 9756
rect 17486 9698 17528 9736
rect 17578 9756 17622 9798
rect 17578 9736 17590 9756
rect 17610 9736 17622 9756
rect 17578 9698 17622 9736
rect 17694 9756 17736 9798
rect 17694 9736 17702 9756
rect 17722 9736 17736 9756
rect 17694 9698 17736 9736
rect 17786 9756 17830 9798
rect 17786 9736 17798 9756
rect 17818 9736 17830 9756
rect 17786 9698 17830 9736
rect 17907 9756 17949 9798
rect 17907 9736 17915 9756
rect 17935 9736 17949 9756
rect 17907 9698 17949 9736
rect 17999 9756 18043 9798
rect 17999 9736 18011 9756
rect 18031 9736 18043 9756
rect 17999 9698 18043 9736
rect 19814 9753 19858 9795
rect 19814 9733 19826 9753
rect 19846 9733 19858 9753
rect 19814 9726 19858 9733
rect 19813 9695 19858 9726
rect 19908 9753 19950 9795
rect 19908 9733 19922 9753
rect 19942 9733 19950 9753
rect 19908 9695 19950 9733
rect 20024 9753 20066 9795
rect 20024 9733 20032 9753
rect 20052 9733 20066 9753
rect 20024 9695 20066 9733
rect 20116 9753 20160 9795
rect 20116 9733 20128 9753
rect 20148 9733 20160 9753
rect 20116 9695 20160 9733
rect 20232 9753 20274 9795
rect 20232 9733 20240 9753
rect 20260 9733 20274 9753
rect 20232 9695 20274 9733
rect 20324 9753 20368 9795
rect 20324 9733 20336 9753
rect 20356 9733 20368 9753
rect 20324 9695 20368 9733
rect 20445 9753 20487 9795
rect 20445 9733 20453 9753
rect 20473 9733 20487 9753
rect 20445 9695 20487 9733
rect 20537 9753 20581 9795
rect 20537 9733 20549 9753
rect 20569 9733 20581 9753
rect 20537 9695 20581 9733
rect 816 9251 860 9289
rect 816 9231 828 9251
rect 848 9231 860 9251
rect 816 9189 860 9231
rect 910 9251 952 9289
rect 910 9231 924 9251
rect 944 9231 952 9251
rect 910 9189 952 9231
rect 1029 9251 1073 9289
rect 1029 9231 1041 9251
rect 1061 9231 1073 9251
rect 1029 9189 1073 9231
rect 1123 9251 1165 9289
rect 1123 9231 1137 9251
rect 1157 9231 1165 9251
rect 1123 9189 1165 9231
rect 1237 9251 1281 9289
rect 1237 9231 1249 9251
rect 1269 9231 1281 9251
rect 1237 9189 1281 9231
rect 1331 9251 1373 9289
rect 1331 9231 1345 9251
rect 1365 9231 1373 9251
rect 1331 9189 1373 9231
rect 1447 9251 1489 9289
rect 1447 9231 1455 9251
rect 1475 9231 1489 9251
rect 1447 9189 1489 9231
rect 1539 9258 1584 9289
rect 1539 9251 1583 9258
rect 1539 9231 1551 9251
rect 1571 9231 1583 9251
rect 1539 9189 1583 9231
rect 3311 9246 3355 9284
rect 3311 9226 3323 9246
rect 3343 9226 3355 9246
rect 3311 9184 3355 9226
rect 3405 9246 3447 9284
rect 3405 9226 3419 9246
rect 3439 9226 3447 9246
rect 3405 9184 3447 9226
rect 3524 9246 3568 9284
rect 3524 9226 3536 9246
rect 3556 9226 3568 9246
rect 3524 9184 3568 9226
rect 3618 9246 3660 9284
rect 3618 9226 3632 9246
rect 3652 9226 3660 9246
rect 3618 9184 3660 9226
rect 3732 9246 3776 9284
rect 3732 9226 3744 9246
rect 3764 9226 3776 9246
rect 3732 9184 3776 9226
rect 3826 9246 3868 9284
rect 3826 9226 3840 9246
rect 3860 9226 3868 9246
rect 3826 9184 3868 9226
rect 3942 9246 3984 9284
rect 3942 9226 3950 9246
rect 3970 9226 3984 9246
rect 3942 9184 3984 9226
rect 4034 9253 4079 9284
rect 4034 9246 4078 9253
rect 4034 9226 4046 9246
rect 4066 9226 4078 9246
rect 4034 9184 4078 9226
rect 11524 9245 11568 9283
rect 11524 9225 11536 9245
rect 11556 9225 11568 9245
rect 8058 9084 8102 9126
rect 8058 9064 8070 9084
rect 8090 9064 8102 9084
rect 8058 9057 8102 9064
rect 8057 9026 8102 9057
rect 8152 9084 8194 9126
rect 8152 9064 8166 9084
rect 8186 9064 8194 9084
rect 8152 9026 8194 9064
rect 8268 9084 8310 9126
rect 8268 9064 8276 9084
rect 8296 9064 8310 9084
rect 8268 9026 8310 9064
rect 8360 9084 8404 9126
rect 8360 9064 8372 9084
rect 8392 9064 8404 9084
rect 8360 9026 8404 9064
rect 8476 9084 8518 9126
rect 8476 9064 8484 9084
rect 8504 9064 8518 9084
rect 8476 9026 8518 9064
rect 8568 9084 8612 9126
rect 8568 9064 8580 9084
rect 8600 9064 8612 9084
rect 8568 9026 8612 9064
rect 8689 9084 8731 9126
rect 8689 9064 8697 9084
rect 8717 9064 8731 9084
rect 8689 9026 8731 9064
rect 8781 9084 8825 9126
rect 11524 9183 11568 9225
rect 11618 9245 11660 9283
rect 11618 9225 11632 9245
rect 11652 9225 11660 9245
rect 11618 9183 11660 9225
rect 11737 9245 11781 9283
rect 11737 9225 11749 9245
rect 11769 9225 11781 9245
rect 11737 9183 11781 9225
rect 11831 9245 11873 9283
rect 11831 9225 11845 9245
rect 11865 9225 11873 9245
rect 11831 9183 11873 9225
rect 11945 9245 11989 9283
rect 11945 9225 11957 9245
rect 11977 9225 11989 9245
rect 11945 9183 11989 9225
rect 12039 9245 12081 9283
rect 12039 9225 12053 9245
rect 12073 9225 12081 9245
rect 12039 9183 12081 9225
rect 12155 9245 12197 9283
rect 12155 9225 12163 9245
rect 12183 9225 12197 9245
rect 12155 9183 12197 9225
rect 12247 9252 12292 9283
rect 12247 9245 12291 9252
rect 12247 9225 12259 9245
rect 12279 9225 12291 9245
rect 12247 9183 12291 9225
rect 14019 9240 14063 9278
rect 14019 9220 14031 9240
rect 14051 9220 14063 9240
rect 8781 9064 8793 9084
rect 8813 9064 8825 9084
rect 8781 9026 8825 9064
rect 9106 9080 9150 9122
rect 9106 9060 9118 9080
rect 9138 9060 9150 9080
rect 9106 9053 9150 9060
rect 9105 9022 9150 9053
rect 9200 9080 9242 9122
rect 9200 9060 9214 9080
rect 9234 9060 9242 9080
rect 9200 9022 9242 9060
rect 9316 9080 9358 9122
rect 9316 9060 9324 9080
rect 9344 9060 9358 9080
rect 9316 9022 9358 9060
rect 9408 9080 9452 9122
rect 9408 9060 9420 9080
rect 9440 9060 9452 9080
rect 9408 9022 9452 9060
rect 9524 9080 9566 9122
rect 9524 9060 9532 9080
rect 9552 9060 9566 9080
rect 9524 9022 9566 9060
rect 9616 9080 9660 9122
rect 9616 9060 9628 9080
rect 9648 9060 9660 9080
rect 9616 9022 9660 9060
rect 9737 9080 9779 9122
rect 9737 9060 9745 9080
rect 9765 9060 9779 9080
rect 9737 9022 9779 9060
rect 9829 9080 9873 9122
rect 9829 9060 9841 9080
rect 9861 9060 9873 9080
rect 14019 9178 14063 9220
rect 14113 9240 14155 9278
rect 14113 9220 14127 9240
rect 14147 9220 14155 9240
rect 14113 9178 14155 9220
rect 14232 9240 14276 9278
rect 14232 9220 14244 9240
rect 14264 9220 14276 9240
rect 14232 9178 14276 9220
rect 14326 9240 14368 9278
rect 14326 9220 14340 9240
rect 14360 9220 14368 9240
rect 14326 9178 14368 9220
rect 14440 9240 14484 9278
rect 14440 9220 14452 9240
rect 14472 9220 14484 9240
rect 14440 9178 14484 9220
rect 14534 9240 14576 9278
rect 14534 9220 14548 9240
rect 14568 9220 14576 9240
rect 14534 9178 14576 9220
rect 14650 9240 14692 9278
rect 14650 9220 14658 9240
rect 14678 9220 14692 9240
rect 14650 9178 14692 9220
rect 14742 9247 14787 9278
rect 14742 9240 14786 9247
rect 14742 9220 14754 9240
rect 14774 9220 14786 9240
rect 14742 9178 14786 9220
rect 9829 9022 9873 9060
rect 18766 9078 18810 9120
rect 18766 9058 18778 9078
rect 18798 9058 18810 9078
rect 18766 9051 18810 9058
rect 18765 9020 18810 9051
rect 18860 9078 18902 9120
rect 18860 9058 18874 9078
rect 18894 9058 18902 9078
rect 18860 9020 18902 9058
rect 18976 9078 19018 9120
rect 18976 9058 18984 9078
rect 19004 9058 19018 9078
rect 18976 9020 19018 9058
rect 19068 9078 19112 9120
rect 19068 9058 19080 9078
rect 19100 9058 19112 9078
rect 19068 9020 19112 9058
rect 19184 9078 19226 9120
rect 19184 9058 19192 9078
rect 19212 9058 19226 9078
rect 19184 9020 19226 9058
rect 19276 9078 19320 9120
rect 19276 9058 19288 9078
rect 19308 9058 19320 9078
rect 19276 9020 19320 9058
rect 19397 9078 19439 9120
rect 19397 9058 19405 9078
rect 19425 9058 19439 9078
rect 19397 9020 19439 9058
rect 19489 9078 19533 9120
rect 19489 9058 19501 9078
rect 19521 9058 19533 9078
rect 19489 9020 19533 9058
rect 19814 9074 19858 9116
rect 19814 9054 19826 9074
rect 19846 9054 19858 9074
rect 19814 9047 19858 9054
rect 19813 9016 19858 9047
rect 19908 9074 19950 9116
rect 19908 9054 19922 9074
rect 19942 9054 19950 9074
rect 19908 9016 19950 9054
rect 20024 9074 20066 9116
rect 20024 9054 20032 9074
rect 20052 9054 20066 9074
rect 20024 9016 20066 9054
rect 20116 9074 20160 9116
rect 20116 9054 20128 9074
rect 20148 9054 20160 9074
rect 20116 9016 20160 9054
rect 20232 9074 20274 9116
rect 20232 9054 20240 9074
rect 20260 9054 20274 9074
rect 20232 9016 20274 9054
rect 20324 9074 20368 9116
rect 20324 9054 20336 9074
rect 20356 9054 20368 9074
rect 20324 9016 20368 9054
rect 20445 9074 20487 9116
rect 20445 9054 20453 9074
rect 20473 9054 20487 9074
rect 20445 9016 20487 9054
rect 20537 9074 20581 9116
rect 20537 9054 20549 9074
rect 20569 9054 20581 9074
rect 20537 9016 20581 9054
rect 816 8483 860 8521
rect 816 8463 828 8483
rect 848 8463 860 8483
rect 816 8421 860 8463
rect 910 8483 952 8521
rect 910 8463 924 8483
rect 944 8463 952 8483
rect 910 8421 952 8463
rect 1029 8483 1073 8521
rect 1029 8463 1041 8483
rect 1061 8463 1073 8483
rect 1029 8421 1073 8463
rect 1123 8483 1165 8521
rect 1123 8463 1137 8483
rect 1157 8463 1165 8483
rect 1123 8421 1165 8463
rect 1237 8483 1281 8521
rect 1237 8463 1249 8483
rect 1269 8463 1281 8483
rect 1237 8421 1281 8463
rect 1331 8483 1373 8521
rect 1331 8463 1345 8483
rect 1365 8463 1373 8483
rect 1331 8421 1373 8463
rect 1447 8483 1489 8521
rect 1447 8463 1455 8483
rect 1475 8463 1489 8483
rect 1447 8421 1489 8463
rect 1539 8490 1584 8521
rect 1539 8483 1583 8490
rect 1539 8463 1551 8483
rect 1571 8463 1583 8483
rect 1539 8421 1583 8463
rect 1864 8479 1908 8517
rect 1864 8459 1876 8479
rect 1896 8459 1908 8479
rect 1864 8417 1908 8459
rect 1958 8479 2000 8517
rect 1958 8459 1972 8479
rect 1992 8459 2000 8479
rect 1958 8417 2000 8459
rect 2077 8479 2121 8517
rect 2077 8459 2089 8479
rect 2109 8459 2121 8479
rect 2077 8417 2121 8459
rect 2171 8479 2213 8517
rect 2171 8459 2185 8479
rect 2205 8459 2213 8479
rect 2171 8417 2213 8459
rect 2285 8479 2329 8517
rect 2285 8459 2297 8479
rect 2317 8459 2329 8479
rect 2285 8417 2329 8459
rect 2379 8479 2421 8517
rect 2379 8459 2393 8479
rect 2413 8459 2421 8479
rect 2379 8417 2421 8459
rect 2495 8479 2537 8517
rect 2495 8459 2503 8479
rect 2523 8459 2537 8479
rect 2495 8417 2537 8459
rect 2587 8486 2632 8517
rect 2587 8479 2631 8486
rect 2587 8459 2599 8479
rect 2619 8459 2631 8479
rect 2587 8417 2631 8459
rect 11524 8477 11568 8515
rect 6611 8317 6655 8359
rect 6611 8297 6623 8317
rect 6643 8297 6655 8317
rect 6611 8290 6655 8297
rect 6610 8259 6655 8290
rect 6705 8317 6747 8359
rect 6705 8297 6719 8317
rect 6739 8297 6747 8317
rect 6705 8259 6747 8297
rect 6821 8317 6863 8359
rect 6821 8297 6829 8317
rect 6849 8297 6863 8317
rect 6821 8259 6863 8297
rect 6913 8317 6957 8359
rect 6913 8297 6925 8317
rect 6945 8297 6957 8317
rect 6913 8259 6957 8297
rect 7029 8317 7071 8359
rect 7029 8297 7037 8317
rect 7057 8297 7071 8317
rect 7029 8259 7071 8297
rect 7121 8317 7165 8359
rect 7121 8297 7133 8317
rect 7153 8297 7165 8317
rect 7121 8259 7165 8297
rect 7242 8317 7284 8359
rect 7242 8297 7250 8317
rect 7270 8297 7284 8317
rect 7242 8259 7284 8297
rect 7334 8317 7378 8359
rect 11524 8457 11536 8477
rect 11556 8457 11568 8477
rect 11524 8415 11568 8457
rect 11618 8477 11660 8515
rect 11618 8457 11632 8477
rect 11652 8457 11660 8477
rect 11618 8415 11660 8457
rect 11737 8477 11781 8515
rect 11737 8457 11749 8477
rect 11769 8457 11781 8477
rect 11737 8415 11781 8457
rect 11831 8477 11873 8515
rect 11831 8457 11845 8477
rect 11865 8457 11873 8477
rect 11831 8415 11873 8457
rect 11945 8477 11989 8515
rect 11945 8457 11957 8477
rect 11977 8457 11989 8477
rect 11945 8415 11989 8457
rect 12039 8477 12081 8515
rect 12039 8457 12053 8477
rect 12073 8457 12081 8477
rect 12039 8415 12081 8457
rect 12155 8477 12197 8515
rect 12155 8457 12163 8477
rect 12183 8457 12197 8477
rect 12155 8415 12197 8457
rect 12247 8484 12292 8515
rect 12247 8477 12291 8484
rect 12247 8457 12259 8477
rect 12279 8457 12291 8477
rect 12247 8415 12291 8457
rect 12572 8473 12616 8511
rect 12572 8453 12584 8473
rect 12604 8453 12616 8473
rect 7334 8297 7346 8317
rect 7366 8297 7378 8317
rect 7334 8259 7378 8297
rect 9106 8312 9150 8354
rect 9106 8292 9118 8312
rect 9138 8292 9150 8312
rect 9106 8285 9150 8292
rect 9105 8254 9150 8285
rect 9200 8312 9242 8354
rect 9200 8292 9214 8312
rect 9234 8292 9242 8312
rect 9200 8254 9242 8292
rect 9316 8312 9358 8354
rect 9316 8292 9324 8312
rect 9344 8292 9358 8312
rect 9316 8254 9358 8292
rect 9408 8312 9452 8354
rect 9408 8292 9420 8312
rect 9440 8292 9452 8312
rect 9408 8254 9452 8292
rect 9524 8312 9566 8354
rect 9524 8292 9532 8312
rect 9552 8292 9566 8312
rect 9524 8254 9566 8292
rect 9616 8312 9660 8354
rect 9616 8292 9628 8312
rect 9648 8292 9660 8312
rect 9616 8254 9660 8292
rect 9737 8312 9779 8354
rect 9737 8292 9745 8312
rect 9765 8292 9779 8312
rect 9737 8254 9779 8292
rect 9829 8312 9873 8354
rect 12572 8411 12616 8453
rect 12666 8473 12708 8511
rect 12666 8453 12680 8473
rect 12700 8453 12708 8473
rect 12666 8411 12708 8453
rect 12785 8473 12829 8511
rect 12785 8453 12797 8473
rect 12817 8453 12829 8473
rect 12785 8411 12829 8453
rect 12879 8473 12921 8511
rect 12879 8453 12893 8473
rect 12913 8453 12921 8473
rect 12879 8411 12921 8453
rect 12993 8473 13037 8511
rect 12993 8453 13005 8473
rect 13025 8453 13037 8473
rect 12993 8411 13037 8453
rect 13087 8473 13129 8511
rect 13087 8453 13101 8473
rect 13121 8453 13129 8473
rect 13087 8411 13129 8453
rect 13203 8473 13245 8511
rect 13203 8453 13211 8473
rect 13231 8453 13245 8473
rect 13203 8411 13245 8453
rect 13295 8480 13340 8511
rect 13295 8473 13339 8480
rect 13295 8453 13307 8473
rect 13327 8453 13339 8473
rect 13295 8411 13339 8453
rect 9829 8292 9841 8312
rect 9861 8292 9873 8312
rect 9829 8254 9873 8292
rect 17319 8311 17363 8353
rect 17319 8291 17331 8311
rect 17351 8291 17363 8311
rect 17319 8284 17363 8291
rect 17318 8253 17363 8284
rect 17413 8311 17455 8353
rect 17413 8291 17427 8311
rect 17447 8291 17455 8311
rect 17413 8253 17455 8291
rect 17529 8311 17571 8353
rect 17529 8291 17537 8311
rect 17557 8291 17571 8311
rect 17529 8253 17571 8291
rect 17621 8311 17665 8353
rect 17621 8291 17633 8311
rect 17653 8291 17665 8311
rect 17621 8253 17665 8291
rect 17737 8311 17779 8353
rect 17737 8291 17745 8311
rect 17765 8291 17779 8311
rect 17737 8253 17779 8291
rect 17829 8311 17873 8353
rect 17829 8291 17841 8311
rect 17861 8291 17873 8311
rect 17829 8253 17873 8291
rect 17950 8311 17992 8353
rect 17950 8291 17958 8311
rect 17978 8291 17992 8311
rect 17950 8253 17992 8291
rect 18042 8311 18086 8353
rect 18042 8291 18054 8311
rect 18074 8291 18086 8311
rect 18042 8253 18086 8291
rect 19814 8306 19858 8348
rect 19814 8286 19826 8306
rect 19846 8286 19858 8306
rect 19814 8279 19858 8286
rect 19813 8248 19858 8279
rect 19908 8306 19950 8348
rect 19908 8286 19922 8306
rect 19942 8286 19950 8306
rect 19908 8248 19950 8286
rect 20024 8306 20066 8348
rect 20024 8286 20032 8306
rect 20052 8286 20066 8306
rect 20024 8248 20066 8286
rect 20116 8306 20160 8348
rect 20116 8286 20128 8306
rect 20148 8286 20160 8306
rect 20116 8248 20160 8286
rect 20232 8306 20274 8348
rect 20232 8286 20240 8306
rect 20260 8286 20274 8306
rect 20232 8248 20274 8286
rect 20324 8306 20368 8348
rect 20324 8286 20336 8306
rect 20356 8286 20368 8306
rect 20324 8248 20368 8286
rect 20445 8306 20487 8348
rect 20445 8286 20453 8306
rect 20473 8286 20487 8306
rect 20445 8248 20487 8286
rect 20537 8306 20581 8348
rect 20537 8286 20549 8306
rect 20569 8286 20581 8306
rect 20537 8248 20581 8286
rect 816 7804 860 7842
rect 816 7784 828 7804
rect 848 7784 860 7804
rect 816 7742 860 7784
rect 910 7804 952 7842
rect 910 7784 924 7804
rect 944 7784 952 7804
rect 910 7742 952 7784
rect 1029 7804 1073 7842
rect 1029 7784 1041 7804
rect 1061 7784 1073 7804
rect 1029 7742 1073 7784
rect 1123 7804 1165 7842
rect 1123 7784 1137 7804
rect 1157 7784 1165 7804
rect 1123 7742 1165 7784
rect 1237 7804 1281 7842
rect 1237 7784 1249 7804
rect 1269 7784 1281 7804
rect 1237 7742 1281 7784
rect 1331 7804 1373 7842
rect 1331 7784 1345 7804
rect 1365 7784 1373 7804
rect 1331 7742 1373 7784
rect 1447 7804 1489 7842
rect 1447 7784 1455 7804
rect 1475 7784 1489 7804
rect 1447 7742 1489 7784
rect 1539 7811 1584 7842
rect 1539 7804 1583 7811
rect 1539 7784 1551 7804
rect 1571 7784 1583 7804
rect 1539 7742 1583 7784
rect 4419 7795 4463 7833
rect 4419 7775 4431 7795
rect 4451 7775 4463 7795
rect 4419 7733 4463 7775
rect 4513 7795 4555 7833
rect 4513 7775 4527 7795
rect 4547 7775 4555 7795
rect 4513 7733 4555 7775
rect 4632 7795 4676 7833
rect 4632 7775 4644 7795
rect 4664 7775 4676 7795
rect 4632 7733 4676 7775
rect 4726 7795 4768 7833
rect 4726 7775 4740 7795
rect 4760 7775 4768 7795
rect 4726 7733 4768 7775
rect 4840 7795 4884 7833
rect 4840 7775 4852 7795
rect 4872 7775 4884 7795
rect 4840 7733 4884 7775
rect 4934 7795 4976 7833
rect 4934 7775 4948 7795
rect 4968 7775 4976 7795
rect 4934 7733 4976 7775
rect 5050 7795 5092 7833
rect 5050 7775 5058 7795
rect 5078 7775 5092 7795
rect 5050 7733 5092 7775
rect 5142 7802 5187 7833
rect 5142 7795 5186 7802
rect 5142 7775 5154 7795
rect 5174 7775 5186 7795
rect 5142 7733 5186 7775
rect 11524 7798 11568 7836
rect 11524 7778 11536 7798
rect 11556 7778 11568 7798
rect 8058 7637 8102 7679
rect 8058 7617 8070 7637
rect 8090 7617 8102 7637
rect 8058 7610 8102 7617
rect 8057 7579 8102 7610
rect 8152 7637 8194 7679
rect 8152 7617 8166 7637
rect 8186 7617 8194 7637
rect 8152 7579 8194 7617
rect 8268 7637 8310 7679
rect 8268 7617 8276 7637
rect 8296 7617 8310 7637
rect 8268 7579 8310 7617
rect 8360 7637 8404 7679
rect 8360 7617 8372 7637
rect 8392 7617 8404 7637
rect 8360 7579 8404 7617
rect 8476 7637 8518 7679
rect 8476 7617 8484 7637
rect 8504 7617 8518 7637
rect 8476 7579 8518 7617
rect 8568 7637 8612 7679
rect 8568 7617 8580 7637
rect 8600 7617 8612 7637
rect 8568 7579 8612 7617
rect 8689 7637 8731 7679
rect 8689 7617 8697 7637
rect 8717 7617 8731 7637
rect 8689 7579 8731 7617
rect 8781 7637 8825 7679
rect 11524 7736 11568 7778
rect 11618 7798 11660 7836
rect 11618 7778 11632 7798
rect 11652 7778 11660 7798
rect 11618 7736 11660 7778
rect 11737 7798 11781 7836
rect 11737 7778 11749 7798
rect 11769 7778 11781 7798
rect 11737 7736 11781 7778
rect 11831 7798 11873 7836
rect 11831 7778 11845 7798
rect 11865 7778 11873 7798
rect 11831 7736 11873 7778
rect 11945 7798 11989 7836
rect 11945 7778 11957 7798
rect 11977 7778 11989 7798
rect 11945 7736 11989 7778
rect 12039 7798 12081 7836
rect 12039 7778 12053 7798
rect 12073 7778 12081 7798
rect 12039 7736 12081 7778
rect 12155 7798 12197 7836
rect 12155 7778 12163 7798
rect 12183 7778 12197 7798
rect 12155 7736 12197 7778
rect 12247 7805 12292 7836
rect 12247 7798 12291 7805
rect 12247 7778 12259 7798
rect 12279 7778 12291 7798
rect 12247 7736 12291 7778
rect 15127 7789 15171 7827
rect 15127 7769 15139 7789
rect 15159 7769 15171 7789
rect 8781 7617 8793 7637
rect 8813 7617 8825 7637
rect 8781 7579 8825 7617
rect 9106 7633 9150 7675
rect 9106 7613 9118 7633
rect 9138 7613 9150 7633
rect 9106 7606 9150 7613
rect 9105 7575 9150 7606
rect 9200 7633 9242 7675
rect 9200 7613 9214 7633
rect 9234 7613 9242 7633
rect 9200 7575 9242 7613
rect 9316 7633 9358 7675
rect 9316 7613 9324 7633
rect 9344 7613 9358 7633
rect 9316 7575 9358 7613
rect 9408 7633 9452 7675
rect 9408 7613 9420 7633
rect 9440 7613 9452 7633
rect 9408 7575 9452 7613
rect 9524 7633 9566 7675
rect 9524 7613 9532 7633
rect 9552 7613 9566 7633
rect 9524 7575 9566 7613
rect 9616 7633 9660 7675
rect 9616 7613 9628 7633
rect 9648 7613 9660 7633
rect 9616 7575 9660 7613
rect 9737 7633 9779 7675
rect 9737 7613 9745 7633
rect 9765 7613 9779 7633
rect 9737 7575 9779 7613
rect 9829 7633 9873 7675
rect 9829 7613 9841 7633
rect 9861 7613 9873 7633
rect 15127 7727 15171 7769
rect 15221 7789 15263 7827
rect 15221 7769 15235 7789
rect 15255 7769 15263 7789
rect 15221 7727 15263 7769
rect 15340 7789 15384 7827
rect 15340 7769 15352 7789
rect 15372 7769 15384 7789
rect 15340 7727 15384 7769
rect 15434 7789 15476 7827
rect 15434 7769 15448 7789
rect 15468 7769 15476 7789
rect 15434 7727 15476 7769
rect 15548 7789 15592 7827
rect 15548 7769 15560 7789
rect 15580 7769 15592 7789
rect 15548 7727 15592 7769
rect 15642 7789 15684 7827
rect 15642 7769 15656 7789
rect 15676 7769 15684 7789
rect 15642 7727 15684 7769
rect 15758 7789 15800 7827
rect 15758 7769 15766 7789
rect 15786 7769 15800 7789
rect 15758 7727 15800 7769
rect 15850 7796 15895 7827
rect 15850 7789 15894 7796
rect 15850 7769 15862 7789
rect 15882 7769 15894 7789
rect 15850 7727 15894 7769
rect 9829 7575 9873 7613
rect 18766 7631 18810 7673
rect 18766 7611 18778 7631
rect 18798 7611 18810 7631
rect 18766 7604 18810 7611
rect 18765 7573 18810 7604
rect 18860 7631 18902 7673
rect 18860 7611 18874 7631
rect 18894 7611 18902 7631
rect 18860 7573 18902 7611
rect 18976 7631 19018 7673
rect 18976 7611 18984 7631
rect 19004 7611 19018 7631
rect 18976 7573 19018 7611
rect 19068 7631 19112 7673
rect 19068 7611 19080 7631
rect 19100 7611 19112 7631
rect 19068 7573 19112 7611
rect 19184 7631 19226 7673
rect 19184 7611 19192 7631
rect 19212 7611 19226 7631
rect 19184 7573 19226 7611
rect 19276 7631 19320 7673
rect 19276 7611 19288 7631
rect 19308 7611 19320 7631
rect 19276 7573 19320 7611
rect 19397 7631 19439 7673
rect 19397 7611 19405 7631
rect 19425 7611 19439 7631
rect 19397 7573 19439 7611
rect 19489 7631 19533 7673
rect 19489 7611 19501 7631
rect 19521 7611 19533 7631
rect 19489 7573 19533 7611
rect 19814 7627 19858 7669
rect 19814 7607 19826 7627
rect 19846 7607 19858 7627
rect 19814 7600 19858 7607
rect 19813 7569 19858 7600
rect 19908 7627 19950 7669
rect 19908 7607 19922 7627
rect 19942 7607 19950 7627
rect 19908 7569 19950 7607
rect 20024 7627 20066 7669
rect 20024 7607 20032 7627
rect 20052 7607 20066 7627
rect 20024 7569 20066 7607
rect 20116 7627 20160 7669
rect 20116 7607 20128 7627
rect 20148 7607 20160 7627
rect 20116 7569 20160 7607
rect 20232 7627 20274 7669
rect 20232 7607 20240 7627
rect 20260 7607 20274 7627
rect 20232 7569 20274 7607
rect 20324 7627 20368 7669
rect 20324 7607 20336 7627
rect 20356 7607 20368 7627
rect 20324 7569 20368 7607
rect 20445 7627 20487 7669
rect 20445 7607 20453 7627
rect 20473 7607 20487 7627
rect 20445 7569 20487 7607
rect 20537 7627 20581 7669
rect 20537 7607 20549 7627
rect 20569 7607 20581 7627
rect 20537 7569 20581 7607
rect 813 6889 857 6927
rect 813 6869 825 6889
rect 845 6869 857 6889
rect 813 6827 857 6869
rect 907 6889 949 6927
rect 907 6869 921 6889
rect 941 6869 949 6889
rect 907 6827 949 6869
rect 1026 6889 1070 6927
rect 1026 6869 1038 6889
rect 1058 6869 1070 6889
rect 1026 6827 1070 6869
rect 1120 6889 1162 6927
rect 1120 6869 1134 6889
rect 1154 6869 1162 6889
rect 1120 6827 1162 6869
rect 1234 6889 1278 6927
rect 1234 6869 1246 6889
rect 1266 6869 1278 6889
rect 1234 6827 1278 6869
rect 1328 6889 1370 6927
rect 1328 6869 1342 6889
rect 1362 6869 1370 6889
rect 1328 6827 1370 6869
rect 1444 6889 1486 6927
rect 1444 6869 1452 6889
rect 1472 6869 1486 6889
rect 1444 6827 1486 6869
rect 1536 6896 1581 6927
rect 1536 6889 1580 6896
rect 1536 6869 1548 6889
rect 1568 6869 1580 6889
rect 1536 6827 1580 6869
rect 1861 6885 1905 6923
rect 1861 6865 1873 6885
rect 1893 6865 1905 6885
rect 1861 6823 1905 6865
rect 1955 6885 1997 6923
rect 1955 6865 1969 6885
rect 1989 6865 1997 6885
rect 1955 6823 1997 6865
rect 2074 6885 2118 6923
rect 2074 6865 2086 6885
rect 2106 6865 2118 6885
rect 2074 6823 2118 6865
rect 2168 6885 2210 6923
rect 2168 6865 2182 6885
rect 2202 6865 2210 6885
rect 2168 6823 2210 6865
rect 2282 6885 2326 6923
rect 2282 6865 2294 6885
rect 2314 6865 2326 6885
rect 2282 6823 2326 6865
rect 2376 6885 2418 6923
rect 2376 6865 2390 6885
rect 2410 6865 2418 6885
rect 2376 6823 2418 6865
rect 2492 6885 2534 6923
rect 2492 6865 2500 6885
rect 2520 6865 2534 6885
rect 2492 6823 2534 6865
rect 2584 6892 2629 6923
rect 2584 6885 2628 6892
rect 2584 6865 2596 6885
rect 2616 6865 2628 6885
rect 2584 6823 2628 6865
rect 11521 6883 11565 6921
rect 5500 6727 5544 6769
rect 5500 6707 5512 6727
rect 5532 6707 5544 6727
rect 5500 6700 5544 6707
rect 5499 6669 5544 6700
rect 5594 6727 5636 6769
rect 5594 6707 5608 6727
rect 5628 6707 5636 6727
rect 5594 6669 5636 6707
rect 5710 6727 5752 6769
rect 5710 6707 5718 6727
rect 5738 6707 5752 6727
rect 5710 6669 5752 6707
rect 5802 6727 5846 6769
rect 5802 6707 5814 6727
rect 5834 6707 5846 6727
rect 5802 6669 5846 6707
rect 5918 6727 5960 6769
rect 5918 6707 5926 6727
rect 5946 6707 5960 6727
rect 5918 6669 5960 6707
rect 6010 6727 6054 6769
rect 6010 6707 6022 6727
rect 6042 6707 6054 6727
rect 6010 6669 6054 6707
rect 6131 6727 6173 6769
rect 6131 6707 6139 6727
rect 6159 6707 6173 6727
rect 6131 6669 6173 6707
rect 6223 6727 6267 6769
rect 11521 6863 11533 6883
rect 11553 6863 11565 6883
rect 11521 6821 11565 6863
rect 11615 6883 11657 6921
rect 11615 6863 11629 6883
rect 11649 6863 11657 6883
rect 11615 6821 11657 6863
rect 11734 6883 11778 6921
rect 11734 6863 11746 6883
rect 11766 6863 11778 6883
rect 11734 6821 11778 6863
rect 11828 6883 11870 6921
rect 11828 6863 11842 6883
rect 11862 6863 11870 6883
rect 11828 6821 11870 6863
rect 11942 6883 11986 6921
rect 11942 6863 11954 6883
rect 11974 6863 11986 6883
rect 11942 6821 11986 6863
rect 12036 6883 12078 6921
rect 12036 6863 12050 6883
rect 12070 6863 12078 6883
rect 12036 6821 12078 6863
rect 12152 6883 12194 6921
rect 12152 6863 12160 6883
rect 12180 6863 12194 6883
rect 12152 6821 12194 6863
rect 12244 6890 12289 6921
rect 12244 6883 12288 6890
rect 12244 6863 12256 6883
rect 12276 6863 12288 6883
rect 12244 6821 12288 6863
rect 12569 6879 12613 6917
rect 12569 6859 12581 6879
rect 12601 6859 12613 6879
rect 6223 6707 6235 6727
rect 6255 6707 6267 6727
rect 6223 6669 6267 6707
rect 9103 6718 9147 6760
rect 9103 6698 9115 6718
rect 9135 6698 9147 6718
rect 9103 6691 9147 6698
rect 9102 6660 9147 6691
rect 9197 6718 9239 6760
rect 9197 6698 9211 6718
rect 9231 6698 9239 6718
rect 9197 6660 9239 6698
rect 9313 6718 9355 6760
rect 9313 6698 9321 6718
rect 9341 6698 9355 6718
rect 9313 6660 9355 6698
rect 9405 6718 9449 6760
rect 9405 6698 9417 6718
rect 9437 6698 9449 6718
rect 9405 6660 9449 6698
rect 9521 6718 9563 6760
rect 9521 6698 9529 6718
rect 9549 6698 9563 6718
rect 9521 6660 9563 6698
rect 9613 6718 9657 6760
rect 9613 6698 9625 6718
rect 9645 6698 9657 6718
rect 9613 6660 9657 6698
rect 9734 6718 9776 6760
rect 9734 6698 9742 6718
rect 9762 6698 9776 6718
rect 9734 6660 9776 6698
rect 9826 6718 9870 6760
rect 12569 6817 12613 6859
rect 12663 6879 12705 6917
rect 12663 6859 12677 6879
rect 12697 6859 12705 6879
rect 12663 6817 12705 6859
rect 12782 6879 12826 6917
rect 12782 6859 12794 6879
rect 12814 6859 12826 6879
rect 12782 6817 12826 6859
rect 12876 6879 12918 6917
rect 12876 6859 12890 6879
rect 12910 6859 12918 6879
rect 12876 6817 12918 6859
rect 12990 6879 13034 6917
rect 12990 6859 13002 6879
rect 13022 6859 13034 6879
rect 12990 6817 13034 6859
rect 13084 6879 13126 6917
rect 13084 6859 13098 6879
rect 13118 6859 13126 6879
rect 13084 6817 13126 6859
rect 13200 6879 13242 6917
rect 13200 6859 13208 6879
rect 13228 6859 13242 6879
rect 13200 6817 13242 6859
rect 13292 6886 13337 6917
rect 13292 6879 13336 6886
rect 13292 6859 13304 6879
rect 13324 6859 13336 6879
rect 13292 6817 13336 6859
rect 9826 6698 9838 6718
rect 9858 6698 9870 6718
rect 9826 6660 9870 6698
rect 16208 6721 16252 6763
rect 16208 6701 16220 6721
rect 16240 6701 16252 6721
rect 16208 6694 16252 6701
rect 16207 6663 16252 6694
rect 16302 6721 16344 6763
rect 16302 6701 16316 6721
rect 16336 6701 16344 6721
rect 16302 6663 16344 6701
rect 16418 6721 16460 6763
rect 16418 6701 16426 6721
rect 16446 6701 16460 6721
rect 16418 6663 16460 6701
rect 16510 6721 16554 6763
rect 16510 6701 16522 6721
rect 16542 6701 16554 6721
rect 16510 6663 16554 6701
rect 16626 6721 16668 6763
rect 16626 6701 16634 6721
rect 16654 6701 16668 6721
rect 16626 6663 16668 6701
rect 16718 6721 16762 6763
rect 16718 6701 16730 6721
rect 16750 6701 16762 6721
rect 16718 6663 16762 6701
rect 16839 6721 16881 6763
rect 16839 6701 16847 6721
rect 16867 6701 16881 6721
rect 16839 6663 16881 6701
rect 16931 6721 16975 6763
rect 16931 6701 16943 6721
rect 16963 6701 16975 6721
rect 16931 6663 16975 6701
rect 19811 6712 19855 6754
rect 19811 6692 19823 6712
rect 19843 6692 19855 6712
rect 19811 6685 19855 6692
rect 19810 6654 19855 6685
rect 19905 6712 19947 6754
rect 19905 6692 19919 6712
rect 19939 6692 19947 6712
rect 19905 6654 19947 6692
rect 20021 6712 20063 6754
rect 20021 6692 20029 6712
rect 20049 6692 20063 6712
rect 20021 6654 20063 6692
rect 20113 6712 20157 6754
rect 20113 6692 20125 6712
rect 20145 6692 20157 6712
rect 20113 6654 20157 6692
rect 20229 6712 20271 6754
rect 20229 6692 20237 6712
rect 20257 6692 20271 6712
rect 20229 6654 20271 6692
rect 20321 6712 20365 6754
rect 20321 6692 20333 6712
rect 20353 6692 20365 6712
rect 20321 6654 20365 6692
rect 20442 6712 20484 6754
rect 20442 6692 20450 6712
rect 20470 6692 20484 6712
rect 20442 6654 20484 6692
rect 20534 6712 20578 6754
rect 20534 6692 20546 6712
rect 20566 6692 20578 6712
rect 20534 6654 20578 6692
rect 813 6210 857 6248
rect 813 6190 825 6210
rect 845 6190 857 6210
rect 813 6148 857 6190
rect 907 6210 949 6248
rect 907 6190 921 6210
rect 941 6190 949 6210
rect 907 6148 949 6190
rect 1026 6210 1070 6248
rect 1026 6190 1038 6210
rect 1058 6190 1070 6210
rect 1026 6148 1070 6190
rect 1120 6210 1162 6248
rect 1120 6190 1134 6210
rect 1154 6190 1162 6210
rect 1120 6148 1162 6190
rect 1234 6210 1278 6248
rect 1234 6190 1246 6210
rect 1266 6190 1278 6210
rect 1234 6148 1278 6190
rect 1328 6210 1370 6248
rect 1328 6190 1342 6210
rect 1362 6190 1370 6210
rect 1328 6148 1370 6190
rect 1444 6210 1486 6248
rect 1444 6190 1452 6210
rect 1472 6190 1486 6210
rect 1444 6148 1486 6190
rect 1536 6217 1581 6248
rect 1536 6210 1580 6217
rect 1536 6190 1548 6210
rect 1568 6190 1580 6210
rect 1536 6148 1580 6190
rect 3308 6205 3352 6243
rect 3308 6185 3320 6205
rect 3340 6185 3352 6205
rect 3308 6143 3352 6185
rect 3402 6205 3444 6243
rect 3402 6185 3416 6205
rect 3436 6185 3444 6205
rect 3402 6143 3444 6185
rect 3521 6205 3565 6243
rect 3521 6185 3533 6205
rect 3553 6185 3565 6205
rect 3521 6143 3565 6185
rect 3615 6205 3657 6243
rect 3615 6185 3629 6205
rect 3649 6185 3657 6205
rect 3615 6143 3657 6185
rect 3729 6205 3773 6243
rect 3729 6185 3741 6205
rect 3761 6185 3773 6205
rect 3729 6143 3773 6185
rect 3823 6205 3865 6243
rect 3823 6185 3837 6205
rect 3857 6185 3865 6205
rect 3823 6143 3865 6185
rect 3939 6205 3981 6243
rect 3939 6185 3947 6205
rect 3967 6185 3981 6205
rect 3939 6143 3981 6185
rect 4031 6212 4076 6243
rect 4031 6205 4075 6212
rect 4031 6185 4043 6205
rect 4063 6185 4075 6205
rect 4031 6143 4075 6185
rect 11521 6204 11565 6242
rect 11521 6184 11533 6204
rect 11553 6184 11565 6204
rect 8055 6043 8099 6085
rect 8055 6023 8067 6043
rect 8087 6023 8099 6043
rect 8055 6016 8099 6023
rect 8054 5985 8099 6016
rect 8149 6043 8191 6085
rect 8149 6023 8163 6043
rect 8183 6023 8191 6043
rect 8149 5985 8191 6023
rect 8265 6043 8307 6085
rect 8265 6023 8273 6043
rect 8293 6023 8307 6043
rect 8265 5985 8307 6023
rect 8357 6043 8401 6085
rect 8357 6023 8369 6043
rect 8389 6023 8401 6043
rect 8357 5985 8401 6023
rect 8473 6043 8515 6085
rect 8473 6023 8481 6043
rect 8501 6023 8515 6043
rect 8473 5985 8515 6023
rect 8565 6043 8609 6085
rect 8565 6023 8577 6043
rect 8597 6023 8609 6043
rect 8565 5985 8609 6023
rect 8686 6043 8728 6085
rect 8686 6023 8694 6043
rect 8714 6023 8728 6043
rect 8686 5985 8728 6023
rect 8778 6043 8822 6085
rect 11521 6142 11565 6184
rect 11615 6204 11657 6242
rect 11615 6184 11629 6204
rect 11649 6184 11657 6204
rect 11615 6142 11657 6184
rect 11734 6204 11778 6242
rect 11734 6184 11746 6204
rect 11766 6184 11778 6204
rect 11734 6142 11778 6184
rect 11828 6204 11870 6242
rect 11828 6184 11842 6204
rect 11862 6184 11870 6204
rect 11828 6142 11870 6184
rect 11942 6204 11986 6242
rect 11942 6184 11954 6204
rect 11974 6184 11986 6204
rect 11942 6142 11986 6184
rect 12036 6204 12078 6242
rect 12036 6184 12050 6204
rect 12070 6184 12078 6204
rect 12036 6142 12078 6184
rect 12152 6204 12194 6242
rect 12152 6184 12160 6204
rect 12180 6184 12194 6204
rect 12152 6142 12194 6184
rect 12244 6211 12289 6242
rect 12244 6204 12288 6211
rect 12244 6184 12256 6204
rect 12276 6184 12288 6204
rect 12244 6142 12288 6184
rect 14016 6199 14060 6237
rect 14016 6179 14028 6199
rect 14048 6179 14060 6199
rect 8778 6023 8790 6043
rect 8810 6023 8822 6043
rect 8778 5985 8822 6023
rect 9103 6039 9147 6081
rect 9103 6019 9115 6039
rect 9135 6019 9147 6039
rect 9103 6012 9147 6019
rect 9102 5981 9147 6012
rect 9197 6039 9239 6081
rect 9197 6019 9211 6039
rect 9231 6019 9239 6039
rect 9197 5981 9239 6019
rect 9313 6039 9355 6081
rect 9313 6019 9321 6039
rect 9341 6019 9355 6039
rect 9313 5981 9355 6019
rect 9405 6039 9449 6081
rect 9405 6019 9417 6039
rect 9437 6019 9449 6039
rect 9405 5981 9449 6019
rect 9521 6039 9563 6081
rect 9521 6019 9529 6039
rect 9549 6019 9563 6039
rect 9521 5981 9563 6019
rect 9613 6039 9657 6081
rect 9613 6019 9625 6039
rect 9645 6019 9657 6039
rect 9613 5981 9657 6019
rect 9734 6039 9776 6081
rect 9734 6019 9742 6039
rect 9762 6019 9776 6039
rect 9734 5981 9776 6019
rect 9826 6039 9870 6081
rect 9826 6019 9838 6039
rect 9858 6019 9870 6039
rect 14016 6137 14060 6179
rect 14110 6199 14152 6237
rect 14110 6179 14124 6199
rect 14144 6179 14152 6199
rect 14110 6137 14152 6179
rect 14229 6199 14273 6237
rect 14229 6179 14241 6199
rect 14261 6179 14273 6199
rect 14229 6137 14273 6179
rect 14323 6199 14365 6237
rect 14323 6179 14337 6199
rect 14357 6179 14365 6199
rect 14323 6137 14365 6179
rect 14437 6199 14481 6237
rect 14437 6179 14449 6199
rect 14469 6179 14481 6199
rect 14437 6137 14481 6179
rect 14531 6199 14573 6237
rect 14531 6179 14545 6199
rect 14565 6179 14573 6199
rect 14531 6137 14573 6179
rect 14647 6199 14689 6237
rect 14647 6179 14655 6199
rect 14675 6179 14689 6199
rect 14647 6137 14689 6179
rect 14739 6206 14784 6237
rect 14739 6199 14783 6206
rect 14739 6179 14751 6199
rect 14771 6179 14783 6199
rect 14739 6137 14783 6179
rect 9826 5981 9870 6019
rect 18763 6037 18807 6079
rect 18763 6017 18775 6037
rect 18795 6017 18807 6037
rect 18763 6010 18807 6017
rect 18762 5979 18807 6010
rect 18857 6037 18899 6079
rect 18857 6017 18871 6037
rect 18891 6017 18899 6037
rect 18857 5979 18899 6017
rect 18973 6037 19015 6079
rect 18973 6017 18981 6037
rect 19001 6017 19015 6037
rect 18973 5979 19015 6017
rect 19065 6037 19109 6079
rect 19065 6017 19077 6037
rect 19097 6017 19109 6037
rect 19065 5979 19109 6017
rect 19181 6037 19223 6079
rect 19181 6017 19189 6037
rect 19209 6017 19223 6037
rect 19181 5979 19223 6017
rect 19273 6037 19317 6079
rect 19273 6017 19285 6037
rect 19305 6017 19317 6037
rect 19273 5979 19317 6017
rect 19394 6037 19436 6079
rect 19394 6017 19402 6037
rect 19422 6017 19436 6037
rect 19394 5979 19436 6017
rect 19486 6037 19530 6079
rect 19486 6017 19498 6037
rect 19518 6017 19530 6037
rect 19486 5979 19530 6017
rect 19811 6033 19855 6075
rect 19811 6013 19823 6033
rect 19843 6013 19855 6033
rect 19811 6006 19855 6013
rect 19810 5975 19855 6006
rect 19905 6033 19947 6075
rect 19905 6013 19919 6033
rect 19939 6013 19947 6033
rect 19905 5975 19947 6013
rect 20021 6033 20063 6075
rect 20021 6013 20029 6033
rect 20049 6013 20063 6033
rect 20021 5975 20063 6013
rect 20113 6033 20157 6075
rect 20113 6013 20125 6033
rect 20145 6013 20157 6033
rect 20113 5975 20157 6013
rect 20229 6033 20271 6075
rect 20229 6013 20237 6033
rect 20257 6013 20271 6033
rect 20229 5975 20271 6013
rect 20321 6033 20365 6075
rect 20321 6013 20333 6033
rect 20353 6013 20365 6033
rect 20321 5975 20365 6013
rect 20442 6033 20484 6075
rect 20442 6013 20450 6033
rect 20470 6013 20484 6033
rect 20442 5975 20484 6013
rect 20534 6033 20578 6075
rect 20534 6013 20546 6033
rect 20566 6013 20578 6033
rect 20534 5975 20578 6013
rect 813 5442 857 5480
rect 813 5422 825 5442
rect 845 5422 857 5442
rect 813 5380 857 5422
rect 907 5442 949 5480
rect 907 5422 921 5442
rect 941 5422 949 5442
rect 907 5380 949 5422
rect 1026 5442 1070 5480
rect 1026 5422 1038 5442
rect 1058 5422 1070 5442
rect 1026 5380 1070 5422
rect 1120 5442 1162 5480
rect 1120 5422 1134 5442
rect 1154 5422 1162 5442
rect 1120 5380 1162 5422
rect 1234 5442 1278 5480
rect 1234 5422 1246 5442
rect 1266 5422 1278 5442
rect 1234 5380 1278 5422
rect 1328 5442 1370 5480
rect 1328 5422 1342 5442
rect 1362 5422 1370 5442
rect 1328 5380 1370 5422
rect 1444 5442 1486 5480
rect 1444 5422 1452 5442
rect 1472 5422 1486 5442
rect 1444 5380 1486 5422
rect 1536 5449 1581 5480
rect 1536 5442 1580 5449
rect 1536 5422 1548 5442
rect 1568 5422 1580 5442
rect 1536 5380 1580 5422
rect 1861 5438 1905 5476
rect 1861 5418 1873 5438
rect 1893 5418 1905 5438
rect 1861 5376 1905 5418
rect 1955 5438 1997 5476
rect 1955 5418 1969 5438
rect 1989 5418 1997 5438
rect 1955 5376 1997 5418
rect 2074 5438 2118 5476
rect 2074 5418 2086 5438
rect 2106 5418 2118 5438
rect 2074 5376 2118 5418
rect 2168 5438 2210 5476
rect 2168 5418 2182 5438
rect 2202 5418 2210 5438
rect 2168 5376 2210 5418
rect 2282 5438 2326 5476
rect 2282 5418 2294 5438
rect 2314 5418 2326 5438
rect 2282 5376 2326 5418
rect 2376 5438 2418 5476
rect 2376 5418 2390 5438
rect 2410 5418 2418 5438
rect 2376 5376 2418 5418
rect 2492 5438 2534 5476
rect 2492 5418 2500 5438
rect 2520 5418 2534 5438
rect 2492 5376 2534 5418
rect 2584 5445 2629 5476
rect 2584 5438 2628 5445
rect 2584 5418 2596 5438
rect 2616 5418 2628 5438
rect 2584 5376 2628 5418
rect 11521 5436 11565 5474
rect 6608 5276 6652 5318
rect 6608 5256 6620 5276
rect 6640 5256 6652 5276
rect 6608 5249 6652 5256
rect 6607 5218 6652 5249
rect 6702 5276 6744 5318
rect 6702 5256 6716 5276
rect 6736 5256 6744 5276
rect 6702 5218 6744 5256
rect 6818 5276 6860 5318
rect 6818 5256 6826 5276
rect 6846 5256 6860 5276
rect 6818 5218 6860 5256
rect 6910 5276 6954 5318
rect 6910 5256 6922 5276
rect 6942 5256 6954 5276
rect 6910 5218 6954 5256
rect 7026 5276 7068 5318
rect 7026 5256 7034 5276
rect 7054 5256 7068 5276
rect 7026 5218 7068 5256
rect 7118 5276 7162 5318
rect 7118 5256 7130 5276
rect 7150 5256 7162 5276
rect 7118 5218 7162 5256
rect 7239 5276 7281 5318
rect 7239 5256 7247 5276
rect 7267 5256 7281 5276
rect 7239 5218 7281 5256
rect 7331 5276 7375 5318
rect 11521 5416 11533 5436
rect 11553 5416 11565 5436
rect 11521 5374 11565 5416
rect 11615 5436 11657 5474
rect 11615 5416 11629 5436
rect 11649 5416 11657 5436
rect 11615 5374 11657 5416
rect 11734 5436 11778 5474
rect 11734 5416 11746 5436
rect 11766 5416 11778 5436
rect 11734 5374 11778 5416
rect 11828 5436 11870 5474
rect 11828 5416 11842 5436
rect 11862 5416 11870 5436
rect 11828 5374 11870 5416
rect 11942 5436 11986 5474
rect 11942 5416 11954 5436
rect 11974 5416 11986 5436
rect 11942 5374 11986 5416
rect 12036 5436 12078 5474
rect 12036 5416 12050 5436
rect 12070 5416 12078 5436
rect 12036 5374 12078 5416
rect 12152 5436 12194 5474
rect 12152 5416 12160 5436
rect 12180 5416 12194 5436
rect 12152 5374 12194 5416
rect 12244 5443 12289 5474
rect 12244 5436 12288 5443
rect 12244 5416 12256 5436
rect 12276 5416 12288 5436
rect 12244 5374 12288 5416
rect 12569 5432 12613 5470
rect 12569 5412 12581 5432
rect 12601 5412 12613 5432
rect 7331 5256 7343 5276
rect 7363 5256 7375 5276
rect 7331 5218 7375 5256
rect 9103 5271 9147 5313
rect 9103 5251 9115 5271
rect 9135 5251 9147 5271
rect 9103 5244 9147 5251
rect 9102 5213 9147 5244
rect 9197 5271 9239 5313
rect 9197 5251 9211 5271
rect 9231 5251 9239 5271
rect 9197 5213 9239 5251
rect 9313 5271 9355 5313
rect 9313 5251 9321 5271
rect 9341 5251 9355 5271
rect 9313 5213 9355 5251
rect 9405 5271 9449 5313
rect 9405 5251 9417 5271
rect 9437 5251 9449 5271
rect 9405 5213 9449 5251
rect 9521 5271 9563 5313
rect 9521 5251 9529 5271
rect 9549 5251 9563 5271
rect 9521 5213 9563 5251
rect 9613 5271 9657 5313
rect 9613 5251 9625 5271
rect 9645 5251 9657 5271
rect 9613 5213 9657 5251
rect 9734 5271 9776 5313
rect 9734 5251 9742 5271
rect 9762 5251 9776 5271
rect 9734 5213 9776 5251
rect 9826 5271 9870 5313
rect 12569 5370 12613 5412
rect 12663 5432 12705 5470
rect 12663 5412 12677 5432
rect 12697 5412 12705 5432
rect 12663 5370 12705 5412
rect 12782 5432 12826 5470
rect 12782 5412 12794 5432
rect 12814 5412 12826 5432
rect 12782 5370 12826 5412
rect 12876 5432 12918 5470
rect 12876 5412 12890 5432
rect 12910 5412 12918 5432
rect 12876 5370 12918 5412
rect 12990 5432 13034 5470
rect 12990 5412 13002 5432
rect 13022 5412 13034 5432
rect 12990 5370 13034 5412
rect 13084 5432 13126 5470
rect 13084 5412 13098 5432
rect 13118 5412 13126 5432
rect 13084 5370 13126 5412
rect 13200 5432 13242 5470
rect 13200 5412 13208 5432
rect 13228 5412 13242 5432
rect 13200 5370 13242 5412
rect 13292 5439 13337 5470
rect 13292 5432 13336 5439
rect 13292 5412 13304 5432
rect 13324 5412 13336 5432
rect 13292 5370 13336 5412
rect 9826 5251 9838 5271
rect 9858 5251 9870 5271
rect 9826 5213 9870 5251
rect 17316 5270 17360 5312
rect 17316 5250 17328 5270
rect 17348 5250 17360 5270
rect 17316 5243 17360 5250
rect 17315 5212 17360 5243
rect 17410 5270 17452 5312
rect 17410 5250 17424 5270
rect 17444 5250 17452 5270
rect 17410 5212 17452 5250
rect 17526 5270 17568 5312
rect 17526 5250 17534 5270
rect 17554 5250 17568 5270
rect 17526 5212 17568 5250
rect 17618 5270 17662 5312
rect 17618 5250 17630 5270
rect 17650 5250 17662 5270
rect 17618 5212 17662 5250
rect 17734 5270 17776 5312
rect 17734 5250 17742 5270
rect 17762 5250 17776 5270
rect 17734 5212 17776 5250
rect 17826 5270 17870 5312
rect 17826 5250 17838 5270
rect 17858 5250 17870 5270
rect 17826 5212 17870 5250
rect 17947 5270 17989 5312
rect 17947 5250 17955 5270
rect 17975 5250 17989 5270
rect 17947 5212 17989 5250
rect 18039 5270 18083 5312
rect 18039 5250 18051 5270
rect 18071 5250 18083 5270
rect 18039 5212 18083 5250
rect 19811 5265 19855 5307
rect 19811 5245 19823 5265
rect 19843 5245 19855 5265
rect 19811 5238 19855 5245
rect 19810 5207 19855 5238
rect 19905 5265 19947 5307
rect 19905 5245 19919 5265
rect 19939 5245 19947 5265
rect 19905 5207 19947 5245
rect 20021 5265 20063 5307
rect 20021 5245 20029 5265
rect 20049 5245 20063 5265
rect 20021 5207 20063 5245
rect 20113 5265 20157 5307
rect 20113 5245 20125 5265
rect 20145 5245 20157 5265
rect 20113 5207 20157 5245
rect 20229 5265 20271 5307
rect 20229 5245 20237 5265
rect 20257 5245 20271 5265
rect 20229 5207 20271 5245
rect 20321 5265 20365 5307
rect 20321 5245 20333 5265
rect 20353 5245 20365 5265
rect 20321 5207 20365 5245
rect 20442 5265 20484 5307
rect 20442 5245 20450 5265
rect 20470 5245 20484 5265
rect 20442 5207 20484 5245
rect 20534 5265 20578 5307
rect 20534 5245 20546 5265
rect 20566 5245 20578 5265
rect 20534 5207 20578 5245
rect 813 4763 857 4801
rect 813 4743 825 4763
rect 845 4743 857 4763
rect 813 4701 857 4743
rect 907 4763 949 4801
rect 907 4743 921 4763
rect 941 4743 949 4763
rect 907 4701 949 4743
rect 1026 4763 1070 4801
rect 1026 4743 1038 4763
rect 1058 4743 1070 4763
rect 1026 4701 1070 4743
rect 1120 4763 1162 4801
rect 1120 4743 1134 4763
rect 1154 4743 1162 4763
rect 1120 4701 1162 4743
rect 1234 4763 1278 4801
rect 1234 4743 1246 4763
rect 1266 4743 1278 4763
rect 1234 4701 1278 4743
rect 1328 4763 1370 4801
rect 1328 4743 1342 4763
rect 1362 4743 1370 4763
rect 1328 4701 1370 4743
rect 1444 4763 1486 4801
rect 1444 4743 1452 4763
rect 1472 4743 1486 4763
rect 1444 4701 1486 4743
rect 1536 4770 1581 4801
rect 1536 4763 1580 4770
rect 1536 4743 1548 4763
rect 1568 4743 1580 4763
rect 1536 4701 1580 4743
rect 3351 4760 3395 4798
rect 3351 4740 3363 4760
rect 3383 4740 3395 4760
rect 3351 4698 3395 4740
rect 3445 4760 3487 4798
rect 3445 4740 3459 4760
rect 3479 4740 3487 4760
rect 3445 4698 3487 4740
rect 3564 4760 3608 4798
rect 3564 4740 3576 4760
rect 3596 4740 3608 4760
rect 3564 4698 3608 4740
rect 3658 4760 3700 4798
rect 3658 4740 3672 4760
rect 3692 4740 3700 4760
rect 3658 4698 3700 4740
rect 3772 4760 3816 4798
rect 3772 4740 3784 4760
rect 3804 4740 3816 4760
rect 3772 4698 3816 4740
rect 3866 4760 3908 4798
rect 3866 4740 3880 4760
rect 3900 4740 3908 4760
rect 3866 4698 3908 4740
rect 3982 4760 4024 4798
rect 3982 4740 3990 4760
rect 4010 4740 4024 4760
rect 3982 4698 4024 4740
rect 4074 4767 4119 4798
rect 4074 4760 4118 4767
rect 4074 4740 4086 4760
rect 4106 4740 4118 4760
rect 4074 4698 4118 4740
rect 11521 4757 11565 4795
rect 11521 4737 11533 4757
rect 11553 4737 11565 4757
rect 8055 4596 8099 4638
rect 8055 4576 8067 4596
rect 8087 4576 8099 4596
rect 8055 4569 8099 4576
rect 8054 4538 8099 4569
rect 8149 4596 8191 4638
rect 8149 4576 8163 4596
rect 8183 4576 8191 4596
rect 8149 4538 8191 4576
rect 8265 4596 8307 4638
rect 8265 4576 8273 4596
rect 8293 4576 8307 4596
rect 8265 4538 8307 4576
rect 8357 4596 8401 4638
rect 8357 4576 8369 4596
rect 8389 4576 8401 4596
rect 8357 4538 8401 4576
rect 8473 4596 8515 4638
rect 8473 4576 8481 4596
rect 8501 4576 8515 4596
rect 8473 4538 8515 4576
rect 8565 4596 8609 4638
rect 8565 4576 8577 4596
rect 8597 4576 8609 4596
rect 8565 4538 8609 4576
rect 8686 4596 8728 4638
rect 8686 4576 8694 4596
rect 8714 4576 8728 4596
rect 8686 4538 8728 4576
rect 8778 4596 8822 4638
rect 11521 4695 11565 4737
rect 11615 4757 11657 4795
rect 11615 4737 11629 4757
rect 11649 4737 11657 4757
rect 11615 4695 11657 4737
rect 11734 4757 11778 4795
rect 11734 4737 11746 4757
rect 11766 4737 11778 4757
rect 11734 4695 11778 4737
rect 11828 4757 11870 4795
rect 11828 4737 11842 4757
rect 11862 4737 11870 4757
rect 11828 4695 11870 4737
rect 11942 4757 11986 4795
rect 11942 4737 11954 4757
rect 11974 4737 11986 4757
rect 11942 4695 11986 4737
rect 12036 4757 12078 4795
rect 12036 4737 12050 4757
rect 12070 4737 12078 4757
rect 12036 4695 12078 4737
rect 12152 4757 12194 4795
rect 12152 4737 12160 4757
rect 12180 4737 12194 4757
rect 12152 4695 12194 4737
rect 12244 4764 12289 4795
rect 12244 4757 12288 4764
rect 12244 4737 12256 4757
rect 12276 4737 12288 4757
rect 12244 4695 12288 4737
rect 14059 4754 14103 4792
rect 14059 4734 14071 4754
rect 14091 4734 14103 4754
rect 8778 4576 8790 4596
rect 8810 4576 8822 4596
rect 8778 4538 8822 4576
rect 9103 4592 9147 4634
rect 9103 4572 9115 4592
rect 9135 4572 9147 4592
rect 9103 4565 9147 4572
rect 9102 4534 9147 4565
rect 9197 4592 9239 4634
rect 9197 4572 9211 4592
rect 9231 4572 9239 4592
rect 9197 4534 9239 4572
rect 9313 4592 9355 4634
rect 9313 4572 9321 4592
rect 9341 4572 9355 4592
rect 9313 4534 9355 4572
rect 9405 4592 9449 4634
rect 9405 4572 9417 4592
rect 9437 4572 9449 4592
rect 9405 4534 9449 4572
rect 9521 4592 9563 4634
rect 9521 4572 9529 4592
rect 9549 4572 9563 4592
rect 9521 4534 9563 4572
rect 9613 4592 9657 4634
rect 9613 4572 9625 4592
rect 9645 4572 9657 4592
rect 9613 4534 9657 4572
rect 9734 4592 9776 4634
rect 9734 4572 9742 4592
rect 9762 4572 9776 4592
rect 9734 4534 9776 4572
rect 9826 4592 9870 4634
rect 9826 4572 9838 4592
rect 9858 4572 9870 4592
rect 14059 4692 14103 4734
rect 14153 4754 14195 4792
rect 14153 4734 14167 4754
rect 14187 4734 14195 4754
rect 14153 4692 14195 4734
rect 14272 4754 14316 4792
rect 14272 4734 14284 4754
rect 14304 4734 14316 4754
rect 14272 4692 14316 4734
rect 14366 4754 14408 4792
rect 14366 4734 14380 4754
rect 14400 4734 14408 4754
rect 14366 4692 14408 4734
rect 14480 4754 14524 4792
rect 14480 4734 14492 4754
rect 14512 4734 14524 4754
rect 14480 4692 14524 4734
rect 14574 4754 14616 4792
rect 14574 4734 14588 4754
rect 14608 4734 14616 4754
rect 14574 4692 14616 4734
rect 14690 4754 14732 4792
rect 14690 4734 14698 4754
rect 14718 4734 14732 4754
rect 14690 4692 14732 4734
rect 14782 4761 14827 4792
rect 14782 4754 14826 4761
rect 14782 4734 14794 4754
rect 14814 4734 14826 4754
rect 14782 4692 14826 4734
rect 9826 4534 9870 4572
rect 18763 4590 18807 4632
rect 18763 4570 18775 4590
rect 18795 4570 18807 4590
rect 18763 4563 18807 4570
rect 18762 4532 18807 4563
rect 18857 4590 18899 4632
rect 18857 4570 18871 4590
rect 18891 4570 18899 4590
rect 18857 4532 18899 4570
rect 18973 4590 19015 4632
rect 18973 4570 18981 4590
rect 19001 4570 19015 4590
rect 18973 4532 19015 4570
rect 19065 4590 19109 4632
rect 19065 4570 19077 4590
rect 19097 4570 19109 4590
rect 19065 4532 19109 4570
rect 19181 4590 19223 4632
rect 19181 4570 19189 4590
rect 19209 4570 19223 4590
rect 19181 4532 19223 4570
rect 19273 4590 19317 4632
rect 19273 4570 19285 4590
rect 19305 4570 19317 4590
rect 19273 4532 19317 4570
rect 19394 4590 19436 4632
rect 19394 4570 19402 4590
rect 19422 4570 19436 4590
rect 19394 4532 19436 4570
rect 19486 4590 19530 4632
rect 19486 4570 19498 4590
rect 19518 4570 19530 4590
rect 19486 4532 19530 4570
rect 19811 4586 19855 4628
rect 19811 4566 19823 4586
rect 19843 4566 19855 4586
rect 19811 4559 19855 4566
rect 19810 4528 19855 4559
rect 19905 4586 19947 4628
rect 19905 4566 19919 4586
rect 19939 4566 19947 4586
rect 19905 4528 19947 4566
rect 20021 4586 20063 4628
rect 20021 4566 20029 4586
rect 20049 4566 20063 4586
rect 20021 4528 20063 4566
rect 20113 4586 20157 4628
rect 20113 4566 20125 4586
rect 20145 4566 20157 4586
rect 20113 4528 20157 4566
rect 20229 4586 20271 4628
rect 20229 4566 20237 4586
rect 20257 4566 20271 4586
rect 20229 4528 20271 4566
rect 20321 4586 20365 4628
rect 20321 4566 20333 4586
rect 20353 4566 20365 4586
rect 20321 4528 20365 4566
rect 20442 4586 20484 4628
rect 20442 4566 20450 4586
rect 20470 4566 20484 4586
rect 20442 4528 20484 4566
rect 20534 4586 20578 4628
rect 20534 4566 20546 4586
rect 20566 4566 20578 4586
rect 20534 4528 20578 4566
rect 814 3922 858 3960
rect 814 3902 826 3922
rect 846 3902 858 3922
rect 814 3860 858 3902
rect 908 3922 950 3960
rect 908 3902 922 3922
rect 942 3902 950 3922
rect 908 3860 950 3902
rect 1027 3922 1071 3960
rect 1027 3902 1039 3922
rect 1059 3902 1071 3922
rect 1027 3860 1071 3902
rect 1121 3922 1163 3960
rect 1121 3902 1135 3922
rect 1155 3902 1163 3922
rect 1121 3860 1163 3902
rect 1235 3922 1279 3960
rect 1235 3902 1247 3922
rect 1267 3902 1279 3922
rect 1235 3860 1279 3902
rect 1329 3922 1371 3960
rect 1329 3902 1343 3922
rect 1363 3902 1371 3922
rect 1329 3860 1371 3902
rect 1445 3922 1487 3960
rect 1445 3902 1453 3922
rect 1473 3902 1487 3922
rect 1445 3860 1487 3902
rect 1537 3929 1582 3960
rect 1537 3922 1581 3929
rect 1537 3902 1549 3922
rect 1569 3902 1581 3922
rect 1537 3860 1581 3902
rect 1862 3918 1906 3956
rect 1862 3898 1874 3918
rect 1894 3898 1906 3918
rect 1862 3856 1906 3898
rect 1956 3918 1998 3956
rect 1956 3898 1970 3918
rect 1990 3898 1998 3918
rect 1956 3856 1998 3898
rect 2075 3918 2119 3956
rect 2075 3898 2087 3918
rect 2107 3898 2119 3918
rect 2075 3856 2119 3898
rect 2169 3918 2211 3956
rect 2169 3898 2183 3918
rect 2203 3898 2211 3918
rect 2169 3856 2211 3898
rect 2283 3918 2327 3956
rect 2283 3898 2295 3918
rect 2315 3898 2327 3918
rect 2283 3856 2327 3898
rect 2377 3918 2419 3956
rect 2377 3898 2391 3918
rect 2411 3898 2419 3918
rect 2377 3856 2419 3898
rect 2493 3918 2535 3956
rect 2493 3898 2501 3918
rect 2521 3898 2535 3918
rect 2493 3856 2535 3898
rect 2585 3925 2630 3956
rect 2585 3918 2629 3925
rect 2585 3898 2597 3918
rect 2617 3898 2629 3918
rect 2585 3856 2629 3898
rect 4764 3924 4808 3962
rect 4764 3904 4776 3924
rect 4796 3904 4808 3924
rect 4764 3862 4808 3904
rect 4858 3924 4900 3962
rect 4858 3904 4872 3924
rect 4892 3904 4900 3924
rect 4858 3862 4900 3904
rect 4977 3924 5021 3962
rect 4977 3904 4989 3924
rect 5009 3904 5021 3924
rect 4977 3862 5021 3904
rect 5071 3924 5113 3962
rect 5071 3904 5085 3924
rect 5105 3904 5113 3924
rect 5071 3862 5113 3904
rect 5185 3924 5229 3962
rect 5185 3904 5197 3924
rect 5217 3904 5229 3924
rect 5185 3862 5229 3904
rect 5279 3924 5321 3962
rect 5279 3904 5293 3924
rect 5313 3904 5321 3924
rect 5279 3862 5321 3904
rect 5395 3924 5437 3962
rect 5395 3904 5403 3924
rect 5423 3904 5437 3924
rect 5395 3862 5437 3904
rect 5487 3931 5532 3962
rect 5487 3924 5531 3931
rect 5487 3904 5499 3924
rect 5519 3904 5531 3924
rect 5487 3862 5531 3904
rect 11522 3916 11566 3954
rect 6566 3754 6610 3796
rect 6566 3734 6578 3754
rect 6598 3734 6610 3754
rect 6566 3727 6610 3734
rect 6565 3696 6610 3727
rect 6660 3754 6702 3796
rect 6660 3734 6674 3754
rect 6694 3734 6702 3754
rect 6660 3696 6702 3734
rect 6776 3754 6818 3796
rect 6776 3734 6784 3754
rect 6804 3734 6818 3754
rect 6776 3696 6818 3734
rect 6868 3754 6912 3796
rect 6868 3734 6880 3754
rect 6900 3734 6912 3754
rect 6868 3696 6912 3734
rect 6984 3754 7026 3796
rect 6984 3734 6992 3754
rect 7012 3734 7026 3754
rect 6984 3696 7026 3734
rect 7076 3754 7120 3796
rect 7076 3734 7088 3754
rect 7108 3734 7120 3754
rect 7076 3696 7120 3734
rect 7197 3754 7239 3796
rect 7197 3734 7205 3754
rect 7225 3734 7239 3754
rect 7197 3696 7239 3734
rect 7289 3754 7333 3796
rect 11522 3896 11534 3916
rect 11554 3896 11566 3916
rect 11522 3854 11566 3896
rect 11616 3916 11658 3954
rect 11616 3896 11630 3916
rect 11650 3896 11658 3916
rect 11616 3854 11658 3896
rect 11735 3916 11779 3954
rect 11735 3896 11747 3916
rect 11767 3896 11779 3916
rect 11735 3854 11779 3896
rect 11829 3916 11871 3954
rect 11829 3896 11843 3916
rect 11863 3896 11871 3916
rect 11829 3854 11871 3896
rect 11943 3916 11987 3954
rect 11943 3896 11955 3916
rect 11975 3896 11987 3916
rect 11943 3854 11987 3896
rect 12037 3916 12079 3954
rect 12037 3896 12051 3916
rect 12071 3896 12079 3916
rect 12037 3854 12079 3896
rect 12153 3916 12195 3954
rect 12153 3896 12161 3916
rect 12181 3896 12195 3916
rect 12153 3854 12195 3896
rect 12245 3923 12290 3954
rect 12245 3916 12289 3923
rect 12245 3896 12257 3916
rect 12277 3896 12289 3916
rect 12245 3854 12289 3896
rect 12570 3912 12614 3950
rect 12570 3892 12582 3912
rect 12602 3892 12614 3912
rect 7289 3734 7301 3754
rect 7321 3734 7333 3754
rect 7289 3696 7333 3734
rect 9104 3751 9148 3793
rect 9104 3731 9116 3751
rect 9136 3731 9148 3751
rect 9104 3724 9148 3731
rect 9103 3693 9148 3724
rect 9198 3751 9240 3793
rect 9198 3731 9212 3751
rect 9232 3731 9240 3751
rect 9198 3693 9240 3731
rect 9314 3751 9356 3793
rect 9314 3731 9322 3751
rect 9342 3731 9356 3751
rect 9314 3693 9356 3731
rect 9406 3751 9450 3793
rect 9406 3731 9418 3751
rect 9438 3731 9450 3751
rect 9406 3693 9450 3731
rect 9522 3751 9564 3793
rect 9522 3731 9530 3751
rect 9550 3731 9564 3751
rect 9522 3693 9564 3731
rect 9614 3751 9658 3793
rect 9614 3731 9626 3751
rect 9646 3731 9658 3751
rect 9614 3693 9658 3731
rect 9735 3751 9777 3793
rect 9735 3731 9743 3751
rect 9763 3731 9777 3751
rect 9735 3693 9777 3731
rect 9827 3751 9871 3793
rect 12570 3850 12614 3892
rect 12664 3912 12706 3950
rect 12664 3892 12678 3912
rect 12698 3892 12706 3912
rect 12664 3850 12706 3892
rect 12783 3912 12827 3950
rect 12783 3892 12795 3912
rect 12815 3892 12827 3912
rect 12783 3850 12827 3892
rect 12877 3912 12919 3950
rect 12877 3892 12891 3912
rect 12911 3892 12919 3912
rect 12877 3850 12919 3892
rect 12991 3912 13035 3950
rect 12991 3892 13003 3912
rect 13023 3892 13035 3912
rect 12991 3850 13035 3892
rect 13085 3912 13127 3950
rect 13085 3892 13099 3912
rect 13119 3892 13127 3912
rect 13085 3850 13127 3892
rect 13201 3912 13243 3950
rect 13201 3892 13209 3912
rect 13229 3892 13243 3912
rect 13201 3850 13243 3892
rect 13293 3919 13338 3950
rect 13293 3912 13337 3919
rect 13293 3892 13305 3912
rect 13325 3892 13337 3912
rect 13293 3850 13337 3892
rect 15472 3918 15516 3956
rect 15472 3898 15484 3918
rect 15504 3898 15516 3918
rect 15472 3856 15516 3898
rect 15566 3918 15608 3956
rect 15566 3898 15580 3918
rect 15600 3898 15608 3918
rect 15566 3856 15608 3898
rect 15685 3918 15729 3956
rect 15685 3898 15697 3918
rect 15717 3898 15729 3918
rect 15685 3856 15729 3898
rect 15779 3918 15821 3956
rect 15779 3898 15793 3918
rect 15813 3898 15821 3918
rect 15779 3856 15821 3898
rect 15893 3918 15937 3956
rect 15893 3898 15905 3918
rect 15925 3898 15937 3918
rect 15893 3856 15937 3898
rect 15987 3918 16029 3956
rect 15987 3898 16001 3918
rect 16021 3898 16029 3918
rect 15987 3856 16029 3898
rect 16103 3918 16145 3956
rect 16103 3898 16111 3918
rect 16131 3898 16145 3918
rect 16103 3856 16145 3898
rect 16195 3925 16240 3956
rect 16195 3918 16239 3925
rect 16195 3898 16207 3918
rect 16227 3898 16239 3918
rect 16195 3856 16239 3898
rect 9827 3731 9839 3751
rect 9859 3731 9871 3751
rect 9827 3693 9871 3731
rect 17274 3748 17318 3790
rect 17274 3728 17286 3748
rect 17306 3728 17318 3748
rect 17274 3721 17318 3728
rect 17273 3690 17318 3721
rect 17368 3748 17410 3790
rect 17368 3728 17382 3748
rect 17402 3728 17410 3748
rect 17368 3690 17410 3728
rect 17484 3748 17526 3790
rect 17484 3728 17492 3748
rect 17512 3728 17526 3748
rect 17484 3690 17526 3728
rect 17576 3748 17620 3790
rect 17576 3728 17588 3748
rect 17608 3728 17620 3748
rect 17576 3690 17620 3728
rect 17692 3748 17734 3790
rect 17692 3728 17700 3748
rect 17720 3728 17734 3748
rect 17692 3690 17734 3728
rect 17784 3748 17828 3790
rect 17784 3728 17796 3748
rect 17816 3728 17828 3748
rect 17784 3690 17828 3728
rect 17905 3748 17947 3790
rect 17905 3728 17913 3748
rect 17933 3728 17947 3748
rect 17905 3690 17947 3728
rect 17997 3748 18041 3790
rect 17997 3728 18009 3748
rect 18029 3728 18041 3748
rect 17997 3690 18041 3728
rect 19812 3745 19856 3787
rect 19812 3725 19824 3745
rect 19844 3725 19856 3745
rect 19812 3718 19856 3725
rect 19811 3687 19856 3718
rect 19906 3745 19948 3787
rect 19906 3725 19920 3745
rect 19940 3725 19948 3745
rect 19906 3687 19948 3725
rect 20022 3745 20064 3787
rect 20022 3725 20030 3745
rect 20050 3725 20064 3745
rect 20022 3687 20064 3725
rect 20114 3745 20158 3787
rect 20114 3725 20126 3745
rect 20146 3725 20158 3745
rect 20114 3687 20158 3725
rect 20230 3745 20272 3787
rect 20230 3725 20238 3745
rect 20258 3725 20272 3745
rect 20230 3687 20272 3725
rect 20322 3745 20366 3787
rect 20322 3725 20334 3745
rect 20354 3725 20366 3745
rect 20322 3687 20366 3725
rect 20443 3745 20485 3787
rect 20443 3725 20451 3745
rect 20471 3725 20485 3745
rect 20443 3687 20485 3725
rect 20535 3745 20579 3787
rect 20535 3725 20547 3745
rect 20567 3725 20579 3745
rect 20535 3687 20579 3725
rect 814 3243 858 3281
rect 814 3223 826 3243
rect 846 3223 858 3243
rect 814 3181 858 3223
rect 908 3243 950 3281
rect 908 3223 922 3243
rect 942 3223 950 3243
rect 908 3181 950 3223
rect 1027 3243 1071 3281
rect 1027 3223 1039 3243
rect 1059 3223 1071 3243
rect 1027 3181 1071 3223
rect 1121 3243 1163 3281
rect 1121 3223 1135 3243
rect 1155 3223 1163 3243
rect 1121 3181 1163 3223
rect 1235 3243 1279 3281
rect 1235 3223 1247 3243
rect 1267 3223 1279 3243
rect 1235 3181 1279 3223
rect 1329 3243 1371 3281
rect 1329 3223 1343 3243
rect 1363 3223 1371 3243
rect 1329 3181 1371 3223
rect 1445 3243 1487 3281
rect 1445 3223 1453 3243
rect 1473 3223 1487 3243
rect 1445 3181 1487 3223
rect 1537 3250 1582 3281
rect 1537 3243 1581 3250
rect 1537 3223 1549 3243
rect 1569 3223 1581 3243
rect 1537 3181 1581 3223
rect 3309 3238 3353 3276
rect 3309 3218 3321 3238
rect 3341 3218 3353 3238
rect 3309 3176 3353 3218
rect 3403 3238 3445 3276
rect 3403 3218 3417 3238
rect 3437 3218 3445 3238
rect 3403 3176 3445 3218
rect 3522 3238 3566 3276
rect 3522 3218 3534 3238
rect 3554 3218 3566 3238
rect 3522 3176 3566 3218
rect 3616 3238 3658 3276
rect 3616 3218 3630 3238
rect 3650 3218 3658 3238
rect 3616 3176 3658 3218
rect 3730 3238 3774 3276
rect 3730 3218 3742 3238
rect 3762 3218 3774 3238
rect 3730 3176 3774 3218
rect 3824 3238 3866 3276
rect 3824 3218 3838 3238
rect 3858 3218 3866 3238
rect 3824 3176 3866 3218
rect 3940 3238 3982 3276
rect 3940 3218 3948 3238
rect 3968 3218 3982 3238
rect 3940 3176 3982 3218
rect 4032 3245 4077 3276
rect 4032 3238 4076 3245
rect 4032 3218 4044 3238
rect 4064 3218 4076 3238
rect 4032 3176 4076 3218
rect 11522 3237 11566 3275
rect 11522 3217 11534 3237
rect 11554 3217 11566 3237
rect 8056 3076 8100 3118
rect 8056 3056 8068 3076
rect 8088 3056 8100 3076
rect 8056 3049 8100 3056
rect 8055 3018 8100 3049
rect 8150 3076 8192 3118
rect 8150 3056 8164 3076
rect 8184 3056 8192 3076
rect 8150 3018 8192 3056
rect 8266 3076 8308 3118
rect 8266 3056 8274 3076
rect 8294 3056 8308 3076
rect 8266 3018 8308 3056
rect 8358 3076 8402 3118
rect 8358 3056 8370 3076
rect 8390 3056 8402 3076
rect 8358 3018 8402 3056
rect 8474 3076 8516 3118
rect 8474 3056 8482 3076
rect 8502 3056 8516 3076
rect 8474 3018 8516 3056
rect 8566 3076 8610 3118
rect 8566 3056 8578 3076
rect 8598 3056 8610 3076
rect 8566 3018 8610 3056
rect 8687 3076 8729 3118
rect 8687 3056 8695 3076
rect 8715 3056 8729 3076
rect 8687 3018 8729 3056
rect 8779 3076 8823 3118
rect 11522 3175 11566 3217
rect 11616 3237 11658 3275
rect 11616 3217 11630 3237
rect 11650 3217 11658 3237
rect 11616 3175 11658 3217
rect 11735 3237 11779 3275
rect 11735 3217 11747 3237
rect 11767 3217 11779 3237
rect 11735 3175 11779 3217
rect 11829 3237 11871 3275
rect 11829 3217 11843 3237
rect 11863 3217 11871 3237
rect 11829 3175 11871 3217
rect 11943 3237 11987 3275
rect 11943 3217 11955 3237
rect 11975 3217 11987 3237
rect 11943 3175 11987 3217
rect 12037 3237 12079 3275
rect 12037 3217 12051 3237
rect 12071 3217 12079 3237
rect 12037 3175 12079 3217
rect 12153 3237 12195 3275
rect 12153 3217 12161 3237
rect 12181 3217 12195 3237
rect 12153 3175 12195 3217
rect 12245 3244 12290 3275
rect 12245 3237 12289 3244
rect 12245 3217 12257 3237
rect 12277 3217 12289 3237
rect 12245 3175 12289 3217
rect 14017 3232 14061 3270
rect 14017 3212 14029 3232
rect 14049 3212 14061 3232
rect 8779 3056 8791 3076
rect 8811 3056 8823 3076
rect 8779 3018 8823 3056
rect 9104 3072 9148 3114
rect 9104 3052 9116 3072
rect 9136 3052 9148 3072
rect 9104 3045 9148 3052
rect 9103 3014 9148 3045
rect 9198 3072 9240 3114
rect 9198 3052 9212 3072
rect 9232 3052 9240 3072
rect 9198 3014 9240 3052
rect 9314 3072 9356 3114
rect 9314 3052 9322 3072
rect 9342 3052 9356 3072
rect 9314 3014 9356 3052
rect 9406 3072 9450 3114
rect 9406 3052 9418 3072
rect 9438 3052 9450 3072
rect 9406 3014 9450 3052
rect 9522 3072 9564 3114
rect 9522 3052 9530 3072
rect 9550 3052 9564 3072
rect 9522 3014 9564 3052
rect 9614 3072 9658 3114
rect 9614 3052 9626 3072
rect 9646 3052 9658 3072
rect 9614 3014 9658 3052
rect 9735 3072 9777 3114
rect 9735 3052 9743 3072
rect 9763 3052 9777 3072
rect 9735 3014 9777 3052
rect 9827 3072 9871 3114
rect 9827 3052 9839 3072
rect 9859 3052 9871 3072
rect 14017 3170 14061 3212
rect 14111 3232 14153 3270
rect 14111 3212 14125 3232
rect 14145 3212 14153 3232
rect 14111 3170 14153 3212
rect 14230 3232 14274 3270
rect 14230 3212 14242 3232
rect 14262 3212 14274 3232
rect 14230 3170 14274 3212
rect 14324 3232 14366 3270
rect 14324 3212 14338 3232
rect 14358 3212 14366 3232
rect 14324 3170 14366 3212
rect 14438 3232 14482 3270
rect 14438 3212 14450 3232
rect 14470 3212 14482 3232
rect 14438 3170 14482 3212
rect 14532 3232 14574 3270
rect 14532 3212 14546 3232
rect 14566 3212 14574 3232
rect 14532 3170 14574 3212
rect 14648 3232 14690 3270
rect 14648 3212 14656 3232
rect 14676 3212 14690 3232
rect 14648 3170 14690 3212
rect 14740 3239 14785 3270
rect 14740 3232 14784 3239
rect 14740 3212 14752 3232
rect 14772 3212 14784 3232
rect 14740 3170 14784 3212
rect 9827 3014 9871 3052
rect 18764 3070 18808 3112
rect 18764 3050 18776 3070
rect 18796 3050 18808 3070
rect 18764 3043 18808 3050
rect 18763 3012 18808 3043
rect 18858 3070 18900 3112
rect 18858 3050 18872 3070
rect 18892 3050 18900 3070
rect 18858 3012 18900 3050
rect 18974 3070 19016 3112
rect 18974 3050 18982 3070
rect 19002 3050 19016 3070
rect 18974 3012 19016 3050
rect 19066 3070 19110 3112
rect 19066 3050 19078 3070
rect 19098 3050 19110 3070
rect 19066 3012 19110 3050
rect 19182 3070 19224 3112
rect 19182 3050 19190 3070
rect 19210 3050 19224 3070
rect 19182 3012 19224 3050
rect 19274 3070 19318 3112
rect 19274 3050 19286 3070
rect 19306 3050 19318 3070
rect 19274 3012 19318 3050
rect 19395 3070 19437 3112
rect 19395 3050 19403 3070
rect 19423 3050 19437 3070
rect 19395 3012 19437 3050
rect 19487 3070 19531 3112
rect 19487 3050 19499 3070
rect 19519 3050 19531 3070
rect 19487 3012 19531 3050
rect 19812 3066 19856 3108
rect 19812 3046 19824 3066
rect 19844 3046 19856 3066
rect 19812 3039 19856 3046
rect 19811 3008 19856 3039
rect 19906 3066 19948 3108
rect 19906 3046 19920 3066
rect 19940 3046 19948 3066
rect 19906 3008 19948 3046
rect 20022 3066 20064 3108
rect 20022 3046 20030 3066
rect 20050 3046 20064 3066
rect 20022 3008 20064 3046
rect 20114 3066 20158 3108
rect 20114 3046 20126 3066
rect 20146 3046 20158 3066
rect 20114 3008 20158 3046
rect 20230 3066 20272 3108
rect 20230 3046 20238 3066
rect 20258 3046 20272 3066
rect 20230 3008 20272 3046
rect 20322 3066 20366 3108
rect 20322 3046 20334 3066
rect 20354 3046 20366 3066
rect 20322 3008 20366 3046
rect 20443 3066 20485 3108
rect 20443 3046 20451 3066
rect 20471 3046 20485 3066
rect 20443 3008 20485 3046
rect 20535 3066 20579 3108
rect 20535 3046 20547 3066
rect 20567 3046 20579 3066
rect 20535 3008 20579 3046
rect 814 2475 858 2513
rect 814 2455 826 2475
rect 846 2455 858 2475
rect 814 2413 858 2455
rect 908 2475 950 2513
rect 908 2455 922 2475
rect 942 2455 950 2475
rect 908 2413 950 2455
rect 1027 2475 1071 2513
rect 1027 2455 1039 2475
rect 1059 2455 1071 2475
rect 1027 2413 1071 2455
rect 1121 2475 1163 2513
rect 1121 2455 1135 2475
rect 1155 2455 1163 2475
rect 1121 2413 1163 2455
rect 1235 2475 1279 2513
rect 1235 2455 1247 2475
rect 1267 2455 1279 2475
rect 1235 2413 1279 2455
rect 1329 2475 1371 2513
rect 1329 2455 1343 2475
rect 1363 2455 1371 2475
rect 1329 2413 1371 2455
rect 1445 2475 1487 2513
rect 1445 2455 1453 2475
rect 1473 2455 1487 2475
rect 1445 2413 1487 2455
rect 1537 2482 1582 2513
rect 1537 2475 1581 2482
rect 1537 2455 1549 2475
rect 1569 2455 1581 2475
rect 1537 2413 1581 2455
rect 1862 2471 1906 2509
rect 1862 2451 1874 2471
rect 1894 2451 1906 2471
rect 1862 2409 1906 2451
rect 1956 2471 1998 2509
rect 1956 2451 1970 2471
rect 1990 2451 1998 2471
rect 1956 2409 1998 2451
rect 2075 2471 2119 2509
rect 2075 2451 2087 2471
rect 2107 2451 2119 2471
rect 2075 2409 2119 2451
rect 2169 2471 2211 2509
rect 2169 2451 2183 2471
rect 2203 2451 2211 2471
rect 2169 2409 2211 2451
rect 2283 2471 2327 2509
rect 2283 2451 2295 2471
rect 2315 2451 2327 2471
rect 2283 2409 2327 2451
rect 2377 2471 2419 2509
rect 2377 2451 2391 2471
rect 2411 2451 2419 2471
rect 2377 2409 2419 2451
rect 2493 2471 2535 2509
rect 2493 2451 2501 2471
rect 2521 2451 2535 2471
rect 2493 2409 2535 2451
rect 2585 2478 2630 2509
rect 2585 2471 2629 2478
rect 2585 2451 2597 2471
rect 2617 2451 2629 2471
rect 2585 2409 2629 2451
rect 11522 2469 11566 2507
rect 6609 2309 6653 2351
rect 6609 2289 6621 2309
rect 6641 2289 6653 2309
rect 6609 2282 6653 2289
rect 6608 2251 6653 2282
rect 6703 2309 6745 2351
rect 6703 2289 6717 2309
rect 6737 2289 6745 2309
rect 6703 2251 6745 2289
rect 6819 2309 6861 2351
rect 6819 2289 6827 2309
rect 6847 2289 6861 2309
rect 6819 2251 6861 2289
rect 6911 2309 6955 2351
rect 6911 2289 6923 2309
rect 6943 2289 6955 2309
rect 6911 2251 6955 2289
rect 7027 2309 7069 2351
rect 7027 2289 7035 2309
rect 7055 2289 7069 2309
rect 7027 2251 7069 2289
rect 7119 2309 7163 2351
rect 7119 2289 7131 2309
rect 7151 2289 7163 2309
rect 7119 2251 7163 2289
rect 7240 2309 7282 2351
rect 7240 2289 7248 2309
rect 7268 2289 7282 2309
rect 7240 2251 7282 2289
rect 7332 2309 7376 2351
rect 11522 2449 11534 2469
rect 11554 2449 11566 2469
rect 11522 2407 11566 2449
rect 11616 2469 11658 2507
rect 11616 2449 11630 2469
rect 11650 2449 11658 2469
rect 11616 2407 11658 2449
rect 11735 2469 11779 2507
rect 11735 2449 11747 2469
rect 11767 2449 11779 2469
rect 11735 2407 11779 2449
rect 11829 2469 11871 2507
rect 11829 2449 11843 2469
rect 11863 2449 11871 2469
rect 11829 2407 11871 2449
rect 11943 2469 11987 2507
rect 11943 2449 11955 2469
rect 11975 2449 11987 2469
rect 11943 2407 11987 2449
rect 12037 2469 12079 2507
rect 12037 2449 12051 2469
rect 12071 2449 12079 2469
rect 12037 2407 12079 2449
rect 12153 2469 12195 2507
rect 12153 2449 12161 2469
rect 12181 2449 12195 2469
rect 12153 2407 12195 2449
rect 12245 2476 12290 2507
rect 12245 2469 12289 2476
rect 12245 2449 12257 2469
rect 12277 2449 12289 2469
rect 12245 2407 12289 2449
rect 12570 2465 12614 2503
rect 12570 2445 12582 2465
rect 12602 2445 12614 2465
rect 7332 2289 7344 2309
rect 7364 2289 7376 2309
rect 7332 2251 7376 2289
rect 9104 2304 9148 2346
rect 9104 2284 9116 2304
rect 9136 2284 9148 2304
rect 9104 2277 9148 2284
rect 9103 2246 9148 2277
rect 9198 2304 9240 2346
rect 9198 2284 9212 2304
rect 9232 2284 9240 2304
rect 9198 2246 9240 2284
rect 9314 2304 9356 2346
rect 9314 2284 9322 2304
rect 9342 2284 9356 2304
rect 9314 2246 9356 2284
rect 9406 2304 9450 2346
rect 9406 2284 9418 2304
rect 9438 2284 9450 2304
rect 9406 2246 9450 2284
rect 9522 2304 9564 2346
rect 9522 2284 9530 2304
rect 9550 2284 9564 2304
rect 9522 2246 9564 2284
rect 9614 2304 9658 2346
rect 9614 2284 9626 2304
rect 9646 2284 9658 2304
rect 9614 2246 9658 2284
rect 9735 2304 9777 2346
rect 9735 2284 9743 2304
rect 9763 2284 9777 2304
rect 9735 2246 9777 2284
rect 9827 2304 9871 2346
rect 12570 2403 12614 2445
rect 12664 2465 12706 2503
rect 12664 2445 12678 2465
rect 12698 2445 12706 2465
rect 12664 2403 12706 2445
rect 12783 2465 12827 2503
rect 12783 2445 12795 2465
rect 12815 2445 12827 2465
rect 12783 2403 12827 2445
rect 12877 2465 12919 2503
rect 12877 2445 12891 2465
rect 12911 2445 12919 2465
rect 12877 2403 12919 2445
rect 12991 2465 13035 2503
rect 12991 2445 13003 2465
rect 13023 2445 13035 2465
rect 12991 2403 13035 2445
rect 13085 2465 13127 2503
rect 13085 2445 13099 2465
rect 13119 2445 13127 2465
rect 13085 2403 13127 2445
rect 13201 2465 13243 2503
rect 13201 2445 13209 2465
rect 13229 2445 13243 2465
rect 13201 2403 13243 2445
rect 13293 2472 13338 2503
rect 13293 2465 13337 2472
rect 13293 2445 13305 2465
rect 13325 2445 13337 2465
rect 13293 2403 13337 2445
rect 9827 2284 9839 2304
rect 9859 2284 9871 2304
rect 9827 2246 9871 2284
rect 17317 2303 17361 2345
rect 17317 2283 17329 2303
rect 17349 2283 17361 2303
rect 17317 2276 17361 2283
rect 17316 2245 17361 2276
rect 17411 2303 17453 2345
rect 17411 2283 17425 2303
rect 17445 2283 17453 2303
rect 17411 2245 17453 2283
rect 17527 2303 17569 2345
rect 17527 2283 17535 2303
rect 17555 2283 17569 2303
rect 17527 2245 17569 2283
rect 17619 2303 17663 2345
rect 17619 2283 17631 2303
rect 17651 2283 17663 2303
rect 17619 2245 17663 2283
rect 17735 2303 17777 2345
rect 17735 2283 17743 2303
rect 17763 2283 17777 2303
rect 17735 2245 17777 2283
rect 17827 2303 17871 2345
rect 17827 2283 17839 2303
rect 17859 2283 17871 2303
rect 17827 2245 17871 2283
rect 17948 2303 17990 2345
rect 17948 2283 17956 2303
rect 17976 2283 17990 2303
rect 17948 2245 17990 2283
rect 18040 2303 18084 2345
rect 18040 2283 18052 2303
rect 18072 2283 18084 2303
rect 18040 2245 18084 2283
rect 19812 2298 19856 2340
rect 19812 2278 19824 2298
rect 19844 2278 19856 2298
rect 19812 2271 19856 2278
rect 19811 2240 19856 2271
rect 19906 2298 19948 2340
rect 19906 2278 19920 2298
rect 19940 2278 19948 2298
rect 19906 2240 19948 2278
rect 20022 2298 20064 2340
rect 20022 2278 20030 2298
rect 20050 2278 20064 2298
rect 20022 2240 20064 2278
rect 20114 2298 20158 2340
rect 20114 2278 20126 2298
rect 20146 2278 20158 2298
rect 20114 2240 20158 2278
rect 20230 2298 20272 2340
rect 20230 2278 20238 2298
rect 20258 2278 20272 2298
rect 20230 2240 20272 2278
rect 20322 2298 20366 2340
rect 20322 2278 20334 2298
rect 20354 2278 20366 2298
rect 20322 2240 20366 2278
rect 20443 2298 20485 2340
rect 20443 2278 20451 2298
rect 20471 2278 20485 2298
rect 20443 2240 20485 2278
rect 20535 2298 20579 2340
rect 20535 2278 20547 2298
rect 20567 2278 20579 2298
rect 20535 2240 20579 2278
rect 814 1796 858 1834
rect 814 1776 826 1796
rect 846 1776 858 1796
rect 814 1734 858 1776
rect 908 1796 950 1834
rect 908 1776 922 1796
rect 942 1776 950 1796
rect 908 1734 950 1776
rect 1027 1796 1071 1834
rect 1027 1776 1039 1796
rect 1059 1776 1071 1796
rect 1027 1734 1071 1776
rect 1121 1796 1163 1834
rect 1121 1776 1135 1796
rect 1155 1776 1163 1796
rect 1121 1734 1163 1776
rect 1235 1796 1279 1834
rect 1235 1776 1247 1796
rect 1267 1776 1279 1796
rect 1235 1734 1279 1776
rect 1329 1796 1371 1834
rect 1329 1776 1343 1796
rect 1363 1776 1371 1796
rect 1329 1734 1371 1776
rect 1445 1796 1487 1834
rect 1445 1776 1453 1796
rect 1473 1776 1487 1796
rect 1445 1734 1487 1776
rect 1537 1803 1582 1834
rect 1537 1796 1581 1803
rect 1537 1776 1549 1796
rect 1569 1776 1581 1796
rect 1537 1734 1581 1776
rect 11522 1790 11566 1828
rect 11522 1770 11534 1790
rect 11554 1770 11566 1790
rect 8056 1629 8100 1671
rect 8056 1609 8068 1629
rect 8088 1609 8100 1629
rect 8056 1602 8100 1609
rect 8055 1571 8100 1602
rect 8150 1629 8192 1671
rect 8150 1609 8164 1629
rect 8184 1609 8192 1629
rect 8150 1571 8192 1609
rect 8266 1629 8308 1671
rect 8266 1609 8274 1629
rect 8294 1609 8308 1629
rect 8266 1571 8308 1609
rect 8358 1629 8402 1671
rect 8358 1609 8370 1629
rect 8390 1609 8402 1629
rect 8358 1571 8402 1609
rect 8474 1629 8516 1671
rect 8474 1609 8482 1629
rect 8502 1609 8516 1629
rect 8474 1571 8516 1609
rect 8566 1629 8610 1671
rect 8566 1609 8578 1629
rect 8598 1609 8610 1629
rect 8566 1571 8610 1609
rect 8687 1629 8729 1671
rect 8687 1609 8695 1629
rect 8715 1609 8729 1629
rect 8687 1571 8729 1609
rect 8779 1629 8823 1671
rect 11522 1728 11566 1770
rect 11616 1790 11658 1828
rect 11616 1770 11630 1790
rect 11650 1770 11658 1790
rect 11616 1728 11658 1770
rect 11735 1790 11779 1828
rect 11735 1770 11747 1790
rect 11767 1770 11779 1790
rect 11735 1728 11779 1770
rect 11829 1790 11871 1828
rect 11829 1770 11843 1790
rect 11863 1770 11871 1790
rect 11829 1728 11871 1770
rect 11943 1790 11987 1828
rect 11943 1770 11955 1790
rect 11975 1770 11987 1790
rect 11943 1728 11987 1770
rect 12037 1790 12079 1828
rect 12037 1770 12051 1790
rect 12071 1770 12079 1790
rect 12037 1728 12079 1770
rect 12153 1790 12195 1828
rect 12153 1770 12161 1790
rect 12181 1770 12195 1790
rect 12153 1728 12195 1770
rect 12245 1797 12290 1828
rect 12245 1790 12289 1797
rect 12245 1770 12257 1790
rect 12277 1770 12289 1790
rect 12245 1728 12289 1770
rect 8779 1609 8791 1629
rect 8811 1609 8823 1629
rect 8779 1571 8823 1609
rect 9104 1625 9148 1667
rect 9104 1605 9116 1625
rect 9136 1605 9148 1625
rect 9104 1598 9148 1605
rect 9103 1567 9148 1598
rect 9198 1625 9240 1667
rect 9198 1605 9212 1625
rect 9232 1605 9240 1625
rect 9198 1567 9240 1605
rect 9314 1625 9356 1667
rect 9314 1605 9322 1625
rect 9342 1605 9356 1625
rect 9314 1567 9356 1605
rect 9406 1625 9450 1667
rect 9406 1605 9418 1625
rect 9438 1605 9450 1625
rect 9406 1567 9450 1605
rect 9522 1625 9564 1667
rect 9522 1605 9530 1625
rect 9550 1605 9564 1625
rect 9522 1567 9564 1605
rect 9614 1625 9658 1667
rect 9614 1605 9626 1625
rect 9646 1605 9658 1625
rect 9614 1567 9658 1605
rect 9735 1625 9777 1667
rect 9735 1605 9743 1625
rect 9763 1605 9777 1625
rect 9735 1567 9777 1605
rect 9827 1625 9871 1667
rect 9827 1605 9839 1625
rect 9859 1605 9871 1625
rect 9827 1567 9871 1605
rect 18764 1623 18808 1665
rect 18764 1603 18776 1623
rect 18796 1603 18808 1623
rect 18764 1596 18808 1603
rect 18763 1565 18808 1596
rect 18858 1623 18900 1665
rect 18858 1603 18872 1623
rect 18892 1603 18900 1623
rect 18858 1565 18900 1603
rect 18974 1623 19016 1665
rect 18974 1603 18982 1623
rect 19002 1603 19016 1623
rect 18974 1565 19016 1603
rect 19066 1623 19110 1665
rect 19066 1603 19078 1623
rect 19098 1603 19110 1623
rect 19066 1565 19110 1603
rect 19182 1623 19224 1665
rect 19182 1603 19190 1623
rect 19210 1603 19224 1623
rect 19182 1565 19224 1603
rect 19274 1623 19318 1665
rect 19274 1603 19286 1623
rect 19306 1603 19318 1623
rect 19274 1565 19318 1603
rect 19395 1623 19437 1665
rect 19395 1603 19403 1623
rect 19423 1603 19437 1623
rect 19395 1565 19437 1603
rect 19487 1623 19531 1665
rect 19487 1603 19499 1623
rect 19519 1603 19531 1623
rect 19487 1565 19531 1603
rect 19812 1619 19856 1661
rect 19812 1599 19824 1619
rect 19844 1599 19856 1619
rect 19812 1592 19856 1599
rect 19811 1561 19856 1592
rect 19906 1619 19948 1661
rect 19906 1599 19920 1619
rect 19940 1599 19948 1619
rect 19906 1561 19948 1599
rect 20022 1619 20064 1661
rect 20022 1599 20030 1619
rect 20050 1599 20064 1619
rect 20022 1561 20064 1599
rect 20114 1619 20158 1661
rect 20114 1599 20126 1619
rect 20146 1599 20158 1619
rect 20114 1561 20158 1599
rect 20230 1619 20272 1661
rect 20230 1599 20238 1619
rect 20258 1599 20272 1619
rect 20230 1561 20272 1599
rect 20322 1619 20366 1661
rect 20322 1599 20334 1619
rect 20354 1599 20366 1619
rect 20322 1561 20366 1599
rect 20443 1619 20485 1661
rect 20443 1599 20451 1619
rect 20471 1599 20485 1619
rect 20443 1561 20485 1599
rect 20535 1619 20579 1661
rect 20535 1599 20547 1619
rect 20567 1599 20579 1619
rect 20535 1561 20579 1599
rect 10525 -363 10569 -325
rect 10525 -383 10537 -363
rect 10557 -383 10569 -363
rect 10525 -425 10569 -383
rect 10619 -363 10661 -325
rect 10619 -383 10633 -363
rect 10653 -383 10661 -363
rect 10619 -425 10661 -383
rect 10738 -363 10782 -325
rect 10738 -383 10750 -363
rect 10770 -383 10782 -363
rect 10738 -425 10782 -383
rect 10832 -363 10874 -325
rect 10832 -383 10846 -363
rect 10866 -383 10874 -363
rect 10832 -425 10874 -383
rect 10946 -363 10990 -325
rect 10946 -383 10958 -363
rect 10978 -383 10990 -363
rect 10946 -425 10990 -383
rect 11040 -363 11082 -325
rect 11040 -383 11054 -363
rect 11074 -383 11082 -363
rect 11040 -425 11082 -383
rect 11156 -363 11198 -325
rect 11156 -383 11164 -363
rect 11184 -383 11198 -363
rect 11156 -425 11198 -383
rect 11248 -356 11293 -325
rect 11248 -363 11292 -356
rect 11248 -383 11260 -363
rect 11280 -383 11292 -363
rect 11248 -425 11292 -383
<< ndiffc >>
rect 501 13051 519 13069
rect 11209 13045 11227 13063
rect 503 12952 521 12970
rect 11211 12946 11229 12964
rect 501 12795 519 12813
rect 9111 12855 9131 12875
rect 9214 12851 9234 12871
rect 9322 12851 9342 12871
rect 9425 12855 9445 12875
rect 9530 12851 9550 12871
rect 9633 12855 9653 12875
rect 9743 12851 9763 12871
rect 9846 12855 9866 12875
rect 10166 12860 10184 12878
rect 821 12728 841 12748
rect 924 12732 944 12752
rect 1034 12728 1054 12748
rect 1137 12732 1157 12752
rect 1242 12728 1262 12748
rect 1345 12732 1365 12752
rect 1453 12732 1473 12752
rect 1556 12728 1576 12748
rect 1869 12724 1889 12744
rect 503 12696 521 12714
rect 1972 12728 1992 12748
rect 2082 12724 2102 12744
rect 2185 12728 2205 12748
rect 2290 12724 2310 12744
rect 2393 12728 2413 12748
rect 2501 12728 2521 12748
rect 2604 12724 2624 12744
rect 10168 12761 10186 12779
rect 11209 12789 11227 12807
rect 19819 12849 19839 12869
rect 19922 12845 19942 12865
rect 20030 12845 20050 12865
rect 20133 12849 20153 12869
rect 20238 12845 20258 12865
rect 20341 12849 20361 12869
rect 20451 12845 20471 12865
rect 20554 12849 20574 12869
rect 20874 12854 20892 12872
rect 11529 12722 11549 12742
rect 11632 12726 11652 12746
rect 11742 12722 11762 12742
rect 11845 12726 11865 12746
rect 11950 12722 11970 12742
rect 12053 12726 12073 12746
rect 12161 12726 12181 12746
rect 12264 12722 12284 12742
rect 12577 12718 12597 12738
rect 11211 12690 11229 12708
rect 12680 12722 12700 12742
rect 12790 12718 12810 12738
rect 12893 12722 12913 12742
rect 12998 12718 13018 12738
rect 13101 12722 13121 12742
rect 13209 12722 13229 12742
rect 13312 12718 13332 12738
rect 10166 12605 10184 12623
rect 20876 12755 20894 12773
rect 20874 12599 20892 12617
rect 10168 12506 10186 12524
rect 20876 12500 20894 12518
rect 501 12400 519 12418
rect 11209 12394 11227 12412
rect 503 12301 521 12319
rect 501 12145 519 12163
rect 11211 12295 11229 12313
rect 8063 12180 8083 12200
rect 8166 12176 8186 12196
rect 8274 12176 8294 12196
rect 8377 12180 8397 12200
rect 8482 12176 8502 12196
rect 8585 12180 8605 12200
rect 8695 12176 8715 12196
rect 10166 12210 10184 12228
rect 8798 12180 8818 12200
rect 9111 12176 9131 12196
rect 503 12046 521 12064
rect 821 12049 841 12069
rect 924 12053 944 12073
rect 1034 12049 1054 12069
rect 1137 12053 1157 12073
rect 1242 12049 1262 12069
rect 1345 12053 1365 12073
rect 1453 12053 1473 12073
rect 9214 12172 9234 12192
rect 9322 12172 9342 12192
rect 9425 12176 9445 12196
rect 9530 12172 9550 12192
rect 9633 12176 9653 12196
rect 9743 12172 9763 12192
rect 9846 12176 9866 12196
rect 1556 12049 1576 12069
rect 3316 12044 3336 12064
rect 3419 12048 3439 12068
rect 3529 12044 3549 12064
rect 3632 12048 3652 12068
rect 3737 12044 3757 12064
rect 3840 12048 3860 12068
rect 3948 12048 3968 12068
rect 4051 12044 4071 12064
rect 10168 12111 10186 12129
rect 11209 12139 11227 12157
rect 18771 12174 18791 12194
rect 18874 12170 18894 12190
rect 18982 12170 19002 12190
rect 19085 12174 19105 12194
rect 19190 12170 19210 12190
rect 19293 12174 19313 12194
rect 19403 12170 19423 12190
rect 20874 12204 20892 12222
rect 19506 12174 19526 12194
rect 19819 12170 19839 12190
rect 11211 12040 11229 12058
rect 11529 12043 11549 12063
rect 11632 12047 11652 12067
rect 11742 12043 11762 12063
rect 11845 12047 11865 12067
rect 11950 12043 11970 12063
rect 12053 12047 12073 12067
rect 12161 12047 12181 12067
rect 19922 12166 19942 12186
rect 20030 12166 20050 12186
rect 20133 12170 20153 12190
rect 20238 12166 20258 12186
rect 20341 12170 20361 12190
rect 20451 12166 20471 12186
rect 20554 12170 20574 12190
rect 12264 12043 12284 12063
rect 14024 12038 14044 12058
rect 14127 12042 14147 12062
rect 14237 12038 14257 12058
rect 14340 12042 14360 12062
rect 14445 12038 14465 12058
rect 14548 12042 14568 12062
rect 14656 12042 14676 12062
rect 14759 12038 14779 12058
rect 20876 12105 20894 12123
rect 10166 11954 10184 11972
rect 20874 11948 20892 11966
rect 10168 11855 10186 11873
rect 20876 11849 20894 11867
rect 501 11604 519 11622
rect 11209 11598 11227 11616
rect 503 11505 521 11523
rect 11211 11499 11229 11517
rect 501 11348 519 11366
rect 6616 11413 6636 11433
rect 6719 11409 6739 11429
rect 6827 11409 6847 11429
rect 6930 11413 6950 11433
rect 7035 11409 7055 11429
rect 7138 11413 7158 11433
rect 7248 11409 7268 11429
rect 7351 11413 7371 11433
rect 9111 11408 9131 11428
rect 821 11281 841 11301
rect 924 11285 944 11305
rect 1034 11281 1054 11301
rect 1137 11285 1157 11305
rect 1242 11281 1262 11301
rect 1345 11285 1365 11305
rect 1453 11285 1473 11305
rect 9214 11404 9234 11424
rect 9322 11404 9342 11424
rect 9425 11408 9445 11428
rect 9530 11404 9550 11424
rect 9633 11408 9653 11428
rect 9743 11404 9763 11424
rect 9846 11408 9866 11428
rect 10166 11413 10184 11431
rect 1556 11281 1576 11301
rect 1869 11277 1889 11297
rect 503 11249 521 11267
rect 1972 11281 1992 11301
rect 2082 11277 2102 11297
rect 2185 11281 2205 11301
rect 2290 11277 2310 11297
rect 2393 11281 2413 11301
rect 2501 11281 2521 11301
rect 2604 11277 2624 11297
rect 10168 11314 10186 11332
rect 11209 11342 11227 11360
rect 17324 11407 17344 11427
rect 17427 11403 17447 11423
rect 17535 11403 17555 11423
rect 17638 11407 17658 11427
rect 17743 11403 17763 11423
rect 17846 11407 17866 11427
rect 17956 11403 17976 11423
rect 18059 11407 18079 11427
rect 19819 11402 19839 11422
rect 11529 11275 11549 11295
rect 11632 11279 11652 11299
rect 11742 11275 11762 11295
rect 11845 11279 11865 11299
rect 11950 11275 11970 11295
rect 12053 11279 12073 11299
rect 12161 11279 12181 11299
rect 19922 11398 19942 11418
rect 20030 11398 20050 11418
rect 20133 11402 20153 11422
rect 20238 11398 20258 11418
rect 20341 11402 20361 11422
rect 20451 11398 20471 11418
rect 20554 11402 20574 11422
rect 20874 11407 20892 11425
rect 12264 11275 12284 11295
rect 12577 11271 12597 11291
rect 11211 11243 11229 11261
rect 12680 11275 12700 11295
rect 12790 11271 12810 11291
rect 12893 11275 12913 11295
rect 12998 11271 13018 11291
rect 13101 11275 13121 11295
rect 13209 11275 13229 11295
rect 13312 11271 13332 11291
rect 10166 11158 10184 11176
rect 20876 11308 20894 11326
rect 20874 11152 20892 11170
rect 10168 11059 10186 11077
rect 20876 11053 20894 11071
rect 501 10953 519 10971
rect 11209 10947 11227 10965
rect 503 10854 521 10872
rect 501 10698 519 10716
rect 11211 10848 11229 10866
rect 8063 10733 8083 10753
rect 8166 10729 8186 10749
rect 8274 10729 8294 10749
rect 8377 10733 8397 10753
rect 8482 10729 8502 10749
rect 8585 10733 8605 10753
rect 8695 10729 8715 10749
rect 10166 10763 10184 10781
rect 8798 10733 8818 10753
rect 9111 10729 9131 10749
rect 503 10599 521 10617
rect 821 10602 841 10622
rect 924 10606 944 10626
rect 1034 10602 1054 10622
rect 1137 10606 1157 10626
rect 1242 10602 1262 10622
rect 1345 10606 1365 10626
rect 1453 10606 1473 10626
rect 9214 10725 9234 10745
rect 9322 10725 9342 10745
rect 9425 10729 9445 10749
rect 9530 10725 9550 10745
rect 9633 10729 9653 10749
rect 9743 10725 9763 10745
rect 9846 10729 9866 10749
rect 1556 10602 1576 10622
rect 3359 10599 3379 10619
rect 3462 10603 3482 10623
rect 3572 10599 3592 10619
rect 3675 10603 3695 10623
rect 3780 10599 3800 10619
rect 3883 10603 3903 10623
rect 3991 10603 4011 10623
rect 4094 10599 4114 10619
rect 10168 10664 10186 10682
rect 11209 10692 11227 10710
rect 18771 10727 18791 10747
rect 18874 10723 18894 10743
rect 18982 10723 19002 10743
rect 19085 10727 19105 10747
rect 19190 10723 19210 10743
rect 19293 10727 19313 10747
rect 19403 10723 19423 10743
rect 20874 10757 20892 10775
rect 19506 10727 19526 10747
rect 19819 10723 19839 10743
rect 11211 10593 11229 10611
rect 11529 10596 11549 10616
rect 11632 10600 11652 10620
rect 11742 10596 11762 10616
rect 11845 10600 11865 10620
rect 11950 10596 11970 10616
rect 12053 10600 12073 10620
rect 12161 10600 12181 10620
rect 19922 10719 19942 10739
rect 20030 10719 20050 10739
rect 20133 10723 20153 10743
rect 20238 10719 20258 10739
rect 20341 10723 20361 10743
rect 20451 10719 20471 10739
rect 20554 10723 20574 10743
rect 12264 10596 12284 10616
rect 14067 10593 14087 10613
rect 14170 10597 14190 10617
rect 14280 10593 14300 10613
rect 14383 10597 14403 10617
rect 14488 10593 14508 10613
rect 14591 10597 14611 10617
rect 14699 10597 14719 10617
rect 14802 10593 14822 10613
rect 20876 10658 20894 10676
rect 10166 10507 10184 10525
rect 20874 10501 20892 10519
rect 10168 10408 10186 10426
rect 20876 10402 20894 10420
rect 502 10084 520 10102
rect 11210 10078 11228 10096
rect 504 9985 522 10003
rect 11212 9979 11230 9997
rect 502 9828 520 9846
rect 6574 9891 6594 9911
rect 6677 9887 6697 9907
rect 6785 9887 6805 9907
rect 6888 9891 6908 9911
rect 6993 9887 7013 9907
rect 7096 9891 7116 9911
rect 7206 9887 7226 9907
rect 7309 9891 7329 9911
rect 9112 9888 9132 9908
rect 822 9761 842 9781
rect 925 9765 945 9785
rect 1035 9761 1055 9781
rect 1138 9765 1158 9785
rect 1243 9761 1263 9781
rect 1346 9765 1366 9785
rect 1454 9765 1474 9785
rect 9215 9884 9235 9904
rect 9323 9884 9343 9904
rect 9426 9888 9446 9908
rect 9531 9884 9551 9904
rect 9634 9888 9654 9908
rect 9744 9884 9764 9904
rect 9847 9888 9867 9908
rect 10167 9893 10185 9911
rect 1557 9761 1577 9781
rect 1870 9757 1890 9777
rect 504 9729 522 9747
rect 1973 9761 1993 9781
rect 2083 9757 2103 9777
rect 2186 9761 2206 9781
rect 2291 9757 2311 9777
rect 2394 9761 2414 9781
rect 2502 9761 2522 9781
rect 2605 9757 2625 9777
rect 10169 9794 10187 9812
rect 11210 9822 11228 9840
rect 17282 9885 17302 9905
rect 17385 9881 17405 9901
rect 17493 9881 17513 9901
rect 17596 9885 17616 9905
rect 17701 9881 17721 9901
rect 17804 9885 17824 9905
rect 17914 9881 17934 9901
rect 18017 9885 18037 9905
rect 19820 9882 19840 9902
rect 11530 9755 11550 9775
rect 11633 9759 11653 9779
rect 11743 9755 11763 9775
rect 11846 9759 11866 9779
rect 11951 9755 11971 9775
rect 12054 9759 12074 9779
rect 12162 9759 12182 9779
rect 19923 9878 19943 9898
rect 20031 9878 20051 9898
rect 20134 9882 20154 9902
rect 20239 9878 20259 9898
rect 20342 9882 20362 9902
rect 20452 9878 20472 9898
rect 20555 9882 20575 9902
rect 20875 9887 20893 9905
rect 12265 9755 12285 9775
rect 12578 9751 12598 9771
rect 11212 9723 11230 9741
rect 12681 9755 12701 9775
rect 12791 9751 12811 9771
rect 12894 9755 12914 9775
rect 12999 9751 13019 9771
rect 13102 9755 13122 9775
rect 13210 9755 13230 9775
rect 13313 9751 13333 9771
rect 10167 9638 10185 9656
rect 20877 9788 20895 9806
rect 20875 9632 20893 9650
rect 10169 9539 10187 9557
rect 20877 9533 20895 9551
rect 502 9433 520 9451
rect 11210 9427 11228 9445
rect 504 9334 522 9352
rect 502 9178 520 9196
rect 11212 9328 11230 9346
rect 8064 9213 8084 9233
rect 8167 9209 8187 9229
rect 8275 9209 8295 9229
rect 8378 9213 8398 9233
rect 8483 9209 8503 9229
rect 8586 9213 8606 9233
rect 8696 9209 8716 9229
rect 10167 9243 10185 9261
rect 8799 9213 8819 9233
rect 9112 9209 9132 9229
rect 504 9079 522 9097
rect 822 9082 842 9102
rect 925 9086 945 9106
rect 1035 9082 1055 9102
rect 1138 9086 1158 9106
rect 1243 9082 1263 9102
rect 1346 9086 1366 9106
rect 1454 9086 1474 9106
rect 9215 9205 9235 9225
rect 9323 9205 9343 9225
rect 9426 9209 9446 9229
rect 9531 9205 9551 9225
rect 9634 9209 9654 9229
rect 9744 9205 9764 9225
rect 9847 9209 9867 9229
rect 1557 9082 1577 9102
rect 3317 9077 3337 9097
rect 3420 9081 3440 9101
rect 3530 9077 3550 9097
rect 3633 9081 3653 9101
rect 3738 9077 3758 9097
rect 3841 9081 3861 9101
rect 3949 9081 3969 9101
rect 4052 9077 4072 9097
rect 10169 9144 10187 9162
rect 11210 9172 11228 9190
rect 18772 9207 18792 9227
rect 18875 9203 18895 9223
rect 18983 9203 19003 9223
rect 19086 9207 19106 9227
rect 19191 9203 19211 9223
rect 19294 9207 19314 9227
rect 19404 9203 19424 9223
rect 20875 9237 20893 9255
rect 19507 9207 19527 9227
rect 19820 9203 19840 9223
rect 11212 9073 11230 9091
rect 11530 9076 11550 9096
rect 11633 9080 11653 9100
rect 11743 9076 11763 9096
rect 11846 9080 11866 9100
rect 11951 9076 11971 9096
rect 12054 9080 12074 9100
rect 12162 9080 12182 9100
rect 19923 9199 19943 9219
rect 20031 9199 20051 9219
rect 20134 9203 20154 9223
rect 20239 9199 20259 9219
rect 20342 9203 20362 9223
rect 20452 9199 20472 9219
rect 20555 9203 20575 9223
rect 12265 9076 12285 9096
rect 14025 9071 14045 9091
rect 14128 9075 14148 9095
rect 14238 9071 14258 9091
rect 14341 9075 14361 9095
rect 14446 9071 14466 9091
rect 14549 9075 14569 9095
rect 14657 9075 14677 9095
rect 14760 9071 14780 9091
rect 20877 9138 20895 9156
rect 10167 8987 10185 9005
rect 20875 8981 20893 8999
rect 10169 8888 10187 8906
rect 20877 8882 20895 8900
rect 502 8637 520 8655
rect 11210 8631 11228 8649
rect 504 8538 522 8556
rect 11212 8532 11230 8550
rect 502 8381 520 8399
rect 6617 8446 6637 8466
rect 6720 8442 6740 8462
rect 6828 8442 6848 8462
rect 6931 8446 6951 8466
rect 7036 8442 7056 8462
rect 7139 8446 7159 8466
rect 7249 8442 7269 8462
rect 7352 8446 7372 8466
rect 9112 8441 9132 8461
rect 822 8314 842 8334
rect 925 8318 945 8338
rect 1035 8314 1055 8334
rect 1138 8318 1158 8338
rect 1243 8314 1263 8334
rect 1346 8318 1366 8338
rect 1454 8318 1474 8338
rect 9215 8437 9235 8457
rect 9323 8437 9343 8457
rect 9426 8441 9446 8461
rect 9531 8437 9551 8457
rect 9634 8441 9654 8461
rect 9744 8437 9764 8457
rect 9847 8441 9867 8461
rect 10167 8446 10185 8464
rect 1557 8314 1577 8334
rect 1870 8310 1890 8330
rect 504 8282 522 8300
rect 1973 8314 1993 8334
rect 2083 8310 2103 8330
rect 2186 8314 2206 8334
rect 2291 8310 2311 8330
rect 2394 8314 2414 8334
rect 2502 8314 2522 8334
rect 2605 8310 2625 8330
rect 10169 8347 10187 8365
rect 11210 8375 11228 8393
rect 17325 8440 17345 8460
rect 17428 8436 17448 8456
rect 17536 8436 17556 8456
rect 17639 8440 17659 8460
rect 17744 8436 17764 8456
rect 17847 8440 17867 8460
rect 17957 8436 17977 8456
rect 18060 8440 18080 8460
rect 19820 8435 19840 8455
rect 11530 8308 11550 8328
rect 11633 8312 11653 8332
rect 11743 8308 11763 8328
rect 11846 8312 11866 8332
rect 11951 8308 11971 8328
rect 12054 8312 12074 8332
rect 12162 8312 12182 8332
rect 19923 8431 19943 8451
rect 20031 8431 20051 8451
rect 20134 8435 20154 8455
rect 20239 8431 20259 8451
rect 20342 8435 20362 8455
rect 20452 8431 20472 8451
rect 20555 8435 20575 8455
rect 20875 8440 20893 8458
rect 12265 8308 12285 8328
rect 12578 8304 12598 8324
rect 11212 8276 11230 8294
rect 12681 8308 12701 8328
rect 12791 8304 12811 8324
rect 12894 8308 12914 8328
rect 12999 8304 13019 8324
rect 13102 8308 13122 8328
rect 13210 8308 13230 8328
rect 13313 8304 13333 8324
rect 10167 8191 10185 8209
rect 20877 8341 20895 8359
rect 20875 8185 20893 8203
rect 10169 8092 10187 8110
rect 20877 8086 20895 8104
rect 502 7986 520 8004
rect 11210 7980 11228 7998
rect 504 7887 522 7905
rect 502 7731 520 7749
rect 11212 7881 11230 7899
rect 8064 7766 8084 7786
rect 8167 7762 8187 7782
rect 8275 7762 8295 7782
rect 8378 7766 8398 7786
rect 8483 7762 8503 7782
rect 8586 7766 8606 7786
rect 8696 7762 8716 7782
rect 10167 7796 10185 7814
rect 8799 7766 8819 7786
rect 9112 7762 9132 7782
rect 504 7632 522 7650
rect 822 7635 842 7655
rect 925 7639 945 7659
rect 1035 7635 1055 7655
rect 1138 7639 1158 7659
rect 1243 7635 1263 7655
rect 1346 7639 1366 7659
rect 1454 7639 1474 7659
rect 9215 7758 9235 7778
rect 9323 7758 9343 7778
rect 9426 7762 9446 7782
rect 9531 7758 9551 7778
rect 9634 7762 9654 7782
rect 9744 7758 9764 7778
rect 9847 7762 9867 7782
rect 1557 7635 1577 7655
rect 4425 7626 4445 7646
rect 4528 7630 4548 7650
rect 4638 7626 4658 7646
rect 4741 7630 4761 7650
rect 4846 7626 4866 7646
rect 4949 7630 4969 7650
rect 5057 7630 5077 7650
rect 5160 7626 5180 7646
rect 10169 7697 10187 7715
rect 11210 7725 11228 7743
rect 18772 7760 18792 7780
rect 18875 7756 18895 7776
rect 18983 7756 19003 7776
rect 19086 7760 19106 7780
rect 19191 7756 19211 7776
rect 19294 7760 19314 7780
rect 19404 7756 19424 7776
rect 20875 7790 20893 7808
rect 19507 7760 19527 7780
rect 19820 7756 19840 7776
rect 11212 7626 11230 7644
rect 11530 7629 11550 7649
rect 11633 7633 11653 7653
rect 11743 7629 11763 7649
rect 11846 7633 11866 7653
rect 11951 7629 11971 7649
rect 12054 7633 12074 7653
rect 12162 7633 12182 7653
rect 19923 7752 19943 7772
rect 20031 7752 20051 7772
rect 20134 7756 20154 7776
rect 20239 7752 20259 7772
rect 20342 7756 20362 7776
rect 20452 7752 20472 7772
rect 20555 7756 20575 7776
rect 12265 7629 12285 7649
rect 15133 7620 15153 7640
rect 15236 7624 15256 7644
rect 15346 7620 15366 7640
rect 15449 7624 15469 7644
rect 15554 7620 15574 7640
rect 15657 7624 15677 7644
rect 15765 7624 15785 7644
rect 15868 7620 15888 7640
rect 20877 7691 20895 7709
rect 10167 7540 10185 7558
rect 20875 7534 20893 7552
rect 10169 7441 10187 7459
rect 20877 7435 20895 7453
rect 499 7043 517 7061
rect 11207 7037 11225 7055
rect 501 6944 519 6962
rect 11209 6938 11227 6956
rect 499 6787 517 6805
rect 5506 6856 5526 6876
rect 5609 6852 5629 6872
rect 5717 6852 5737 6872
rect 5820 6856 5840 6876
rect 5925 6852 5945 6872
rect 6028 6856 6048 6876
rect 6138 6852 6158 6872
rect 6241 6856 6261 6876
rect 9109 6847 9129 6867
rect 819 6720 839 6740
rect 922 6724 942 6744
rect 1032 6720 1052 6740
rect 1135 6724 1155 6744
rect 1240 6720 1260 6740
rect 1343 6724 1363 6744
rect 1451 6724 1471 6744
rect 9212 6843 9232 6863
rect 9320 6843 9340 6863
rect 9423 6847 9443 6867
rect 9528 6843 9548 6863
rect 9631 6847 9651 6867
rect 9741 6843 9761 6863
rect 9844 6847 9864 6867
rect 10164 6852 10182 6870
rect 1554 6720 1574 6740
rect 1867 6716 1887 6736
rect 501 6688 519 6706
rect 1970 6720 1990 6740
rect 2080 6716 2100 6736
rect 2183 6720 2203 6740
rect 2288 6716 2308 6736
rect 2391 6720 2411 6740
rect 2499 6720 2519 6740
rect 2602 6716 2622 6736
rect 10166 6753 10184 6771
rect 11207 6781 11225 6799
rect 16214 6850 16234 6870
rect 16317 6846 16337 6866
rect 16425 6846 16445 6866
rect 16528 6850 16548 6870
rect 16633 6846 16653 6866
rect 16736 6850 16756 6870
rect 16846 6846 16866 6866
rect 16949 6850 16969 6870
rect 19817 6841 19837 6861
rect 11527 6714 11547 6734
rect 11630 6718 11650 6738
rect 11740 6714 11760 6734
rect 11843 6718 11863 6738
rect 11948 6714 11968 6734
rect 12051 6718 12071 6738
rect 12159 6718 12179 6738
rect 19920 6837 19940 6857
rect 20028 6837 20048 6857
rect 20131 6841 20151 6861
rect 20236 6837 20256 6857
rect 20339 6841 20359 6861
rect 20449 6837 20469 6857
rect 20552 6841 20572 6861
rect 20872 6846 20890 6864
rect 12262 6714 12282 6734
rect 12575 6710 12595 6730
rect 11209 6682 11227 6700
rect 12678 6714 12698 6734
rect 12788 6710 12808 6730
rect 12891 6714 12911 6734
rect 12996 6710 13016 6730
rect 13099 6714 13119 6734
rect 13207 6714 13227 6734
rect 13310 6710 13330 6730
rect 10164 6597 10182 6615
rect 20874 6747 20892 6765
rect 20872 6591 20890 6609
rect 10166 6498 10184 6516
rect 20874 6492 20892 6510
rect 499 6392 517 6410
rect 11207 6386 11225 6404
rect 501 6293 519 6311
rect 499 6137 517 6155
rect 11209 6287 11227 6305
rect 8061 6172 8081 6192
rect 8164 6168 8184 6188
rect 8272 6168 8292 6188
rect 8375 6172 8395 6192
rect 8480 6168 8500 6188
rect 8583 6172 8603 6192
rect 8693 6168 8713 6188
rect 10164 6202 10182 6220
rect 8796 6172 8816 6192
rect 9109 6168 9129 6188
rect 501 6038 519 6056
rect 819 6041 839 6061
rect 922 6045 942 6065
rect 1032 6041 1052 6061
rect 1135 6045 1155 6065
rect 1240 6041 1260 6061
rect 1343 6045 1363 6065
rect 1451 6045 1471 6065
rect 9212 6164 9232 6184
rect 9320 6164 9340 6184
rect 9423 6168 9443 6188
rect 9528 6164 9548 6184
rect 9631 6168 9651 6188
rect 9741 6164 9761 6184
rect 9844 6168 9864 6188
rect 1554 6041 1574 6061
rect 3314 6036 3334 6056
rect 3417 6040 3437 6060
rect 3527 6036 3547 6056
rect 3630 6040 3650 6060
rect 3735 6036 3755 6056
rect 3838 6040 3858 6060
rect 3946 6040 3966 6060
rect 4049 6036 4069 6056
rect 10166 6103 10184 6121
rect 11207 6131 11225 6149
rect 18769 6166 18789 6186
rect 18872 6162 18892 6182
rect 18980 6162 19000 6182
rect 19083 6166 19103 6186
rect 19188 6162 19208 6182
rect 19291 6166 19311 6186
rect 19401 6162 19421 6182
rect 20872 6196 20890 6214
rect 19504 6166 19524 6186
rect 19817 6162 19837 6182
rect 11209 6032 11227 6050
rect 11527 6035 11547 6055
rect 11630 6039 11650 6059
rect 11740 6035 11760 6055
rect 11843 6039 11863 6059
rect 11948 6035 11968 6055
rect 12051 6039 12071 6059
rect 12159 6039 12179 6059
rect 19920 6158 19940 6178
rect 20028 6158 20048 6178
rect 20131 6162 20151 6182
rect 20236 6158 20256 6178
rect 20339 6162 20359 6182
rect 20449 6158 20469 6178
rect 20552 6162 20572 6182
rect 12262 6035 12282 6055
rect 14022 6030 14042 6050
rect 14125 6034 14145 6054
rect 14235 6030 14255 6050
rect 14338 6034 14358 6054
rect 14443 6030 14463 6050
rect 14546 6034 14566 6054
rect 14654 6034 14674 6054
rect 14757 6030 14777 6050
rect 20874 6097 20892 6115
rect 10164 5946 10182 5964
rect 20872 5940 20890 5958
rect 10166 5847 10184 5865
rect 20874 5841 20892 5859
rect 499 5596 517 5614
rect 11207 5590 11225 5608
rect 501 5497 519 5515
rect 11209 5491 11227 5509
rect 499 5340 517 5358
rect 6614 5405 6634 5425
rect 6717 5401 6737 5421
rect 6825 5401 6845 5421
rect 6928 5405 6948 5425
rect 7033 5401 7053 5421
rect 7136 5405 7156 5425
rect 7246 5401 7266 5421
rect 7349 5405 7369 5425
rect 9109 5400 9129 5420
rect 819 5273 839 5293
rect 922 5277 942 5297
rect 1032 5273 1052 5293
rect 1135 5277 1155 5297
rect 1240 5273 1260 5293
rect 1343 5277 1363 5297
rect 1451 5277 1471 5297
rect 9212 5396 9232 5416
rect 9320 5396 9340 5416
rect 9423 5400 9443 5420
rect 9528 5396 9548 5416
rect 9631 5400 9651 5420
rect 9741 5396 9761 5416
rect 9844 5400 9864 5420
rect 10164 5405 10182 5423
rect 1554 5273 1574 5293
rect 1867 5269 1887 5289
rect 501 5241 519 5259
rect 1970 5273 1990 5293
rect 2080 5269 2100 5289
rect 2183 5273 2203 5293
rect 2288 5269 2308 5289
rect 2391 5273 2411 5293
rect 2499 5273 2519 5293
rect 2602 5269 2622 5289
rect 10166 5306 10184 5324
rect 11207 5334 11225 5352
rect 17322 5399 17342 5419
rect 17425 5395 17445 5415
rect 17533 5395 17553 5415
rect 17636 5399 17656 5419
rect 17741 5395 17761 5415
rect 17844 5399 17864 5419
rect 17954 5395 17974 5415
rect 18057 5399 18077 5419
rect 19817 5394 19837 5414
rect 11527 5267 11547 5287
rect 11630 5271 11650 5291
rect 11740 5267 11760 5287
rect 11843 5271 11863 5291
rect 11948 5267 11968 5287
rect 12051 5271 12071 5291
rect 12159 5271 12179 5291
rect 19920 5390 19940 5410
rect 20028 5390 20048 5410
rect 20131 5394 20151 5414
rect 20236 5390 20256 5410
rect 20339 5394 20359 5414
rect 20449 5390 20469 5410
rect 20552 5394 20572 5414
rect 20872 5399 20890 5417
rect 12262 5267 12282 5287
rect 12575 5263 12595 5283
rect 11209 5235 11227 5253
rect 12678 5267 12698 5287
rect 12788 5263 12808 5283
rect 12891 5267 12911 5287
rect 12996 5263 13016 5283
rect 13099 5267 13119 5287
rect 13207 5267 13227 5287
rect 13310 5263 13330 5283
rect 10164 5150 10182 5168
rect 20874 5300 20892 5318
rect 20872 5144 20890 5162
rect 10166 5051 10184 5069
rect 20874 5045 20892 5063
rect 499 4945 517 4963
rect 11207 4939 11225 4957
rect 501 4846 519 4864
rect 499 4690 517 4708
rect 11209 4840 11227 4858
rect 8061 4725 8081 4745
rect 8164 4721 8184 4741
rect 8272 4721 8292 4741
rect 8375 4725 8395 4745
rect 8480 4721 8500 4741
rect 8583 4725 8603 4745
rect 8693 4721 8713 4741
rect 10164 4755 10182 4773
rect 8796 4725 8816 4745
rect 9109 4721 9129 4741
rect 501 4591 519 4609
rect 819 4594 839 4614
rect 922 4598 942 4618
rect 1032 4594 1052 4614
rect 1135 4598 1155 4618
rect 1240 4594 1260 4614
rect 1343 4598 1363 4618
rect 1451 4598 1471 4618
rect 9212 4717 9232 4737
rect 9320 4717 9340 4737
rect 9423 4721 9443 4741
rect 9528 4717 9548 4737
rect 9631 4721 9651 4741
rect 9741 4717 9761 4737
rect 9844 4721 9864 4741
rect 1554 4594 1574 4614
rect 3357 4591 3377 4611
rect 3460 4595 3480 4615
rect 3570 4591 3590 4611
rect 3673 4595 3693 4615
rect 3778 4591 3798 4611
rect 3881 4595 3901 4615
rect 3989 4595 4009 4615
rect 4092 4591 4112 4611
rect 10166 4656 10184 4674
rect 11207 4684 11225 4702
rect 18769 4719 18789 4739
rect 18872 4715 18892 4735
rect 18980 4715 19000 4735
rect 19083 4719 19103 4739
rect 19188 4715 19208 4735
rect 19291 4719 19311 4739
rect 19401 4715 19421 4735
rect 20872 4749 20890 4767
rect 19504 4719 19524 4739
rect 19817 4715 19837 4735
rect 11209 4585 11227 4603
rect 11527 4588 11547 4608
rect 11630 4592 11650 4612
rect 11740 4588 11760 4608
rect 11843 4592 11863 4612
rect 11948 4588 11968 4608
rect 12051 4592 12071 4612
rect 12159 4592 12179 4612
rect 19920 4711 19940 4731
rect 20028 4711 20048 4731
rect 20131 4715 20151 4735
rect 20236 4711 20256 4731
rect 20339 4715 20359 4735
rect 20449 4711 20469 4731
rect 20552 4715 20572 4735
rect 12262 4588 12282 4608
rect 14065 4585 14085 4605
rect 14168 4589 14188 4609
rect 14278 4585 14298 4605
rect 14381 4589 14401 4609
rect 14486 4585 14506 4605
rect 14589 4589 14609 4609
rect 14697 4589 14717 4609
rect 14800 4585 14820 4605
rect 20874 4650 20892 4668
rect 10164 4499 10182 4517
rect 20872 4493 20890 4511
rect 10166 4400 10184 4418
rect 20874 4394 20892 4412
rect 500 4076 518 4094
rect 11208 4070 11226 4088
rect 502 3977 520 3995
rect 500 3820 518 3838
rect 11210 3971 11228 3989
rect 6572 3883 6592 3903
rect 6675 3879 6695 3899
rect 6783 3879 6803 3899
rect 6886 3883 6906 3903
rect 6991 3879 7011 3899
rect 7094 3883 7114 3903
rect 7204 3879 7224 3899
rect 7307 3883 7327 3903
rect 9110 3880 9130 3900
rect 820 3753 840 3773
rect 923 3757 943 3777
rect 1033 3753 1053 3773
rect 1136 3757 1156 3777
rect 1241 3753 1261 3773
rect 1344 3757 1364 3777
rect 1452 3757 1472 3777
rect 9213 3876 9233 3896
rect 9321 3876 9341 3896
rect 9424 3880 9444 3900
rect 9529 3876 9549 3896
rect 9632 3880 9652 3900
rect 9742 3876 9762 3896
rect 9845 3880 9865 3900
rect 10165 3885 10183 3903
rect 1555 3753 1575 3773
rect 1868 3749 1888 3769
rect 502 3721 520 3739
rect 1971 3753 1991 3773
rect 2081 3749 2101 3769
rect 2184 3753 2204 3773
rect 2289 3749 2309 3769
rect 2392 3753 2412 3773
rect 2500 3753 2520 3773
rect 2603 3749 2623 3769
rect 4770 3755 4790 3775
rect 4873 3759 4893 3779
rect 4983 3755 5003 3775
rect 5086 3759 5106 3779
rect 5191 3755 5211 3775
rect 5294 3759 5314 3779
rect 5402 3759 5422 3779
rect 5505 3755 5525 3775
rect 10167 3786 10185 3804
rect 11208 3814 11226 3832
rect 17280 3877 17300 3897
rect 17383 3873 17403 3893
rect 17491 3873 17511 3893
rect 17594 3877 17614 3897
rect 17699 3873 17719 3893
rect 17802 3877 17822 3897
rect 17912 3873 17932 3893
rect 18015 3877 18035 3897
rect 19818 3874 19838 3894
rect 11528 3747 11548 3767
rect 11631 3751 11651 3771
rect 11741 3747 11761 3767
rect 11844 3751 11864 3771
rect 11949 3747 11969 3767
rect 12052 3751 12072 3771
rect 12160 3751 12180 3771
rect 19921 3870 19941 3890
rect 20029 3870 20049 3890
rect 20132 3874 20152 3894
rect 20237 3870 20257 3890
rect 20340 3874 20360 3894
rect 20450 3870 20470 3890
rect 20553 3874 20573 3894
rect 20873 3879 20891 3897
rect 12263 3747 12283 3767
rect 12576 3743 12596 3763
rect 11210 3715 11228 3733
rect 12679 3747 12699 3767
rect 12789 3743 12809 3763
rect 12892 3747 12912 3767
rect 12997 3743 13017 3763
rect 13100 3747 13120 3767
rect 13208 3747 13228 3767
rect 13311 3743 13331 3763
rect 15478 3749 15498 3769
rect 15581 3753 15601 3773
rect 15691 3749 15711 3769
rect 15794 3753 15814 3773
rect 15899 3749 15919 3769
rect 16002 3753 16022 3773
rect 16110 3753 16130 3773
rect 16213 3749 16233 3769
rect 10165 3630 10183 3648
rect 20875 3780 20893 3798
rect 20873 3624 20891 3642
rect 10167 3531 10185 3549
rect 20875 3525 20893 3543
rect 500 3425 518 3443
rect 11208 3419 11226 3437
rect 502 3326 520 3344
rect 500 3170 518 3188
rect 11210 3320 11228 3338
rect 8062 3205 8082 3225
rect 8165 3201 8185 3221
rect 8273 3201 8293 3221
rect 8376 3205 8396 3225
rect 8481 3201 8501 3221
rect 8584 3205 8604 3225
rect 8694 3201 8714 3221
rect 10165 3235 10183 3253
rect 8797 3205 8817 3225
rect 9110 3201 9130 3221
rect 502 3071 520 3089
rect 820 3074 840 3094
rect 923 3078 943 3098
rect 1033 3074 1053 3094
rect 1136 3078 1156 3098
rect 1241 3074 1261 3094
rect 1344 3078 1364 3098
rect 1452 3078 1472 3098
rect 9213 3197 9233 3217
rect 9321 3197 9341 3217
rect 9424 3201 9444 3221
rect 9529 3197 9549 3217
rect 9632 3201 9652 3221
rect 9742 3197 9762 3217
rect 9845 3201 9865 3221
rect 1555 3074 1575 3094
rect 3315 3069 3335 3089
rect 3418 3073 3438 3093
rect 3528 3069 3548 3089
rect 3631 3073 3651 3093
rect 3736 3069 3756 3089
rect 3839 3073 3859 3093
rect 3947 3073 3967 3093
rect 4050 3069 4070 3089
rect 10167 3136 10185 3154
rect 11208 3164 11226 3182
rect 18770 3199 18790 3219
rect 18873 3195 18893 3215
rect 18981 3195 19001 3215
rect 19084 3199 19104 3219
rect 19189 3195 19209 3215
rect 19292 3199 19312 3219
rect 19402 3195 19422 3215
rect 20873 3229 20891 3247
rect 19505 3199 19525 3219
rect 19818 3195 19838 3215
rect 11210 3065 11228 3083
rect 11528 3068 11548 3088
rect 11631 3072 11651 3092
rect 11741 3068 11761 3088
rect 11844 3072 11864 3092
rect 11949 3068 11969 3088
rect 12052 3072 12072 3092
rect 12160 3072 12180 3092
rect 19921 3191 19941 3211
rect 20029 3191 20049 3211
rect 20132 3195 20152 3215
rect 20237 3191 20257 3211
rect 20340 3195 20360 3215
rect 20450 3191 20470 3211
rect 20553 3195 20573 3215
rect 12263 3068 12283 3088
rect 14023 3063 14043 3083
rect 14126 3067 14146 3087
rect 14236 3063 14256 3083
rect 14339 3067 14359 3087
rect 14444 3063 14464 3083
rect 14547 3067 14567 3087
rect 14655 3067 14675 3087
rect 14758 3063 14778 3083
rect 20875 3130 20893 3148
rect 10165 2979 10183 2997
rect 20873 2973 20891 2991
rect 10167 2880 10185 2898
rect 20875 2874 20893 2892
rect 500 2629 518 2647
rect 11208 2623 11226 2641
rect 502 2530 520 2548
rect 11210 2524 11228 2542
rect 500 2373 518 2391
rect 6615 2438 6635 2458
rect 6718 2434 6738 2454
rect 6826 2434 6846 2454
rect 6929 2438 6949 2458
rect 7034 2434 7054 2454
rect 7137 2438 7157 2458
rect 7247 2434 7267 2454
rect 7350 2438 7370 2458
rect 9110 2433 9130 2453
rect 820 2306 840 2326
rect 923 2310 943 2330
rect 1033 2306 1053 2326
rect 1136 2310 1156 2330
rect 1241 2306 1261 2326
rect 1344 2310 1364 2330
rect 1452 2310 1472 2330
rect 9213 2429 9233 2449
rect 9321 2429 9341 2449
rect 9424 2433 9444 2453
rect 9529 2429 9549 2449
rect 9632 2433 9652 2453
rect 9742 2429 9762 2449
rect 9845 2433 9865 2453
rect 10165 2438 10183 2456
rect 1555 2306 1575 2326
rect 1868 2302 1888 2322
rect 502 2274 520 2292
rect 1971 2306 1991 2326
rect 2081 2302 2101 2322
rect 2184 2306 2204 2326
rect 2289 2302 2309 2322
rect 2392 2306 2412 2326
rect 2500 2306 2520 2326
rect 2603 2302 2623 2322
rect 10167 2339 10185 2357
rect 11208 2367 11226 2385
rect 17323 2432 17343 2452
rect 17426 2428 17446 2448
rect 17534 2428 17554 2448
rect 17637 2432 17657 2452
rect 17742 2428 17762 2448
rect 17845 2432 17865 2452
rect 17955 2428 17975 2448
rect 18058 2432 18078 2452
rect 19818 2427 19838 2447
rect 11528 2300 11548 2320
rect 11631 2304 11651 2324
rect 11741 2300 11761 2320
rect 11844 2304 11864 2324
rect 11949 2300 11969 2320
rect 12052 2304 12072 2324
rect 12160 2304 12180 2324
rect 19921 2423 19941 2443
rect 20029 2423 20049 2443
rect 20132 2427 20152 2447
rect 20237 2423 20257 2443
rect 20340 2427 20360 2447
rect 20450 2423 20470 2443
rect 20553 2427 20573 2447
rect 20873 2432 20891 2450
rect 12263 2300 12283 2320
rect 12576 2296 12596 2316
rect 11210 2268 11228 2286
rect 12679 2300 12699 2320
rect 12789 2296 12809 2316
rect 12892 2300 12912 2320
rect 12997 2296 13017 2316
rect 13100 2300 13120 2320
rect 13208 2300 13228 2320
rect 13311 2296 13331 2316
rect 10165 2183 10183 2201
rect 20875 2333 20893 2351
rect 20873 2177 20891 2195
rect 10167 2084 10185 2102
rect 20875 2078 20893 2096
rect 500 1978 518 1996
rect 11208 1972 11226 1990
rect 502 1879 520 1897
rect 500 1723 518 1741
rect 11210 1873 11228 1891
rect 8062 1758 8082 1778
rect 8165 1754 8185 1774
rect 8273 1754 8293 1774
rect 8376 1758 8396 1778
rect 8481 1754 8501 1774
rect 8584 1758 8604 1778
rect 8694 1754 8714 1774
rect 10165 1788 10183 1806
rect 8797 1758 8817 1778
rect 9110 1754 9130 1774
rect 9213 1750 9233 1770
rect 9321 1750 9341 1770
rect 9424 1754 9444 1774
rect 9529 1750 9549 1770
rect 9632 1754 9652 1774
rect 9742 1750 9762 1770
rect 9845 1754 9865 1774
rect 502 1624 520 1642
rect 820 1627 840 1647
rect 923 1631 943 1651
rect 1033 1627 1053 1647
rect 1136 1631 1156 1651
rect 1241 1627 1261 1647
rect 1344 1631 1364 1651
rect 1452 1631 1472 1651
rect 1555 1627 1575 1647
rect 10167 1689 10185 1707
rect 11208 1717 11226 1735
rect 18770 1752 18790 1772
rect 18873 1748 18893 1768
rect 18981 1748 19001 1768
rect 19084 1752 19104 1772
rect 19189 1748 19209 1768
rect 19292 1752 19312 1772
rect 19402 1748 19422 1768
rect 20873 1782 20891 1800
rect 19505 1752 19525 1772
rect 19818 1748 19838 1768
rect 19921 1744 19941 1764
rect 20029 1744 20049 1764
rect 20132 1748 20152 1768
rect 20237 1744 20257 1764
rect 20340 1748 20360 1768
rect 20450 1744 20470 1764
rect 20553 1748 20573 1768
rect 11210 1618 11228 1636
rect 11528 1621 11548 1641
rect 11631 1625 11651 1645
rect 11741 1621 11761 1641
rect 11844 1625 11864 1645
rect 11949 1621 11969 1641
rect 12052 1625 12072 1645
rect 12160 1625 12180 1645
rect 12263 1621 12283 1641
rect 20875 1683 20893 1701
rect 10165 1532 10183 1550
rect 20873 1526 20891 1544
rect 10167 1433 10185 1451
rect 20875 1427 20893 1445
rect 10531 -532 10551 -512
rect 10634 -528 10654 -508
rect 10744 -532 10764 -512
rect 10847 -528 10867 -508
rect 10952 -532 10972 -512
rect 11055 -528 11075 -508
rect 11163 -528 11183 -508
rect 11266 -532 11286 -512
<< pdiffc >>
rect 827 12877 847 12897
rect 923 12877 943 12897
rect 1040 12877 1060 12897
rect 1136 12877 1156 12897
rect 1248 12877 1268 12897
rect 1344 12877 1364 12897
rect 1454 12877 1474 12897
rect 1550 12877 1570 12897
rect 1875 12873 1895 12893
rect 1971 12873 1991 12893
rect 2088 12873 2108 12893
rect 2184 12873 2204 12893
rect 2296 12873 2316 12893
rect 2392 12873 2412 12893
rect 2502 12873 2522 12893
rect 2598 12873 2618 12893
rect 11535 12871 11555 12891
rect 11631 12871 11651 12891
rect 11748 12871 11768 12891
rect 11844 12871 11864 12891
rect 11956 12871 11976 12891
rect 12052 12871 12072 12891
rect 12162 12871 12182 12891
rect 12258 12871 12278 12891
rect 12583 12867 12603 12887
rect 9117 12706 9137 12726
rect 9213 12706 9233 12726
rect 9323 12706 9343 12726
rect 9419 12706 9439 12726
rect 9531 12706 9551 12726
rect 9627 12706 9647 12726
rect 9744 12706 9764 12726
rect 12679 12867 12699 12887
rect 12796 12867 12816 12887
rect 12892 12867 12912 12887
rect 13004 12867 13024 12887
rect 13100 12867 13120 12887
rect 13210 12867 13230 12887
rect 13306 12867 13326 12887
rect 9840 12706 9860 12726
rect 19825 12700 19845 12720
rect 19921 12700 19941 12720
rect 20031 12700 20051 12720
rect 20127 12700 20147 12720
rect 20239 12700 20259 12720
rect 20335 12700 20355 12720
rect 20452 12700 20472 12720
rect 20548 12700 20568 12720
rect 827 12198 847 12218
rect 923 12198 943 12218
rect 1040 12198 1060 12218
rect 1136 12198 1156 12218
rect 1248 12198 1268 12218
rect 1344 12198 1364 12218
rect 1454 12198 1474 12218
rect 1550 12198 1570 12218
rect 3322 12193 3342 12213
rect 3418 12193 3438 12213
rect 3535 12193 3555 12213
rect 3631 12193 3651 12213
rect 3743 12193 3763 12213
rect 3839 12193 3859 12213
rect 3949 12193 3969 12213
rect 4045 12193 4065 12213
rect 11535 12192 11555 12212
rect 8069 12031 8089 12051
rect 8165 12031 8185 12051
rect 8275 12031 8295 12051
rect 8371 12031 8391 12051
rect 8483 12031 8503 12051
rect 8579 12031 8599 12051
rect 8696 12031 8716 12051
rect 11631 12192 11651 12212
rect 11748 12192 11768 12212
rect 11844 12192 11864 12212
rect 11956 12192 11976 12212
rect 12052 12192 12072 12212
rect 12162 12192 12182 12212
rect 12258 12192 12278 12212
rect 14030 12187 14050 12207
rect 8792 12031 8812 12051
rect 9117 12027 9137 12047
rect 9213 12027 9233 12047
rect 9323 12027 9343 12047
rect 9419 12027 9439 12047
rect 9531 12027 9551 12047
rect 9627 12027 9647 12047
rect 9744 12027 9764 12047
rect 9840 12027 9860 12047
rect 14126 12187 14146 12207
rect 14243 12187 14263 12207
rect 14339 12187 14359 12207
rect 14451 12187 14471 12207
rect 14547 12187 14567 12207
rect 14657 12187 14677 12207
rect 14753 12187 14773 12207
rect 18777 12025 18797 12045
rect 18873 12025 18893 12045
rect 18983 12025 19003 12045
rect 19079 12025 19099 12045
rect 19191 12025 19211 12045
rect 19287 12025 19307 12045
rect 19404 12025 19424 12045
rect 19500 12025 19520 12045
rect 19825 12021 19845 12041
rect 19921 12021 19941 12041
rect 20031 12021 20051 12041
rect 20127 12021 20147 12041
rect 20239 12021 20259 12041
rect 20335 12021 20355 12041
rect 20452 12021 20472 12041
rect 20548 12021 20568 12041
rect 827 11430 847 11450
rect 923 11430 943 11450
rect 1040 11430 1060 11450
rect 1136 11430 1156 11450
rect 1248 11430 1268 11450
rect 1344 11430 1364 11450
rect 1454 11430 1474 11450
rect 1550 11430 1570 11450
rect 1875 11426 1895 11446
rect 1971 11426 1991 11446
rect 2088 11426 2108 11446
rect 2184 11426 2204 11446
rect 2296 11426 2316 11446
rect 2392 11426 2412 11446
rect 2502 11426 2522 11446
rect 2598 11426 2618 11446
rect 6622 11264 6642 11284
rect 6718 11264 6738 11284
rect 6828 11264 6848 11284
rect 6924 11264 6944 11284
rect 7036 11264 7056 11284
rect 7132 11264 7152 11284
rect 7249 11264 7269 11284
rect 11535 11424 11555 11444
rect 11631 11424 11651 11444
rect 11748 11424 11768 11444
rect 11844 11424 11864 11444
rect 11956 11424 11976 11444
rect 12052 11424 12072 11444
rect 12162 11424 12182 11444
rect 12258 11424 12278 11444
rect 12583 11420 12603 11440
rect 7345 11264 7365 11284
rect 9117 11259 9137 11279
rect 9213 11259 9233 11279
rect 9323 11259 9343 11279
rect 9419 11259 9439 11279
rect 9531 11259 9551 11279
rect 9627 11259 9647 11279
rect 9744 11259 9764 11279
rect 12679 11420 12699 11440
rect 12796 11420 12816 11440
rect 12892 11420 12912 11440
rect 13004 11420 13024 11440
rect 13100 11420 13120 11440
rect 13210 11420 13230 11440
rect 13306 11420 13326 11440
rect 9840 11259 9860 11279
rect 17330 11258 17350 11278
rect 17426 11258 17446 11278
rect 17536 11258 17556 11278
rect 17632 11258 17652 11278
rect 17744 11258 17764 11278
rect 17840 11258 17860 11278
rect 17957 11258 17977 11278
rect 18053 11258 18073 11278
rect 19825 11253 19845 11273
rect 19921 11253 19941 11273
rect 20031 11253 20051 11273
rect 20127 11253 20147 11273
rect 20239 11253 20259 11273
rect 20335 11253 20355 11273
rect 20452 11253 20472 11273
rect 20548 11253 20568 11273
rect 827 10751 847 10771
rect 923 10751 943 10771
rect 1040 10751 1060 10771
rect 1136 10751 1156 10771
rect 1248 10751 1268 10771
rect 1344 10751 1364 10771
rect 1454 10751 1474 10771
rect 1550 10751 1570 10771
rect 3365 10748 3385 10768
rect 3461 10748 3481 10768
rect 3578 10748 3598 10768
rect 3674 10748 3694 10768
rect 3786 10748 3806 10768
rect 3882 10748 3902 10768
rect 3992 10748 4012 10768
rect 4088 10748 4108 10768
rect 11535 10745 11555 10765
rect 8069 10584 8089 10604
rect 8165 10584 8185 10604
rect 8275 10584 8295 10604
rect 8371 10584 8391 10604
rect 8483 10584 8503 10604
rect 8579 10584 8599 10604
rect 8696 10584 8716 10604
rect 11631 10745 11651 10765
rect 11748 10745 11768 10765
rect 11844 10745 11864 10765
rect 11956 10745 11976 10765
rect 12052 10745 12072 10765
rect 12162 10745 12182 10765
rect 12258 10745 12278 10765
rect 14073 10742 14093 10762
rect 8792 10584 8812 10604
rect 9117 10580 9137 10600
rect 9213 10580 9233 10600
rect 9323 10580 9343 10600
rect 9419 10580 9439 10600
rect 9531 10580 9551 10600
rect 9627 10580 9647 10600
rect 9744 10580 9764 10600
rect 9840 10580 9860 10600
rect 14169 10742 14189 10762
rect 14286 10742 14306 10762
rect 14382 10742 14402 10762
rect 14494 10742 14514 10762
rect 14590 10742 14610 10762
rect 14700 10742 14720 10762
rect 14796 10742 14816 10762
rect 18777 10578 18797 10598
rect 18873 10578 18893 10598
rect 18983 10578 19003 10598
rect 19079 10578 19099 10598
rect 19191 10578 19211 10598
rect 19287 10578 19307 10598
rect 19404 10578 19424 10598
rect 19500 10578 19520 10598
rect 19825 10574 19845 10594
rect 19921 10574 19941 10594
rect 20031 10574 20051 10594
rect 20127 10574 20147 10594
rect 20239 10574 20259 10594
rect 20335 10574 20355 10594
rect 20452 10574 20472 10594
rect 20548 10574 20568 10594
rect 828 9910 848 9930
rect 924 9910 944 9930
rect 1041 9910 1061 9930
rect 1137 9910 1157 9930
rect 1249 9910 1269 9930
rect 1345 9910 1365 9930
rect 1455 9910 1475 9930
rect 1551 9910 1571 9930
rect 1876 9906 1896 9926
rect 1972 9906 1992 9926
rect 2089 9906 2109 9926
rect 2185 9906 2205 9926
rect 2297 9906 2317 9926
rect 2393 9906 2413 9926
rect 2503 9906 2523 9926
rect 2599 9906 2619 9926
rect 6580 9742 6600 9762
rect 6676 9742 6696 9762
rect 6786 9742 6806 9762
rect 6882 9742 6902 9762
rect 6994 9742 7014 9762
rect 7090 9742 7110 9762
rect 7207 9742 7227 9762
rect 11536 9904 11556 9924
rect 11632 9904 11652 9924
rect 11749 9904 11769 9924
rect 11845 9904 11865 9924
rect 11957 9904 11977 9924
rect 12053 9904 12073 9924
rect 12163 9904 12183 9924
rect 12259 9904 12279 9924
rect 12584 9900 12604 9920
rect 7303 9742 7323 9762
rect 9118 9739 9138 9759
rect 9214 9739 9234 9759
rect 9324 9739 9344 9759
rect 9420 9739 9440 9759
rect 9532 9739 9552 9759
rect 9628 9739 9648 9759
rect 9745 9739 9765 9759
rect 12680 9900 12700 9920
rect 12797 9900 12817 9920
rect 12893 9900 12913 9920
rect 13005 9900 13025 9920
rect 13101 9900 13121 9920
rect 13211 9900 13231 9920
rect 13307 9900 13327 9920
rect 9841 9739 9861 9759
rect 17288 9736 17308 9756
rect 17384 9736 17404 9756
rect 17494 9736 17514 9756
rect 17590 9736 17610 9756
rect 17702 9736 17722 9756
rect 17798 9736 17818 9756
rect 17915 9736 17935 9756
rect 18011 9736 18031 9756
rect 19826 9733 19846 9753
rect 19922 9733 19942 9753
rect 20032 9733 20052 9753
rect 20128 9733 20148 9753
rect 20240 9733 20260 9753
rect 20336 9733 20356 9753
rect 20453 9733 20473 9753
rect 20549 9733 20569 9753
rect 828 9231 848 9251
rect 924 9231 944 9251
rect 1041 9231 1061 9251
rect 1137 9231 1157 9251
rect 1249 9231 1269 9251
rect 1345 9231 1365 9251
rect 1455 9231 1475 9251
rect 1551 9231 1571 9251
rect 3323 9226 3343 9246
rect 3419 9226 3439 9246
rect 3536 9226 3556 9246
rect 3632 9226 3652 9246
rect 3744 9226 3764 9246
rect 3840 9226 3860 9246
rect 3950 9226 3970 9246
rect 4046 9226 4066 9246
rect 11536 9225 11556 9245
rect 8070 9064 8090 9084
rect 8166 9064 8186 9084
rect 8276 9064 8296 9084
rect 8372 9064 8392 9084
rect 8484 9064 8504 9084
rect 8580 9064 8600 9084
rect 8697 9064 8717 9084
rect 11632 9225 11652 9245
rect 11749 9225 11769 9245
rect 11845 9225 11865 9245
rect 11957 9225 11977 9245
rect 12053 9225 12073 9245
rect 12163 9225 12183 9245
rect 12259 9225 12279 9245
rect 14031 9220 14051 9240
rect 8793 9064 8813 9084
rect 9118 9060 9138 9080
rect 9214 9060 9234 9080
rect 9324 9060 9344 9080
rect 9420 9060 9440 9080
rect 9532 9060 9552 9080
rect 9628 9060 9648 9080
rect 9745 9060 9765 9080
rect 9841 9060 9861 9080
rect 14127 9220 14147 9240
rect 14244 9220 14264 9240
rect 14340 9220 14360 9240
rect 14452 9220 14472 9240
rect 14548 9220 14568 9240
rect 14658 9220 14678 9240
rect 14754 9220 14774 9240
rect 18778 9058 18798 9078
rect 18874 9058 18894 9078
rect 18984 9058 19004 9078
rect 19080 9058 19100 9078
rect 19192 9058 19212 9078
rect 19288 9058 19308 9078
rect 19405 9058 19425 9078
rect 19501 9058 19521 9078
rect 19826 9054 19846 9074
rect 19922 9054 19942 9074
rect 20032 9054 20052 9074
rect 20128 9054 20148 9074
rect 20240 9054 20260 9074
rect 20336 9054 20356 9074
rect 20453 9054 20473 9074
rect 20549 9054 20569 9074
rect 828 8463 848 8483
rect 924 8463 944 8483
rect 1041 8463 1061 8483
rect 1137 8463 1157 8483
rect 1249 8463 1269 8483
rect 1345 8463 1365 8483
rect 1455 8463 1475 8483
rect 1551 8463 1571 8483
rect 1876 8459 1896 8479
rect 1972 8459 1992 8479
rect 2089 8459 2109 8479
rect 2185 8459 2205 8479
rect 2297 8459 2317 8479
rect 2393 8459 2413 8479
rect 2503 8459 2523 8479
rect 2599 8459 2619 8479
rect 6623 8297 6643 8317
rect 6719 8297 6739 8317
rect 6829 8297 6849 8317
rect 6925 8297 6945 8317
rect 7037 8297 7057 8317
rect 7133 8297 7153 8317
rect 7250 8297 7270 8317
rect 11536 8457 11556 8477
rect 11632 8457 11652 8477
rect 11749 8457 11769 8477
rect 11845 8457 11865 8477
rect 11957 8457 11977 8477
rect 12053 8457 12073 8477
rect 12163 8457 12183 8477
rect 12259 8457 12279 8477
rect 12584 8453 12604 8473
rect 7346 8297 7366 8317
rect 9118 8292 9138 8312
rect 9214 8292 9234 8312
rect 9324 8292 9344 8312
rect 9420 8292 9440 8312
rect 9532 8292 9552 8312
rect 9628 8292 9648 8312
rect 9745 8292 9765 8312
rect 12680 8453 12700 8473
rect 12797 8453 12817 8473
rect 12893 8453 12913 8473
rect 13005 8453 13025 8473
rect 13101 8453 13121 8473
rect 13211 8453 13231 8473
rect 13307 8453 13327 8473
rect 9841 8292 9861 8312
rect 17331 8291 17351 8311
rect 17427 8291 17447 8311
rect 17537 8291 17557 8311
rect 17633 8291 17653 8311
rect 17745 8291 17765 8311
rect 17841 8291 17861 8311
rect 17958 8291 17978 8311
rect 18054 8291 18074 8311
rect 19826 8286 19846 8306
rect 19922 8286 19942 8306
rect 20032 8286 20052 8306
rect 20128 8286 20148 8306
rect 20240 8286 20260 8306
rect 20336 8286 20356 8306
rect 20453 8286 20473 8306
rect 20549 8286 20569 8306
rect 828 7784 848 7804
rect 924 7784 944 7804
rect 1041 7784 1061 7804
rect 1137 7784 1157 7804
rect 1249 7784 1269 7804
rect 1345 7784 1365 7804
rect 1455 7784 1475 7804
rect 1551 7784 1571 7804
rect 4431 7775 4451 7795
rect 4527 7775 4547 7795
rect 4644 7775 4664 7795
rect 4740 7775 4760 7795
rect 4852 7775 4872 7795
rect 4948 7775 4968 7795
rect 5058 7775 5078 7795
rect 5154 7775 5174 7795
rect 11536 7778 11556 7798
rect 8070 7617 8090 7637
rect 8166 7617 8186 7637
rect 8276 7617 8296 7637
rect 8372 7617 8392 7637
rect 8484 7617 8504 7637
rect 8580 7617 8600 7637
rect 8697 7617 8717 7637
rect 11632 7778 11652 7798
rect 11749 7778 11769 7798
rect 11845 7778 11865 7798
rect 11957 7778 11977 7798
rect 12053 7778 12073 7798
rect 12163 7778 12183 7798
rect 12259 7778 12279 7798
rect 15139 7769 15159 7789
rect 8793 7617 8813 7637
rect 9118 7613 9138 7633
rect 9214 7613 9234 7633
rect 9324 7613 9344 7633
rect 9420 7613 9440 7633
rect 9532 7613 9552 7633
rect 9628 7613 9648 7633
rect 9745 7613 9765 7633
rect 9841 7613 9861 7633
rect 15235 7769 15255 7789
rect 15352 7769 15372 7789
rect 15448 7769 15468 7789
rect 15560 7769 15580 7789
rect 15656 7769 15676 7789
rect 15766 7769 15786 7789
rect 15862 7769 15882 7789
rect 18778 7611 18798 7631
rect 18874 7611 18894 7631
rect 18984 7611 19004 7631
rect 19080 7611 19100 7631
rect 19192 7611 19212 7631
rect 19288 7611 19308 7631
rect 19405 7611 19425 7631
rect 19501 7611 19521 7631
rect 19826 7607 19846 7627
rect 19922 7607 19942 7627
rect 20032 7607 20052 7627
rect 20128 7607 20148 7627
rect 20240 7607 20260 7627
rect 20336 7607 20356 7627
rect 20453 7607 20473 7627
rect 20549 7607 20569 7627
rect 825 6869 845 6889
rect 921 6869 941 6889
rect 1038 6869 1058 6889
rect 1134 6869 1154 6889
rect 1246 6869 1266 6889
rect 1342 6869 1362 6889
rect 1452 6869 1472 6889
rect 1548 6869 1568 6889
rect 1873 6865 1893 6885
rect 1969 6865 1989 6885
rect 2086 6865 2106 6885
rect 2182 6865 2202 6885
rect 2294 6865 2314 6885
rect 2390 6865 2410 6885
rect 2500 6865 2520 6885
rect 2596 6865 2616 6885
rect 5512 6707 5532 6727
rect 5608 6707 5628 6727
rect 5718 6707 5738 6727
rect 5814 6707 5834 6727
rect 5926 6707 5946 6727
rect 6022 6707 6042 6727
rect 6139 6707 6159 6727
rect 11533 6863 11553 6883
rect 11629 6863 11649 6883
rect 11746 6863 11766 6883
rect 11842 6863 11862 6883
rect 11954 6863 11974 6883
rect 12050 6863 12070 6883
rect 12160 6863 12180 6883
rect 12256 6863 12276 6883
rect 12581 6859 12601 6879
rect 6235 6707 6255 6727
rect 9115 6698 9135 6718
rect 9211 6698 9231 6718
rect 9321 6698 9341 6718
rect 9417 6698 9437 6718
rect 9529 6698 9549 6718
rect 9625 6698 9645 6718
rect 9742 6698 9762 6718
rect 12677 6859 12697 6879
rect 12794 6859 12814 6879
rect 12890 6859 12910 6879
rect 13002 6859 13022 6879
rect 13098 6859 13118 6879
rect 13208 6859 13228 6879
rect 13304 6859 13324 6879
rect 9838 6698 9858 6718
rect 16220 6701 16240 6721
rect 16316 6701 16336 6721
rect 16426 6701 16446 6721
rect 16522 6701 16542 6721
rect 16634 6701 16654 6721
rect 16730 6701 16750 6721
rect 16847 6701 16867 6721
rect 16943 6701 16963 6721
rect 19823 6692 19843 6712
rect 19919 6692 19939 6712
rect 20029 6692 20049 6712
rect 20125 6692 20145 6712
rect 20237 6692 20257 6712
rect 20333 6692 20353 6712
rect 20450 6692 20470 6712
rect 20546 6692 20566 6712
rect 825 6190 845 6210
rect 921 6190 941 6210
rect 1038 6190 1058 6210
rect 1134 6190 1154 6210
rect 1246 6190 1266 6210
rect 1342 6190 1362 6210
rect 1452 6190 1472 6210
rect 1548 6190 1568 6210
rect 3320 6185 3340 6205
rect 3416 6185 3436 6205
rect 3533 6185 3553 6205
rect 3629 6185 3649 6205
rect 3741 6185 3761 6205
rect 3837 6185 3857 6205
rect 3947 6185 3967 6205
rect 4043 6185 4063 6205
rect 11533 6184 11553 6204
rect 8067 6023 8087 6043
rect 8163 6023 8183 6043
rect 8273 6023 8293 6043
rect 8369 6023 8389 6043
rect 8481 6023 8501 6043
rect 8577 6023 8597 6043
rect 8694 6023 8714 6043
rect 11629 6184 11649 6204
rect 11746 6184 11766 6204
rect 11842 6184 11862 6204
rect 11954 6184 11974 6204
rect 12050 6184 12070 6204
rect 12160 6184 12180 6204
rect 12256 6184 12276 6204
rect 14028 6179 14048 6199
rect 8790 6023 8810 6043
rect 9115 6019 9135 6039
rect 9211 6019 9231 6039
rect 9321 6019 9341 6039
rect 9417 6019 9437 6039
rect 9529 6019 9549 6039
rect 9625 6019 9645 6039
rect 9742 6019 9762 6039
rect 9838 6019 9858 6039
rect 14124 6179 14144 6199
rect 14241 6179 14261 6199
rect 14337 6179 14357 6199
rect 14449 6179 14469 6199
rect 14545 6179 14565 6199
rect 14655 6179 14675 6199
rect 14751 6179 14771 6199
rect 18775 6017 18795 6037
rect 18871 6017 18891 6037
rect 18981 6017 19001 6037
rect 19077 6017 19097 6037
rect 19189 6017 19209 6037
rect 19285 6017 19305 6037
rect 19402 6017 19422 6037
rect 19498 6017 19518 6037
rect 19823 6013 19843 6033
rect 19919 6013 19939 6033
rect 20029 6013 20049 6033
rect 20125 6013 20145 6033
rect 20237 6013 20257 6033
rect 20333 6013 20353 6033
rect 20450 6013 20470 6033
rect 20546 6013 20566 6033
rect 825 5422 845 5442
rect 921 5422 941 5442
rect 1038 5422 1058 5442
rect 1134 5422 1154 5442
rect 1246 5422 1266 5442
rect 1342 5422 1362 5442
rect 1452 5422 1472 5442
rect 1548 5422 1568 5442
rect 1873 5418 1893 5438
rect 1969 5418 1989 5438
rect 2086 5418 2106 5438
rect 2182 5418 2202 5438
rect 2294 5418 2314 5438
rect 2390 5418 2410 5438
rect 2500 5418 2520 5438
rect 2596 5418 2616 5438
rect 6620 5256 6640 5276
rect 6716 5256 6736 5276
rect 6826 5256 6846 5276
rect 6922 5256 6942 5276
rect 7034 5256 7054 5276
rect 7130 5256 7150 5276
rect 7247 5256 7267 5276
rect 11533 5416 11553 5436
rect 11629 5416 11649 5436
rect 11746 5416 11766 5436
rect 11842 5416 11862 5436
rect 11954 5416 11974 5436
rect 12050 5416 12070 5436
rect 12160 5416 12180 5436
rect 12256 5416 12276 5436
rect 12581 5412 12601 5432
rect 7343 5256 7363 5276
rect 9115 5251 9135 5271
rect 9211 5251 9231 5271
rect 9321 5251 9341 5271
rect 9417 5251 9437 5271
rect 9529 5251 9549 5271
rect 9625 5251 9645 5271
rect 9742 5251 9762 5271
rect 12677 5412 12697 5432
rect 12794 5412 12814 5432
rect 12890 5412 12910 5432
rect 13002 5412 13022 5432
rect 13098 5412 13118 5432
rect 13208 5412 13228 5432
rect 13304 5412 13324 5432
rect 9838 5251 9858 5271
rect 17328 5250 17348 5270
rect 17424 5250 17444 5270
rect 17534 5250 17554 5270
rect 17630 5250 17650 5270
rect 17742 5250 17762 5270
rect 17838 5250 17858 5270
rect 17955 5250 17975 5270
rect 18051 5250 18071 5270
rect 19823 5245 19843 5265
rect 19919 5245 19939 5265
rect 20029 5245 20049 5265
rect 20125 5245 20145 5265
rect 20237 5245 20257 5265
rect 20333 5245 20353 5265
rect 20450 5245 20470 5265
rect 20546 5245 20566 5265
rect 825 4743 845 4763
rect 921 4743 941 4763
rect 1038 4743 1058 4763
rect 1134 4743 1154 4763
rect 1246 4743 1266 4763
rect 1342 4743 1362 4763
rect 1452 4743 1472 4763
rect 1548 4743 1568 4763
rect 3363 4740 3383 4760
rect 3459 4740 3479 4760
rect 3576 4740 3596 4760
rect 3672 4740 3692 4760
rect 3784 4740 3804 4760
rect 3880 4740 3900 4760
rect 3990 4740 4010 4760
rect 4086 4740 4106 4760
rect 11533 4737 11553 4757
rect 8067 4576 8087 4596
rect 8163 4576 8183 4596
rect 8273 4576 8293 4596
rect 8369 4576 8389 4596
rect 8481 4576 8501 4596
rect 8577 4576 8597 4596
rect 8694 4576 8714 4596
rect 11629 4737 11649 4757
rect 11746 4737 11766 4757
rect 11842 4737 11862 4757
rect 11954 4737 11974 4757
rect 12050 4737 12070 4757
rect 12160 4737 12180 4757
rect 12256 4737 12276 4757
rect 14071 4734 14091 4754
rect 8790 4576 8810 4596
rect 9115 4572 9135 4592
rect 9211 4572 9231 4592
rect 9321 4572 9341 4592
rect 9417 4572 9437 4592
rect 9529 4572 9549 4592
rect 9625 4572 9645 4592
rect 9742 4572 9762 4592
rect 9838 4572 9858 4592
rect 14167 4734 14187 4754
rect 14284 4734 14304 4754
rect 14380 4734 14400 4754
rect 14492 4734 14512 4754
rect 14588 4734 14608 4754
rect 14698 4734 14718 4754
rect 14794 4734 14814 4754
rect 18775 4570 18795 4590
rect 18871 4570 18891 4590
rect 18981 4570 19001 4590
rect 19077 4570 19097 4590
rect 19189 4570 19209 4590
rect 19285 4570 19305 4590
rect 19402 4570 19422 4590
rect 19498 4570 19518 4590
rect 19823 4566 19843 4586
rect 19919 4566 19939 4586
rect 20029 4566 20049 4586
rect 20125 4566 20145 4586
rect 20237 4566 20257 4586
rect 20333 4566 20353 4586
rect 20450 4566 20470 4586
rect 20546 4566 20566 4586
rect 826 3902 846 3922
rect 922 3902 942 3922
rect 1039 3902 1059 3922
rect 1135 3902 1155 3922
rect 1247 3902 1267 3922
rect 1343 3902 1363 3922
rect 1453 3902 1473 3922
rect 1549 3902 1569 3922
rect 1874 3898 1894 3918
rect 1970 3898 1990 3918
rect 2087 3898 2107 3918
rect 2183 3898 2203 3918
rect 2295 3898 2315 3918
rect 2391 3898 2411 3918
rect 2501 3898 2521 3918
rect 2597 3898 2617 3918
rect 4776 3904 4796 3924
rect 4872 3904 4892 3924
rect 4989 3904 5009 3924
rect 5085 3904 5105 3924
rect 5197 3904 5217 3924
rect 5293 3904 5313 3924
rect 5403 3904 5423 3924
rect 5499 3904 5519 3924
rect 6578 3734 6598 3754
rect 6674 3734 6694 3754
rect 6784 3734 6804 3754
rect 6880 3734 6900 3754
rect 6992 3734 7012 3754
rect 7088 3734 7108 3754
rect 7205 3734 7225 3754
rect 11534 3896 11554 3916
rect 11630 3896 11650 3916
rect 11747 3896 11767 3916
rect 11843 3896 11863 3916
rect 11955 3896 11975 3916
rect 12051 3896 12071 3916
rect 12161 3896 12181 3916
rect 12257 3896 12277 3916
rect 12582 3892 12602 3912
rect 7301 3734 7321 3754
rect 9116 3731 9136 3751
rect 9212 3731 9232 3751
rect 9322 3731 9342 3751
rect 9418 3731 9438 3751
rect 9530 3731 9550 3751
rect 9626 3731 9646 3751
rect 9743 3731 9763 3751
rect 12678 3892 12698 3912
rect 12795 3892 12815 3912
rect 12891 3892 12911 3912
rect 13003 3892 13023 3912
rect 13099 3892 13119 3912
rect 13209 3892 13229 3912
rect 13305 3892 13325 3912
rect 15484 3898 15504 3918
rect 15580 3898 15600 3918
rect 15697 3898 15717 3918
rect 15793 3898 15813 3918
rect 15905 3898 15925 3918
rect 16001 3898 16021 3918
rect 16111 3898 16131 3918
rect 16207 3898 16227 3918
rect 9839 3731 9859 3751
rect 17286 3728 17306 3748
rect 17382 3728 17402 3748
rect 17492 3728 17512 3748
rect 17588 3728 17608 3748
rect 17700 3728 17720 3748
rect 17796 3728 17816 3748
rect 17913 3728 17933 3748
rect 18009 3728 18029 3748
rect 19824 3725 19844 3745
rect 19920 3725 19940 3745
rect 20030 3725 20050 3745
rect 20126 3725 20146 3745
rect 20238 3725 20258 3745
rect 20334 3725 20354 3745
rect 20451 3725 20471 3745
rect 20547 3725 20567 3745
rect 826 3223 846 3243
rect 922 3223 942 3243
rect 1039 3223 1059 3243
rect 1135 3223 1155 3243
rect 1247 3223 1267 3243
rect 1343 3223 1363 3243
rect 1453 3223 1473 3243
rect 1549 3223 1569 3243
rect 3321 3218 3341 3238
rect 3417 3218 3437 3238
rect 3534 3218 3554 3238
rect 3630 3218 3650 3238
rect 3742 3218 3762 3238
rect 3838 3218 3858 3238
rect 3948 3218 3968 3238
rect 4044 3218 4064 3238
rect 11534 3217 11554 3237
rect 8068 3056 8088 3076
rect 8164 3056 8184 3076
rect 8274 3056 8294 3076
rect 8370 3056 8390 3076
rect 8482 3056 8502 3076
rect 8578 3056 8598 3076
rect 8695 3056 8715 3076
rect 11630 3217 11650 3237
rect 11747 3217 11767 3237
rect 11843 3217 11863 3237
rect 11955 3217 11975 3237
rect 12051 3217 12071 3237
rect 12161 3217 12181 3237
rect 12257 3217 12277 3237
rect 14029 3212 14049 3232
rect 8791 3056 8811 3076
rect 9116 3052 9136 3072
rect 9212 3052 9232 3072
rect 9322 3052 9342 3072
rect 9418 3052 9438 3072
rect 9530 3052 9550 3072
rect 9626 3052 9646 3072
rect 9743 3052 9763 3072
rect 9839 3052 9859 3072
rect 14125 3212 14145 3232
rect 14242 3212 14262 3232
rect 14338 3212 14358 3232
rect 14450 3212 14470 3232
rect 14546 3212 14566 3232
rect 14656 3212 14676 3232
rect 14752 3212 14772 3232
rect 18776 3050 18796 3070
rect 18872 3050 18892 3070
rect 18982 3050 19002 3070
rect 19078 3050 19098 3070
rect 19190 3050 19210 3070
rect 19286 3050 19306 3070
rect 19403 3050 19423 3070
rect 19499 3050 19519 3070
rect 19824 3046 19844 3066
rect 19920 3046 19940 3066
rect 20030 3046 20050 3066
rect 20126 3046 20146 3066
rect 20238 3046 20258 3066
rect 20334 3046 20354 3066
rect 20451 3046 20471 3066
rect 20547 3046 20567 3066
rect 826 2455 846 2475
rect 922 2455 942 2475
rect 1039 2455 1059 2475
rect 1135 2455 1155 2475
rect 1247 2455 1267 2475
rect 1343 2455 1363 2475
rect 1453 2455 1473 2475
rect 1549 2455 1569 2475
rect 1874 2451 1894 2471
rect 1970 2451 1990 2471
rect 2087 2451 2107 2471
rect 2183 2451 2203 2471
rect 2295 2451 2315 2471
rect 2391 2451 2411 2471
rect 2501 2451 2521 2471
rect 2597 2451 2617 2471
rect 6621 2289 6641 2309
rect 6717 2289 6737 2309
rect 6827 2289 6847 2309
rect 6923 2289 6943 2309
rect 7035 2289 7055 2309
rect 7131 2289 7151 2309
rect 7248 2289 7268 2309
rect 11534 2449 11554 2469
rect 11630 2449 11650 2469
rect 11747 2449 11767 2469
rect 11843 2449 11863 2469
rect 11955 2449 11975 2469
rect 12051 2449 12071 2469
rect 12161 2449 12181 2469
rect 12257 2449 12277 2469
rect 12582 2445 12602 2465
rect 7344 2289 7364 2309
rect 9116 2284 9136 2304
rect 9212 2284 9232 2304
rect 9322 2284 9342 2304
rect 9418 2284 9438 2304
rect 9530 2284 9550 2304
rect 9626 2284 9646 2304
rect 9743 2284 9763 2304
rect 12678 2445 12698 2465
rect 12795 2445 12815 2465
rect 12891 2445 12911 2465
rect 13003 2445 13023 2465
rect 13099 2445 13119 2465
rect 13209 2445 13229 2465
rect 13305 2445 13325 2465
rect 9839 2284 9859 2304
rect 17329 2283 17349 2303
rect 17425 2283 17445 2303
rect 17535 2283 17555 2303
rect 17631 2283 17651 2303
rect 17743 2283 17763 2303
rect 17839 2283 17859 2303
rect 17956 2283 17976 2303
rect 18052 2283 18072 2303
rect 19824 2278 19844 2298
rect 19920 2278 19940 2298
rect 20030 2278 20050 2298
rect 20126 2278 20146 2298
rect 20238 2278 20258 2298
rect 20334 2278 20354 2298
rect 20451 2278 20471 2298
rect 20547 2278 20567 2298
rect 826 1776 846 1796
rect 922 1776 942 1796
rect 1039 1776 1059 1796
rect 1135 1776 1155 1796
rect 1247 1776 1267 1796
rect 1343 1776 1363 1796
rect 1453 1776 1473 1796
rect 1549 1776 1569 1796
rect 11534 1770 11554 1790
rect 8068 1609 8088 1629
rect 8164 1609 8184 1629
rect 8274 1609 8294 1629
rect 8370 1609 8390 1629
rect 8482 1609 8502 1629
rect 8578 1609 8598 1629
rect 8695 1609 8715 1629
rect 11630 1770 11650 1790
rect 11747 1770 11767 1790
rect 11843 1770 11863 1790
rect 11955 1770 11975 1790
rect 12051 1770 12071 1790
rect 12161 1770 12181 1790
rect 12257 1770 12277 1790
rect 8791 1609 8811 1629
rect 9116 1605 9136 1625
rect 9212 1605 9232 1625
rect 9322 1605 9342 1625
rect 9418 1605 9438 1625
rect 9530 1605 9550 1625
rect 9626 1605 9646 1625
rect 9743 1605 9763 1625
rect 9839 1605 9859 1625
rect 18776 1603 18796 1623
rect 18872 1603 18892 1623
rect 18982 1603 19002 1623
rect 19078 1603 19098 1623
rect 19190 1603 19210 1623
rect 19286 1603 19306 1623
rect 19403 1603 19423 1623
rect 19499 1603 19519 1623
rect 19824 1599 19844 1619
rect 19920 1599 19940 1619
rect 20030 1599 20050 1619
rect 20126 1599 20146 1619
rect 20238 1599 20258 1619
rect 20334 1599 20354 1619
rect 20451 1599 20471 1619
rect 20547 1599 20567 1619
rect 10537 -383 10557 -363
rect 10633 -383 10653 -363
rect 10750 -383 10770 -363
rect 10846 -383 10866 -363
rect 10958 -383 10978 -363
rect 11054 -383 11074 -363
rect 11164 -383 11184 -363
rect 11260 -383 11280 -363
<< psubdiff >>
rect 9681 12972 9792 12983
rect 9681 12942 9723 12972
rect 9751 12942 9792 12972
rect 20389 12966 20500 12981
rect 9681 12928 9792 12942
rect 20389 12936 20431 12966
rect 20459 12936 20500 12966
rect 895 12661 1006 12675
rect 895 12631 936 12661
rect 964 12631 1006 12661
rect 895 12616 1006 12631
rect 1943 12657 2054 12671
rect 20389 12922 20500 12936
rect 1943 12627 1984 12657
rect 2012 12627 2054 12657
rect 11603 12655 11714 12669
rect 1943 12612 2054 12627
rect 11603 12625 11644 12655
rect 11672 12625 11714 12655
rect 11603 12610 11714 12625
rect 12651 12651 12762 12665
rect 12651 12621 12692 12651
rect 12720 12621 12762 12651
rect 12651 12606 12762 12621
rect 8633 12297 8744 12312
rect 8633 12267 8675 12297
rect 8703 12267 8744 12297
rect 8633 12253 8744 12267
rect 9681 12293 9792 12308
rect 9681 12263 9723 12293
rect 9751 12263 9792 12293
rect 19341 12291 19452 12306
rect 9681 12249 9792 12263
rect 19341 12261 19383 12291
rect 19411 12261 19452 12291
rect 895 11982 1006 11996
rect 19341 12247 19452 12261
rect 20389 12287 20500 12302
rect 20389 12257 20431 12287
rect 20459 12257 20500 12287
rect 895 11952 936 11982
rect 964 11952 1006 11982
rect 895 11939 1006 11952
rect 3390 11977 3501 11991
rect 20389 12243 20500 12257
rect 3390 11947 3431 11977
rect 3459 11947 3501 11977
rect 11603 11976 11714 11990
rect 3390 11932 3501 11947
rect 11603 11946 11644 11976
rect 11672 11946 11714 11976
rect 11603 11933 11714 11946
rect 14098 11971 14209 11985
rect 14098 11941 14139 11971
rect 14167 11941 14209 11971
rect 14098 11926 14209 11941
rect 7186 11530 7297 11545
rect 7186 11500 7228 11530
rect 7256 11500 7297 11530
rect 7186 11486 7297 11500
rect 9681 11525 9792 11538
rect 9681 11495 9723 11525
rect 9751 11495 9792 11525
rect 17894 11524 18005 11539
rect 9681 11481 9792 11495
rect 17894 11494 17936 11524
rect 17964 11494 18005 11524
rect 895 11214 1006 11228
rect 17894 11480 18005 11494
rect 20389 11519 20500 11532
rect 20389 11489 20431 11519
rect 20459 11489 20500 11519
rect 895 11184 936 11214
rect 964 11184 1006 11214
rect 895 11169 1006 11184
rect 1943 11210 2054 11224
rect 20389 11475 20500 11489
rect 1943 11180 1984 11210
rect 2012 11180 2054 11210
rect 11603 11208 11714 11222
rect 1943 11165 2054 11180
rect 11603 11178 11644 11208
rect 11672 11178 11714 11208
rect 11603 11163 11714 11178
rect 12651 11204 12762 11218
rect 12651 11174 12692 11204
rect 12720 11174 12762 11204
rect 12651 11159 12762 11174
rect 8633 10850 8744 10865
rect 8633 10820 8675 10850
rect 8703 10820 8744 10850
rect 8633 10806 8744 10820
rect 9681 10846 9792 10861
rect 9681 10816 9723 10846
rect 9751 10816 9792 10846
rect 19341 10844 19452 10859
rect 9681 10802 9792 10816
rect 19341 10814 19383 10844
rect 19411 10814 19452 10844
rect 895 10535 1006 10549
rect 19341 10800 19452 10814
rect 20389 10840 20500 10855
rect 20389 10810 20431 10840
rect 20459 10810 20500 10840
rect 895 10505 936 10535
rect 964 10505 1006 10535
rect 895 10490 1006 10505
rect 3433 10532 3544 10546
rect 20389 10796 20500 10810
rect 3433 10502 3474 10532
rect 3502 10502 3544 10532
rect 11603 10529 11714 10543
rect 3433 10487 3544 10502
rect 11603 10499 11644 10529
rect 11672 10499 11714 10529
rect 11603 10484 11714 10499
rect 14141 10526 14252 10540
rect 14141 10496 14182 10526
rect 14210 10496 14252 10526
rect 14141 10481 14252 10496
rect 7144 10008 7255 10023
rect 7144 9978 7186 10008
rect 7214 9978 7255 10008
rect 7144 9964 7255 9978
rect 9682 10005 9793 10020
rect 9682 9975 9724 10005
rect 9752 9975 9793 10005
rect 17852 10002 17963 10017
rect 9682 9961 9793 9975
rect 17852 9972 17894 10002
rect 17922 9972 17963 10002
rect 896 9694 1007 9708
rect 17852 9958 17963 9972
rect 20390 9999 20501 10014
rect 20390 9969 20432 9999
rect 20460 9969 20501 9999
rect 896 9664 937 9694
rect 965 9664 1007 9694
rect 896 9649 1007 9664
rect 1944 9690 2055 9704
rect 20390 9955 20501 9969
rect 1944 9660 1985 9690
rect 2013 9660 2055 9690
rect 11604 9688 11715 9702
rect 1944 9645 2055 9660
rect 11604 9658 11645 9688
rect 11673 9658 11715 9688
rect 11604 9643 11715 9658
rect 12652 9684 12763 9698
rect 12652 9654 12693 9684
rect 12721 9654 12763 9684
rect 12652 9639 12763 9654
rect 8634 9330 8745 9345
rect 8634 9300 8676 9330
rect 8704 9300 8745 9330
rect 8634 9286 8745 9300
rect 9682 9326 9793 9341
rect 9682 9296 9724 9326
rect 9752 9296 9793 9326
rect 19342 9324 19453 9339
rect 9682 9282 9793 9296
rect 19342 9294 19384 9324
rect 19412 9294 19453 9324
rect 896 9015 1007 9029
rect 19342 9280 19453 9294
rect 20390 9320 20501 9335
rect 20390 9290 20432 9320
rect 20460 9290 20501 9320
rect 896 8985 937 9015
rect 965 8985 1007 9015
rect 896 8972 1007 8985
rect 3391 9010 3502 9024
rect 20390 9276 20501 9290
rect 3391 8980 3432 9010
rect 3460 8980 3502 9010
rect 11604 9009 11715 9023
rect 3391 8965 3502 8980
rect 11604 8979 11645 9009
rect 11673 8979 11715 9009
rect 11604 8966 11715 8979
rect 14099 9004 14210 9018
rect 14099 8974 14140 9004
rect 14168 8974 14210 9004
rect 14099 8959 14210 8974
rect 7187 8563 7298 8578
rect 7187 8533 7229 8563
rect 7257 8533 7298 8563
rect 7187 8519 7298 8533
rect 9682 8558 9793 8571
rect 9682 8528 9724 8558
rect 9752 8528 9793 8558
rect 17895 8557 18006 8572
rect 9682 8514 9793 8528
rect 17895 8527 17937 8557
rect 17965 8527 18006 8557
rect 896 8247 1007 8261
rect 17895 8513 18006 8527
rect 20390 8552 20501 8565
rect 20390 8522 20432 8552
rect 20460 8522 20501 8552
rect 896 8217 937 8247
rect 965 8217 1007 8247
rect 896 8202 1007 8217
rect 1944 8243 2055 8257
rect 20390 8508 20501 8522
rect 1944 8213 1985 8243
rect 2013 8213 2055 8243
rect 11604 8241 11715 8255
rect 1944 8198 2055 8213
rect 11604 8211 11645 8241
rect 11673 8211 11715 8241
rect 11604 8196 11715 8211
rect 12652 8237 12763 8251
rect 12652 8207 12693 8237
rect 12721 8207 12763 8237
rect 12652 8192 12763 8207
rect 8634 7883 8745 7898
rect 8634 7853 8676 7883
rect 8704 7853 8745 7883
rect 8634 7839 8745 7853
rect 9682 7879 9793 7894
rect 9682 7849 9724 7879
rect 9752 7849 9793 7879
rect 19342 7877 19453 7892
rect 9682 7835 9793 7849
rect 19342 7847 19384 7877
rect 19412 7847 19453 7877
rect 896 7568 1007 7582
rect 19342 7833 19453 7847
rect 20390 7873 20501 7888
rect 20390 7843 20432 7873
rect 20460 7843 20501 7873
rect 20390 7829 20501 7843
rect 896 7538 937 7568
rect 965 7538 1007 7568
rect 896 7523 1007 7538
rect 4499 7559 4610 7573
rect 11604 7562 11715 7576
rect 4499 7529 4540 7559
rect 4568 7529 4610 7559
rect 4499 7514 4610 7529
rect 11604 7532 11645 7562
rect 11673 7532 11715 7562
rect 11604 7517 11715 7532
rect 15207 7553 15318 7567
rect 15207 7523 15248 7553
rect 15276 7523 15318 7553
rect 15207 7508 15318 7523
rect 6076 6973 6187 6988
rect 6076 6943 6118 6973
rect 6146 6943 6187 6973
rect 6076 6929 6187 6943
rect 9679 6964 9790 6979
rect 9679 6934 9721 6964
rect 9749 6934 9790 6964
rect 16784 6967 16895 6982
rect 16784 6937 16826 6967
rect 16854 6937 16895 6967
rect 9679 6920 9790 6934
rect 16784 6923 16895 6937
rect 20387 6958 20498 6973
rect 20387 6928 20429 6958
rect 20457 6928 20498 6958
rect 893 6653 1004 6667
rect 893 6623 934 6653
rect 962 6623 1004 6653
rect 893 6608 1004 6623
rect 1941 6649 2052 6663
rect 20387 6914 20498 6928
rect 1941 6619 1982 6649
rect 2010 6619 2052 6649
rect 11601 6647 11712 6661
rect 1941 6604 2052 6619
rect 11601 6617 11642 6647
rect 11670 6617 11712 6647
rect 11601 6602 11712 6617
rect 12649 6643 12760 6657
rect 12649 6613 12690 6643
rect 12718 6613 12760 6643
rect 12649 6598 12760 6613
rect 8631 6289 8742 6304
rect 8631 6259 8673 6289
rect 8701 6259 8742 6289
rect 8631 6245 8742 6259
rect 9679 6285 9790 6300
rect 9679 6255 9721 6285
rect 9749 6255 9790 6285
rect 19339 6283 19450 6298
rect 9679 6241 9790 6255
rect 19339 6253 19381 6283
rect 19409 6253 19450 6283
rect 893 5974 1004 5988
rect 19339 6239 19450 6253
rect 20387 6279 20498 6294
rect 20387 6249 20429 6279
rect 20457 6249 20498 6279
rect 893 5944 934 5974
rect 962 5944 1004 5974
rect 893 5931 1004 5944
rect 3388 5969 3499 5983
rect 20387 6235 20498 6249
rect 3388 5939 3429 5969
rect 3457 5939 3499 5969
rect 11601 5968 11712 5982
rect 3388 5924 3499 5939
rect 11601 5938 11642 5968
rect 11670 5938 11712 5968
rect 11601 5925 11712 5938
rect 14096 5963 14207 5977
rect 14096 5933 14137 5963
rect 14165 5933 14207 5963
rect 14096 5918 14207 5933
rect 7184 5522 7295 5537
rect 7184 5492 7226 5522
rect 7254 5492 7295 5522
rect 7184 5478 7295 5492
rect 9679 5517 9790 5530
rect 9679 5487 9721 5517
rect 9749 5487 9790 5517
rect 17892 5516 18003 5531
rect 9679 5473 9790 5487
rect 17892 5486 17934 5516
rect 17962 5486 18003 5516
rect 893 5206 1004 5220
rect 17892 5472 18003 5486
rect 20387 5511 20498 5524
rect 20387 5481 20429 5511
rect 20457 5481 20498 5511
rect 893 5176 934 5206
rect 962 5176 1004 5206
rect 893 5161 1004 5176
rect 1941 5202 2052 5216
rect 20387 5467 20498 5481
rect 1941 5172 1982 5202
rect 2010 5172 2052 5202
rect 11601 5200 11712 5214
rect 1941 5157 2052 5172
rect 11601 5170 11642 5200
rect 11670 5170 11712 5200
rect 11601 5155 11712 5170
rect 12649 5196 12760 5210
rect 12649 5166 12690 5196
rect 12718 5166 12760 5196
rect 12649 5151 12760 5166
rect 8631 4842 8742 4857
rect 8631 4812 8673 4842
rect 8701 4812 8742 4842
rect 8631 4798 8742 4812
rect 9679 4838 9790 4853
rect 9679 4808 9721 4838
rect 9749 4808 9790 4838
rect 19339 4836 19450 4851
rect 9679 4794 9790 4808
rect 19339 4806 19381 4836
rect 19409 4806 19450 4836
rect 893 4527 1004 4541
rect 19339 4792 19450 4806
rect 20387 4832 20498 4847
rect 20387 4802 20429 4832
rect 20457 4802 20498 4832
rect 893 4497 934 4527
rect 962 4497 1004 4527
rect 893 4482 1004 4497
rect 3431 4524 3542 4538
rect 20387 4788 20498 4802
rect 3431 4494 3472 4524
rect 3500 4494 3542 4524
rect 11601 4521 11712 4535
rect 3431 4479 3542 4494
rect 11601 4491 11642 4521
rect 11670 4491 11712 4521
rect 11601 4476 11712 4491
rect 14139 4518 14250 4532
rect 14139 4488 14180 4518
rect 14208 4488 14250 4518
rect 14139 4473 14250 4488
rect 7142 4000 7253 4015
rect 7142 3970 7184 4000
rect 7212 3970 7253 4000
rect 7142 3956 7253 3970
rect 9680 3997 9791 4012
rect 9680 3967 9722 3997
rect 9750 3967 9791 3997
rect 17850 3994 17961 4009
rect 9680 3953 9791 3967
rect 894 3686 1005 3700
rect 894 3656 935 3686
rect 963 3656 1005 3686
rect 894 3641 1005 3656
rect 1942 3682 2053 3696
rect 1942 3652 1983 3682
rect 2011 3652 2053 3682
rect 1942 3637 2053 3652
rect 4844 3688 4955 3702
rect 17850 3964 17892 3994
rect 17920 3964 17961 3994
rect 4844 3658 4885 3688
rect 4913 3658 4955 3688
rect 17850 3950 17961 3964
rect 20388 3991 20499 4006
rect 20388 3961 20430 3991
rect 20458 3961 20499 3991
rect 20388 3947 20499 3961
rect 11602 3680 11713 3694
rect 4844 3643 4955 3658
rect 11602 3650 11643 3680
rect 11671 3650 11713 3680
rect 11602 3635 11713 3650
rect 12650 3676 12761 3690
rect 12650 3646 12691 3676
rect 12719 3646 12761 3676
rect 12650 3631 12761 3646
rect 15552 3682 15663 3696
rect 15552 3652 15593 3682
rect 15621 3652 15663 3682
rect 15552 3637 15663 3652
rect 8632 3322 8743 3337
rect 8632 3292 8674 3322
rect 8702 3292 8743 3322
rect 8632 3278 8743 3292
rect 9680 3318 9791 3333
rect 9680 3288 9722 3318
rect 9750 3288 9791 3318
rect 19340 3316 19451 3331
rect 9680 3274 9791 3288
rect 19340 3286 19382 3316
rect 19410 3286 19451 3316
rect 894 3007 1005 3021
rect 19340 3272 19451 3286
rect 20388 3312 20499 3327
rect 20388 3282 20430 3312
rect 20458 3282 20499 3312
rect 894 2977 935 3007
rect 963 2977 1005 3007
rect 894 2964 1005 2977
rect 3389 3002 3500 3016
rect 20388 3268 20499 3282
rect 3389 2972 3430 3002
rect 3458 2972 3500 3002
rect 11602 3001 11713 3015
rect 3389 2957 3500 2972
rect 11602 2971 11643 3001
rect 11671 2971 11713 3001
rect 11602 2958 11713 2971
rect 14097 2996 14208 3010
rect 14097 2966 14138 2996
rect 14166 2966 14208 2996
rect 14097 2951 14208 2966
rect 7185 2555 7296 2570
rect 7185 2525 7227 2555
rect 7255 2525 7296 2555
rect 7185 2511 7296 2525
rect 9680 2550 9791 2563
rect 9680 2520 9722 2550
rect 9750 2520 9791 2550
rect 17893 2549 18004 2564
rect 9680 2506 9791 2520
rect 17893 2519 17935 2549
rect 17963 2519 18004 2549
rect 894 2239 1005 2253
rect 17893 2505 18004 2519
rect 20388 2544 20499 2557
rect 20388 2514 20430 2544
rect 20458 2514 20499 2544
rect 894 2209 935 2239
rect 963 2209 1005 2239
rect 894 2194 1005 2209
rect 1942 2235 2053 2249
rect 20388 2500 20499 2514
rect 1942 2205 1983 2235
rect 2011 2205 2053 2235
rect 11602 2233 11713 2247
rect 1942 2190 2053 2205
rect 11602 2203 11643 2233
rect 11671 2203 11713 2233
rect 11602 2188 11713 2203
rect 12650 2229 12761 2243
rect 12650 2199 12691 2229
rect 12719 2199 12761 2229
rect 12650 2184 12761 2199
rect 8632 1875 8743 1890
rect 8632 1845 8674 1875
rect 8702 1845 8743 1875
rect 8632 1831 8743 1845
rect 9680 1871 9791 1886
rect 9680 1841 9722 1871
rect 9750 1841 9791 1871
rect 19340 1869 19451 1884
rect 9680 1827 9791 1841
rect 19340 1839 19382 1869
rect 19410 1839 19451 1869
rect 894 1560 1005 1574
rect 19340 1825 19451 1839
rect 20388 1865 20499 1880
rect 20388 1835 20430 1865
rect 20458 1835 20499 1865
rect 20388 1821 20499 1835
rect 894 1530 935 1560
rect 963 1530 1005 1560
rect 11602 1554 11713 1568
rect 894 1515 1005 1530
rect 11602 1524 11643 1554
rect 11671 1524 11713 1554
rect 11602 1509 11713 1524
rect 10605 -599 10716 -585
rect 10605 -629 10646 -599
rect 10674 -629 10716 -599
rect 10605 -644 10716 -629
<< nsubdiff >>
rect 896 13008 1006 13022
rect 896 12978 939 13008
rect 967 12978 1006 13008
rect 896 12963 1006 12978
rect 1944 13004 2054 13018
rect 1944 12974 1987 13004
rect 2015 12974 2054 13004
rect 11604 13002 11714 13016
rect 1944 12959 2054 12974
rect 11604 12972 11647 13002
rect 11675 12972 11714 13002
rect 11604 12957 11714 12972
rect 12652 12998 12762 13012
rect 12652 12968 12695 12998
rect 12723 12968 12762 12998
rect 12652 12953 12762 12968
rect 9681 12625 9791 12640
rect 9681 12595 9720 12625
rect 9748 12595 9791 12625
rect 9681 12581 9791 12595
rect 20389 12619 20499 12634
rect 20389 12589 20428 12619
rect 20456 12589 20499 12619
rect 20389 12575 20499 12589
rect 896 12329 1006 12343
rect 896 12299 939 12329
rect 967 12299 1006 12329
rect 896 12284 1006 12299
rect 3391 12324 3501 12338
rect 3391 12294 3434 12324
rect 3462 12294 3501 12324
rect 3391 12279 3501 12294
rect 11604 12323 11714 12337
rect 11604 12293 11647 12323
rect 11675 12293 11714 12323
rect 11604 12278 11714 12293
rect 14099 12318 14209 12332
rect 14099 12288 14142 12318
rect 14170 12288 14209 12318
rect 14099 12273 14209 12288
rect 8633 11950 8743 11965
rect 8633 11920 8672 11950
rect 8700 11920 8743 11950
rect 8633 11906 8743 11920
rect 9681 11946 9791 11961
rect 9681 11916 9720 11946
rect 9748 11916 9791 11946
rect 9681 11902 9791 11916
rect 19341 11944 19451 11959
rect 19341 11914 19380 11944
rect 19408 11914 19451 11944
rect 19341 11900 19451 11914
rect 20389 11940 20499 11955
rect 20389 11910 20428 11940
rect 20456 11910 20499 11940
rect 20389 11896 20499 11910
rect 896 11561 1006 11575
rect 896 11531 939 11561
rect 967 11531 1006 11561
rect 896 11516 1006 11531
rect 1944 11557 2054 11571
rect 1944 11527 1987 11557
rect 2015 11527 2054 11557
rect 1944 11512 2054 11527
rect 11604 11555 11714 11569
rect 11604 11525 11647 11555
rect 11675 11525 11714 11555
rect 11604 11510 11714 11525
rect 12652 11551 12762 11565
rect 12652 11521 12695 11551
rect 12723 11521 12762 11551
rect 12652 11506 12762 11521
rect 7186 11183 7296 11198
rect 7186 11153 7225 11183
rect 7253 11153 7296 11183
rect 7186 11139 7296 11153
rect 9681 11178 9791 11193
rect 9681 11148 9720 11178
rect 9748 11148 9791 11178
rect 9681 11134 9791 11148
rect 17894 11177 18004 11192
rect 17894 11147 17933 11177
rect 17961 11147 18004 11177
rect 17894 11133 18004 11147
rect 20389 11172 20499 11187
rect 20389 11142 20428 11172
rect 20456 11142 20499 11172
rect 20389 11128 20499 11142
rect 896 10882 1006 10896
rect 896 10852 939 10882
rect 967 10852 1006 10882
rect 896 10837 1006 10852
rect 3434 10879 3544 10893
rect 3434 10849 3477 10879
rect 3505 10849 3544 10879
rect 3434 10834 3544 10849
rect 11604 10876 11714 10890
rect 11604 10846 11647 10876
rect 11675 10846 11714 10876
rect 11604 10831 11714 10846
rect 14142 10873 14252 10887
rect 14142 10843 14185 10873
rect 14213 10843 14252 10873
rect 14142 10828 14252 10843
rect 8633 10503 8743 10518
rect 8633 10473 8672 10503
rect 8700 10473 8743 10503
rect 8633 10459 8743 10473
rect 9681 10499 9791 10514
rect 9681 10469 9720 10499
rect 9748 10469 9791 10499
rect 9681 10455 9791 10469
rect 19341 10497 19451 10512
rect 19341 10467 19380 10497
rect 19408 10467 19451 10497
rect 19341 10453 19451 10467
rect 20389 10493 20499 10508
rect 20389 10463 20428 10493
rect 20456 10463 20499 10493
rect 20389 10449 20499 10463
rect 897 10041 1007 10055
rect 897 10011 940 10041
rect 968 10011 1007 10041
rect 897 9996 1007 10011
rect 1945 10037 2055 10051
rect 1945 10007 1988 10037
rect 2016 10007 2055 10037
rect 1945 9992 2055 10007
rect 11605 10035 11715 10049
rect 11605 10005 11648 10035
rect 11676 10005 11715 10035
rect 11605 9990 11715 10005
rect 12653 10031 12763 10045
rect 12653 10001 12696 10031
rect 12724 10001 12763 10031
rect 12653 9986 12763 10001
rect 7144 9661 7254 9676
rect 7144 9631 7183 9661
rect 7211 9631 7254 9661
rect 7144 9617 7254 9631
rect 9682 9658 9792 9673
rect 9682 9628 9721 9658
rect 9749 9628 9792 9658
rect 9682 9614 9792 9628
rect 17852 9655 17962 9670
rect 17852 9625 17891 9655
rect 17919 9625 17962 9655
rect 17852 9611 17962 9625
rect 20390 9652 20500 9667
rect 20390 9622 20429 9652
rect 20457 9622 20500 9652
rect 20390 9608 20500 9622
rect 897 9362 1007 9376
rect 897 9332 940 9362
rect 968 9332 1007 9362
rect 897 9317 1007 9332
rect 3392 9357 3502 9371
rect 3392 9327 3435 9357
rect 3463 9327 3502 9357
rect 3392 9312 3502 9327
rect 11605 9356 11715 9370
rect 11605 9326 11648 9356
rect 11676 9326 11715 9356
rect 11605 9311 11715 9326
rect 14100 9351 14210 9365
rect 14100 9321 14143 9351
rect 14171 9321 14210 9351
rect 14100 9306 14210 9321
rect 8634 8983 8744 8998
rect 8634 8953 8673 8983
rect 8701 8953 8744 8983
rect 8634 8939 8744 8953
rect 9682 8979 9792 8994
rect 9682 8949 9721 8979
rect 9749 8949 9792 8979
rect 9682 8935 9792 8949
rect 19342 8977 19452 8992
rect 19342 8947 19381 8977
rect 19409 8947 19452 8977
rect 19342 8933 19452 8947
rect 20390 8973 20500 8988
rect 20390 8943 20429 8973
rect 20457 8943 20500 8973
rect 20390 8929 20500 8943
rect 897 8594 1007 8608
rect 897 8564 940 8594
rect 968 8564 1007 8594
rect 897 8549 1007 8564
rect 1945 8590 2055 8604
rect 1945 8560 1988 8590
rect 2016 8560 2055 8590
rect 1945 8545 2055 8560
rect 11605 8588 11715 8602
rect 11605 8558 11648 8588
rect 11676 8558 11715 8588
rect 11605 8543 11715 8558
rect 12653 8584 12763 8598
rect 12653 8554 12696 8584
rect 12724 8554 12763 8584
rect 12653 8539 12763 8554
rect 7187 8216 7297 8231
rect 7187 8186 7226 8216
rect 7254 8186 7297 8216
rect 7187 8172 7297 8186
rect 9682 8211 9792 8226
rect 9682 8181 9721 8211
rect 9749 8181 9792 8211
rect 9682 8167 9792 8181
rect 17895 8210 18005 8225
rect 17895 8180 17934 8210
rect 17962 8180 18005 8210
rect 17895 8166 18005 8180
rect 20390 8205 20500 8220
rect 20390 8175 20429 8205
rect 20457 8175 20500 8205
rect 20390 8161 20500 8175
rect 897 7915 1007 7929
rect 897 7885 940 7915
rect 968 7885 1007 7915
rect 897 7870 1007 7885
rect 4500 7906 4610 7920
rect 4500 7876 4543 7906
rect 4571 7876 4610 7906
rect 4500 7861 4610 7876
rect 11605 7909 11715 7923
rect 11605 7879 11648 7909
rect 11676 7879 11715 7909
rect 11605 7864 11715 7879
rect 15208 7900 15318 7914
rect 15208 7870 15251 7900
rect 15279 7870 15318 7900
rect 15208 7855 15318 7870
rect 8634 7536 8744 7551
rect 8634 7506 8673 7536
rect 8701 7506 8744 7536
rect 8634 7492 8744 7506
rect 9682 7532 9792 7547
rect 9682 7502 9721 7532
rect 9749 7502 9792 7532
rect 9682 7488 9792 7502
rect 19342 7530 19452 7545
rect 19342 7500 19381 7530
rect 19409 7500 19452 7530
rect 19342 7486 19452 7500
rect 20390 7526 20500 7541
rect 20390 7496 20429 7526
rect 20457 7496 20500 7526
rect 20390 7482 20500 7496
rect 894 7000 1004 7014
rect 894 6970 937 7000
rect 965 6970 1004 7000
rect 894 6955 1004 6970
rect 1942 6996 2052 7010
rect 1942 6966 1985 6996
rect 2013 6966 2052 6996
rect 1942 6951 2052 6966
rect 11602 6994 11712 7008
rect 11602 6964 11645 6994
rect 11673 6964 11712 6994
rect 11602 6949 11712 6964
rect 12650 6990 12760 7004
rect 12650 6960 12693 6990
rect 12721 6960 12760 6990
rect 12650 6945 12760 6960
rect 6076 6626 6186 6641
rect 6076 6596 6115 6626
rect 6143 6596 6186 6626
rect 6076 6582 6186 6596
rect 9679 6617 9789 6632
rect 9679 6587 9718 6617
rect 9746 6587 9789 6617
rect 9679 6573 9789 6587
rect 16784 6620 16894 6635
rect 16784 6590 16823 6620
rect 16851 6590 16894 6620
rect 16784 6576 16894 6590
rect 20387 6611 20497 6626
rect 20387 6581 20426 6611
rect 20454 6581 20497 6611
rect 20387 6567 20497 6581
rect 894 6321 1004 6335
rect 894 6291 937 6321
rect 965 6291 1004 6321
rect 894 6276 1004 6291
rect 3389 6316 3499 6330
rect 3389 6286 3432 6316
rect 3460 6286 3499 6316
rect 3389 6271 3499 6286
rect 11602 6315 11712 6329
rect 11602 6285 11645 6315
rect 11673 6285 11712 6315
rect 11602 6270 11712 6285
rect 14097 6310 14207 6324
rect 14097 6280 14140 6310
rect 14168 6280 14207 6310
rect 14097 6265 14207 6280
rect 8631 5942 8741 5957
rect 8631 5912 8670 5942
rect 8698 5912 8741 5942
rect 8631 5898 8741 5912
rect 9679 5938 9789 5953
rect 9679 5908 9718 5938
rect 9746 5908 9789 5938
rect 9679 5894 9789 5908
rect 19339 5936 19449 5951
rect 19339 5906 19378 5936
rect 19406 5906 19449 5936
rect 19339 5892 19449 5906
rect 20387 5932 20497 5947
rect 20387 5902 20426 5932
rect 20454 5902 20497 5932
rect 20387 5888 20497 5902
rect 894 5553 1004 5567
rect 894 5523 937 5553
rect 965 5523 1004 5553
rect 894 5508 1004 5523
rect 1942 5549 2052 5563
rect 1942 5519 1985 5549
rect 2013 5519 2052 5549
rect 1942 5504 2052 5519
rect 11602 5547 11712 5561
rect 11602 5517 11645 5547
rect 11673 5517 11712 5547
rect 11602 5502 11712 5517
rect 12650 5543 12760 5557
rect 12650 5513 12693 5543
rect 12721 5513 12760 5543
rect 12650 5498 12760 5513
rect 7184 5175 7294 5190
rect 7184 5145 7223 5175
rect 7251 5145 7294 5175
rect 7184 5131 7294 5145
rect 9679 5170 9789 5185
rect 9679 5140 9718 5170
rect 9746 5140 9789 5170
rect 9679 5126 9789 5140
rect 17892 5169 18002 5184
rect 17892 5139 17931 5169
rect 17959 5139 18002 5169
rect 17892 5125 18002 5139
rect 20387 5164 20497 5179
rect 20387 5134 20426 5164
rect 20454 5134 20497 5164
rect 20387 5120 20497 5134
rect 894 4874 1004 4888
rect 894 4844 937 4874
rect 965 4844 1004 4874
rect 894 4829 1004 4844
rect 3432 4871 3542 4885
rect 3432 4841 3475 4871
rect 3503 4841 3542 4871
rect 3432 4826 3542 4841
rect 11602 4868 11712 4882
rect 11602 4838 11645 4868
rect 11673 4838 11712 4868
rect 11602 4823 11712 4838
rect 14140 4865 14250 4879
rect 14140 4835 14183 4865
rect 14211 4835 14250 4865
rect 14140 4820 14250 4835
rect 8631 4495 8741 4510
rect 8631 4465 8670 4495
rect 8698 4465 8741 4495
rect 8631 4451 8741 4465
rect 9679 4491 9789 4506
rect 9679 4461 9718 4491
rect 9746 4461 9789 4491
rect 9679 4447 9789 4461
rect 19339 4489 19449 4504
rect 19339 4459 19378 4489
rect 19406 4459 19449 4489
rect 19339 4445 19449 4459
rect 20387 4485 20497 4500
rect 20387 4455 20426 4485
rect 20454 4455 20497 4485
rect 20387 4441 20497 4455
rect 895 4033 1005 4047
rect 895 4003 938 4033
rect 966 4003 1005 4033
rect 895 3988 1005 4003
rect 1943 4029 2053 4043
rect 1943 3999 1986 4029
rect 2014 3999 2053 4029
rect 1943 3984 2053 3999
rect 4845 4035 4955 4049
rect 4845 4005 4888 4035
rect 4916 4005 4955 4035
rect 4845 3990 4955 4005
rect 11603 4027 11713 4041
rect 11603 3997 11646 4027
rect 11674 3997 11713 4027
rect 11603 3982 11713 3997
rect 12651 4023 12761 4037
rect 12651 3993 12694 4023
rect 12722 3993 12761 4023
rect 12651 3978 12761 3993
rect 15553 4029 15663 4043
rect 15553 3999 15596 4029
rect 15624 3999 15663 4029
rect 15553 3984 15663 3999
rect 7142 3653 7252 3668
rect 7142 3623 7181 3653
rect 7209 3623 7252 3653
rect 7142 3609 7252 3623
rect 9680 3650 9790 3665
rect 9680 3620 9719 3650
rect 9747 3620 9790 3650
rect 9680 3606 9790 3620
rect 17850 3647 17960 3662
rect 17850 3617 17889 3647
rect 17917 3617 17960 3647
rect 17850 3603 17960 3617
rect 20388 3644 20498 3659
rect 20388 3614 20427 3644
rect 20455 3614 20498 3644
rect 20388 3600 20498 3614
rect 895 3354 1005 3368
rect 895 3324 938 3354
rect 966 3324 1005 3354
rect 895 3309 1005 3324
rect 3390 3349 3500 3363
rect 3390 3319 3433 3349
rect 3461 3319 3500 3349
rect 3390 3304 3500 3319
rect 11603 3348 11713 3362
rect 11603 3318 11646 3348
rect 11674 3318 11713 3348
rect 11603 3303 11713 3318
rect 14098 3343 14208 3357
rect 14098 3313 14141 3343
rect 14169 3313 14208 3343
rect 14098 3298 14208 3313
rect 8632 2975 8742 2990
rect 8632 2945 8671 2975
rect 8699 2945 8742 2975
rect 8632 2931 8742 2945
rect 9680 2971 9790 2986
rect 9680 2941 9719 2971
rect 9747 2941 9790 2971
rect 9680 2927 9790 2941
rect 19340 2969 19450 2984
rect 19340 2939 19379 2969
rect 19407 2939 19450 2969
rect 19340 2925 19450 2939
rect 20388 2965 20498 2980
rect 20388 2935 20427 2965
rect 20455 2935 20498 2965
rect 20388 2921 20498 2935
rect 895 2586 1005 2600
rect 895 2556 938 2586
rect 966 2556 1005 2586
rect 895 2541 1005 2556
rect 1943 2582 2053 2596
rect 1943 2552 1986 2582
rect 2014 2552 2053 2582
rect 1943 2537 2053 2552
rect 11603 2580 11713 2594
rect 11603 2550 11646 2580
rect 11674 2550 11713 2580
rect 11603 2535 11713 2550
rect 12651 2576 12761 2590
rect 12651 2546 12694 2576
rect 12722 2546 12761 2576
rect 12651 2531 12761 2546
rect 7185 2208 7295 2223
rect 7185 2178 7224 2208
rect 7252 2178 7295 2208
rect 7185 2164 7295 2178
rect 9680 2203 9790 2218
rect 9680 2173 9719 2203
rect 9747 2173 9790 2203
rect 9680 2159 9790 2173
rect 17893 2202 18003 2217
rect 17893 2172 17932 2202
rect 17960 2172 18003 2202
rect 17893 2158 18003 2172
rect 20388 2197 20498 2212
rect 20388 2167 20427 2197
rect 20455 2167 20498 2197
rect 20388 2153 20498 2167
rect 895 1907 1005 1921
rect 895 1877 938 1907
rect 966 1877 1005 1907
rect 895 1862 1005 1877
rect 11603 1901 11713 1915
rect 11603 1871 11646 1901
rect 11674 1871 11713 1901
rect 11603 1856 11713 1871
rect 8632 1528 8742 1543
rect 8632 1498 8671 1528
rect 8699 1498 8742 1528
rect 8632 1484 8742 1498
rect 9680 1524 9790 1539
rect 9680 1494 9719 1524
rect 9747 1494 9790 1524
rect 9680 1480 9790 1494
rect 19340 1522 19450 1537
rect 19340 1492 19379 1522
rect 19407 1492 19450 1522
rect 19340 1478 19450 1492
rect 20388 1518 20498 1533
rect 20388 1488 20427 1518
rect 20455 1488 20498 1518
rect 20388 1474 20498 1488
rect 10606 -252 10716 -238
rect 10606 -282 10649 -252
rect 10677 -282 10716 -252
rect 10606 -297 10716 -282
<< psubdiffcont >>
rect 9723 12942 9751 12972
rect 20431 12936 20459 12966
rect 936 12631 964 12661
rect 1984 12627 2012 12657
rect 11644 12625 11672 12655
rect 12692 12621 12720 12651
rect 8675 12267 8703 12297
rect 9723 12263 9751 12293
rect 19383 12261 19411 12291
rect 20431 12257 20459 12287
rect 936 11952 964 11982
rect 3431 11947 3459 11977
rect 11644 11946 11672 11976
rect 14139 11941 14167 11971
rect 7228 11500 7256 11530
rect 9723 11495 9751 11525
rect 17936 11494 17964 11524
rect 20431 11489 20459 11519
rect 936 11184 964 11214
rect 1984 11180 2012 11210
rect 11644 11178 11672 11208
rect 12692 11174 12720 11204
rect 8675 10820 8703 10850
rect 9723 10816 9751 10846
rect 19383 10814 19411 10844
rect 20431 10810 20459 10840
rect 936 10505 964 10535
rect 3474 10502 3502 10532
rect 11644 10499 11672 10529
rect 14182 10496 14210 10526
rect 7186 9978 7214 10008
rect 9724 9975 9752 10005
rect 17894 9972 17922 10002
rect 20432 9969 20460 9999
rect 937 9664 965 9694
rect 1985 9660 2013 9690
rect 11645 9658 11673 9688
rect 12693 9654 12721 9684
rect 8676 9300 8704 9330
rect 9724 9296 9752 9326
rect 19384 9294 19412 9324
rect 20432 9290 20460 9320
rect 937 8985 965 9015
rect 3432 8980 3460 9010
rect 11645 8979 11673 9009
rect 14140 8974 14168 9004
rect 7229 8533 7257 8563
rect 9724 8528 9752 8558
rect 17937 8527 17965 8557
rect 20432 8522 20460 8552
rect 937 8217 965 8247
rect 1985 8213 2013 8243
rect 11645 8211 11673 8241
rect 12693 8207 12721 8237
rect 8676 7853 8704 7883
rect 9724 7849 9752 7879
rect 19384 7847 19412 7877
rect 20432 7843 20460 7873
rect 937 7538 965 7568
rect 4540 7529 4568 7559
rect 11645 7532 11673 7562
rect 15248 7523 15276 7553
rect 6118 6943 6146 6973
rect 9721 6934 9749 6964
rect 16826 6937 16854 6967
rect 20429 6928 20457 6958
rect 934 6623 962 6653
rect 1982 6619 2010 6649
rect 11642 6617 11670 6647
rect 12690 6613 12718 6643
rect 8673 6259 8701 6289
rect 9721 6255 9749 6285
rect 19381 6253 19409 6283
rect 20429 6249 20457 6279
rect 934 5944 962 5974
rect 3429 5939 3457 5969
rect 11642 5938 11670 5968
rect 14137 5933 14165 5963
rect 7226 5492 7254 5522
rect 9721 5487 9749 5517
rect 17934 5486 17962 5516
rect 20429 5481 20457 5511
rect 934 5176 962 5206
rect 1982 5172 2010 5202
rect 11642 5170 11670 5200
rect 12690 5166 12718 5196
rect 8673 4812 8701 4842
rect 9721 4808 9749 4838
rect 19381 4806 19409 4836
rect 20429 4802 20457 4832
rect 934 4497 962 4527
rect 3472 4494 3500 4524
rect 11642 4491 11670 4521
rect 14180 4488 14208 4518
rect 7184 3970 7212 4000
rect 9722 3967 9750 3997
rect 935 3656 963 3686
rect 1983 3652 2011 3682
rect 17892 3964 17920 3994
rect 4885 3658 4913 3688
rect 20430 3961 20458 3991
rect 11643 3650 11671 3680
rect 12691 3646 12719 3676
rect 15593 3652 15621 3682
rect 8674 3292 8702 3322
rect 9722 3288 9750 3318
rect 19382 3286 19410 3316
rect 20430 3282 20458 3312
rect 935 2977 963 3007
rect 3430 2972 3458 3002
rect 11643 2971 11671 3001
rect 14138 2966 14166 2996
rect 7227 2525 7255 2555
rect 9722 2520 9750 2550
rect 17935 2519 17963 2549
rect 20430 2514 20458 2544
rect 935 2209 963 2239
rect 1983 2205 2011 2235
rect 11643 2203 11671 2233
rect 12691 2199 12719 2229
rect 8674 1845 8702 1875
rect 9722 1841 9750 1871
rect 19382 1839 19410 1869
rect 20430 1835 20458 1865
rect 935 1530 963 1560
rect 11643 1524 11671 1554
rect 10646 -629 10674 -599
<< nsubdiffcont >>
rect 939 12978 967 13008
rect 1987 12974 2015 13004
rect 11647 12972 11675 13002
rect 12695 12968 12723 12998
rect 9720 12595 9748 12625
rect 20428 12589 20456 12619
rect 939 12299 967 12329
rect 3434 12294 3462 12324
rect 11647 12293 11675 12323
rect 14142 12288 14170 12318
rect 8672 11920 8700 11950
rect 9720 11916 9748 11946
rect 19380 11914 19408 11944
rect 20428 11910 20456 11940
rect 939 11531 967 11561
rect 1987 11527 2015 11557
rect 11647 11525 11675 11555
rect 12695 11521 12723 11551
rect 7225 11153 7253 11183
rect 9720 11148 9748 11178
rect 17933 11147 17961 11177
rect 20428 11142 20456 11172
rect 939 10852 967 10882
rect 3477 10849 3505 10879
rect 11647 10846 11675 10876
rect 14185 10843 14213 10873
rect 8672 10473 8700 10503
rect 9720 10469 9748 10499
rect 19380 10467 19408 10497
rect 20428 10463 20456 10493
rect 940 10011 968 10041
rect 1988 10007 2016 10037
rect 11648 10005 11676 10035
rect 12696 10001 12724 10031
rect 7183 9631 7211 9661
rect 9721 9628 9749 9658
rect 17891 9625 17919 9655
rect 20429 9622 20457 9652
rect 940 9332 968 9362
rect 3435 9327 3463 9357
rect 11648 9326 11676 9356
rect 14143 9321 14171 9351
rect 8673 8953 8701 8983
rect 9721 8949 9749 8979
rect 19381 8947 19409 8977
rect 20429 8943 20457 8973
rect 940 8564 968 8594
rect 1988 8560 2016 8590
rect 11648 8558 11676 8588
rect 12696 8554 12724 8584
rect 7226 8186 7254 8216
rect 9721 8181 9749 8211
rect 17934 8180 17962 8210
rect 20429 8175 20457 8205
rect 940 7885 968 7915
rect 4543 7876 4571 7906
rect 11648 7879 11676 7909
rect 15251 7870 15279 7900
rect 8673 7506 8701 7536
rect 9721 7502 9749 7532
rect 19381 7500 19409 7530
rect 20429 7496 20457 7526
rect 937 6970 965 7000
rect 1985 6966 2013 6996
rect 11645 6964 11673 6994
rect 12693 6960 12721 6990
rect 6115 6596 6143 6626
rect 9718 6587 9746 6617
rect 16823 6590 16851 6620
rect 20426 6581 20454 6611
rect 937 6291 965 6321
rect 3432 6286 3460 6316
rect 11645 6285 11673 6315
rect 14140 6280 14168 6310
rect 8670 5912 8698 5942
rect 9718 5908 9746 5938
rect 19378 5906 19406 5936
rect 20426 5902 20454 5932
rect 937 5523 965 5553
rect 1985 5519 2013 5549
rect 11645 5517 11673 5547
rect 12693 5513 12721 5543
rect 7223 5145 7251 5175
rect 9718 5140 9746 5170
rect 17931 5139 17959 5169
rect 20426 5134 20454 5164
rect 937 4844 965 4874
rect 3475 4841 3503 4871
rect 11645 4838 11673 4868
rect 14183 4835 14211 4865
rect 8670 4465 8698 4495
rect 9718 4461 9746 4491
rect 19378 4459 19406 4489
rect 20426 4455 20454 4485
rect 938 4003 966 4033
rect 1986 3999 2014 4029
rect 4888 4005 4916 4035
rect 11646 3997 11674 4027
rect 12694 3993 12722 4023
rect 15596 3999 15624 4029
rect 7181 3623 7209 3653
rect 9719 3620 9747 3650
rect 17889 3617 17917 3647
rect 20427 3614 20455 3644
rect 938 3324 966 3354
rect 3433 3319 3461 3349
rect 11646 3318 11674 3348
rect 14141 3313 14169 3343
rect 8671 2945 8699 2975
rect 9719 2941 9747 2971
rect 19379 2939 19407 2969
rect 20427 2935 20455 2965
rect 938 2556 966 2586
rect 1986 2552 2014 2582
rect 11646 2550 11674 2580
rect 12694 2546 12722 2576
rect 7224 2178 7252 2208
rect 9719 2173 9747 2203
rect 17932 2172 17960 2202
rect 20427 2167 20455 2197
rect 938 1877 966 1907
rect 11646 1871 11674 1901
rect 8671 1498 8699 1528
rect 9719 1494 9747 1524
rect 19379 1492 19407 1522
rect 20427 1488 20455 1518
rect 10649 -282 10677 -252
<< poly >>
rect 859 12935 909 12948
rect 1072 12935 1122 12948
rect 1280 12935 1330 12948
rect 1488 12935 1538 12948
rect 1907 12931 1957 12944
rect 2120 12931 2170 12944
rect 2328 12931 2378 12944
rect 2536 12931 2586 12944
rect 859 12807 909 12835
rect 859 12787 872 12807
rect 892 12787 909 12807
rect 859 12758 909 12787
rect 1072 12806 1122 12835
rect 1072 12782 1083 12806
rect 1107 12782 1122 12806
rect 1072 12758 1122 12782
rect 1280 12811 1330 12835
rect 1280 12787 1292 12811
rect 1316 12787 1330 12811
rect 1280 12758 1330 12787
rect 1488 12809 1538 12835
rect 11567 12929 11617 12942
rect 11780 12929 11830 12942
rect 11988 12929 12038 12942
rect 12196 12929 12246 12942
rect 9149 12887 9199 12903
rect 9357 12887 9407 12903
rect 9565 12887 9615 12903
rect 9778 12887 9828 12903
rect 1488 12783 1506 12809
rect 1532 12783 1538 12809
rect 1488 12758 1538 12783
rect 1907 12803 1957 12831
rect 1907 12783 1920 12803
rect 1940 12783 1957 12803
rect 1907 12754 1957 12783
rect 2120 12802 2170 12831
rect 2120 12778 2131 12802
rect 2155 12778 2170 12802
rect 2120 12754 2170 12778
rect 2328 12807 2378 12831
rect 2328 12783 2340 12807
rect 2364 12783 2378 12807
rect 2328 12754 2378 12783
rect 2536 12805 2586 12831
rect 2536 12779 2554 12805
rect 2580 12779 2586 12805
rect 2536 12754 2586 12779
rect 9149 12820 9199 12845
rect 9149 12794 9155 12820
rect 9181 12794 9199 12820
rect 9149 12768 9199 12794
rect 9357 12816 9407 12845
rect 9357 12792 9371 12816
rect 9395 12792 9407 12816
rect 9357 12768 9407 12792
rect 9565 12821 9615 12845
rect 9565 12797 9580 12821
rect 9604 12797 9615 12821
rect 9565 12768 9615 12797
rect 9778 12816 9828 12845
rect 9778 12796 9795 12816
rect 9815 12796 9828 12816
rect 12615 12925 12665 12938
rect 12828 12925 12878 12938
rect 13036 12925 13086 12938
rect 13244 12925 13294 12938
rect 9778 12768 9828 12796
rect 859 12700 909 12716
rect 1072 12700 1122 12716
rect 1280 12700 1330 12716
rect 1488 12700 1538 12716
rect 1907 12696 1957 12712
rect 2120 12696 2170 12712
rect 2328 12696 2378 12712
rect 2536 12696 2586 12712
rect 11567 12801 11617 12829
rect 11567 12781 11580 12801
rect 11600 12781 11617 12801
rect 11567 12752 11617 12781
rect 11780 12800 11830 12829
rect 11780 12776 11791 12800
rect 11815 12776 11830 12800
rect 11780 12752 11830 12776
rect 11988 12805 12038 12829
rect 11988 12781 12000 12805
rect 12024 12781 12038 12805
rect 11988 12752 12038 12781
rect 12196 12803 12246 12829
rect 19857 12881 19907 12897
rect 20065 12881 20115 12897
rect 20273 12881 20323 12897
rect 20486 12881 20536 12897
rect 12196 12777 12214 12803
rect 12240 12777 12246 12803
rect 12196 12752 12246 12777
rect 12615 12797 12665 12825
rect 12615 12777 12628 12797
rect 12648 12777 12665 12797
rect 12615 12748 12665 12777
rect 12828 12796 12878 12825
rect 12828 12772 12839 12796
rect 12863 12772 12878 12796
rect 12828 12748 12878 12772
rect 13036 12801 13086 12825
rect 13036 12777 13048 12801
rect 13072 12777 13086 12801
rect 13036 12748 13086 12777
rect 13244 12799 13294 12825
rect 13244 12773 13262 12799
rect 13288 12773 13294 12799
rect 13244 12748 13294 12773
rect 19857 12814 19907 12839
rect 19857 12788 19863 12814
rect 19889 12788 19907 12814
rect 19857 12762 19907 12788
rect 20065 12810 20115 12839
rect 20065 12786 20079 12810
rect 20103 12786 20115 12810
rect 20065 12762 20115 12786
rect 20273 12815 20323 12839
rect 20273 12791 20288 12815
rect 20312 12791 20323 12815
rect 20273 12762 20323 12791
rect 20486 12810 20536 12839
rect 20486 12790 20503 12810
rect 20523 12790 20536 12810
rect 20486 12762 20536 12790
rect 11567 12694 11617 12710
rect 11780 12694 11830 12710
rect 11988 12694 12038 12710
rect 12196 12694 12246 12710
rect 12615 12690 12665 12706
rect 12828 12690 12878 12706
rect 13036 12690 13086 12706
rect 13244 12690 13294 12706
rect 9149 12655 9199 12668
rect 9357 12655 9407 12668
rect 9565 12655 9615 12668
rect 9778 12655 9828 12668
rect 19857 12649 19907 12662
rect 20065 12649 20115 12662
rect 20273 12649 20323 12662
rect 20486 12649 20536 12662
rect 859 12256 909 12269
rect 1072 12256 1122 12269
rect 1280 12256 1330 12269
rect 1488 12256 1538 12269
rect 3354 12251 3404 12264
rect 3567 12251 3617 12264
rect 3775 12251 3825 12264
rect 3983 12251 4033 12264
rect 859 12128 909 12156
rect 859 12108 872 12128
rect 892 12108 909 12128
rect 859 12079 909 12108
rect 1072 12127 1122 12156
rect 1072 12103 1083 12127
rect 1107 12103 1122 12127
rect 1072 12079 1122 12103
rect 1280 12132 1330 12156
rect 1280 12108 1292 12132
rect 1316 12108 1330 12132
rect 1280 12079 1330 12108
rect 1488 12130 1538 12156
rect 11567 12250 11617 12263
rect 11780 12250 11830 12263
rect 11988 12250 12038 12263
rect 12196 12250 12246 12263
rect 8101 12212 8151 12228
rect 8309 12212 8359 12228
rect 8517 12212 8567 12228
rect 8730 12212 8780 12228
rect 9149 12208 9199 12224
rect 9357 12208 9407 12224
rect 9565 12208 9615 12224
rect 9778 12208 9828 12224
rect 1488 12104 1506 12130
rect 1532 12104 1538 12130
rect 1488 12079 1538 12104
rect 3354 12123 3404 12151
rect 3354 12103 3367 12123
rect 3387 12103 3404 12123
rect 3354 12074 3404 12103
rect 3567 12122 3617 12151
rect 3567 12098 3578 12122
rect 3602 12098 3617 12122
rect 3567 12074 3617 12098
rect 3775 12127 3825 12151
rect 3775 12103 3787 12127
rect 3811 12103 3825 12127
rect 3775 12074 3825 12103
rect 3983 12125 4033 12151
rect 3983 12099 4001 12125
rect 4027 12099 4033 12125
rect 3983 12074 4033 12099
rect 8101 12145 8151 12170
rect 8101 12119 8107 12145
rect 8133 12119 8151 12145
rect 8101 12093 8151 12119
rect 8309 12141 8359 12170
rect 8309 12117 8323 12141
rect 8347 12117 8359 12141
rect 8309 12093 8359 12117
rect 8517 12146 8567 12170
rect 8517 12122 8532 12146
rect 8556 12122 8567 12146
rect 8517 12093 8567 12122
rect 8730 12141 8780 12170
rect 8730 12121 8747 12141
rect 8767 12121 8780 12141
rect 8730 12093 8780 12121
rect 9149 12141 9199 12166
rect 9149 12115 9155 12141
rect 9181 12115 9199 12141
rect 859 12021 909 12037
rect 1072 12021 1122 12037
rect 1280 12021 1330 12037
rect 1488 12021 1538 12037
rect 3354 12016 3404 12032
rect 3567 12016 3617 12032
rect 3775 12016 3825 12032
rect 3983 12016 4033 12032
rect 9149 12089 9199 12115
rect 9357 12137 9407 12166
rect 9357 12113 9371 12137
rect 9395 12113 9407 12137
rect 9357 12089 9407 12113
rect 9565 12142 9615 12166
rect 9565 12118 9580 12142
rect 9604 12118 9615 12142
rect 9565 12089 9615 12118
rect 9778 12137 9828 12166
rect 9778 12117 9795 12137
rect 9815 12117 9828 12137
rect 9778 12089 9828 12117
rect 14062 12245 14112 12258
rect 14275 12245 14325 12258
rect 14483 12245 14533 12258
rect 14691 12245 14741 12258
rect 11567 12122 11617 12150
rect 8101 11980 8151 11993
rect 8309 11980 8359 11993
rect 8517 11980 8567 11993
rect 8730 11980 8780 11993
rect 11567 12102 11580 12122
rect 11600 12102 11617 12122
rect 11567 12073 11617 12102
rect 11780 12121 11830 12150
rect 11780 12097 11791 12121
rect 11815 12097 11830 12121
rect 11780 12073 11830 12097
rect 11988 12126 12038 12150
rect 11988 12102 12000 12126
rect 12024 12102 12038 12126
rect 11988 12073 12038 12102
rect 12196 12124 12246 12150
rect 18809 12206 18859 12222
rect 19017 12206 19067 12222
rect 19225 12206 19275 12222
rect 19438 12206 19488 12222
rect 19857 12202 19907 12218
rect 20065 12202 20115 12218
rect 20273 12202 20323 12218
rect 20486 12202 20536 12218
rect 12196 12098 12214 12124
rect 12240 12098 12246 12124
rect 12196 12073 12246 12098
rect 14062 12117 14112 12145
rect 14062 12097 14075 12117
rect 14095 12097 14112 12117
rect 14062 12068 14112 12097
rect 14275 12116 14325 12145
rect 14275 12092 14286 12116
rect 14310 12092 14325 12116
rect 14275 12068 14325 12092
rect 14483 12121 14533 12145
rect 14483 12097 14495 12121
rect 14519 12097 14533 12121
rect 14483 12068 14533 12097
rect 14691 12119 14741 12145
rect 14691 12093 14709 12119
rect 14735 12093 14741 12119
rect 14691 12068 14741 12093
rect 18809 12139 18859 12164
rect 18809 12113 18815 12139
rect 18841 12113 18859 12139
rect 18809 12087 18859 12113
rect 19017 12135 19067 12164
rect 19017 12111 19031 12135
rect 19055 12111 19067 12135
rect 19017 12087 19067 12111
rect 19225 12140 19275 12164
rect 19225 12116 19240 12140
rect 19264 12116 19275 12140
rect 19225 12087 19275 12116
rect 19438 12135 19488 12164
rect 19438 12115 19455 12135
rect 19475 12115 19488 12135
rect 19438 12087 19488 12115
rect 19857 12135 19907 12160
rect 19857 12109 19863 12135
rect 19889 12109 19907 12135
rect 11567 12015 11617 12031
rect 11780 12015 11830 12031
rect 11988 12015 12038 12031
rect 12196 12015 12246 12031
rect 14062 12010 14112 12026
rect 14275 12010 14325 12026
rect 14483 12010 14533 12026
rect 14691 12010 14741 12026
rect 9149 11976 9199 11989
rect 9357 11976 9407 11989
rect 9565 11976 9615 11989
rect 9778 11976 9828 11989
rect 19857 12083 19907 12109
rect 20065 12131 20115 12160
rect 20065 12107 20079 12131
rect 20103 12107 20115 12131
rect 20065 12083 20115 12107
rect 20273 12136 20323 12160
rect 20273 12112 20288 12136
rect 20312 12112 20323 12136
rect 20273 12083 20323 12112
rect 20486 12131 20536 12160
rect 20486 12111 20503 12131
rect 20523 12111 20536 12131
rect 20486 12083 20536 12111
rect 18809 11974 18859 11987
rect 19017 11974 19067 11987
rect 19225 11974 19275 11987
rect 19438 11974 19488 11987
rect 19857 11970 19907 11983
rect 20065 11970 20115 11983
rect 20273 11970 20323 11983
rect 20486 11970 20536 11983
rect 859 11488 909 11501
rect 1072 11488 1122 11501
rect 1280 11488 1330 11501
rect 1488 11488 1538 11501
rect 1907 11484 1957 11497
rect 2120 11484 2170 11497
rect 2328 11484 2378 11497
rect 2536 11484 2586 11497
rect 859 11360 909 11388
rect 859 11340 872 11360
rect 892 11340 909 11360
rect 859 11311 909 11340
rect 1072 11359 1122 11388
rect 1072 11335 1083 11359
rect 1107 11335 1122 11359
rect 1072 11311 1122 11335
rect 1280 11364 1330 11388
rect 1280 11340 1292 11364
rect 1316 11340 1330 11364
rect 1280 11311 1330 11340
rect 1488 11362 1538 11388
rect 11567 11482 11617 11495
rect 11780 11482 11830 11495
rect 11988 11482 12038 11495
rect 12196 11482 12246 11495
rect 6654 11445 6704 11461
rect 6862 11445 6912 11461
rect 7070 11445 7120 11461
rect 7283 11445 7333 11461
rect 9149 11440 9199 11456
rect 9357 11440 9407 11456
rect 9565 11440 9615 11456
rect 9778 11440 9828 11456
rect 1488 11336 1506 11362
rect 1532 11336 1538 11362
rect 1488 11311 1538 11336
rect 1907 11356 1957 11384
rect 1907 11336 1920 11356
rect 1940 11336 1957 11356
rect 1907 11307 1957 11336
rect 2120 11355 2170 11384
rect 2120 11331 2131 11355
rect 2155 11331 2170 11355
rect 2120 11307 2170 11331
rect 2328 11360 2378 11384
rect 2328 11336 2340 11360
rect 2364 11336 2378 11360
rect 2328 11307 2378 11336
rect 2536 11358 2586 11384
rect 2536 11332 2554 11358
rect 2580 11332 2586 11358
rect 2536 11307 2586 11332
rect 6654 11378 6704 11403
rect 6654 11352 6660 11378
rect 6686 11352 6704 11378
rect 6654 11326 6704 11352
rect 6862 11374 6912 11403
rect 6862 11350 6876 11374
rect 6900 11350 6912 11374
rect 6862 11326 6912 11350
rect 7070 11379 7120 11403
rect 7070 11355 7085 11379
rect 7109 11355 7120 11379
rect 7070 11326 7120 11355
rect 7283 11374 7333 11403
rect 7283 11354 7300 11374
rect 7320 11354 7333 11374
rect 7283 11326 7333 11354
rect 9149 11373 9199 11398
rect 9149 11347 9155 11373
rect 9181 11347 9199 11373
rect 859 11253 909 11269
rect 1072 11253 1122 11269
rect 1280 11253 1330 11269
rect 1488 11253 1538 11269
rect 1907 11249 1957 11265
rect 2120 11249 2170 11265
rect 2328 11249 2378 11265
rect 2536 11249 2586 11265
rect 9149 11321 9199 11347
rect 9357 11369 9407 11398
rect 9357 11345 9371 11369
rect 9395 11345 9407 11369
rect 9357 11321 9407 11345
rect 9565 11374 9615 11398
rect 9565 11350 9580 11374
rect 9604 11350 9615 11374
rect 9565 11321 9615 11350
rect 9778 11369 9828 11398
rect 9778 11349 9795 11369
rect 9815 11349 9828 11369
rect 12615 11478 12665 11491
rect 12828 11478 12878 11491
rect 13036 11478 13086 11491
rect 13244 11478 13294 11491
rect 9778 11321 9828 11349
rect 6654 11213 6704 11226
rect 6862 11213 6912 11226
rect 7070 11213 7120 11226
rect 7283 11213 7333 11226
rect 11567 11354 11617 11382
rect 11567 11334 11580 11354
rect 11600 11334 11617 11354
rect 11567 11305 11617 11334
rect 11780 11353 11830 11382
rect 11780 11329 11791 11353
rect 11815 11329 11830 11353
rect 11780 11305 11830 11329
rect 11988 11358 12038 11382
rect 11988 11334 12000 11358
rect 12024 11334 12038 11358
rect 11988 11305 12038 11334
rect 12196 11356 12246 11382
rect 17362 11439 17412 11455
rect 17570 11439 17620 11455
rect 17778 11439 17828 11455
rect 17991 11439 18041 11455
rect 19857 11434 19907 11450
rect 20065 11434 20115 11450
rect 20273 11434 20323 11450
rect 20486 11434 20536 11450
rect 12196 11330 12214 11356
rect 12240 11330 12246 11356
rect 12196 11305 12246 11330
rect 12615 11350 12665 11378
rect 12615 11330 12628 11350
rect 12648 11330 12665 11350
rect 12615 11301 12665 11330
rect 12828 11349 12878 11378
rect 12828 11325 12839 11349
rect 12863 11325 12878 11349
rect 12828 11301 12878 11325
rect 13036 11354 13086 11378
rect 13036 11330 13048 11354
rect 13072 11330 13086 11354
rect 13036 11301 13086 11330
rect 13244 11352 13294 11378
rect 13244 11326 13262 11352
rect 13288 11326 13294 11352
rect 13244 11301 13294 11326
rect 17362 11372 17412 11397
rect 17362 11346 17368 11372
rect 17394 11346 17412 11372
rect 17362 11320 17412 11346
rect 17570 11368 17620 11397
rect 17570 11344 17584 11368
rect 17608 11344 17620 11368
rect 17570 11320 17620 11344
rect 17778 11373 17828 11397
rect 17778 11349 17793 11373
rect 17817 11349 17828 11373
rect 17778 11320 17828 11349
rect 17991 11368 18041 11397
rect 17991 11348 18008 11368
rect 18028 11348 18041 11368
rect 17991 11320 18041 11348
rect 19857 11367 19907 11392
rect 19857 11341 19863 11367
rect 19889 11341 19907 11367
rect 11567 11247 11617 11263
rect 11780 11247 11830 11263
rect 11988 11247 12038 11263
rect 12196 11247 12246 11263
rect 12615 11243 12665 11259
rect 12828 11243 12878 11259
rect 13036 11243 13086 11259
rect 13244 11243 13294 11259
rect 9149 11208 9199 11221
rect 9357 11208 9407 11221
rect 9565 11208 9615 11221
rect 9778 11208 9828 11221
rect 19857 11315 19907 11341
rect 20065 11363 20115 11392
rect 20065 11339 20079 11363
rect 20103 11339 20115 11363
rect 20065 11315 20115 11339
rect 20273 11368 20323 11392
rect 20273 11344 20288 11368
rect 20312 11344 20323 11368
rect 20273 11315 20323 11344
rect 20486 11363 20536 11392
rect 20486 11343 20503 11363
rect 20523 11343 20536 11363
rect 20486 11315 20536 11343
rect 17362 11207 17412 11220
rect 17570 11207 17620 11220
rect 17778 11207 17828 11220
rect 17991 11207 18041 11220
rect 19857 11202 19907 11215
rect 20065 11202 20115 11215
rect 20273 11202 20323 11215
rect 20486 11202 20536 11215
rect 859 10809 909 10822
rect 1072 10809 1122 10822
rect 1280 10809 1330 10822
rect 1488 10809 1538 10822
rect 3397 10806 3447 10819
rect 3610 10806 3660 10819
rect 3818 10806 3868 10819
rect 4026 10806 4076 10819
rect 859 10681 909 10709
rect 859 10661 872 10681
rect 892 10661 909 10681
rect 859 10632 909 10661
rect 1072 10680 1122 10709
rect 1072 10656 1083 10680
rect 1107 10656 1122 10680
rect 1072 10632 1122 10656
rect 1280 10685 1330 10709
rect 1280 10661 1292 10685
rect 1316 10661 1330 10685
rect 1280 10632 1330 10661
rect 1488 10683 1538 10709
rect 11567 10803 11617 10816
rect 11780 10803 11830 10816
rect 11988 10803 12038 10816
rect 12196 10803 12246 10816
rect 8101 10765 8151 10781
rect 8309 10765 8359 10781
rect 8517 10765 8567 10781
rect 8730 10765 8780 10781
rect 9149 10761 9199 10777
rect 9357 10761 9407 10777
rect 9565 10761 9615 10777
rect 9778 10761 9828 10777
rect 1488 10657 1506 10683
rect 1532 10657 1538 10683
rect 1488 10632 1538 10657
rect 3397 10678 3447 10706
rect 3397 10658 3410 10678
rect 3430 10658 3447 10678
rect 3397 10629 3447 10658
rect 3610 10677 3660 10706
rect 3610 10653 3621 10677
rect 3645 10653 3660 10677
rect 3610 10629 3660 10653
rect 3818 10682 3868 10706
rect 3818 10658 3830 10682
rect 3854 10658 3868 10682
rect 3818 10629 3868 10658
rect 4026 10680 4076 10706
rect 4026 10654 4044 10680
rect 4070 10654 4076 10680
rect 4026 10629 4076 10654
rect 8101 10698 8151 10723
rect 8101 10672 8107 10698
rect 8133 10672 8151 10698
rect 8101 10646 8151 10672
rect 8309 10694 8359 10723
rect 8309 10670 8323 10694
rect 8347 10670 8359 10694
rect 8309 10646 8359 10670
rect 8517 10699 8567 10723
rect 8517 10675 8532 10699
rect 8556 10675 8567 10699
rect 8517 10646 8567 10675
rect 8730 10694 8780 10723
rect 8730 10674 8747 10694
rect 8767 10674 8780 10694
rect 8730 10646 8780 10674
rect 9149 10694 9199 10719
rect 9149 10668 9155 10694
rect 9181 10668 9199 10694
rect 859 10574 909 10590
rect 1072 10574 1122 10590
rect 1280 10574 1330 10590
rect 1488 10574 1538 10590
rect 3397 10571 3447 10587
rect 3610 10571 3660 10587
rect 3818 10571 3868 10587
rect 4026 10571 4076 10587
rect 9149 10642 9199 10668
rect 9357 10690 9407 10719
rect 9357 10666 9371 10690
rect 9395 10666 9407 10690
rect 9357 10642 9407 10666
rect 9565 10695 9615 10719
rect 9565 10671 9580 10695
rect 9604 10671 9615 10695
rect 9565 10642 9615 10671
rect 9778 10690 9828 10719
rect 9778 10670 9795 10690
rect 9815 10670 9828 10690
rect 9778 10642 9828 10670
rect 14105 10800 14155 10813
rect 14318 10800 14368 10813
rect 14526 10800 14576 10813
rect 14734 10800 14784 10813
rect 11567 10675 11617 10703
rect 8101 10533 8151 10546
rect 8309 10533 8359 10546
rect 8517 10533 8567 10546
rect 8730 10533 8780 10546
rect 11567 10655 11580 10675
rect 11600 10655 11617 10675
rect 11567 10626 11617 10655
rect 11780 10674 11830 10703
rect 11780 10650 11791 10674
rect 11815 10650 11830 10674
rect 11780 10626 11830 10650
rect 11988 10679 12038 10703
rect 11988 10655 12000 10679
rect 12024 10655 12038 10679
rect 11988 10626 12038 10655
rect 12196 10677 12246 10703
rect 18809 10759 18859 10775
rect 19017 10759 19067 10775
rect 19225 10759 19275 10775
rect 19438 10759 19488 10775
rect 19857 10755 19907 10771
rect 20065 10755 20115 10771
rect 20273 10755 20323 10771
rect 20486 10755 20536 10771
rect 12196 10651 12214 10677
rect 12240 10651 12246 10677
rect 12196 10626 12246 10651
rect 14105 10672 14155 10700
rect 14105 10652 14118 10672
rect 14138 10652 14155 10672
rect 14105 10623 14155 10652
rect 14318 10671 14368 10700
rect 14318 10647 14329 10671
rect 14353 10647 14368 10671
rect 14318 10623 14368 10647
rect 14526 10676 14576 10700
rect 14526 10652 14538 10676
rect 14562 10652 14576 10676
rect 14526 10623 14576 10652
rect 14734 10674 14784 10700
rect 14734 10648 14752 10674
rect 14778 10648 14784 10674
rect 14734 10623 14784 10648
rect 18809 10692 18859 10717
rect 18809 10666 18815 10692
rect 18841 10666 18859 10692
rect 18809 10640 18859 10666
rect 19017 10688 19067 10717
rect 19017 10664 19031 10688
rect 19055 10664 19067 10688
rect 19017 10640 19067 10664
rect 19225 10693 19275 10717
rect 19225 10669 19240 10693
rect 19264 10669 19275 10693
rect 19225 10640 19275 10669
rect 19438 10688 19488 10717
rect 19438 10668 19455 10688
rect 19475 10668 19488 10688
rect 19438 10640 19488 10668
rect 19857 10688 19907 10713
rect 19857 10662 19863 10688
rect 19889 10662 19907 10688
rect 11567 10568 11617 10584
rect 11780 10568 11830 10584
rect 11988 10568 12038 10584
rect 12196 10568 12246 10584
rect 14105 10565 14155 10581
rect 14318 10565 14368 10581
rect 14526 10565 14576 10581
rect 14734 10565 14784 10581
rect 9149 10529 9199 10542
rect 9357 10529 9407 10542
rect 9565 10529 9615 10542
rect 9778 10529 9828 10542
rect 19857 10636 19907 10662
rect 20065 10684 20115 10713
rect 20065 10660 20079 10684
rect 20103 10660 20115 10684
rect 20065 10636 20115 10660
rect 20273 10689 20323 10713
rect 20273 10665 20288 10689
rect 20312 10665 20323 10689
rect 20273 10636 20323 10665
rect 20486 10684 20536 10713
rect 20486 10664 20503 10684
rect 20523 10664 20536 10684
rect 20486 10636 20536 10664
rect 18809 10527 18859 10540
rect 19017 10527 19067 10540
rect 19225 10527 19275 10540
rect 19438 10527 19488 10540
rect 19857 10523 19907 10536
rect 20065 10523 20115 10536
rect 20273 10523 20323 10536
rect 20486 10523 20536 10536
rect 860 9968 910 9981
rect 1073 9968 1123 9981
rect 1281 9968 1331 9981
rect 1489 9968 1539 9981
rect 1908 9964 1958 9977
rect 2121 9964 2171 9977
rect 2329 9964 2379 9977
rect 2537 9964 2587 9977
rect 860 9840 910 9868
rect 860 9820 873 9840
rect 893 9820 910 9840
rect 860 9791 910 9820
rect 1073 9839 1123 9868
rect 1073 9815 1084 9839
rect 1108 9815 1123 9839
rect 1073 9791 1123 9815
rect 1281 9844 1331 9868
rect 1281 9820 1293 9844
rect 1317 9820 1331 9844
rect 1281 9791 1331 9820
rect 1489 9842 1539 9868
rect 11568 9962 11618 9975
rect 11781 9962 11831 9975
rect 11989 9962 12039 9975
rect 12197 9962 12247 9975
rect 6612 9923 6662 9939
rect 6820 9923 6870 9939
rect 7028 9923 7078 9939
rect 7241 9923 7291 9939
rect 9150 9920 9200 9936
rect 9358 9920 9408 9936
rect 9566 9920 9616 9936
rect 9779 9920 9829 9936
rect 1489 9816 1507 9842
rect 1533 9816 1539 9842
rect 1489 9791 1539 9816
rect 1908 9836 1958 9864
rect 1908 9816 1921 9836
rect 1941 9816 1958 9836
rect 1908 9787 1958 9816
rect 2121 9835 2171 9864
rect 2121 9811 2132 9835
rect 2156 9811 2171 9835
rect 2121 9787 2171 9811
rect 2329 9840 2379 9864
rect 2329 9816 2341 9840
rect 2365 9816 2379 9840
rect 2329 9787 2379 9816
rect 2537 9838 2587 9864
rect 2537 9812 2555 9838
rect 2581 9812 2587 9838
rect 2537 9787 2587 9812
rect 6612 9856 6662 9881
rect 6612 9830 6618 9856
rect 6644 9830 6662 9856
rect 6612 9804 6662 9830
rect 6820 9852 6870 9881
rect 6820 9828 6834 9852
rect 6858 9828 6870 9852
rect 6820 9804 6870 9828
rect 7028 9857 7078 9881
rect 7028 9833 7043 9857
rect 7067 9833 7078 9857
rect 7028 9804 7078 9833
rect 7241 9852 7291 9881
rect 7241 9832 7258 9852
rect 7278 9832 7291 9852
rect 7241 9804 7291 9832
rect 9150 9853 9200 9878
rect 9150 9827 9156 9853
rect 9182 9827 9200 9853
rect 860 9733 910 9749
rect 1073 9733 1123 9749
rect 1281 9733 1331 9749
rect 1489 9733 1539 9749
rect 1908 9729 1958 9745
rect 2121 9729 2171 9745
rect 2329 9729 2379 9745
rect 2537 9729 2587 9745
rect 9150 9801 9200 9827
rect 9358 9849 9408 9878
rect 9358 9825 9372 9849
rect 9396 9825 9408 9849
rect 9358 9801 9408 9825
rect 9566 9854 9616 9878
rect 9566 9830 9581 9854
rect 9605 9830 9616 9854
rect 9566 9801 9616 9830
rect 9779 9849 9829 9878
rect 9779 9829 9796 9849
rect 9816 9829 9829 9849
rect 12616 9958 12666 9971
rect 12829 9958 12879 9971
rect 13037 9958 13087 9971
rect 13245 9958 13295 9971
rect 9779 9801 9829 9829
rect 6612 9691 6662 9704
rect 6820 9691 6870 9704
rect 7028 9691 7078 9704
rect 7241 9691 7291 9704
rect 11568 9834 11618 9862
rect 11568 9814 11581 9834
rect 11601 9814 11618 9834
rect 11568 9785 11618 9814
rect 11781 9833 11831 9862
rect 11781 9809 11792 9833
rect 11816 9809 11831 9833
rect 11781 9785 11831 9809
rect 11989 9838 12039 9862
rect 11989 9814 12001 9838
rect 12025 9814 12039 9838
rect 11989 9785 12039 9814
rect 12197 9836 12247 9862
rect 17320 9917 17370 9933
rect 17528 9917 17578 9933
rect 17736 9917 17786 9933
rect 17949 9917 17999 9933
rect 19858 9914 19908 9930
rect 20066 9914 20116 9930
rect 20274 9914 20324 9930
rect 20487 9914 20537 9930
rect 12197 9810 12215 9836
rect 12241 9810 12247 9836
rect 12197 9785 12247 9810
rect 12616 9830 12666 9858
rect 12616 9810 12629 9830
rect 12649 9810 12666 9830
rect 12616 9781 12666 9810
rect 12829 9829 12879 9858
rect 12829 9805 12840 9829
rect 12864 9805 12879 9829
rect 12829 9781 12879 9805
rect 13037 9834 13087 9858
rect 13037 9810 13049 9834
rect 13073 9810 13087 9834
rect 13037 9781 13087 9810
rect 13245 9832 13295 9858
rect 13245 9806 13263 9832
rect 13289 9806 13295 9832
rect 13245 9781 13295 9806
rect 17320 9850 17370 9875
rect 17320 9824 17326 9850
rect 17352 9824 17370 9850
rect 17320 9798 17370 9824
rect 17528 9846 17578 9875
rect 17528 9822 17542 9846
rect 17566 9822 17578 9846
rect 17528 9798 17578 9822
rect 17736 9851 17786 9875
rect 17736 9827 17751 9851
rect 17775 9827 17786 9851
rect 17736 9798 17786 9827
rect 17949 9846 17999 9875
rect 17949 9826 17966 9846
rect 17986 9826 17999 9846
rect 17949 9798 17999 9826
rect 19858 9847 19908 9872
rect 19858 9821 19864 9847
rect 19890 9821 19908 9847
rect 11568 9727 11618 9743
rect 11781 9727 11831 9743
rect 11989 9727 12039 9743
rect 12197 9727 12247 9743
rect 12616 9723 12666 9739
rect 12829 9723 12879 9739
rect 13037 9723 13087 9739
rect 13245 9723 13295 9739
rect 9150 9688 9200 9701
rect 9358 9688 9408 9701
rect 9566 9688 9616 9701
rect 9779 9688 9829 9701
rect 19858 9795 19908 9821
rect 20066 9843 20116 9872
rect 20066 9819 20080 9843
rect 20104 9819 20116 9843
rect 20066 9795 20116 9819
rect 20274 9848 20324 9872
rect 20274 9824 20289 9848
rect 20313 9824 20324 9848
rect 20274 9795 20324 9824
rect 20487 9843 20537 9872
rect 20487 9823 20504 9843
rect 20524 9823 20537 9843
rect 20487 9795 20537 9823
rect 17320 9685 17370 9698
rect 17528 9685 17578 9698
rect 17736 9685 17786 9698
rect 17949 9685 17999 9698
rect 19858 9682 19908 9695
rect 20066 9682 20116 9695
rect 20274 9682 20324 9695
rect 20487 9682 20537 9695
rect 860 9289 910 9302
rect 1073 9289 1123 9302
rect 1281 9289 1331 9302
rect 1489 9289 1539 9302
rect 3355 9284 3405 9297
rect 3568 9284 3618 9297
rect 3776 9284 3826 9297
rect 3984 9284 4034 9297
rect 860 9161 910 9189
rect 860 9141 873 9161
rect 893 9141 910 9161
rect 860 9112 910 9141
rect 1073 9160 1123 9189
rect 1073 9136 1084 9160
rect 1108 9136 1123 9160
rect 1073 9112 1123 9136
rect 1281 9165 1331 9189
rect 1281 9141 1293 9165
rect 1317 9141 1331 9165
rect 1281 9112 1331 9141
rect 1489 9163 1539 9189
rect 11568 9283 11618 9296
rect 11781 9283 11831 9296
rect 11989 9283 12039 9296
rect 12197 9283 12247 9296
rect 8102 9245 8152 9261
rect 8310 9245 8360 9261
rect 8518 9245 8568 9261
rect 8731 9245 8781 9261
rect 9150 9241 9200 9257
rect 9358 9241 9408 9257
rect 9566 9241 9616 9257
rect 9779 9241 9829 9257
rect 1489 9137 1507 9163
rect 1533 9137 1539 9163
rect 1489 9112 1539 9137
rect 3355 9156 3405 9184
rect 3355 9136 3368 9156
rect 3388 9136 3405 9156
rect 3355 9107 3405 9136
rect 3568 9155 3618 9184
rect 3568 9131 3579 9155
rect 3603 9131 3618 9155
rect 3568 9107 3618 9131
rect 3776 9160 3826 9184
rect 3776 9136 3788 9160
rect 3812 9136 3826 9160
rect 3776 9107 3826 9136
rect 3984 9158 4034 9184
rect 3984 9132 4002 9158
rect 4028 9132 4034 9158
rect 3984 9107 4034 9132
rect 8102 9178 8152 9203
rect 8102 9152 8108 9178
rect 8134 9152 8152 9178
rect 8102 9126 8152 9152
rect 8310 9174 8360 9203
rect 8310 9150 8324 9174
rect 8348 9150 8360 9174
rect 8310 9126 8360 9150
rect 8518 9179 8568 9203
rect 8518 9155 8533 9179
rect 8557 9155 8568 9179
rect 8518 9126 8568 9155
rect 8731 9174 8781 9203
rect 8731 9154 8748 9174
rect 8768 9154 8781 9174
rect 8731 9126 8781 9154
rect 9150 9174 9200 9199
rect 9150 9148 9156 9174
rect 9182 9148 9200 9174
rect 860 9054 910 9070
rect 1073 9054 1123 9070
rect 1281 9054 1331 9070
rect 1489 9054 1539 9070
rect 3355 9049 3405 9065
rect 3568 9049 3618 9065
rect 3776 9049 3826 9065
rect 3984 9049 4034 9065
rect 9150 9122 9200 9148
rect 9358 9170 9408 9199
rect 9358 9146 9372 9170
rect 9396 9146 9408 9170
rect 9358 9122 9408 9146
rect 9566 9175 9616 9199
rect 9566 9151 9581 9175
rect 9605 9151 9616 9175
rect 9566 9122 9616 9151
rect 9779 9170 9829 9199
rect 9779 9150 9796 9170
rect 9816 9150 9829 9170
rect 9779 9122 9829 9150
rect 14063 9278 14113 9291
rect 14276 9278 14326 9291
rect 14484 9278 14534 9291
rect 14692 9278 14742 9291
rect 11568 9155 11618 9183
rect 8102 9013 8152 9026
rect 8310 9013 8360 9026
rect 8518 9013 8568 9026
rect 8731 9013 8781 9026
rect 11568 9135 11581 9155
rect 11601 9135 11618 9155
rect 11568 9106 11618 9135
rect 11781 9154 11831 9183
rect 11781 9130 11792 9154
rect 11816 9130 11831 9154
rect 11781 9106 11831 9130
rect 11989 9159 12039 9183
rect 11989 9135 12001 9159
rect 12025 9135 12039 9159
rect 11989 9106 12039 9135
rect 12197 9157 12247 9183
rect 18810 9239 18860 9255
rect 19018 9239 19068 9255
rect 19226 9239 19276 9255
rect 19439 9239 19489 9255
rect 19858 9235 19908 9251
rect 20066 9235 20116 9251
rect 20274 9235 20324 9251
rect 20487 9235 20537 9251
rect 12197 9131 12215 9157
rect 12241 9131 12247 9157
rect 12197 9106 12247 9131
rect 14063 9150 14113 9178
rect 14063 9130 14076 9150
rect 14096 9130 14113 9150
rect 14063 9101 14113 9130
rect 14276 9149 14326 9178
rect 14276 9125 14287 9149
rect 14311 9125 14326 9149
rect 14276 9101 14326 9125
rect 14484 9154 14534 9178
rect 14484 9130 14496 9154
rect 14520 9130 14534 9154
rect 14484 9101 14534 9130
rect 14692 9152 14742 9178
rect 14692 9126 14710 9152
rect 14736 9126 14742 9152
rect 14692 9101 14742 9126
rect 18810 9172 18860 9197
rect 18810 9146 18816 9172
rect 18842 9146 18860 9172
rect 18810 9120 18860 9146
rect 19018 9168 19068 9197
rect 19018 9144 19032 9168
rect 19056 9144 19068 9168
rect 19018 9120 19068 9144
rect 19226 9173 19276 9197
rect 19226 9149 19241 9173
rect 19265 9149 19276 9173
rect 19226 9120 19276 9149
rect 19439 9168 19489 9197
rect 19439 9148 19456 9168
rect 19476 9148 19489 9168
rect 19439 9120 19489 9148
rect 19858 9168 19908 9193
rect 19858 9142 19864 9168
rect 19890 9142 19908 9168
rect 11568 9048 11618 9064
rect 11781 9048 11831 9064
rect 11989 9048 12039 9064
rect 12197 9048 12247 9064
rect 14063 9043 14113 9059
rect 14276 9043 14326 9059
rect 14484 9043 14534 9059
rect 14692 9043 14742 9059
rect 9150 9009 9200 9022
rect 9358 9009 9408 9022
rect 9566 9009 9616 9022
rect 9779 9009 9829 9022
rect 19858 9116 19908 9142
rect 20066 9164 20116 9193
rect 20066 9140 20080 9164
rect 20104 9140 20116 9164
rect 20066 9116 20116 9140
rect 20274 9169 20324 9193
rect 20274 9145 20289 9169
rect 20313 9145 20324 9169
rect 20274 9116 20324 9145
rect 20487 9164 20537 9193
rect 20487 9144 20504 9164
rect 20524 9144 20537 9164
rect 20487 9116 20537 9144
rect 18810 9007 18860 9020
rect 19018 9007 19068 9020
rect 19226 9007 19276 9020
rect 19439 9007 19489 9020
rect 19858 9003 19908 9016
rect 20066 9003 20116 9016
rect 20274 9003 20324 9016
rect 20487 9003 20537 9016
rect 860 8521 910 8534
rect 1073 8521 1123 8534
rect 1281 8521 1331 8534
rect 1489 8521 1539 8534
rect 1908 8517 1958 8530
rect 2121 8517 2171 8530
rect 2329 8517 2379 8530
rect 2537 8517 2587 8530
rect 860 8393 910 8421
rect 860 8373 873 8393
rect 893 8373 910 8393
rect 860 8344 910 8373
rect 1073 8392 1123 8421
rect 1073 8368 1084 8392
rect 1108 8368 1123 8392
rect 1073 8344 1123 8368
rect 1281 8397 1331 8421
rect 1281 8373 1293 8397
rect 1317 8373 1331 8397
rect 1281 8344 1331 8373
rect 1489 8395 1539 8421
rect 11568 8515 11618 8528
rect 11781 8515 11831 8528
rect 11989 8515 12039 8528
rect 12197 8515 12247 8528
rect 6655 8478 6705 8494
rect 6863 8478 6913 8494
rect 7071 8478 7121 8494
rect 7284 8478 7334 8494
rect 9150 8473 9200 8489
rect 9358 8473 9408 8489
rect 9566 8473 9616 8489
rect 9779 8473 9829 8489
rect 1489 8369 1507 8395
rect 1533 8369 1539 8395
rect 1489 8344 1539 8369
rect 1908 8389 1958 8417
rect 1908 8369 1921 8389
rect 1941 8369 1958 8389
rect 1908 8340 1958 8369
rect 2121 8388 2171 8417
rect 2121 8364 2132 8388
rect 2156 8364 2171 8388
rect 2121 8340 2171 8364
rect 2329 8393 2379 8417
rect 2329 8369 2341 8393
rect 2365 8369 2379 8393
rect 2329 8340 2379 8369
rect 2537 8391 2587 8417
rect 2537 8365 2555 8391
rect 2581 8365 2587 8391
rect 2537 8340 2587 8365
rect 6655 8411 6705 8436
rect 6655 8385 6661 8411
rect 6687 8385 6705 8411
rect 6655 8359 6705 8385
rect 6863 8407 6913 8436
rect 6863 8383 6877 8407
rect 6901 8383 6913 8407
rect 6863 8359 6913 8383
rect 7071 8412 7121 8436
rect 7071 8388 7086 8412
rect 7110 8388 7121 8412
rect 7071 8359 7121 8388
rect 7284 8407 7334 8436
rect 7284 8387 7301 8407
rect 7321 8387 7334 8407
rect 7284 8359 7334 8387
rect 9150 8406 9200 8431
rect 9150 8380 9156 8406
rect 9182 8380 9200 8406
rect 860 8286 910 8302
rect 1073 8286 1123 8302
rect 1281 8286 1331 8302
rect 1489 8286 1539 8302
rect 1908 8282 1958 8298
rect 2121 8282 2171 8298
rect 2329 8282 2379 8298
rect 2537 8282 2587 8298
rect 9150 8354 9200 8380
rect 9358 8402 9408 8431
rect 9358 8378 9372 8402
rect 9396 8378 9408 8402
rect 9358 8354 9408 8378
rect 9566 8407 9616 8431
rect 9566 8383 9581 8407
rect 9605 8383 9616 8407
rect 9566 8354 9616 8383
rect 9779 8402 9829 8431
rect 9779 8382 9796 8402
rect 9816 8382 9829 8402
rect 12616 8511 12666 8524
rect 12829 8511 12879 8524
rect 13037 8511 13087 8524
rect 13245 8511 13295 8524
rect 9779 8354 9829 8382
rect 6655 8246 6705 8259
rect 6863 8246 6913 8259
rect 7071 8246 7121 8259
rect 7284 8246 7334 8259
rect 11568 8387 11618 8415
rect 11568 8367 11581 8387
rect 11601 8367 11618 8387
rect 11568 8338 11618 8367
rect 11781 8386 11831 8415
rect 11781 8362 11792 8386
rect 11816 8362 11831 8386
rect 11781 8338 11831 8362
rect 11989 8391 12039 8415
rect 11989 8367 12001 8391
rect 12025 8367 12039 8391
rect 11989 8338 12039 8367
rect 12197 8389 12247 8415
rect 17363 8472 17413 8488
rect 17571 8472 17621 8488
rect 17779 8472 17829 8488
rect 17992 8472 18042 8488
rect 19858 8467 19908 8483
rect 20066 8467 20116 8483
rect 20274 8467 20324 8483
rect 20487 8467 20537 8483
rect 12197 8363 12215 8389
rect 12241 8363 12247 8389
rect 12197 8338 12247 8363
rect 12616 8383 12666 8411
rect 12616 8363 12629 8383
rect 12649 8363 12666 8383
rect 12616 8334 12666 8363
rect 12829 8382 12879 8411
rect 12829 8358 12840 8382
rect 12864 8358 12879 8382
rect 12829 8334 12879 8358
rect 13037 8387 13087 8411
rect 13037 8363 13049 8387
rect 13073 8363 13087 8387
rect 13037 8334 13087 8363
rect 13245 8385 13295 8411
rect 13245 8359 13263 8385
rect 13289 8359 13295 8385
rect 13245 8334 13295 8359
rect 17363 8405 17413 8430
rect 17363 8379 17369 8405
rect 17395 8379 17413 8405
rect 17363 8353 17413 8379
rect 17571 8401 17621 8430
rect 17571 8377 17585 8401
rect 17609 8377 17621 8401
rect 17571 8353 17621 8377
rect 17779 8406 17829 8430
rect 17779 8382 17794 8406
rect 17818 8382 17829 8406
rect 17779 8353 17829 8382
rect 17992 8401 18042 8430
rect 17992 8381 18009 8401
rect 18029 8381 18042 8401
rect 17992 8353 18042 8381
rect 19858 8400 19908 8425
rect 19858 8374 19864 8400
rect 19890 8374 19908 8400
rect 11568 8280 11618 8296
rect 11781 8280 11831 8296
rect 11989 8280 12039 8296
rect 12197 8280 12247 8296
rect 12616 8276 12666 8292
rect 12829 8276 12879 8292
rect 13037 8276 13087 8292
rect 13245 8276 13295 8292
rect 9150 8241 9200 8254
rect 9358 8241 9408 8254
rect 9566 8241 9616 8254
rect 9779 8241 9829 8254
rect 19858 8348 19908 8374
rect 20066 8396 20116 8425
rect 20066 8372 20080 8396
rect 20104 8372 20116 8396
rect 20066 8348 20116 8372
rect 20274 8401 20324 8425
rect 20274 8377 20289 8401
rect 20313 8377 20324 8401
rect 20274 8348 20324 8377
rect 20487 8396 20537 8425
rect 20487 8376 20504 8396
rect 20524 8376 20537 8396
rect 20487 8348 20537 8376
rect 17363 8240 17413 8253
rect 17571 8240 17621 8253
rect 17779 8240 17829 8253
rect 17992 8240 18042 8253
rect 19858 8235 19908 8248
rect 20066 8235 20116 8248
rect 20274 8235 20324 8248
rect 20487 8235 20537 8248
rect 860 7842 910 7855
rect 1073 7842 1123 7855
rect 1281 7842 1331 7855
rect 1489 7842 1539 7855
rect 4463 7833 4513 7846
rect 4676 7833 4726 7846
rect 4884 7833 4934 7846
rect 5092 7833 5142 7846
rect 11568 7836 11618 7849
rect 11781 7836 11831 7849
rect 11989 7836 12039 7849
rect 12197 7836 12247 7849
rect 860 7714 910 7742
rect 860 7694 873 7714
rect 893 7694 910 7714
rect 860 7665 910 7694
rect 1073 7713 1123 7742
rect 1073 7689 1084 7713
rect 1108 7689 1123 7713
rect 1073 7665 1123 7689
rect 1281 7718 1331 7742
rect 1281 7694 1293 7718
rect 1317 7694 1331 7718
rect 1281 7665 1331 7694
rect 1489 7716 1539 7742
rect 8102 7798 8152 7814
rect 8310 7798 8360 7814
rect 8518 7798 8568 7814
rect 8731 7798 8781 7814
rect 9150 7794 9200 7810
rect 9358 7794 9408 7810
rect 9566 7794 9616 7810
rect 9779 7794 9829 7810
rect 1489 7690 1507 7716
rect 1533 7690 1539 7716
rect 1489 7665 1539 7690
rect 4463 7705 4513 7733
rect 4463 7685 4476 7705
rect 4496 7685 4513 7705
rect 4463 7656 4513 7685
rect 4676 7704 4726 7733
rect 4676 7680 4687 7704
rect 4711 7680 4726 7704
rect 4676 7656 4726 7680
rect 4884 7709 4934 7733
rect 4884 7685 4896 7709
rect 4920 7685 4934 7709
rect 4884 7656 4934 7685
rect 5092 7707 5142 7733
rect 5092 7681 5110 7707
rect 5136 7681 5142 7707
rect 5092 7656 5142 7681
rect 8102 7731 8152 7756
rect 8102 7705 8108 7731
rect 8134 7705 8152 7731
rect 8102 7679 8152 7705
rect 8310 7727 8360 7756
rect 8310 7703 8324 7727
rect 8348 7703 8360 7727
rect 8310 7679 8360 7703
rect 8518 7732 8568 7756
rect 8518 7708 8533 7732
rect 8557 7708 8568 7732
rect 8518 7679 8568 7708
rect 8731 7727 8781 7756
rect 8731 7707 8748 7727
rect 8768 7707 8781 7727
rect 8731 7679 8781 7707
rect 9150 7727 9200 7752
rect 9150 7701 9156 7727
rect 9182 7701 9200 7727
rect 860 7607 910 7623
rect 1073 7607 1123 7623
rect 1281 7607 1331 7623
rect 1489 7607 1539 7623
rect 4463 7598 4513 7614
rect 4676 7598 4726 7614
rect 4884 7598 4934 7614
rect 5092 7598 5142 7614
rect 9150 7675 9200 7701
rect 9358 7723 9408 7752
rect 9358 7699 9372 7723
rect 9396 7699 9408 7723
rect 9358 7675 9408 7699
rect 9566 7728 9616 7752
rect 9566 7704 9581 7728
rect 9605 7704 9616 7728
rect 9566 7675 9616 7704
rect 9779 7723 9829 7752
rect 9779 7703 9796 7723
rect 9816 7703 9829 7723
rect 9779 7675 9829 7703
rect 15171 7827 15221 7840
rect 15384 7827 15434 7840
rect 15592 7827 15642 7840
rect 15800 7827 15850 7840
rect 11568 7708 11618 7736
rect 8102 7566 8152 7579
rect 8310 7566 8360 7579
rect 8518 7566 8568 7579
rect 8731 7566 8781 7579
rect 11568 7688 11581 7708
rect 11601 7688 11618 7708
rect 11568 7659 11618 7688
rect 11781 7707 11831 7736
rect 11781 7683 11792 7707
rect 11816 7683 11831 7707
rect 11781 7659 11831 7683
rect 11989 7712 12039 7736
rect 11989 7688 12001 7712
rect 12025 7688 12039 7712
rect 11989 7659 12039 7688
rect 12197 7710 12247 7736
rect 18810 7792 18860 7808
rect 19018 7792 19068 7808
rect 19226 7792 19276 7808
rect 19439 7792 19489 7808
rect 19858 7788 19908 7804
rect 20066 7788 20116 7804
rect 20274 7788 20324 7804
rect 20487 7788 20537 7804
rect 12197 7684 12215 7710
rect 12241 7684 12247 7710
rect 12197 7659 12247 7684
rect 15171 7699 15221 7727
rect 15171 7679 15184 7699
rect 15204 7679 15221 7699
rect 15171 7650 15221 7679
rect 15384 7698 15434 7727
rect 15384 7674 15395 7698
rect 15419 7674 15434 7698
rect 15384 7650 15434 7674
rect 15592 7703 15642 7727
rect 15592 7679 15604 7703
rect 15628 7679 15642 7703
rect 15592 7650 15642 7679
rect 15800 7701 15850 7727
rect 15800 7675 15818 7701
rect 15844 7675 15850 7701
rect 15800 7650 15850 7675
rect 18810 7725 18860 7750
rect 18810 7699 18816 7725
rect 18842 7699 18860 7725
rect 18810 7673 18860 7699
rect 19018 7721 19068 7750
rect 19018 7697 19032 7721
rect 19056 7697 19068 7721
rect 19018 7673 19068 7697
rect 19226 7726 19276 7750
rect 19226 7702 19241 7726
rect 19265 7702 19276 7726
rect 19226 7673 19276 7702
rect 19439 7721 19489 7750
rect 19439 7701 19456 7721
rect 19476 7701 19489 7721
rect 19439 7673 19489 7701
rect 19858 7721 19908 7746
rect 19858 7695 19864 7721
rect 19890 7695 19908 7721
rect 11568 7601 11618 7617
rect 11781 7601 11831 7617
rect 11989 7601 12039 7617
rect 12197 7601 12247 7617
rect 15171 7592 15221 7608
rect 15384 7592 15434 7608
rect 15592 7592 15642 7608
rect 15800 7592 15850 7608
rect 9150 7562 9200 7575
rect 9358 7562 9408 7575
rect 9566 7562 9616 7575
rect 9779 7562 9829 7575
rect 19858 7669 19908 7695
rect 20066 7717 20116 7746
rect 20066 7693 20080 7717
rect 20104 7693 20116 7717
rect 20066 7669 20116 7693
rect 20274 7722 20324 7746
rect 20274 7698 20289 7722
rect 20313 7698 20324 7722
rect 20274 7669 20324 7698
rect 20487 7717 20537 7746
rect 20487 7697 20504 7717
rect 20524 7697 20537 7717
rect 20487 7669 20537 7697
rect 18810 7560 18860 7573
rect 19018 7560 19068 7573
rect 19226 7560 19276 7573
rect 19439 7560 19489 7573
rect 19858 7556 19908 7569
rect 20066 7556 20116 7569
rect 20274 7556 20324 7569
rect 20487 7556 20537 7569
rect 857 6927 907 6940
rect 1070 6927 1120 6940
rect 1278 6927 1328 6940
rect 1486 6927 1536 6940
rect 1905 6923 1955 6936
rect 2118 6923 2168 6936
rect 2326 6923 2376 6936
rect 2534 6923 2584 6936
rect 857 6799 907 6827
rect 857 6779 870 6799
rect 890 6779 907 6799
rect 857 6750 907 6779
rect 1070 6798 1120 6827
rect 1070 6774 1081 6798
rect 1105 6774 1120 6798
rect 1070 6750 1120 6774
rect 1278 6803 1328 6827
rect 1278 6779 1290 6803
rect 1314 6779 1328 6803
rect 1278 6750 1328 6779
rect 1486 6801 1536 6827
rect 11565 6921 11615 6934
rect 11778 6921 11828 6934
rect 11986 6921 12036 6934
rect 12194 6921 12244 6934
rect 5544 6888 5594 6904
rect 5752 6888 5802 6904
rect 5960 6888 6010 6904
rect 6173 6888 6223 6904
rect 9147 6879 9197 6895
rect 9355 6879 9405 6895
rect 9563 6879 9613 6895
rect 9776 6879 9826 6895
rect 1486 6775 1504 6801
rect 1530 6775 1536 6801
rect 1486 6750 1536 6775
rect 1905 6795 1955 6823
rect 1905 6775 1918 6795
rect 1938 6775 1955 6795
rect 1905 6746 1955 6775
rect 2118 6794 2168 6823
rect 2118 6770 2129 6794
rect 2153 6770 2168 6794
rect 2118 6746 2168 6770
rect 2326 6799 2376 6823
rect 2326 6775 2338 6799
rect 2362 6775 2376 6799
rect 2326 6746 2376 6775
rect 2534 6797 2584 6823
rect 2534 6771 2552 6797
rect 2578 6771 2584 6797
rect 2534 6746 2584 6771
rect 5544 6821 5594 6846
rect 5544 6795 5550 6821
rect 5576 6795 5594 6821
rect 5544 6769 5594 6795
rect 5752 6817 5802 6846
rect 5752 6793 5766 6817
rect 5790 6793 5802 6817
rect 5752 6769 5802 6793
rect 5960 6822 6010 6846
rect 5960 6798 5975 6822
rect 5999 6798 6010 6822
rect 5960 6769 6010 6798
rect 6173 6817 6223 6846
rect 6173 6797 6190 6817
rect 6210 6797 6223 6817
rect 6173 6769 6223 6797
rect 9147 6812 9197 6837
rect 9147 6786 9153 6812
rect 9179 6786 9197 6812
rect 857 6692 907 6708
rect 1070 6692 1120 6708
rect 1278 6692 1328 6708
rect 1486 6692 1536 6708
rect 1905 6688 1955 6704
rect 2118 6688 2168 6704
rect 2326 6688 2376 6704
rect 2534 6688 2584 6704
rect 9147 6760 9197 6786
rect 9355 6808 9405 6837
rect 9355 6784 9369 6808
rect 9393 6784 9405 6808
rect 9355 6760 9405 6784
rect 9563 6813 9613 6837
rect 9563 6789 9578 6813
rect 9602 6789 9613 6813
rect 9563 6760 9613 6789
rect 9776 6808 9826 6837
rect 9776 6788 9793 6808
rect 9813 6788 9826 6808
rect 12613 6917 12663 6930
rect 12826 6917 12876 6930
rect 13034 6917 13084 6930
rect 13242 6917 13292 6930
rect 9776 6760 9826 6788
rect 5544 6656 5594 6669
rect 5752 6656 5802 6669
rect 5960 6656 6010 6669
rect 6173 6656 6223 6669
rect 11565 6793 11615 6821
rect 11565 6773 11578 6793
rect 11598 6773 11615 6793
rect 11565 6744 11615 6773
rect 11778 6792 11828 6821
rect 11778 6768 11789 6792
rect 11813 6768 11828 6792
rect 11778 6744 11828 6768
rect 11986 6797 12036 6821
rect 11986 6773 11998 6797
rect 12022 6773 12036 6797
rect 11986 6744 12036 6773
rect 12194 6795 12244 6821
rect 16252 6882 16302 6898
rect 16460 6882 16510 6898
rect 16668 6882 16718 6898
rect 16881 6882 16931 6898
rect 19855 6873 19905 6889
rect 20063 6873 20113 6889
rect 20271 6873 20321 6889
rect 20484 6873 20534 6889
rect 12194 6769 12212 6795
rect 12238 6769 12244 6795
rect 12194 6744 12244 6769
rect 12613 6789 12663 6817
rect 12613 6769 12626 6789
rect 12646 6769 12663 6789
rect 12613 6740 12663 6769
rect 12826 6788 12876 6817
rect 12826 6764 12837 6788
rect 12861 6764 12876 6788
rect 12826 6740 12876 6764
rect 13034 6793 13084 6817
rect 13034 6769 13046 6793
rect 13070 6769 13084 6793
rect 13034 6740 13084 6769
rect 13242 6791 13292 6817
rect 13242 6765 13260 6791
rect 13286 6765 13292 6791
rect 13242 6740 13292 6765
rect 16252 6815 16302 6840
rect 16252 6789 16258 6815
rect 16284 6789 16302 6815
rect 16252 6763 16302 6789
rect 16460 6811 16510 6840
rect 16460 6787 16474 6811
rect 16498 6787 16510 6811
rect 16460 6763 16510 6787
rect 16668 6816 16718 6840
rect 16668 6792 16683 6816
rect 16707 6792 16718 6816
rect 16668 6763 16718 6792
rect 16881 6811 16931 6840
rect 16881 6791 16898 6811
rect 16918 6791 16931 6811
rect 16881 6763 16931 6791
rect 19855 6806 19905 6831
rect 19855 6780 19861 6806
rect 19887 6780 19905 6806
rect 11565 6686 11615 6702
rect 11778 6686 11828 6702
rect 11986 6686 12036 6702
rect 12194 6686 12244 6702
rect 12613 6682 12663 6698
rect 12826 6682 12876 6698
rect 13034 6682 13084 6698
rect 13242 6682 13292 6698
rect 19855 6754 19905 6780
rect 20063 6802 20113 6831
rect 20063 6778 20077 6802
rect 20101 6778 20113 6802
rect 20063 6754 20113 6778
rect 20271 6807 20321 6831
rect 20271 6783 20286 6807
rect 20310 6783 20321 6807
rect 20271 6754 20321 6783
rect 20484 6802 20534 6831
rect 20484 6782 20501 6802
rect 20521 6782 20534 6802
rect 20484 6754 20534 6782
rect 9147 6647 9197 6660
rect 9355 6647 9405 6660
rect 9563 6647 9613 6660
rect 9776 6647 9826 6660
rect 16252 6650 16302 6663
rect 16460 6650 16510 6663
rect 16668 6650 16718 6663
rect 16881 6650 16931 6663
rect 19855 6641 19905 6654
rect 20063 6641 20113 6654
rect 20271 6641 20321 6654
rect 20484 6641 20534 6654
rect 857 6248 907 6261
rect 1070 6248 1120 6261
rect 1278 6248 1328 6261
rect 1486 6248 1536 6261
rect 3352 6243 3402 6256
rect 3565 6243 3615 6256
rect 3773 6243 3823 6256
rect 3981 6243 4031 6256
rect 857 6120 907 6148
rect 857 6100 870 6120
rect 890 6100 907 6120
rect 857 6071 907 6100
rect 1070 6119 1120 6148
rect 1070 6095 1081 6119
rect 1105 6095 1120 6119
rect 1070 6071 1120 6095
rect 1278 6124 1328 6148
rect 1278 6100 1290 6124
rect 1314 6100 1328 6124
rect 1278 6071 1328 6100
rect 1486 6122 1536 6148
rect 11565 6242 11615 6255
rect 11778 6242 11828 6255
rect 11986 6242 12036 6255
rect 12194 6242 12244 6255
rect 8099 6204 8149 6220
rect 8307 6204 8357 6220
rect 8515 6204 8565 6220
rect 8728 6204 8778 6220
rect 9147 6200 9197 6216
rect 9355 6200 9405 6216
rect 9563 6200 9613 6216
rect 9776 6200 9826 6216
rect 1486 6096 1504 6122
rect 1530 6096 1536 6122
rect 1486 6071 1536 6096
rect 3352 6115 3402 6143
rect 3352 6095 3365 6115
rect 3385 6095 3402 6115
rect 3352 6066 3402 6095
rect 3565 6114 3615 6143
rect 3565 6090 3576 6114
rect 3600 6090 3615 6114
rect 3565 6066 3615 6090
rect 3773 6119 3823 6143
rect 3773 6095 3785 6119
rect 3809 6095 3823 6119
rect 3773 6066 3823 6095
rect 3981 6117 4031 6143
rect 3981 6091 3999 6117
rect 4025 6091 4031 6117
rect 3981 6066 4031 6091
rect 8099 6137 8149 6162
rect 8099 6111 8105 6137
rect 8131 6111 8149 6137
rect 8099 6085 8149 6111
rect 8307 6133 8357 6162
rect 8307 6109 8321 6133
rect 8345 6109 8357 6133
rect 8307 6085 8357 6109
rect 8515 6138 8565 6162
rect 8515 6114 8530 6138
rect 8554 6114 8565 6138
rect 8515 6085 8565 6114
rect 8728 6133 8778 6162
rect 8728 6113 8745 6133
rect 8765 6113 8778 6133
rect 8728 6085 8778 6113
rect 9147 6133 9197 6158
rect 9147 6107 9153 6133
rect 9179 6107 9197 6133
rect 857 6013 907 6029
rect 1070 6013 1120 6029
rect 1278 6013 1328 6029
rect 1486 6013 1536 6029
rect 3352 6008 3402 6024
rect 3565 6008 3615 6024
rect 3773 6008 3823 6024
rect 3981 6008 4031 6024
rect 9147 6081 9197 6107
rect 9355 6129 9405 6158
rect 9355 6105 9369 6129
rect 9393 6105 9405 6129
rect 9355 6081 9405 6105
rect 9563 6134 9613 6158
rect 9563 6110 9578 6134
rect 9602 6110 9613 6134
rect 9563 6081 9613 6110
rect 9776 6129 9826 6158
rect 9776 6109 9793 6129
rect 9813 6109 9826 6129
rect 9776 6081 9826 6109
rect 14060 6237 14110 6250
rect 14273 6237 14323 6250
rect 14481 6237 14531 6250
rect 14689 6237 14739 6250
rect 11565 6114 11615 6142
rect 8099 5972 8149 5985
rect 8307 5972 8357 5985
rect 8515 5972 8565 5985
rect 8728 5972 8778 5985
rect 11565 6094 11578 6114
rect 11598 6094 11615 6114
rect 11565 6065 11615 6094
rect 11778 6113 11828 6142
rect 11778 6089 11789 6113
rect 11813 6089 11828 6113
rect 11778 6065 11828 6089
rect 11986 6118 12036 6142
rect 11986 6094 11998 6118
rect 12022 6094 12036 6118
rect 11986 6065 12036 6094
rect 12194 6116 12244 6142
rect 18807 6198 18857 6214
rect 19015 6198 19065 6214
rect 19223 6198 19273 6214
rect 19436 6198 19486 6214
rect 19855 6194 19905 6210
rect 20063 6194 20113 6210
rect 20271 6194 20321 6210
rect 20484 6194 20534 6210
rect 12194 6090 12212 6116
rect 12238 6090 12244 6116
rect 12194 6065 12244 6090
rect 14060 6109 14110 6137
rect 14060 6089 14073 6109
rect 14093 6089 14110 6109
rect 14060 6060 14110 6089
rect 14273 6108 14323 6137
rect 14273 6084 14284 6108
rect 14308 6084 14323 6108
rect 14273 6060 14323 6084
rect 14481 6113 14531 6137
rect 14481 6089 14493 6113
rect 14517 6089 14531 6113
rect 14481 6060 14531 6089
rect 14689 6111 14739 6137
rect 14689 6085 14707 6111
rect 14733 6085 14739 6111
rect 14689 6060 14739 6085
rect 18807 6131 18857 6156
rect 18807 6105 18813 6131
rect 18839 6105 18857 6131
rect 18807 6079 18857 6105
rect 19015 6127 19065 6156
rect 19015 6103 19029 6127
rect 19053 6103 19065 6127
rect 19015 6079 19065 6103
rect 19223 6132 19273 6156
rect 19223 6108 19238 6132
rect 19262 6108 19273 6132
rect 19223 6079 19273 6108
rect 19436 6127 19486 6156
rect 19436 6107 19453 6127
rect 19473 6107 19486 6127
rect 19436 6079 19486 6107
rect 19855 6127 19905 6152
rect 19855 6101 19861 6127
rect 19887 6101 19905 6127
rect 11565 6007 11615 6023
rect 11778 6007 11828 6023
rect 11986 6007 12036 6023
rect 12194 6007 12244 6023
rect 14060 6002 14110 6018
rect 14273 6002 14323 6018
rect 14481 6002 14531 6018
rect 14689 6002 14739 6018
rect 9147 5968 9197 5981
rect 9355 5968 9405 5981
rect 9563 5968 9613 5981
rect 9776 5968 9826 5981
rect 19855 6075 19905 6101
rect 20063 6123 20113 6152
rect 20063 6099 20077 6123
rect 20101 6099 20113 6123
rect 20063 6075 20113 6099
rect 20271 6128 20321 6152
rect 20271 6104 20286 6128
rect 20310 6104 20321 6128
rect 20271 6075 20321 6104
rect 20484 6123 20534 6152
rect 20484 6103 20501 6123
rect 20521 6103 20534 6123
rect 20484 6075 20534 6103
rect 18807 5966 18857 5979
rect 19015 5966 19065 5979
rect 19223 5966 19273 5979
rect 19436 5966 19486 5979
rect 19855 5962 19905 5975
rect 20063 5962 20113 5975
rect 20271 5962 20321 5975
rect 20484 5962 20534 5975
rect 857 5480 907 5493
rect 1070 5480 1120 5493
rect 1278 5480 1328 5493
rect 1486 5480 1536 5493
rect 1905 5476 1955 5489
rect 2118 5476 2168 5489
rect 2326 5476 2376 5489
rect 2534 5476 2584 5489
rect 857 5352 907 5380
rect 857 5332 870 5352
rect 890 5332 907 5352
rect 857 5303 907 5332
rect 1070 5351 1120 5380
rect 1070 5327 1081 5351
rect 1105 5327 1120 5351
rect 1070 5303 1120 5327
rect 1278 5356 1328 5380
rect 1278 5332 1290 5356
rect 1314 5332 1328 5356
rect 1278 5303 1328 5332
rect 1486 5354 1536 5380
rect 11565 5474 11615 5487
rect 11778 5474 11828 5487
rect 11986 5474 12036 5487
rect 12194 5474 12244 5487
rect 6652 5437 6702 5453
rect 6860 5437 6910 5453
rect 7068 5437 7118 5453
rect 7281 5437 7331 5453
rect 9147 5432 9197 5448
rect 9355 5432 9405 5448
rect 9563 5432 9613 5448
rect 9776 5432 9826 5448
rect 1486 5328 1504 5354
rect 1530 5328 1536 5354
rect 1486 5303 1536 5328
rect 1905 5348 1955 5376
rect 1905 5328 1918 5348
rect 1938 5328 1955 5348
rect 1905 5299 1955 5328
rect 2118 5347 2168 5376
rect 2118 5323 2129 5347
rect 2153 5323 2168 5347
rect 2118 5299 2168 5323
rect 2326 5352 2376 5376
rect 2326 5328 2338 5352
rect 2362 5328 2376 5352
rect 2326 5299 2376 5328
rect 2534 5350 2584 5376
rect 2534 5324 2552 5350
rect 2578 5324 2584 5350
rect 2534 5299 2584 5324
rect 6652 5370 6702 5395
rect 6652 5344 6658 5370
rect 6684 5344 6702 5370
rect 6652 5318 6702 5344
rect 6860 5366 6910 5395
rect 6860 5342 6874 5366
rect 6898 5342 6910 5366
rect 6860 5318 6910 5342
rect 7068 5371 7118 5395
rect 7068 5347 7083 5371
rect 7107 5347 7118 5371
rect 7068 5318 7118 5347
rect 7281 5366 7331 5395
rect 7281 5346 7298 5366
rect 7318 5346 7331 5366
rect 7281 5318 7331 5346
rect 9147 5365 9197 5390
rect 9147 5339 9153 5365
rect 9179 5339 9197 5365
rect 857 5245 907 5261
rect 1070 5245 1120 5261
rect 1278 5245 1328 5261
rect 1486 5245 1536 5261
rect 1905 5241 1955 5257
rect 2118 5241 2168 5257
rect 2326 5241 2376 5257
rect 2534 5241 2584 5257
rect 9147 5313 9197 5339
rect 9355 5361 9405 5390
rect 9355 5337 9369 5361
rect 9393 5337 9405 5361
rect 9355 5313 9405 5337
rect 9563 5366 9613 5390
rect 9563 5342 9578 5366
rect 9602 5342 9613 5366
rect 9563 5313 9613 5342
rect 9776 5361 9826 5390
rect 9776 5341 9793 5361
rect 9813 5341 9826 5361
rect 12613 5470 12663 5483
rect 12826 5470 12876 5483
rect 13034 5470 13084 5483
rect 13242 5470 13292 5483
rect 9776 5313 9826 5341
rect 6652 5205 6702 5218
rect 6860 5205 6910 5218
rect 7068 5205 7118 5218
rect 7281 5205 7331 5218
rect 11565 5346 11615 5374
rect 11565 5326 11578 5346
rect 11598 5326 11615 5346
rect 11565 5297 11615 5326
rect 11778 5345 11828 5374
rect 11778 5321 11789 5345
rect 11813 5321 11828 5345
rect 11778 5297 11828 5321
rect 11986 5350 12036 5374
rect 11986 5326 11998 5350
rect 12022 5326 12036 5350
rect 11986 5297 12036 5326
rect 12194 5348 12244 5374
rect 17360 5431 17410 5447
rect 17568 5431 17618 5447
rect 17776 5431 17826 5447
rect 17989 5431 18039 5447
rect 19855 5426 19905 5442
rect 20063 5426 20113 5442
rect 20271 5426 20321 5442
rect 20484 5426 20534 5442
rect 12194 5322 12212 5348
rect 12238 5322 12244 5348
rect 12194 5297 12244 5322
rect 12613 5342 12663 5370
rect 12613 5322 12626 5342
rect 12646 5322 12663 5342
rect 12613 5293 12663 5322
rect 12826 5341 12876 5370
rect 12826 5317 12837 5341
rect 12861 5317 12876 5341
rect 12826 5293 12876 5317
rect 13034 5346 13084 5370
rect 13034 5322 13046 5346
rect 13070 5322 13084 5346
rect 13034 5293 13084 5322
rect 13242 5344 13292 5370
rect 13242 5318 13260 5344
rect 13286 5318 13292 5344
rect 13242 5293 13292 5318
rect 17360 5364 17410 5389
rect 17360 5338 17366 5364
rect 17392 5338 17410 5364
rect 17360 5312 17410 5338
rect 17568 5360 17618 5389
rect 17568 5336 17582 5360
rect 17606 5336 17618 5360
rect 17568 5312 17618 5336
rect 17776 5365 17826 5389
rect 17776 5341 17791 5365
rect 17815 5341 17826 5365
rect 17776 5312 17826 5341
rect 17989 5360 18039 5389
rect 17989 5340 18006 5360
rect 18026 5340 18039 5360
rect 17989 5312 18039 5340
rect 19855 5359 19905 5384
rect 19855 5333 19861 5359
rect 19887 5333 19905 5359
rect 11565 5239 11615 5255
rect 11778 5239 11828 5255
rect 11986 5239 12036 5255
rect 12194 5239 12244 5255
rect 12613 5235 12663 5251
rect 12826 5235 12876 5251
rect 13034 5235 13084 5251
rect 13242 5235 13292 5251
rect 9147 5200 9197 5213
rect 9355 5200 9405 5213
rect 9563 5200 9613 5213
rect 9776 5200 9826 5213
rect 19855 5307 19905 5333
rect 20063 5355 20113 5384
rect 20063 5331 20077 5355
rect 20101 5331 20113 5355
rect 20063 5307 20113 5331
rect 20271 5360 20321 5384
rect 20271 5336 20286 5360
rect 20310 5336 20321 5360
rect 20271 5307 20321 5336
rect 20484 5355 20534 5384
rect 20484 5335 20501 5355
rect 20521 5335 20534 5355
rect 20484 5307 20534 5335
rect 17360 5199 17410 5212
rect 17568 5199 17618 5212
rect 17776 5199 17826 5212
rect 17989 5199 18039 5212
rect 19855 5194 19905 5207
rect 20063 5194 20113 5207
rect 20271 5194 20321 5207
rect 20484 5194 20534 5207
rect 857 4801 907 4814
rect 1070 4801 1120 4814
rect 1278 4801 1328 4814
rect 1486 4801 1536 4814
rect 3395 4798 3445 4811
rect 3608 4798 3658 4811
rect 3816 4798 3866 4811
rect 4024 4798 4074 4811
rect 857 4673 907 4701
rect 857 4653 870 4673
rect 890 4653 907 4673
rect 857 4624 907 4653
rect 1070 4672 1120 4701
rect 1070 4648 1081 4672
rect 1105 4648 1120 4672
rect 1070 4624 1120 4648
rect 1278 4677 1328 4701
rect 1278 4653 1290 4677
rect 1314 4653 1328 4677
rect 1278 4624 1328 4653
rect 1486 4675 1536 4701
rect 11565 4795 11615 4808
rect 11778 4795 11828 4808
rect 11986 4795 12036 4808
rect 12194 4795 12244 4808
rect 8099 4757 8149 4773
rect 8307 4757 8357 4773
rect 8515 4757 8565 4773
rect 8728 4757 8778 4773
rect 9147 4753 9197 4769
rect 9355 4753 9405 4769
rect 9563 4753 9613 4769
rect 9776 4753 9826 4769
rect 1486 4649 1504 4675
rect 1530 4649 1536 4675
rect 1486 4624 1536 4649
rect 3395 4670 3445 4698
rect 3395 4650 3408 4670
rect 3428 4650 3445 4670
rect 3395 4621 3445 4650
rect 3608 4669 3658 4698
rect 3608 4645 3619 4669
rect 3643 4645 3658 4669
rect 3608 4621 3658 4645
rect 3816 4674 3866 4698
rect 3816 4650 3828 4674
rect 3852 4650 3866 4674
rect 3816 4621 3866 4650
rect 4024 4672 4074 4698
rect 4024 4646 4042 4672
rect 4068 4646 4074 4672
rect 4024 4621 4074 4646
rect 8099 4690 8149 4715
rect 8099 4664 8105 4690
rect 8131 4664 8149 4690
rect 8099 4638 8149 4664
rect 8307 4686 8357 4715
rect 8307 4662 8321 4686
rect 8345 4662 8357 4686
rect 8307 4638 8357 4662
rect 8515 4691 8565 4715
rect 8515 4667 8530 4691
rect 8554 4667 8565 4691
rect 8515 4638 8565 4667
rect 8728 4686 8778 4715
rect 8728 4666 8745 4686
rect 8765 4666 8778 4686
rect 8728 4638 8778 4666
rect 9147 4686 9197 4711
rect 9147 4660 9153 4686
rect 9179 4660 9197 4686
rect 857 4566 907 4582
rect 1070 4566 1120 4582
rect 1278 4566 1328 4582
rect 1486 4566 1536 4582
rect 3395 4563 3445 4579
rect 3608 4563 3658 4579
rect 3816 4563 3866 4579
rect 4024 4563 4074 4579
rect 9147 4634 9197 4660
rect 9355 4682 9405 4711
rect 9355 4658 9369 4682
rect 9393 4658 9405 4682
rect 9355 4634 9405 4658
rect 9563 4687 9613 4711
rect 9563 4663 9578 4687
rect 9602 4663 9613 4687
rect 9563 4634 9613 4663
rect 9776 4682 9826 4711
rect 9776 4662 9793 4682
rect 9813 4662 9826 4682
rect 9776 4634 9826 4662
rect 14103 4792 14153 4805
rect 14316 4792 14366 4805
rect 14524 4792 14574 4805
rect 14732 4792 14782 4805
rect 11565 4667 11615 4695
rect 8099 4525 8149 4538
rect 8307 4525 8357 4538
rect 8515 4525 8565 4538
rect 8728 4525 8778 4538
rect 11565 4647 11578 4667
rect 11598 4647 11615 4667
rect 11565 4618 11615 4647
rect 11778 4666 11828 4695
rect 11778 4642 11789 4666
rect 11813 4642 11828 4666
rect 11778 4618 11828 4642
rect 11986 4671 12036 4695
rect 11986 4647 11998 4671
rect 12022 4647 12036 4671
rect 11986 4618 12036 4647
rect 12194 4669 12244 4695
rect 18807 4751 18857 4767
rect 19015 4751 19065 4767
rect 19223 4751 19273 4767
rect 19436 4751 19486 4767
rect 19855 4747 19905 4763
rect 20063 4747 20113 4763
rect 20271 4747 20321 4763
rect 20484 4747 20534 4763
rect 12194 4643 12212 4669
rect 12238 4643 12244 4669
rect 12194 4618 12244 4643
rect 14103 4664 14153 4692
rect 14103 4644 14116 4664
rect 14136 4644 14153 4664
rect 14103 4615 14153 4644
rect 14316 4663 14366 4692
rect 14316 4639 14327 4663
rect 14351 4639 14366 4663
rect 14316 4615 14366 4639
rect 14524 4668 14574 4692
rect 14524 4644 14536 4668
rect 14560 4644 14574 4668
rect 14524 4615 14574 4644
rect 14732 4666 14782 4692
rect 14732 4640 14750 4666
rect 14776 4640 14782 4666
rect 14732 4615 14782 4640
rect 18807 4684 18857 4709
rect 18807 4658 18813 4684
rect 18839 4658 18857 4684
rect 18807 4632 18857 4658
rect 19015 4680 19065 4709
rect 19015 4656 19029 4680
rect 19053 4656 19065 4680
rect 19015 4632 19065 4656
rect 19223 4685 19273 4709
rect 19223 4661 19238 4685
rect 19262 4661 19273 4685
rect 19223 4632 19273 4661
rect 19436 4680 19486 4709
rect 19436 4660 19453 4680
rect 19473 4660 19486 4680
rect 19436 4632 19486 4660
rect 19855 4680 19905 4705
rect 19855 4654 19861 4680
rect 19887 4654 19905 4680
rect 11565 4560 11615 4576
rect 11778 4560 11828 4576
rect 11986 4560 12036 4576
rect 12194 4560 12244 4576
rect 14103 4557 14153 4573
rect 14316 4557 14366 4573
rect 14524 4557 14574 4573
rect 14732 4557 14782 4573
rect 9147 4521 9197 4534
rect 9355 4521 9405 4534
rect 9563 4521 9613 4534
rect 9776 4521 9826 4534
rect 19855 4628 19905 4654
rect 20063 4676 20113 4705
rect 20063 4652 20077 4676
rect 20101 4652 20113 4676
rect 20063 4628 20113 4652
rect 20271 4681 20321 4705
rect 20271 4657 20286 4681
rect 20310 4657 20321 4681
rect 20271 4628 20321 4657
rect 20484 4676 20534 4705
rect 20484 4656 20501 4676
rect 20521 4656 20534 4676
rect 20484 4628 20534 4656
rect 18807 4519 18857 4532
rect 19015 4519 19065 4532
rect 19223 4519 19273 4532
rect 19436 4519 19486 4532
rect 19855 4515 19905 4528
rect 20063 4515 20113 4528
rect 20271 4515 20321 4528
rect 20484 4515 20534 4528
rect 858 3960 908 3973
rect 1071 3960 1121 3973
rect 1279 3960 1329 3973
rect 1487 3960 1537 3973
rect 1906 3956 1956 3969
rect 2119 3956 2169 3969
rect 2327 3956 2377 3969
rect 2535 3956 2585 3969
rect 4808 3962 4858 3975
rect 5021 3962 5071 3975
rect 5229 3962 5279 3975
rect 5437 3962 5487 3975
rect 858 3832 908 3860
rect 858 3812 871 3832
rect 891 3812 908 3832
rect 858 3783 908 3812
rect 1071 3831 1121 3860
rect 1071 3807 1082 3831
rect 1106 3807 1121 3831
rect 1071 3783 1121 3807
rect 1279 3836 1329 3860
rect 1279 3812 1291 3836
rect 1315 3812 1329 3836
rect 1279 3783 1329 3812
rect 1487 3834 1537 3860
rect 11566 3954 11616 3967
rect 11779 3954 11829 3967
rect 11987 3954 12037 3967
rect 12195 3954 12245 3967
rect 6610 3915 6660 3931
rect 6818 3915 6868 3931
rect 7026 3915 7076 3931
rect 7239 3915 7289 3931
rect 9148 3912 9198 3928
rect 9356 3912 9406 3928
rect 9564 3912 9614 3928
rect 9777 3912 9827 3928
rect 1487 3808 1505 3834
rect 1531 3808 1537 3834
rect 1487 3783 1537 3808
rect 1906 3828 1956 3856
rect 1906 3808 1919 3828
rect 1939 3808 1956 3828
rect 1906 3779 1956 3808
rect 2119 3827 2169 3856
rect 2119 3803 2130 3827
rect 2154 3803 2169 3827
rect 2119 3779 2169 3803
rect 2327 3832 2377 3856
rect 2327 3808 2339 3832
rect 2363 3808 2377 3832
rect 2327 3779 2377 3808
rect 2535 3830 2585 3856
rect 2535 3804 2553 3830
rect 2579 3804 2585 3830
rect 2535 3779 2585 3804
rect 4808 3834 4858 3862
rect 4808 3814 4821 3834
rect 4841 3814 4858 3834
rect 4808 3785 4858 3814
rect 5021 3833 5071 3862
rect 5021 3809 5032 3833
rect 5056 3809 5071 3833
rect 5021 3785 5071 3809
rect 5229 3838 5279 3862
rect 5229 3814 5241 3838
rect 5265 3814 5279 3838
rect 5229 3785 5279 3814
rect 5437 3836 5487 3862
rect 5437 3810 5455 3836
rect 5481 3810 5487 3836
rect 5437 3785 5487 3810
rect 6610 3848 6660 3873
rect 6610 3822 6616 3848
rect 6642 3822 6660 3848
rect 6610 3796 6660 3822
rect 6818 3844 6868 3873
rect 6818 3820 6832 3844
rect 6856 3820 6868 3844
rect 6818 3796 6868 3820
rect 7026 3849 7076 3873
rect 7026 3825 7041 3849
rect 7065 3825 7076 3849
rect 7026 3796 7076 3825
rect 7239 3844 7289 3873
rect 7239 3824 7256 3844
rect 7276 3824 7289 3844
rect 7239 3796 7289 3824
rect 9148 3845 9198 3870
rect 9148 3819 9154 3845
rect 9180 3819 9198 3845
rect 858 3725 908 3741
rect 1071 3725 1121 3741
rect 1279 3725 1329 3741
rect 1487 3725 1537 3741
rect 1906 3721 1956 3737
rect 2119 3721 2169 3737
rect 2327 3721 2377 3737
rect 2535 3721 2585 3737
rect 4808 3727 4858 3743
rect 5021 3727 5071 3743
rect 5229 3727 5279 3743
rect 5437 3727 5487 3743
rect 9148 3793 9198 3819
rect 9356 3841 9406 3870
rect 9356 3817 9370 3841
rect 9394 3817 9406 3841
rect 9356 3793 9406 3817
rect 9564 3846 9614 3870
rect 9564 3822 9579 3846
rect 9603 3822 9614 3846
rect 9564 3793 9614 3822
rect 9777 3841 9827 3870
rect 9777 3821 9794 3841
rect 9814 3821 9827 3841
rect 12614 3950 12664 3963
rect 12827 3950 12877 3963
rect 13035 3950 13085 3963
rect 13243 3950 13293 3963
rect 15516 3956 15566 3969
rect 15729 3956 15779 3969
rect 15937 3956 15987 3969
rect 16145 3956 16195 3969
rect 9777 3793 9827 3821
rect 6610 3683 6660 3696
rect 6818 3683 6868 3696
rect 7026 3683 7076 3696
rect 7239 3683 7289 3696
rect 11566 3826 11616 3854
rect 11566 3806 11579 3826
rect 11599 3806 11616 3826
rect 11566 3777 11616 3806
rect 11779 3825 11829 3854
rect 11779 3801 11790 3825
rect 11814 3801 11829 3825
rect 11779 3777 11829 3801
rect 11987 3830 12037 3854
rect 11987 3806 11999 3830
rect 12023 3806 12037 3830
rect 11987 3777 12037 3806
rect 12195 3828 12245 3854
rect 17318 3909 17368 3925
rect 17526 3909 17576 3925
rect 17734 3909 17784 3925
rect 17947 3909 17997 3925
rect 19856 3906 19906 3922
rect 20064 3906 20114 3922
rect 20272 3906 20322 3922
rect 20485 3906 20535 3922
rect 12195 3802 12213 3828
rect 12239 3802 12245 3828
rect 12195 3777 12245 3802
rect 12614 3822 12664 3850
rect 12614 3802 12627 3822
rect 12647 3802 12664 3822
rect 12614 3773 12664 3802
rect 12827 3821 12877 3850
rect 12827 3797 12838 3821
rect 12862 3797 12877 3821
rect 12827 3773 12877 3797
rect 13035 3826 13085 3850
rect 13035 3802 13047 3826
rect 13071 3802 13085 3826
rect 13035 3773 13085 3802
rect 13243 3824 13293 3850
rect 13243 3798 13261 3824
rect 13287 3798 13293 3824
rect 13243 3773 13293 3798
rect 15516 3828 15566 3856
rect 15516 3808 15529 3828
rect 15549 3808 15566 3828
rect 15516 3779 15566 3808
rect 15729 3827 15779 3856
rect 15729 3803 15740 3827
rect 15764 3803 15779 3827
rect 15729 3779 15779 3803
rect 15937 3832 15987 3856
rect 15937 3808 15949 3832
rect 15973 3808 15987 3832
rect 15937 3779 15987 3808
rect 16145 3830 16195 3856
rect 16145 3804 16163 3830
rect 16189 3804 16195 3830
rect 16145 3779 16195 3804
rect 17318 3842 17368 3867
rect 17318 3816 17324 3842
rect 17350 3816 17368 3842
rect 17318 3790 17368 3816
rect 17526 3838 17576 3867
rect 17526 3814 17540 3838
rect 17564 3814 17576 3838
rect 17526 3790 17576 3814
rect 17734 3843 17784 3867
rect 17734 3819 17749 3843
rect 17773 3819 17784 3843
rect 17734 3790 17784 3819
rect 17947 3838 17997 3867
rect 17947 3818 17964 3838
rect 17984 3818 17997 3838
rect 17947 3790 17997 3818
rect 19856 3839 19906 3864
rect 19856 3813 19862 3839
rect 19888 3813 19906 3839
rect 11566 3719 11616 3735
rect 11779 3719 11829 3735
rect 11987 3719 12037 3735
rect 12195 3719 12245 3735
rect 12614 3715 12664 3731
rect 12827 3715 12877 3731
rect 13035 3715 13085 3731
rect 13243 3715 13293 3731
rect 15516 3721 15566 3737
rect 15729 3721 15779 3737
rect 15937 3721 15987 3737
rect 16145 3721 16195 3737
rect 9148 3680 9198 3693
rect 9356 3680 9406 3693
rect 9564 3680 9614 3693
rect 9777 3680 9827 3693
rect 19856 3787 19906 3813
rect 20064 3835 20114 3864
rect 20064 3811 20078 3835
rect 20102 3811 20114 3835
rect 20064 3787 20114 3811
rect 20272 3840 20322 3864
rect 20272 3816 20287 3840
rect 20311 3816 20322 3840
rect 20272 3787 20322 3816
rect 20485 3835 20535 3864
rect 20485 3815 20502 3835
rect 20522 3815 20535 3835
rect 20485 3787 20535 3815
rect 17318 3677 17368 3690
rect 17526 3677 17576 3690
rect 17734 3677 17784 3690
rect 17947 3677 17997 3690
rect 19856 3674 19906 3687
rect 20064 3674 20114 3687
rect 20272 3674 20322 3687
rect 20485 3674 20535 3687
rect 858 3281 908 3294
rect 1071 3281 1121 3294
rect 1279 3281 1329 3294
rect 1487 3281 1537 3294
rect 3353 3276 3403 3289
rect 3566 3276 3616 3289
rect 3774 3276 3824 3289
rect 3982 3276 4032 3289
rect 858 3153 908 3181
rect 858 3133 871 3153
rect 891 3133 908 3153
rect 858 3104 908 3133
rect 1071 3152 1121 3181
rect 1071 3128 1082 3152
rect 1106 3128 1121 3152
rect 1071 3104 1121 3128
rect 1279 3157 1329 3181
rect 1279 3133 1291 3157
rect 1315 3133 1329 3157
rect 1279 3104 1329 3133
rect 1487 3155 1537 3181
rect 11566 3275 11616 3288
rect 11779 3275 11829 3288
rect 11987 3275 12037 3288
rect 12195 3275 12245 3288
rect 8100 3237 8150 3253
rect 8308 3237 8358 3253
rect 8516 3237 8566 3253
rect 8729 3237 8779 3253
rect 9148 3233 9198 3249
rect 9356 3233 9406 3249
rect 9564 3233 9614 3249
rect 9777 3233 9827 3249
rect 1487 3129 1505 3155
rect 1531 3129 1537 3155
rect 1487 3104 1537 3129
rect 3353 3148 3403 3176
rect 3353 3128 3366 3148
rect 3386 3128 3403 3148
rect 3353 3099 3403 3128
rect 3566 3147 3616 3176
rect 3566 3123 3577 3147
rect 3601 3123 3616 3147
rect 3566 3099 3616 3123
rect 3774 3152 3824 3176
rect 3774 3128 3786 3152
rect 3810 3128 3824 3152
rect 3774 3099 3824 3128
rect 3982 3150 4032 3176
rect 3982 3124 4000 3150
rect 4026 3124 4032 3150
rect 3982 3099 4032 3124
rect 8100 3170 8150 3195
rect 8100 3144 8106 3170
rect 8132 3144 8150 3170
rect 8100 3118 8150 3144
rect 8308 3166 8358 3195
rect 8308 3142 8322 3166
rect 8346 3142 8358 3166
rect 8308 3118 8358 3142
rect 8516 3171 8566 3195
rect 8516 3147 8531 3171
rect 8555 3147 8566 3171
rect 8516 3118 8566 3147
rect 8729 3166 8779 3195
rect 8729 3146 8746 3166
rect 8766 3146 8779 3166
rect 8729 3118 8779 3146
rect 9148 3166 9198 3191
rect 9148 3140 9154 3166
rect 9180 3140 9198 3166
rect 858 3046 908 3062
rect 1071 3046 1121 3062
rect 1279 3046 1329 3062
rect 1487 3046 1537 3062
rect 3353 3041 3403 3057
rect 3566 3041 3616 3057
rect 3774 3041 3824 3057
rect 3982 3041 4032 3057
rect 9148 3114 9198 3140
rect 9356 3162 9406 3191
rect 9356 3138 9370 3162
rect 9394 3138 9406 3162
rect 9356 3114 9406 3138
rect 9564 3167 9614 3191
rect 9564 3143 9579 3167
rect 9603 3143 9614 3167
rect 9564 3114 9614 3143
rect 9777 3162 9827 3191
rect 9777 3142 9794 3162
rect 9814 3142 9827 3162
rect 9777 3114 9827 3142
rect 14061 3270 14111 3283
rect 14274 3270 14324 3283
rect 14482 3270 14532 3283
rect 14690 3270 14740 3283
rect 11566 3147 11616 3175
rect 8100 3005 8150 3018
rect 8308 3005 8358 3018
rect 8516 3005 8566 3018
rect 8729 3005 8779 3018
rect 11566 3127 11579 3147
rect 11599 3127 11616 3147
rect 11566 3098 11616 3127
rect 11779 3146 11829 3175
rect 11779 3122 11790 3146
rect 11814 3122 11829 3146
rect 11779 3098 11829 3122
rect 11987 3151 12037 3175
rect 11987 3127 11999 3151
rect 12023 3127 12037 3151
rect 11987 3098 12037 3127
rect 12195 3149 12245 3175
rect 18808 3231 18858 3247
rect 19016 3231 19066 3247
rect 19224 3231 19274 3247
rect 19437 3231 19487 3247
rect 19856 3227 19906 3243
rect 20064 3227 20114 3243
rect 20272 3227 20322 3243
rect 20485 3227 20535 3243
rect 12195 3123 12213 3149
rect 12239 3123 12245 3149
rect 12195 3098 12245 3123
rect 14061 3142 14111 3170
rect 14061 3122 14074 3142
rect 14094 3122 14111 3142
rect 14061 3093 14111 3122
rect 14274 3141 14324 3170
rect 14274 3117 14285 3141
rect 14309 3117 14324 3141
rect 14274 3093 14324 3117
rect 14482 3146 14532 3170
rect 14482 3122 14494 3146
rect 14518 3122 14532 3146
rect 14482 3093 14532 3122
rect 14690 3144 14740 3170
rect 14690 3118 14708 3144
rect 14734 3118 14740 3144
rect 14690 3093 14740 3118
rect 18808 3164 18858 3189
rect 18808 3138 18814 3164
rect 18840 3138 18858 3164
rect 18808 3112 18858 3138
rect 19016 3160 19066 3189
rect 19016 3136 19030 3160
rect 19054 3136 19066 3160
rect 19016 3112 19066 3136
rect 19224 3165 19274 3189
rect 19224 3141 19239 3165
rect 19263 3141 19274 3165
rect 19224 3112 19274 3141
rect 19437 3160 19487 3189
rect 19437 3140 19454 3160
rect 19474 3140 19487 3160
rect 19437 3112 19487 3140
rect 19856 3160 19906 3185
rect 19856 3134 19862 3160
rect 19888 3134 19906 3160
rect 11566 3040 11616 3056
rect 11779 3040 11829 3056
rect 11987 3040 12037 3056
rect 12195 3040 12245 3056
rect 14061 3035 14111 3051
rect 14274 3035 14324 3051
rect 14482 3035 14532 3051
rect 14690 3035 14740 3051
rect 9148 3001 9198 3014
rect 9356 3001 9406 3014
rect 9564 3001 9614 3014
rect 9777 3001 9827 3014
rect 19856 3108 19906 3134
rect 20064 3156 20114 3185
rect 20064 3132 20078 3156
rect 20102 3132 20114 3156
rect 20064 3108 20114 3132
rect 20272 3161 20322 3185
rect 20272 3137 20287 3161
rect 20311 3137 20322 3161
rect 20272 3108 20322 3137
rect 20485 3156 20535 3185
rect 20485 3136 20502 3156
rect 20522 3136 20535 3156
rect 20485 3108 20535 3136
rect 18808 2999 18858 3012
rect 19016 2999 19066 3012
rect 19224 2999 19274 3012
rect 19437 2999 19487 3012
rect 19856 2995 19906 3008
rect 20064 2995 20114 3008
rect 20272 2995 20322 3008
rect 20485 2995 20535 3008
rect 858 2513 908 2526
rect 1071 2513 1121 2526
rect 1279 2513 1329 2526
rect 1487 2513 1537 2526
rect 1906 2509 1956 2522
rect 2119 2509 2169 2522
rect 2327 2509 2377 2522
rect 2535 2509 2585 2522
rect 858 2385 908 2413
rect 858 2365 871 2385
rect 891 2365 908 2385
rect 858 2336 908 2365
rect 1071 2384 1121 2413
rect 1071 2360 1082 2384
rect 1106 2360 1121 2384
rect 1071 2336 1121 2360
rect 1279 2389 1329 2413
rect 1279 2365 1291 2389
rect 1315 2365 1329 2389
rect 1279 2336 1329 2365
rect 1487 2387 1537 2413
rect 11566 2507 11616 2520
rect 11779 2507 11829 2520
rect 11987 2507 12037 2520
rect 12195 2507 12245 2520
rect 6653 2470 6703 2486
rect 6861 2470 6911 2486
rect 7069 2470 7119 2486
rect 7282 2470 7332 2486
rect 9148 2465 9198 2481
rect 9356 2465 9406 2481
rect 9564 2465 9614 2481
rect 9777 2465 9827 2481
rect 1487 2361 1505 2387
rect 1531 2361 1537 2387
rect 1487 2336 1537 2361
rect 1906 2381 1956 2409
rect 1906 2361 1919 2381
rect 1939 2361 1956 2381
rect 1906 2332 1956 2361
rect 2119 2380 2169 2409
rect 2119 2356 2130 2380
rect 2154 2356 2169 2380
rect 2119 2332 2169 2356
rect 2327 2385 2377 2409
rect 2327 2361 2339 2385
rect 2363 2361 2377 2385
rect 2327 2332 2377 2361
rect 2535 2383 2585 2409
rect 2535 2357 2553 2383
rect 2579 2357 2585 2383
rect 2535 2332 2585 2357
rect 6653 2403 6703 2428
rect 6653 2377 6659 2403
rect 6685 2377 6703 2403
rect 6653 2351 6703 2377
rect 6861 2399 6911 2428
rect 6861 2375 6875 2399
rect 6899 2375 6911 2399
rect 6861 2351 6911 2375
rect 7069 2404 7119 2428
rect 7069 2380 7084 2404
rect 7108 2380 7119 2404
rect 7069 2351 7119 2380
rect 7282 2399 7332 2428
rect 7282 2379 7299 2399
rect 7319 2379 7332 2399
rect 7282 2351 7332 2379
rect 9148 2398 9198 2423
rect 9148 2372 9154 2398
rect 9180 2372 9198 2398
rect 858 2278 908 2294
rect 1071 2278 1121 2294
rect 1279 2278 1329 2294
rect 1487 2278 1537 2294
rect 1906 2274 1956 2290
rect 2119 2274 2169 2290
rect 2327 2274 2377 2290
rect 2535 2274 2585 2290
rect 9148 2346 9198 2372
rect 9356 2394 9406 2423
rect 9356 2370 9370 2394
rect 9394 2370 9406 2394
rect 9356 2346 9406 2370
rect 9564 2399 9614 2423
rect 9564 2375 9579 2399
rect 9603 2375 9614 2399
rect 9564 2346 9614 2375
rect 9777 2394 9827 2423
rect 9777 2374 9794 2394
rect 9814 2374 9827 2394
rect 12614 2503 12664 2516
rect 12827 2503 12877 2516
rect 13035 2503 13085 2516
rect 13243 2503 13293 2516
rect 9777 2346 9827 2374
rect 6653 2238 6703 2251
rect 6861 2238 6911 2251
rect 7069 2238 7119 2251
rect 7282 2238 7332 2251
rect 11566 2379 11616 2407
rect 11566 2359 11579 2379
rect 11599 2359 11616 2379
rect 11566 2330 11616 2359
rect 11779 2378 11829 2407
rect 11779 2354 11790 2378
rect 11814 2354 11829 2378
rect 11779 2330 11829 2354
rect 11987 2383 12037 2407
rect 11987 2359 11999 2383
rect 12023 2359 12037 2383
rect 11987 2330 12037 2359
rect 12195 2381 12245 2407
rect 17361 2464 17411 2480
rect 17569 2464 17619 2480
rect 17777 2464 17827 2480
rect 17990 2464 18040 2480
rect 19856 2459 19906 2475
rect 20064 2459 20114 2475
rect 20272 2459 20322 2475
rect 20485 2459 20535 2475
rect 12195 2355 12213 2381
rect 12239 2355 12245 2381
rect 12195 2330 12245 2355
rect 12614 2375 12664 2403
rect 12614 2355 12627 2375
rect 12647 2355 12664 2375
rect 12614 2326 12664 2355
rect 12827 2374 12877 2403
rect 12827 2350 12838 2374
rect 12862 2350 12877 2374
rect 12827 2326 12877 2350
rect 13035 2379 13085 2403
rect 13035 2355 13047 2379
rect 13071 2355 13085 2379
rect 13035 2326 13085 2355
rect 13243 2377 13293 2403
rect 13243 2351 13261 2377
rect 13287 2351 13293 2377
rect 13243 2326 13293 2351
rect 17361 2397 17411 2422
rect 17361 2371 17367 2397
rect 17393 2371 17411 2397
rect 17361 2345 17411 2371
rect 17569 2393 17619 2422
rect 17569 2369 17583 2393
rect 17607 2369 17619 2393
rect 17569 2345 17619 2369
rect 17777 2398 17827 2422
rect 17777 2374 17792 2398
rect 17816 2374 17827 2398
rect 17777 2345 17827 2374
rect 17990 2393 18040 2422
rect 17990 2373 18007 2393
rect 18027 2373 18040 2393
rect 17990 2345 18040 2373
rect 19856 2392 19906 2417
rect 19856 2366 19862 2392
rect 19888 2366 19906 2392
rect 11566 2272 11616 2288
rect 11779 2272 11829 2288
rect 11987 2272 12037 2288
rect 12195 2272 12245 2288
rect 12614 2268 12664 2284
rect 12827 2268 12877 2284
rect 13035 2268 13085 2284
rect 13243 2268 13293 2284
rect 9148 2233 9198 2246
rect 9356 2233 9406 2246
rect 9564 2233 9614 2246
rect 9777 2233 9827 2246
rect 19856 2340 19906 2366
rect 20064 2388 20114 2417
rect 20064 2364 20078 2388
rect 20102 2364 20114 2388
rect 20064 2340 20114 2364
rect 20272 2393 20322 2417
rect 20272 2369 20287 2393
rect 20311 2369 20322 2393
rect 20272 2340 20322 2369
rect 20485 2388 20535 2417
rect 20485 2368 20502 2388
rect 20522 2368 20535 2388
rect 20485 2340 20535 2368
rect 17361 2232 17411 2245
rect 17569 2232 17619 2245
rect 17777 2232 17827 2245
rect 17990 2232 18040 2245
rect 19856 2227 19906 2240
rect 20064 2227 20114 2240
rect 20272 2227 20322 2240
rect 20485 2227 20535 2240
rect 858 1834 908 1847
rect 1071 1834 1121 1847
rect 1279 1834 1329 1847
rect 1487 1834 1537 1847
rect 11566 1828 11616 1841
rect 11779 1828 11829 1841
rect 11987 1828 12037 1841
rect 12195 1828 12245 1841
rect 8100 1790 8150 1806
rect 8308 1790 8358 1806
rect 8516 1790 8566 1806
rect 8729 1790 8779 1806
rect 9148 1786 9198 1802
rect 9356 1786 9406 1802
rect 9564 1786 9614 1802
rect 9777 1786 9827 1802
rect 858 1706 908 1734
rect 858 1686 871 1706
rect 891 1686 908 1706
rect 858 1657 908 1686
rect 1071 1705 1121 1734
rect 1071 1681 1082 1705
rect 1106 1681 1121 1705
rect 1071 1657 1121 1681
rect 1279 1710 1329 1734
rect 1279 1686 1291 1710
rect 1315 1686 1329 1710
rect 1279 1657 1329 1686
rect 1487 1708 1537 1734
rect 1487 1682 1505 1708
rect 1531 1682 1537 1708
rect 1487 1657 1537 1682
rect 8100 1723 8150 1748
rect 8100 1697 8106 1723
rect 8132 1697 8150 1723
rect 8100 1671 8150 1697
rect 8308 1719 8358 1748
rect 8308 1695 8322 1719
rect 8346 1695 8358 1719
rect 8308 1671 8358 1695
rect 8516 1724 8566 1748
rect 8516 1700 8531 1724
rect 8555 1700 8566 1724
rect 8516 1671 8566 1700
rect 8729 1719 8779 1748
rect 8729 1699 8746 1719
rect 8766 1699 8779 1719
rect 8729 1671 8779 1699
rect 9148 1719 9198 1744
rect 9148 1693 9154 1719
rect 9180 1693 9198 1719
rect 858 1599 908 1615
rect 1071 1599 1121 1615
rect 1279 1599 1329 1615
rect 1487 1599 1537 1615
rect 9148 1667 9198 1693
rect 9356 1715 9406 1744
rect 9356 1691 9370 1715
rect 9394 1691 9406 1715
rect 9356 1667 9406 1691
rect 9564 1720 9614 1744
rect 9564 1696 9579 1720
rect 9603 1696 9614 1720
rect 9564 1667 9614 1696
rect 9777 1715 9827 1744
rect 9777 1695 9794 1715
rect 9814 1695 9827 1715
rect 9777 1667 9827 1695
rect 18808 1784 18858 1800
rect 19016 1784 19066 1800
rect 19224 1784 19274 1800
rect 19437 1784 19487 1800
rect 19856 1780 19906 1796
rect 20064 1780 20114 1796
rect 20272 1780 20322 1796
rect 20485 1780 20535 1796
rect 11566 1700 11616 1728
rect 8100 1558 8150 1571
rect 8308 1558 8358 1571
rect 8516 1558 8566 1571
rect 8729 1558 8779 1571
rect 11566 1680 11579 1700
rect 11599 1680 11616 1700
rect 11566 1651 11616 1680
rect 11779 1699 11829 1728
rect 11779 1675 11790 1699
rect 11814 1675 11829 1699
rect 11779 1651 11829 1675
rect 11987 1704 12037 1728
rect 11987 1680 11999 1704
rect 12023 1680 12037 1704
rect 11987 1651 12037 1680
rect 12195 1702 12245 1728
rect 12195 1676 12213 1702
rect 12239 1676 12245 1702
rect 12195 1651 12245 1676
rect 18808 1717 18858 1742
rect 18808 1691 18814 1717
rect 18840 1691 18858 1717
rect 18808 1665 18858 1691
rect 19016 1713 19066 1742
rect 19016 1689 19030 1713
rect 19054 1689 19066 1713
rect 19016 1665 19066 1689
rect 19224 1718 19274 1742
rect 19224 1694 19239 1718
rect 19263 1694 19274 1718
rect 19224 1665 19274 1694
rect 19437 1713 19487 1742
rect 19437 1693 19454 1713
rect 19474 1693 19487 1713
rect 19437 1665 19487 1693
rect 19856 1713 19906 1738
rect 19856 1687 19862 1713
rect 19888 1687 19906 1713
rect 11566 1593 11616 1609
rect 11779 1593 11829 1609
rect 11987 1593 12037 1609
rect 12195 1593 12245 1609
rect 9148 1554 9198 1567
rect 9356 1554 9406 1567
rect 9564 1554 9614 1567
rect 9777 1554 9827 1567
rect 19856 1661 19906 1687
rect 20064 1709 20114 1738
rect 20064 1685 20078 1709
rect 20102 1685 20114 1709
rect 20064 1661 20114 1685
rect 20272 1714 20322 1738
rect 20272 1690 20287 1714
rect 20311 1690 20322 1714
rect 20272 1661 20322 1690
rect 20485 1709 20535 1738
rect 20485 1689 20502 1709
rect 20522 1689 20535 1709
rect 20485 1661 20535 1689
rect 18808 1552 18858 1565
rect 19016 1552 19066 1565
rect 19224 1552 19274 1565
rect 19437 1552 19487 1565
rect 19856 1548 19906 1561
rect 20064 1548 20114 1561
rect 20272 1548 20322 1561
rect 20485 1548 20535 1561
rect 10569 -325 10619 -312
rect 10782 -325 10832 -312
rect 10990 -325 11040 -312
rect 11198 -325 11248 -312
rect 10569 -453 10619 -425
rect 10569 -473 10582 -453
rect 10602 -473 10619 -453
rect 10569 -502 10619 -473
rect 10782 -454 10832 -425
rect 10782 -478 10793 -454
rect 10817 -478 10832 -454
rect 10782 -502 10832 -478
rect 10990 -449 11040 -425
rect 10990 -473 11002 -449
rect 11026 -473 11040 -449
rect 10990 -502 11040 -473
rect 11198 -451 11248 -425
rect 11198 -477 11216 -451
rect 11242 -477 11248 -451
rect 11198 -502 11248 -477
rect 10569 -560 10619 -544
rect 10782 -560 10832 -544
rect 10990 -560 11040 -544
rect 11198 -560 11248 -544
<< polycont >>
rect 872 12787 892 12807
rect 1083 12782 1107 12806
rect 1292 12787 1316 12811
rect 1506 12783 1532 12809
rect 1920 12783 1940 12803
rect 2131 12778 2155 12802
rect 2340 12783 2364 12807
rect 2554 12779 2580 12805
rect 9155 12794 9181 12820
rect 9371 12792 9395 12816
rect 9580 12797 9604 12821
rect 9795 12796 9815 12816
rect 11580 12781 11600 12801
rect 11791 12776 11815 12800
rect 12000 12781 12024 12805
rect 12214 12777 12240 12803
rect 12628 12777 12648 12797
rect 12839 12772 12863 12796
rect 13048 12777 13072 12801
rect 13262 12773 13288 12799
rect 19863 12788 19889 12814
rect 20079 12786 20103 12810
rect 20288 12791 20312 12815
rect 20503 12790 20523 12810
rect 872 12108 892 12128
rect 1083 12103 1107 12127
rect 1292 12108 1316 12132
rect 1506 12104 1532 12130
rect 3367 12103 3387 12123
rect 3578 12098 3602 12122
rect 3787 12103 3811 12127
rect 4001 12099 4027 12125
rect 8107 12119 8133 12145
rect 8323 12117 8347 12141
rect 8532 12122 8556 12146
rect 8747 12121 8767 12141
rect 9155 12115 9181 12141
rect 9371 12113 9395 12137
rect 9580 12118 9604 12142
rect 9795 12117 9815 12137
rect 11580 12102 11600 12122
rect 11791 12097 11815 12121
rect 12000 12102 12024 12126
rect 12214 12098 12240 12124
rect 14075 12097 14095 12117
rect 14286 12092 14310 12116
rect 14495 12097 14519 12121
rect 14709 12093 14735 12119
rect 18815 12113 18841 12139
rect 19031 12111 19055 12135
rect 19240 12116 19264 12140
rect 19455 12115 19475 12135
rect 19863 12109 19889 12135
rect 20079 12107 20103 12131
rect 20288 12112 20312 12136
rect 20503 12111 20523 12131
rect 872 11340 892 11360
rect 1083 11335 1107 11359
rect 1292 11340 1316 11364
rect 1506 11336 1532 11362
rect 1920 11336 1940 11356
rect 2131 11331 2155 11355
rect 2340 11336 2364 11360
rect 2554 11332 2580 11358
rect 6660 11352 6686 11378
rect 6876 11350 6900 11374
rect 7085 11355 7109 11379
rect 7300 11354 7320 11374
rect 9155 11347 9181 11373
rect 9371 11345 9395 11369
rect 9580 11350 9604 11374
rect 9795 11349 9815 11369
rect 11580 11334 11600 11354
rect 11791 11329 11815 11353
rect 12000 11334 12024 11358
rect 12214 11330 12240 11356
rect 12628 11330 12648 11350
rect 12839 11325 12863 11349
rect 13048 11330 13072 11354
rect 13262 11326 13288 11352
rect 17368 11346 17394 11372
rect 17584 11344 17608 11368
rect 17793 11349 17817 11373
rect 18008 11348 18028 11368
rect 19863 11341 19889 11367
rect 20079 11339 20103 11363
rect 20288 11344 20312 11368
rect 20503 11343 20523 11363
rect 872 10661 892 10681
rect 1083 10656 1107 10680
rect 1292 10661 1316 10685
rect 1506 10657 1532 10683
rect 3410 10658 3430 10678
rect 3621 10653 3645 10677
rect 3830 10658 3854 10682
rect 4044 10654 4070 10680
rect 8107 10672 8133 10698
rect 8323 10670 8347 10694
rect 8532 10675 8556 10699
rect 8747 10674 8767 10694
rect 9155 10668 9181 10694
rect 9371 10666 9395 10690
rect 9580 10671 9604 10695
rect 9795 10670 9815 10690
rect 11580 10655 11600 10675
rect 11791 10650 11815 10674
rect 12000 10655 12024 10679
rect 12214 10651 12240 10677
rect 14118 10652 14138 10672
rect 14329 10647 14353 10671
rect 14538 10652 14562 10676
rect 14752 10648 14778 10674
rect 18815 10666 18841 10692
rect 19031 10664 19055 10688
rect 19240 10669 19264 10693
rect 19455 10668 19475 10688
rect 19863 10662 19889 10688
rect 20079 10660 20103 10684
rect 20288 10665 20312 10689
rect 20503 10664 20523 10684
rect 873 9820 893 9840
rect 1084 9815 1108 9839
rect 1293 9820 1317 9844
rect 1507 9816 1533 9842
rect 1921 9816 1941 9836
rect 2132 9811 2156 9835
rect 2341 9816 2365 9840
rect 2555 9812 2581 9838
rect 6618 9830 6644 9856
rect 6834 9828 6858 9852
rect 7043 9833 7067 9857
rect 7258 9832 7278 9852
rect 9156 9827 9182 9853
rect 9372 9825 9396 9849
rect 9581 9830 9605 9854
rect 9796 9829 9816 9849
rect 11581 9814 11601 9834
rect 11792 9809 11816 9833
rect 12001 9814 12025 9838
rect 12215 9810 12241 9836
rect 12629 9810 12649 9830
rect 12840 9805 12864 9829
rect 13049 9810 13073 9834
rect 13263 9806 13289 9832
rect 17326 9824 17352 9850
rect 17542 9822 17566 9846
rect 17751 9827 17775 9851
rect 17966 9826 17986 9846
rect 19864 9821 19890 9847
rect 20080 9819 20104 9843
rect 20289 9824 20313 9848
rect 20504 9823 20524 9843
rect 873 9141 893 9161
rect 1084 9136 1108 9160
rect 1293 9141 1317 9165
rect 1507 9137 1533 9163
rect 3368 9136 3388 9156
rect 3579 9131 3603 9155
rect 3788 9136 3812 9160
rect 4002 9132 4028 9158
rect 8108 9152 8134 9178
rect 8324 9150 8348 9174
rect 8533 9155 8557 9179
rect 8748 9154 8768 9174
rect 9156 9148 9182 9174
rect 9372 9146 9396 9170
rect 9581 9151 9605 9175
rect 9796 9150 9816 9170
rect 11581 9135 11601 9155
rect 11792 9130 11816 9154
rect 12001 9135 12025 9159
rect 12215 9131 12241 9157
rect 14076 9130 14096 9150
rect 14287 9125 14311 9149
rect 14496 9130 14520 9154
rect 14710 9126 14736 9152
rect 18816 9146 18842 9172
rect 19032 9144 19056 9168
rect 19241 9149 19265 9173
rect 19456 9148 19476 9168
rect 19864 9142 19890 9168
rect 20080 9140 20104 9164
rect 20289 9145 20313 9169
rect 20504 9144 20524 9164
rect 873 8373 893 8393
rect 1084 8368 1108 8392
rect 1293 8373 1317 8397
rect 1507 8369 1533 8395
rect 1921 8369 1941 8389
rect 2132 8364 2156 8388
rect 2341 8369 2365 8393
rect 2555 8365 2581 8391
rect 6661 8385 6687 8411
rect 6877 8383 6901 8407
rect 7086 8388 7110 8412
rect 7301 8387 7321 8407
rect 9156 8380 9182 8406
rect 9372 8378 9396 8402
rect 9581 8383 9605 8407
rect 9796 8382 9816 8402
rect 11581 8367 11601 8387
rect 11792 8362 11816 8386
rect 12001 8367 12025 8391
rect 12215 8363 12241 8389
rect 12629 8363 12649 8383
rect 12840 8358 12864 8382
rect 13049 8363 13073 8387
rect 13263 8359 13289 8385
rect 17369 8379 17395 8405
rect 17585 8377 17609 8401
rect 17794 8382 17818 8406
rect 18009 8381 18029 8401
rect 19864 8374 19890 8400
rect 20080 8372 20104 8396
rect 20289 8377 20313 8401
rect 20504 8376 20524 8396
rect 873 7694 893 7714
rect 1084 7689 1108 7713
rect 1293 7694 1317 7718
rect 1507 7690 1533 7716
rect 4476 7685 4496 7705
rect 4687 7680 4711 7704
rect 4896 7685 4920 7709
rect 5110 7681 5136 7707
rect 8108 7705 8134 7731
rect 8324 7703 8348 7727
rect 8533 7708 8557 7732
rect 8748 7707 8768 7727
rect 9156 7701 9182 7727
rect 9372 7699 9396 7723
rect 9581 7704 9605 7728
rect 9796 7703 9816 7723
rect 11581 7688 11601 7708
rect 11792 7683 11816 7707
rect 12001 7688 12025 7712
rect 12215 7684 12241 7710
rect 15184 7679 15204 7699
rect 15395 7674 15419 7698
rect 15604 7679 15628 7703
rect 15818 7675 15844 7701
rect 18816 7699 18842 7725
rect 19032 7697 19056 7721
rect 19241 7702 19265 7726
rect 19456 7701 19476 7721
rect 19864 7695 19890 7721
rect 20080 7693 20104 7717
rect 20289 7698 20313 7722
rect 20504 7697 20524 7717
rect 870 6779 890 6799
rect 1081 6774 1105 6798
rect 1290 6779 1314 6803
rect 1504 6775 1530 6801
rect 1918 6775 1938 6795
rect 2129 6770 2153 6794
rect 2338 6775 2362 6799
rect 2552 6771 2578 6797
rect 5550 6795 5576 6821
rect 5766 6793 5790 6817
rect 5975 6798 5999 6822
rect 6190 6797 6210 6817
rect 9153 6786 9179 6812
rect 9369 6784 9393 6808
rect 9578 6789 9602 6813
rect 9793 6788 9813 6808
rect 11578 6773 11598 6793
rect 11789 6768 11813 6792
rect 11998 6773 12022 6797
rect 12212 6769 12238 6795
rect 12626 6769 12646 6789
rect 12837 6764 12861 6788
rect 13046 6769 13070 6793
rect 13260 6765 13286 6791
rect 16258 6789 16284 6815
rect 16474 6787 16498 6811
rect 16683 6792 16707 6816
rect 16898 6791 16918 6811
rect 19861 6780 19887 6806
rect 20077 6778 20101 6802
rect 20286 6783 20310 6807
rect 20501 6782 20521 6802
rect 870 6100 890 6120
rect 1081 6095 1105 6119
rect 1290 6100 1314 6124
rect 1504 6096 1530 6122
rect 3365 6095 3385 6115
rect 3576 6090 3600 6114
rect 3785 6095 3809 6119
rect 3999 6091 4025 6117
rect 8105 6111 8131 6137
rect 8321 6109 8345 6133
rect 8530 6114 8554 6138
rect 8745 6113 8765 6133
rect 9153 6107 9179 6133
rect 9369 6105 9393 6129
rect 9578 6110 9602 6134
rect 9793 6109 9813 6129
rect 11578 6094 11598 6114
rect 11789 6089 11813 6113
rect 11998 6094 12022 6118
rect 12212 6090 12238 6116
rect 14073 6089 14093 6109
rect 14284 6084 14308 6108
rect 14493 6089 14517 6113
rect 14707 6085 14733 6111
rect 18813 6105 18839 6131
rect 19029 6103 19053 6127
rect 19238 6108 19262 6132
rect 19453 6107 19473 6127
rect 19861 6101 19887 6127
rect 20077 6099 20101 6123
rect 20286 6104 20310 6128
rect 20501 6103 20521 6123
rect 870 5332 890 5352
rect 1081 5327 1105 5351
rect 1290 5332 1314 5356
rect 1504 5328 1530 5354
rect 1918 5328 1938 5348
rect 2129 5323 2153 5347
rect 2338 5328 2362 5352
rect 2552 5324 2578 5350
rect 6658 5344 6684 5370
rect 6874 5342 6898 5366
rect 7083 5347 7107 5371
rect 7298 5346 7318 5366
rect 9153 5339 9179 5365
rect 9369 5337 9393 5361
rect 9578 5342 9602 5366
rect 9793 5341 9813 5361
rect 11578 5326 11598 5346
rect 11789 5321 11813 5345
rect 11998 5326 12022 5350
rect 12212 5322 12238 5348
rect 12626 5322 12646 5342
rect 12837 5317 12861 5341
rect 13046 5322 13070 5346
rect 13260 5318 13286 5344
rect 17366 5338 17392 5364
rect 17582 5336 17606 5360
rect 17791 5341 17815 5365
rect 18006 5340 18026 5360
rect 19861 5333 19887 5359
rect 20077 5331 20101 5355
rect 20286 5336 20310 5360
rect 20501 5335 20521 5355
rect 870 4653 890 4673
rect 1081 4648 1105 4672
rect 1290 4653 1314 4677
rect 1504 4649 1530 4675
rect 3408 4650 3428 4670
rect 3619 4645 3643 4669
rect 3828 4650 3852 4674
rect 4042 4646 4068 4672
rect 8105 4664 8131 4690
rect 8321 4662 8345 4686
rect 8530 4667 8554 4691
rect 8745 4666 8765 4686
rect 9153 4660 9179 4686
rect 9369 4658 9393 4682
rect 9578 4663 9602 4687
rect 9793 4662 9813 4682
rect 11578 4647 11598 4667
rect 11789 4642 11813 4666
rect 11998 4647 12022 4671
rect 12212 4643 12238 4669
rect 14116 4644 14136 4664
rect 14327 4639 14351 4663
rect 14536 4644 14560 4668
rect 14750 4640 14776 4666
rect 18813 4658 18839 4684
rect 19029 4656 19053 4680
rect 19238 4661 19262 4685
rect 19453 4660 19473 4680
rect 19861 4654 19887 4680
rect 20077 4652 20101 4676
rect 20286 4657 20310 4681
rect 20501 4656 20521 4676
rect 871 3812 891 3832
rect 1082 3807 1106 3831
rect 1291 3812 1315 3836
rect 1505 3808 1531 3834
rect 1919 3808 1939 3828
rect 2130 3803 2154 3827
rect 2339 3808 2363 3832
rect 2553 3804 2579 3830
rect 4821 3814 4841 3834
rect 5032 3809 5056 3833
rect 5241 3814 5265 3838
rect 5455 3810 5481 3836
rect 6616 3822 6642 3848
rect 6832 3820 6856 3844
rect 7041 3825 7065 3849
rect 7256 3824 7276 3844
rect 9154 3819 9180 3845
rect 9370 3817 9394 3841
rect 9579 3822 9603 3846
rect 9794 3821 9814 3841
rect 11579 3806 11599 3826
rect 11790 3801 11814 3825
rect 11999 3806 12023 3830
rect 12213 3802 12239 3828
rect 12627 3802 12647 3822
rect 12838 3797 12862 3821
rect 13047 3802 13071 3826
rect 13261 3798 13287 3824
rect 15529 3808 15549 3828
rect 15740 3803 15764 3827
rect 15949 3808 15973 3832
rect 16163 3804 16189 3830
rect 17324 3816 17350 3842
rect 17540 3814 17564 3838
rect 17749 3819 17773 3843
rect 17964 3818 17984 3838
rect 19862 3813 19888 3839
rect 20078 3811 20102 3835
rect 20287 3816 20311 3840
rect 20502 3815 20522 3835
rect 871 3133 891 3153
rect 1082 3128 1106 3152
rect 1291 3133 1315 3157
rect 1505 3129 1531 3155
rect 3366 3128 3386 3148
rect 3577 3123 3601 3147
rect 3786 3128 3810 3152
rect 4000 3124 4026 3150
rect 8106 3144 8132 3170
rect 8322 3142 8346 3166
rect 8531 3147 8555 3171
rect 8746 3146 8766 3166
rect 9154 3140 9180 3166
rect 9370 3138 9394 3162
rect 9579 3143 9603 3167
rect 9794 3142 9814 3162
rect 11579 3127 11599 3147
rect 11790 3122 11814 3146
rect 11999 3127 12023 3151
rect 12213 3123 12239 3149
rect 14074 3122 14094 3142
rect 14285 3117 14309 3141
rect 14494 3122 14518 3146
rect 14708 3118 14734 3144
rect 18814 3138 18840 3164
rect 19030 3136 19054 3160
rect 19239 3141 19263 3165
rect 19454 3140 19474 3160
rect 19862 3134 19888 3160
rect 20078 3132 20102 3156
rect 20287 3137 20311 3161
rect 20502 3136 20522 3156
rect 871 2365 891 2385
rect 1082 2360 1106 2384
rect 1291 2365 1315 2389
rect 1505 2361 1531 2387
rect 1919 2361 1939 2381
rect 2130 2356 2154 2380
rect 2339 2361 2363 2385
rect 2553 2357 2579 2383
rect 6659 2377 6685 2403
rect 6875 2375 6899 2399
rect 7084 2380 7108 2404
rect 7299 2379 7319 2399
rect 9154 2372 9180 2398
rect 9370 2370 9394 2394
rect 9579 2375 9603 2399
rect 9794 2374 9814 2394
rect 11579 2359 11599 2379
rect 11790 2354 11814 2378
rect 11999 2359 12023 2383
rect 12213 2355 12239 2381
rect 12627 2355 12647 2375
rect 12838 2350 12862 2374
rect 13047 2355 13071 2379
rect 13261 2351 13287 2377
rect 17367 2371 17393 2397
rect 17583 2369 17607 2393
rect 17792 2374 17816 2398
rect 18007 2373 18027 2393
rect 19862 2366 19888 2392
rect 20078 2364 20102 2388
rect 20287 2369 20311 2393
rect 20502 2368 20522 2388
rect 871 1686 891 1706
rect 1082 1681 1106 1705
rect 1291 1686 1315 1710
rect 1505 1682 1531 1708
rect 8106 1697 8132 1723
rect 8322 1695 8346 1719
rect 8531 1700 8555 1724
rect 8746 1699 8766 1719
rect 9154 1693 9180 1719
rect 9370 1691 9394 1715
rect 9579 1696 9603 1720
rect 9794 1695 9814 1715
rect 11579 1680 11599 1700
rect 11790 1675 11814 1699
rect 11999 1680 12023 1704
rect 12213 1676 12239 1702
rect 18814 1691 18840 1717
rect 19030 1689 19054 1713
rect 19239 1694 19263 1718
rect 19454 1693 19474 1713
rect 19862 1687 19888 1713
rect 20078 1685 20102 1709
rect 20287 1690 20311 1714
rect 20502 1689 20522 1709
rect 10582 -473 10602 -453
rect 10793 -478 10817 -454
rect 11002 -473 11026 -449
rect 11216 -477 11242 -451
<< ndiffres >>
rect 480 13069 537 13088
rect 480 13066 501 13069
rect 386 13051 501 13066
rect 519 13051 537 13069
rect 11188 13063 11245 13082
rect 11188 13060 11209 13063
rect 386 13028 537 13051
rect 11094 13045 11209 13060
rect 11227 13045 11245 13063
rect 386 12992 428 13028
rect 11094 13022 11245 13045
rect 385 12991 485 12992
rect 385 12970 541 12991
rect 385 12952 503 12970
rect 521 12952 541 12970
rect 11094 12986 11136 13022
rect 11093 12985 11193 12986
rect 385 12948 541 12952
rect 480 12932 541 12948
rect 11093 12964 11249 12985
rect 11093 12946 11211 12964
rect 11229 12946 11249 12964
rect 11093 12942 11249 12946
rect 480 12813 537 12832
rect 480 12810 501 12813
rect 386 12795 501 12810
rect 519 12795 537 12813
rect 386 12772 537 12795
rect 386 12736 428 12772
rect 11188 12926 11249 12942
rect 10146 12882 10207 12898
rect 10146 12878 10302 12882
rect 10146 12860 10166 12878
rect 10184 12860 10302 12878
rect 385 12735 485 12736
rect 385 12714 541 12735
rect 10146 12839 10302 12860
rect 10202 12838 10302 12839
rect 10259 12802 10301 12838
rect 11188 12807 11245 12826
rect 11188 12804 11209 12807
rect 10150 12779 10301 12802
rect 385 12696 503 12714
rect 521 12696 541 12714
rect 385 12692 541 12696
rect 480 12676 541 12692
rect 10150 12761 10168 12779
rect 10186 12764 10301 12779
rect 11094 12789 11209 12804
rect 11227 12789 11245 12807
rect 11094 12766 11245 12789
rect 10186 12761 10207 12764
rect 10150 12742 10207 12761
rect 11094 12730 11136 12766
rect 20854 12876 20915 12892
rect 20854 12872 21010 12876
rect 20854 12854 20874 12872
rect 20892 12854 21010 12872
rect 11093 12729 11193 12730
rect 11093 12708 11249 12729
rect 20854 12833 21010 12854
rect 20910 12832 21010 12833
rect 20967 12796 21009 12832
rect 20858 12773 21009 12796
rect 11093 12690 11211 12708
rect 11229 12690 11249 12708
rect 11093 12686 11249 12690
rect 11188 12670 11249 12686
rect 10146 12627 10207 12643
rect 10146 12623 10302 12627
rect 10146 12605 10166 12623
rect 10184 12605 10302 12623
rect 20858 12755 20876 12773
rect 20894 12758 21009 12773
rect 20894 12755 20915 12758
rect 20858 12736 20915 12755
rect 10146 12584 10302 12605
rect 10202 12583 10302 12584
rect 10259 12547 10301 12583
rect 20854 12621 20915 12637
rect 20854 12617 21010 12621
rect 20854 12599 20874 12617
rect 20892 12599 21010 12617
rect 20854 12578 21010 12599
rect 20910 12577 21010 12578
rect 10150 12524 10301 12547
rect 20967 12541 21009 12577
rect 10150 12506 10168 12524
rect 10186 12509 10301 12524
rect 20858 12518 21009 12541
rect 10186 12506 10207 12509
rect 10150 12487 10207 12506
rect 20858 12500 20876 12518
rect 20894 12503 21009 12518
rect 20894 12500 20915 12503
rect 20858 12481 20915 12500
rect 480 12418 537 12437
rect 480 12415 501 12418
rect 386 12400 501 12415
rect 519 12400 537 12418
rect 11188 12412 11245 12431
rect 11188 12409 11209 12412
rect 386 12377 537 12400
rect 11094 12394 11209 12409
rect 11227 12394 11245 12412
rect 386 12341 428 12377
rect 11094 12371 11245 12394
rect 385 12340 485 12341
rect 385 12319 541 12340
rect 385 12301 503 12319
rect 521 12301 541 12319
rect 385 12297 541 12301
rect 480 12281 541 12297
rect 11094 12335 11136 12371
rect 11093 12334 11193 12335
rect 11093 12313 11249 12334
rect 480 12163 537 12182
rect 480 12160 501 12163
rect 386 12145 501 12160
rect 519 12145 537 12163
rect 11093 12295 11211 12313
rect 11229 12295 11249 12313
rect 11093 12291 11249 12295
rect 11188 12275 11249 12291
rect 386 12122 537 12145
rect 386 12086 428 12122
rect 385 12085 485 12086
rect 385 12064 541 12085
rect 10146 12232 10207 12248
rect 10146 12228 10302 12232
rect 10146 12210 10166 12228
rect 10184 12210 10302 12228
rect 385 12046 503 12064
rect 521 12046 541 12064
rect 385 12042 541 12046
rect 480 12026 541 12042
rect 10146 12189 10302 12210
rect 10202 12188 10302 12189
rect 10259 12152 10301 12188
rect 11188 12157 11245 12176
rect 11188 12154 11209 12157
rect 10150 12129 10301 12152
rect 10150 12111 10168 12129
rect 10186 12114 10301 12129
rect 11094 12139 11209 12154
rect 11227 12139 11245 12157
rect 11094 12116 11245 12139
rect 10186 12111 10207 12114
rect 10150 12092 10207 12111
rect 11094 12080 11136 12116
rect 11093 12079 11193 12080
rect 11093 12058 11249 12079
rect 20854 12226 20915 12242
rect 20854 12222 21010 12226
rect 20854 12204 20874 12222
rect 20892 12204 21010 12222
rect 11093 12040 11211 12058
rect 11229 12040 11249 12058
rect 11093 12036 11249 12040
rect 11188 12020 11249 12036
rect 20854 12183 21010 12204
rect 20910 12182 21010 12183
rect 10146 11976 10207 11992
rect 20967 12146 21009 12182
rect 20858 12123 21009 12146
rect 20858 12105 20876 12123
rect 20894 12108 21009 12123
rect 20894 12105 20915 12108
rect 20858 12086 20915 12105
rect 10146 11972 10302 11976
rect 10146 11954 10166 11972
rect 10184 11954 10302 11972
rect 10146 11933 10302 11954
rect 20854 11970 20915 11986
rect 20854 11966 21010 11970
rect 10202 11932 10302 11933
rect 10259 11896 10301 11932
rect 20854 11948 20874 11966
rect 20892 11948 21010 11966
rect 20854 11927 21010 11948
rect 20910 11926 21010 11927
rect 10150 11873 10301 11896
rect 20967 11890 21009 11926
rect 10150 11855 10168 11873
rect 10186 11858 10301 11873
rect 20858 11867 21009 11890
rect 10186 11855 10207 11858
rect 10150 11836 10207 11855
rect 20858 11849 20876 11867
rect 20894 11852 21009 11867
rect 20894 11849 20915 11852
rect 20858 11830 20915 11849
rect 480 11622 537 11641
rect 480 11619 501 11622
rect 386 11604 501 11619
rect 519 11604 537 11622
rect 11188 11616 11245 11635
rect 11188 11613 11209 11616
rect 386 11581 537 11604
rect 11094 11598 11209 11613
rect 11227 11598 11245 11616
rect 386 11545 428 11581
rect 11094 11575 11245 11598
rect 385 11544 485 11545
rect 385 11523 541 11544
rect 385 11505 503 11523
rect 521 11505 541 11523
rect 11094 11539 11136 11575
rect 11093 11538 11193 11539
rect 385 11501 541 11505
rect 480 11485 541 11501
rect 11093 11517 11249 11538
rect 11093 11499 11211 11517
rect 11229 11499 11249 11517
rect 11093 11495 11249 11499
rect 480 11366 537 11385
rect 480 11363 501 11366
rect 386 11348 501 11363
rect 519 11348 537 11366
rect 386 11325 537 11348
rect 386 11289 428 11325
rect 11188 11479 11249 11495
rect 385 11288 485 11289
rect 385 11267 541 11288
rect 10146 11435 10207 11451
rect 10146 11431 10302 11435
rect 10146 11413 10166 11431
rect 10184 11413 10302 11431
rect 385 11249 503 11267
rect 521 11249 541 11267
rect 385 11245 541 11249
rect 480 11229 541 11245
rect 10146 11392 10302 11413
rect 10202 11391 10302 11392
rect 10259 11355 10301 11391
rect 11188 11360 11245 11379
rect 11188 11357 11209 11360
rect 10150 11332 10301 11355
rect 10150 11314 10168 11332
rect 10186 11317 10301 11332
rect 11094 11342 11209 11357
rect 11227 11342 11245 11360
rect 11094 11319 11245 11342
rect 10186 11314 10207 11317
rect 10150 11295 10207 11314
rect 11094 11283 11136 11319
rect 11093 11282 11193 11283
rect 11093 11261 11249 11282
rect 20854 11429 20915 11445
rect 20854 11425 21010 11429
rect 20854 11407 20874 11425
rect 20892 11407 21010 11425
rect 11093 11243 11211 11261
rect 11229 11243 11249 11261
rect 11093 11239 11249 11243
rect 11188 11223 11249 11239
rect 20854 11386 21010 11407
rect 20910 11385 21010 11386
rect 20967 11349 21009 11385
rect 20858 11326 21009 11349
rect 10146 11180 10207 11196
rect 10146 11176 10302 11180
rect 10146 11158 10166 11176
rect 10184 11158 10302 11176
rect 20858 11308 20876 11326
rect 20894 11311 21009 11326
rect 20894 11308 20915 11311
rect 20858 11289 20915 11308
rect 10146 11137 10302 11158
rect 10202 11136 10302 11137
rect 10259 11100 10301 11136
rect 20854 11174 20915 11190
rect 20854 11170 21010 11174
rect 20854 11152 20874 11170
rect 20892 11152 21010 11170
rect 20854 11131 21010 11152
rect 20910 11130 21010 11131
rect 10150 11077 10301 11100
rect 20967 11094 21009 11130
rect 10150 11059 10168 11077
rect 10186 11062 10301 11077
rect 20858 11071 21009 11094
rect 10186 11059 10207 11062
rect 10150 11040 10207 11059
rect 20858 11053 20876 11071
rect 20894 11056 21009 11071
rect 20894 11053 20915 11056
rect 20858 11034 20915 11053
rect 480 10971 537 10990
rect 480 10968 501 10971
rect 386 10953 501 10968
rect 519 10953 537 10971
rect 11188 10965 11245 10984
rect 11188 10962 11209 10965
rect 386 10930 537 10953
rect 11094 10947 11209 10962
rect 11227 10947 11245 10965
rect 386 10894 428 10930
rect 11094 10924 11245 10947
rect 385 10893 485 10894
rect 385 10872 541 10893
rect 385 10854 503 10872
rect 521 10854 541 10872
rect 385 10850 541 10854
rect 480 10834 541 10850
rect 11094 10888 11136 10924
rect 11093 10887 11193 10888
rect 11093 10866 11249 10887
rect 480 10716 537 10735
rect 480 10713 501 10716
rect 386 10698 501 10713
rect 519 10698 537 10716
rect 11093 10848 11211 10866
rect 11229 10848 11249 10866
rect 11093 10844 11249 10848
rect 11188 10828 11249 10844
rect 386 10675 537 10698
rect 386 10639 428 10675
rect 385 10638 485 10639
rect 385 10617 541 10638
rect 10146 10785 10207 10801
rect 10146 10781 10302 10785
rect 10146 10763 10166 10781
rect 10184 10763 10302 10781
rect 385 10599 503 10617
rect 521 10599 541 10617
rect 385 10595 541 10599
rect 480 10579 541 10595
rect 10146 10742 10302 10763
rect 10202 10741 10302 10742
rect 10259 10705 10301 10741
rect 11188 10710 11245 10729
rect 11188 10707 11209 10710
rect 10150 10682 10301 10705
rect 10150 10664 10168 10682
rect 10186 10667 10301 10682
rect 11094 10692 11209 10707
rect 11227 10692 11245 10710
rect 11094 10669 11245 10692
rect 10186 10664 10207 10667
rect 10150 10645 10207 10664
rect 11094 10633 11136 10669
rect 11093 10632 11193 10633
rect 11093 10611 11249 10632
rect 20854 10779 20915 10795
rect 20854 10775 21010 10779
rect 20854 10757 20874 10775
rect 20892 10757 21010 10775
rect 11093 10593 11211 10611
rect 11229 10593 11249 10611
rect 11093 10589 11249 10593
rect 11188 10573 11249 10589
rect 20854 10736 21010 10757
rect 20910 10735 21010 10736
rect 10146 10529 10207 10545
rect 20967 10699 21009 10735
rect 20858 10676 21009 10699
rect 20858 10658 20876 10676
rect 20894 10661 21009 10676
rect 20894 10658 20915 10661
rect 20858 10639 20915 10658
rect 10146 10525 10302 10529
rect 10146 10507 10166 10525
rect 10184 10507 10302 10525
rect 10146 10486 10302 10507
rect 10202 10485 10302 10486
rect 10259 10449 10301 10485
rect 20854 10523 20915 10539
rect 20854 10519 21010 10523
rect 20854 10501 20874 10519
rect 20892 10501 21010 10519
rect 20854 10480 21010 10501
rect 20910 10479 21010 10480
rect 10150 10426 10301 10449
rect 20967 10443 21009 10479
rect 10150 10408 10168 10426
rect 10186 10411 10301 10426
rect 20858 10420 21009 10443
rect 10186 10408 10207 10411
rect 10150 10389 10207 10408
rect 20858 10402 20876 10420
rect 20894 10405 21009 10420
rect 20894 10402 20915 10405
rect 20858 10383 20915 10402
rect 481 10102 538 10121
rect 481 10099 502 10102
rect 387 10084 502 10099
rect 520 10084 538 10102
rect 11189 10096 11246 10115
rect 11189 10093 11210 10096
rect 387 10061 538 10084
rect 11095 10078 11210 10093
rect 11228 10078 11246 10096
rect 387 10025 429 10061
rect 11095 10055 11246 10078
rect 386 10024 486 10025
rect 386 10003 542 10024
rect 386 9985 504 10003
rect 522 9985 542 10003
rect 386 9981 542 9985
rect 481 9965 542 9981
rect 11095 10019 11137 10055
rect 11094 10018 11194 10019
rect 11094 9997 11250 10018
rect 11094 9979 11212 9997
rect 11230 9979 11250 9997
rect 11094 9975 11250 9979
rect 481 9846 538 9865
rect 481 9843 502 9846
rect 387 9828 502 9843
rect 520 9828 538 9846
rect 387 9805 538 9828
rect 387 9769 429 9805
rect 11189 9959 11250 9975
rect 386 9768 486 9769
rect 386 9747 542 9768
rect 10147 9915 10208 9931
rect 10147 9911 10303 9915
rect 10147 9893 10167 9911
rect 10185 9893 10303 9911
rect 386 9729 504 9747
rect 522 9729 542 9747
rect 386 9725 542 9729
rect 481 9709 542 9725
rect 10147 9872 10303 9893
rect 10203 9871 10303 9872
rect 10260 9835 10302 9871
rect 11189 9840 11246 9859
rect 11189 9837 11210 9840
rect 10151 9812 10302 9835
rect 10151 9794 10169 9812
rect 10187 9797 10302 9812
rect 11095 9822 11210 9837
rect 11228 9822 11246 9840
rect 11095 9799 11246 9822
rect 10187 9794 10208 9797
rect 10151 9775 10208 9794
rect 11095 9763 11137 9799
rect 11094 9762 11194 9763
rect 11094 9741 11250 9762
rect 20855 9909 20916 9925
rect 20855 9905 21011 9909
rect 20855 9887 20875 9905
rect 20893 9887 21011 9905
rect 11094 9723 11212 9741
rect 11230 9723 11250 9741
rect 11094 9719 11250 9723
rect 11189 9703 11250 9719
rect 20855 9866 21011 9887
rect 20911 9865 21011 9866
rect 20968 9829 21010 9865
rect 20859 9806 21010 9829
rect 10147 9660 10208 9676
rect 10147 9656 10303 9660
rect 10147 9638 10167 9656
rect 10185 9638 10303 9656
rect 20859 9788 20877 9806
rect 20895 9791 21010 9806
rect 20895 9788 20916 9791
rect 20859 9769 20916 9788
rect 10147 9617 10303 9638
rect 10203 9616 10303 9617
rect 10260 9580 10302 9616
rect 20855 9654 20916 9670
rect 20855 9650 21011 9654
rect 20855 9632 20875 9650
rect 20893 9632 21011 9650
rect 20855 9611 21011 9632
rect 20911 9610 21011 9611
rect 10151 9557 10302 9580
rect 20968 9574 21010 9610
rect 10151 9539 10169 9557
rect 10187 9542 10302 9557
rect 20859 9551 21010 9574
rect 10187 9539 10208 9542
rect 10151 9520 10208 9539
rect 20859 9533 20877 9551
rect 20895 9536 21010 9551
rect 20895 9533 20916 9536
rect 20859 9514 20916 9533
rect 481 9451 538 9470
rect 481 9448 502 9451
rect 387 9433 502 9448
rect 520 9433 538 9451
rect 11189 9445 11246 9464
rect 11189 9442 11210 9445
rect 387 9410 538 9433
rect 11095 9427 11210 9442
rect 11228 9427 11246 9445
rect 387 9374 429 9410
rect 11095 9404 11246 9427
rect 386 9373 486 9374
rect 386 9352 542 9373
rect 386 9334 504 9352
rect 522 9334 542 9352
rect 386 9330 542 9334
rect 481 9314 542 9330
rect 11095 9368 11137 9404
rect 11094 9367 11194 9368
rect 11094 9346 11250 9367
rect 481 9196 538 9215
rect 481 9193 502 9196
rect 387 9178 502 9193
rect 520 9178 538 9196
rect 11094 9328 11212 9346
rect 11230 9328 11250 9346
rect 11094 9324 11250 9328
rect 11189 9308 11250 9324
rect 387 9155 538 9178
rect 387 9119 429 9155
rect 386 9118 486 9119
rect 386 9097 542 9118
rect 10147 9265 10208 9281
rect 10147 9261 10303 9265
rect 10147 9243 10167 9261
rect 10185 9243 10303 9261
rect 386 9079 504 9097
rect 522 9079 542 9097
rect 386 9075 542 9079
rect 481 9059 542 9075
rect 10147 9222 10303 9243
rect 10203 9221 10303 9222
rect 10260 9185 10302 9221
rect 11189 9190 11246 9209
rect 11189 9187 11210 9190
rect 10151 9162 10302 9185
rect 10151 9144 10169 9162
rect 10187 9147 10302 9162
rect 11095 9172 11210 9187
rect 11228 9172 11246 9190
rect 11095 9149 11246 9172
rect 10187 9144 10208 9147
rect 10151 9125 10208 9144
rect 11095 9113 11137 9149
rect 11094 9112 11194 9113
rect 11094 9091 11250 9112
rect 20855 9259 20916 9275
rect 20855 9255 21011 9259
rect 20855 9237 20875 9255
rect 20893 9237 21011 9255
rect 11094 9073 11212 9091
rect 11230 9073 11250 9091
rect 11094 9069 11250 9073
rect 11189 9053 11250 9069
rect 20855 9216 21011 9237
rect 20911 9215 21011 9216
rect 10147 9009 10208 9025
rect 20968 9179 21010 9215
rect 20859 9156 21010 9179
rect 20859 9138 20877 9156
rect 20895 9141 21010 9156
rect 20895 9138 20916 9141
rect 20859 9119 20916 9138
rect 10147 9005 10303 9009
rect 10147 8987 10167 9005
rect 10185 8987 10303 9005
rect 10147 8966 10303 8987
rect 20855 9003 20916 9019
rect 20855 8999 21011 9003
rect 10203 8965 10303 8966
rect 10260 8929 10302 8965
rect 20855 8981 20875 8999
rect 20893 8981 21011 8999
rect 20855 8960 21011 8981
rect 20911 8959 21011 8960
rect 10151 8906 10302 8929
rect 20968 8923 21010 8959
rect 10151 8888 10169 8906
rect 10187 8891 10302 8906
rect 20859 8900 21010 8923
rect 10187 8888 10208 8891
rect 10151 8869 10208 8888
rect 20859 8882 20877 8900
rect 20895 8885 21010 8900
rect 20895 8882 20916 8885
rect 20859 8863 20916 8882
rect 481 8655 538 8674
rect 481 8652 502 8655
rect 387 8637 502 8652
rect 520 8637 538 8655
rect 11189 8649 11246 8668
rect 11189 8646 11210 8649
rect 387 8614 538 8637
rect 11095 8631 11210 8646
rect 11228 8631 11246 8649
rect 387 8578 429 8614
rect 11095 8608 11246 8631
rect 386 8577 486 8578
rect 386 8556 542 8577
rect 386 8538 504 8556
rect 522 8538 542 8556
rect 11095 8572 11137 8608
rect 11094 8571 11194 8572
rect 386 8534 542 8538
rect 481 8518 542 8534
rect 11094 8550 11250 8571
rect 11094 8532 11212 8550
rect 11230 8532 11250 8550
rect 11094 8528 11250 8532
rect 481 8399 538 8418
rect 481 8396 502 8399
rect 387 8381 502 8396
rect 520 8381 538 8399
rect 387 8358 538 8381
rect 387 8322 429 8358
rect 11189 8512 11250 8528
rect 386 8321 486 8322
rect 386 8300 542 8321
rect 10147 8468 10208 8484
rect 10147 8464 10303 8468
rect 10147 8446 10167 8464
rect 10185 8446 10303 8464
rect 386 8282 504 8300
rect 522 8282 542 8300
rect 386 8278 542 8282
rect 481 8262 542 8278
rect 10147 8425 10303 8446
rect 10203 8424 10303 8425
rect 10260 8388 10302 8424
rect 11189 8393 11246 8412
rect 11189 8390 11210 8393
rect 10151 8365 10302 8388
rect 10151 8347 10169 8365
rect 10187 8350 10302 8365
rect 11095 8375 11210 8390
rect 11228 8375 11246 8393
rect 11095 8352 11246 8375
rect 10187 8347 10208 8350
rect 10151 8328 10208 8347
rect 11095 8316 11137 8352
rect 11094 8315 11194 8316
rect 11094 8294 11250 8315
rect 20855 8462 20916 8478
rect 20855 8458 21011 8462
rect 20855 8440 20875 8458
rect 20893 8440 21011 8458
rect 11094 8276 11212 8294
rect 11230 8276 11250 8294
rect 11094 8272 11250 8276
rect 11189 8256 11250 8272
rect 20855 8419 21011 8440
rect 20911 8418 21011 8419
rect 20968 8382 21010 8418
rect 20859 8359 21010 8382
rect 10147 8213 10208 8229
rect 10147 8209 10303 8213
rect 10147 8191 10167 8209
rect 10185 8191 10303 8209
rect 20859 8341 20877 8359
rect 20895 8344 21010 8359
rect 20895 8341 20916 8344
rect 20859 8322 20916 8341
rect 10147 8170 10303 8191
rect 10203 8169 10303 8170
rect 10260 8133 10302 8169
rect 20855 8207 20916 8223
rect 20855 8203 21011 8207
rect 20855 8185 20875 8203
rect 20893 8185 21011 8203
rect 20855 8164 21011 8185
rect 20911 8163 21011 8164
rect 10151 8110 10302 8133
rect 20968 8127 21010 8163
rect 10151 8092 10169 8110
rect 10187 8095 10302 8110
rect 20859 8104 21010 8127
rect 10187 8092 10208 8095
rect 10151 8073 10208 8092
rect 20859 8086 20877 8104
rect 20895 8089 21010 8104
rect 20895 8086 20916 8089
rect 20859 8067 20916 8086
rect 481 8004 538 8023
rect 481 8001 502 8004
rect 387 7986 502 8001
rect 520 7986 538 8004
rect 11189 7998 11246 8017
rect 11189 7995 11210 7998
rect 387 7963 538 7986
rect 11095 7980 11210 7995
rect 11228 7980 11246 7998
rect 387 7927 429 7963
rect 11095 7957 11246 7980
rect 386 7926 486 7927
rect 386 7905 542 7926
rect 386 7887 504 7905
rect 522 7887 542 7905
rect 386 7883 542 7887
rect 481 7867 542 7883
rect 11095 7921 11137 7957
rect 11094 7920 11194 7921
rect 11094 7899 11250 7920
rect 481 7749 538 7768
rect 481 7746 502 7749
rect 387 7731 502 7746
rect 520 7731 538 7749
rect 11094 7881 11212 7899
rect 11230 7881 11250 7899
rect 11094 7877 11250 7881
rect 11189 7861 11250 7877
rect 387 7708 538 7731
rect 387 7672 429 7708
rect 386 7671 486 7672
rect 386 7650 542 7671
rect 10147 7818 10208 7834
rect 10147 7814 10303 7818
rect 10147 7796 10167 7814
rect 10185 7796 10303 7814
rect 386 7632 504 7650
rect 522 7632 542 7650
rect 386 7628 542 7632
rect 481 7612 542 7628
rect 10147 7775 10303 7796
rect 10203 7774 10303 7775
rect 10260 7738 10302 7774
rect 11189 7743 11246 7762
rect 11189 7740 11210 7743
rect 10151 7715 10302 7738
rect 10151 7697 10169 7715
rect 10187 7700 10302 7715
rect 11095 7725 11210 7740
rect 11228 7725 11246 7743
rect 11095 7702 11246 7725
rect 10187 7697 10208 7700
rect 10151 7678 10208 7697
rect 11095 7666 11137 7702
rect 11094 7665 11194 7666
rect 11094 7644 11250 7665
rect 20855 7812 20916 7828
rect 20855 7808 21011 7812
rect 20855 7790 20875 7808
rect 20893 7790 21011 7808
rect 11094 7626 11212 7644
rect 11230 7626 11250 7644
rect 11094 7622 11250 7626
rect 11189 7606 11250 7622
rect 20855 7769 21011 7790
rect 20911 7768 21011 7769
rect 10147 7562 10208 7578
rect 20968 7732 21010 7768
rect 20859 7709 21010 7732
rect 20859 7691 20877 7709
rect 20895 7694 21010 7709
rect 20895 7691 20916 7694
rect 20859 7672 20916 7691
rect 10147 7558 10303 7562
rect 10147 7540 10167 7558
rect 10185 7540 10303 7558
rect 10147 7519 10303 7540
rect 10203 7518 10303 7519
rect 10260 7482 10302 7518
rect 20855 7556 20916 7572
rect 20855 7552 21011 7556
rect 20855 7534 20875 7552
rect 20893 7534 21011 7552
rect 20855 7513 21011 7534
rect 20911 7512 21011 7513
rect 10151 7459 10302 7482
rect 20968 7476 21010 7512
rect 10151 7441 10169 7459
rect 10187 7444 10302 7459
rect 20859 7453 21010 7476
rect 10187 7441 10208 7444
rect 10151 7422 10208 7441
rect 20859 7435 20877 7453
rect 20895 7438 21010 7453
rect 20895 7435 20916 7438
rect 20859 7416 20916 7435
rect 478 7061 535 7080
rect 478 7058 499 7061
rect 384 7043 499 7058
rect 517 7043 535 7061
rect 11186 7055 11243 7074
rect 11186 7052 11207 7055
rect 384 7020 535 7043
rect 11092 7037 11207 7052
rect 11225 7037 11243 7055
rect 384 6984 426 7020
rect 11092 7014 11243 7037
rect 383 6983 483 6984
rect 383 6962 539 6983
rect 383 6944 501 6962
rect 519 6944 539 6962
rect 383 6940 539 6944
rect 478 6924 539 6940
rect 11092 6978 11134 7014
rect 11091 6977 11191 6978
rect 11091 6956 11247 6977
rect 11091 6938 11209 6956
rect 11227 6938 11247 6956
rect 11091 6934 11247 6938
rect 478 6805 535 6824
rect 478 6802 499 6805
rect 384 6787 499 6802
rect 517 6787 535 6805
rect 384 6764 535 6787
rect 384 6728 426 6764
rect 11186 6918 11247 6934
rect 383 6727 483 6728
rect 383 6706 539 6727
rect 10144 6874 10205 6890
rect 10144 6870 10300 6874
rect 10144 6852 10164 6870
rect 10182 6852 10300 6870
rect 383 6688 501 6706
rect 519 6688 539 6706
rect 383 6684 539 6688
rect 478 6668 539 6684
rect 10144 6831 10300 6852
rect 10200 6830 10300 6831
rect 10257 6794 10299 6830
rect 11186 6799 11243 6818
rect 11186 6796 11207 6799
rect 10148 6771 10299 6794
rect 10148 6753 10166 6771
rect 10184 6756 10299 6771
rect 11092 6781 11207 6796
rect 11225 6781 11243 6799
rect 11092 6758 11243 6781
rect 10184 6753 10205 6756
rect 10148 6734 10205 6753
rect 11092 6722 11134 6758
rect 11091 6721 11191 6722
rect 11091 6700 11247 6721
rect 20852 6868 20913 6884
rect 20852 6864 21008 6868
rect 20852 6846 20872 6864
rect 20890 6846 21008 6864
rect 11091 6682 11209 6700
rect 11227 6682 11247 6700
rect 11091 6678 11247 6682
rect 11186 6662 11247 6678
rect 20852 6825 21008 6846
rect 20908 6824 21008 6825
rect 20965 6788 21007 6824
rect 20856 6765 21007 6788
rect 10144 6619 10205 6635
rect 10144 6615 10300 6619
rect 10144 6597 10164 6615
rect 10182 6597 10300 6615
rect 20856 6747 20874 6765
rect 20892 6750 21007 6765
rect 20892 6747 20913 6750
rect 20856 6728 20913 6747
rect 10144 6576 10300 6597
rect 10200 6575 10300 6576
rect 10257 6539 10299 6575
rect 20852 6613 20913 6629
rect 20852 6609 21008 6613
rect 20852 6591 20872 6609
rect 20890 6591 21008 6609
rect 20852 6570 21008 6591
rect 20908 6569 21008 6570
rect 10148 6516 10299 6539
rect 20965 6533 21007 6569
rect 10148 6498 10166 6516
rect 10184 6501 10299 6516
rect 20856 6510 21007 6533
rect 10184 6498 10205 6501
rect 10148 6479 10205 6498
rect 20856 6492 20874 6510
rect 20892 6495 21007 6510
rect 20892 6492 20913 6495
rect 20856 6473 20913 6492
rect 478 6410 535 6429
rect 478 6407 499 6410
rect 384 6392 499 6407
rect 517 6392 535 6410
rect 11186 6404 11243 6423
rect 11186 6401 11207 6404
rect 384 6369 535 6392
rect 11092 6386 11207 6401
rect 11225 6386 11243 6404
rect 384 6333 426 6369
rect 11092 6363 11243 6386
rect 383 6332 483 6333
rect 383 6311 539 6332
rect 383 6293 501 6311
rect 519 6293 539 6311
rect 383 6289 539 6293
rect 478 6273 539 6289
rect 11092 6327 11134 6363
rect 11091 6326 11191 6327
rect 11091 6305 11247 6326
rect 478 6155 535 6174
rect 478 6152 499 6155
rect 384 6137 499 6152
rect 517 6137 535 6155
rect 11091 6287 11209 6305
rect 11227 6287 11247 6305
rect 11091 6283 11247 6287
rect 11186 6267 11247 6283
rect 384 6114 535 6137
rect 384 6078 426 6114
rect 383 6077 483 6078
rect 383 6056 539 6077
rect 10144 6224 10205 6240
rect 10144 6220 10300 6224
rect 10144 6202 10164 6220
rect 10182 6202 10300 6220
rect 383 6038 501 6056
rect 519 6038 539 6056
rect 383 6034 539 6038
rect 478 6018 539 6034
rect 10144 6181 10300 6202
rect 10200 6180 10300 6181
rect 10257 6144 10299 6180
rect 11186 6149 11243 6168
rect 11186 6146 11207 6149
rect 10148 6121 10299 6144
rect 10148 6103 10166 6121
rect 10184 6106 10299 6121
rect 11092 6131 11207 6146
rect 11225 6131 11243 6149
rect 11092 6108 11243 6131
rect 10184 6103 10205 6106
rect 10148 6084 10205 6103
rect 11092 6072 11134 6108
rect 11091 6071 11191 6072
rect 11091 6050 11247 6071
rect 20852 6218 20913 6234
rect 20852 6214 21008 6218
rect 20852 6196 20872 6214
rect 20890 6196 21008 6214
rect 11091 6032 11209 6050
rect 11227 6032 11247 6050
rect 11091 6028 11247 6032
rect 11186 6012 11247 6028
rect 20852 6175 21008 6196
rect 20908 6174 21008 6175
rect 10144 5968 10205 5984
rect 20965 6138 21007 6174
rect 20856 6115 21007 6138
rect 20856 6097 20874 6115
rect 20892 6100 21007 6115
rect 20892 6097 20913 6100
rect 20856 6078 20913 6097
rect 10144 5964 10300 5968
rect 10144 5946 10164 5964
rect 10182 5946 10300 5964
rect 10144 5925 10300 5946
rect 20852 5962 20913 5978
rect 20852 5958 21008 5962
rect 10200 5924 10300 5925
rect 10257 5888 10299 5924
rect 20852 5940 20872 5958
rect 20890 5940 21008 5958
rect 20852 5919 21008 5940
rect 20908 5918 21008 5919
rect 10148 5865 10299 5888
rect 20965 5882 21007 5918
rect 10148 5847 10166 5865
rect 10184 5850 10299 5865
rect 20856 5859 21007 5882
rect 10184 5847 10205 5850
rect 10148 5828 10205 5847
rect 20856 5841 20874 5859
rect 20892 5844 21007 5859
rect 20892 5841 20913 5844
rect 20856 5822 20913 5841
rect 478 5614 535 5633
rect 478 5611 499 5614
rect 384 5596 499 5611
rect 517 5596 535 5614
rect 11186 5608 11243 5627
rect 11186 5605 11207 5608
rect 384 5573 535 5596
rect 11092 5590 11207 5605
rect 11225 5590 11243 5608
rect 384 5537 426 5573
rect 11092 5567 11243 5590
rect 383 5536 483 5537
rect 383 5515 539 5536
rect 383 5497 501 5515
rect 519 5497 539 5515
rect 11092 5531 11134 5567
rect 11091 5530 11191 5531
rect 383 5493 539 5497
rect 478 5477 539 5493
rect 11091 5509 11247 5530
rect 11091 5491 11209 5509
rect 11227 5491 11247 5509
rect 11091 5487 11247 5491
rect 478 5358 535 5377
rect 478 5355 499 5358
rect 384 5340 499 5355
rect 517 5340 535 5358
rect 384 5317 535 5340
rect 384 5281 426 5317
rect 11186 5471 11247 5487
rect 383 5280 483 5281
rect 383 5259 539 5280
rect 10144 5427 10205 5443
rect 10144 5423 10300 5427
rect 10144 5405 10164 5423
rect 10182 5405 10300 5423
rect 383 5241 501 5259
rect 519 5241 539 5259
rect 383 5237 539 5241
rect 478 5221 539 5237
rect 10144 5384 10300 5405
rect 10200 5383 10300 5384
rect 10257 5347 10299 5383
rect 11186 5352 11243 5371
rect 11186 5349 11207 5352
rect 10148 5324 10299 5347
rect 10148 5306 10166 5324
rect 10184 5309 10299 5324
rect 11092 5334 11207 5349
rect 11225 5334 11243 5352
rect 11092 5311 11243 5334
rect 10184 5306 10205 5309
rect 10148 5287 10205 5306
rect 11092 5275 11134 5311
rect 11091 5274 11191 5275
rect 11091 5253 11247 5274
rect 20852 5421 20913 5437
rect 20852 5417 21008 5421
rect 20852 5399 20872 5417
rect 20890 5399 21008 5417
rect 11091 5235 11209 5253
rect 11227 5235 11247 5253
rect 11091 5231 11247 5235
rect 11186 5215 11247 5231
rect 20852 5378 21008 5399
rect 20908 5377 21008 5378
rect 20965 5341 21007 5377
rect 20856 5318 21007 5341
rect 10144 5172 10205 5188
rect 10144 5168 10300 5172
rect 10144 5150 10164 5168
rect 10182 5150 10300 5168
rect 20856 5300 20874 5318
rect 20892 5303 21007 5318
rect 20892 5300 20913 5303
rect 20856 5281 20913 5300
rect 10144 5129 10300 5150
rect 10200 5128 10300 5129
rect 10257 5092 10299 5128
rect 20852 5166 20913 5182
rect 20852 5162 21008 5166
rect 20852 5144 20872 5162
rect 20890 5144 21008 5162
rect 20852 5123 21008 5144
rect 20908 5122 21008 5123
rect 10148 5069 10299 5092
rect 20965 5086 21007 5122
rect 10148 5051 10166 5069
rect 10184 5054 10299 5069
rect 20856 5063 21007 5086
rect 10184 5051 10205 5054
rect 10148 5032 10205 5051
rect 20856 5045 20874 5063
rect 20892 5048 21007 5063
rect 20892 5045 20913 5048
rect 20856 5026 20913 5045
rect 478 4963 535 4982
rect 478 4960 499 4963
rect 384 4945 499 4960
rect 517 4945 535 4963
rect 11186 4957 11243 4976
rect 11186 4954 11207 4957
rect 384 4922 535 4945
rect 11092 4939 11207 4954
rect 11225 4939 11243 4957
rect 384 4886 426 4922
rect 11092 4916 11243 4939
rect 383 4885 483 4886
rect 383 4864 539 4885
rect 383 4846 501 4864
rect 519 4846 539 4864
rect 383 4842 539 4846
rect 478 4826 539 4842
rect 11092 4880 11134 4916
rect 11091 4879 11191 4880
rect 11091 4858 11247 4879
rect 478 4708 535 4727
rect 478 4705 499 4708
rect 384 4690 499 4705
rect 517 4690 535 4708
rect 11091 4840 11209 4858
rect 11227 4840 11247 4858
rect 11091 4836 11247 4840
rect 11186 4820 11247 4836
rect 384 4667 535 4690
rect 384 4631 426 4667
rect 383 4630 483 4631
rect 383 4609 539 4630
rect 10144 4777 10205 4793
rect 10144 4773 10300 4777
rect 10144 4755 10164 4773
rect 10182 4755 10300 4773
rect 383 4591 501 4609
rect 519 4591 539 4609
rect 383 4587 539 4591
rect 478 4571 539 4587
rect 10144 4734 10300 4755
rect 10200 4733 10300 4734
rect 10257 4697 10299 4733
rect 11186 4702 11243 4721
rect 11186 4699 11207 4702
rect 10148 4674 10299 4697
rect 10148 4656 10166 4674
rect 10184 4659 10299 4674
rect 11092 4684 11207 4699
rect 11225 4684 11243 4702
rect 11092 4661 11243 4684
rect 10184 4656 10205 4659
rect 10148 4637 10205 4656
rect 11092 4625 11134 4661
rect 11091 4624 11191 4625
rect 11091 4603 11247 4624
rect 20852 4771 20913 4787
rect 20852 4767 21008 4771
rect 20852 4749 20872 4767
rect 20890 4749 21008 4767
rect 11091 4585 11209 4603
rect 11227 4585 11247 4603
rect 11091 4581 11247 4585
rect 11186 4565 11247 4581
rect 20852 4728 21008 4749
rect 20908 4727 21008 4728
rect 10144 4521 10205 4537
rect 20965 4691 21007 4727
rect 20856 4668 21007 4691
rect 20856 4650 20874 4668
rect 20892 4653 21007 4668
rect 20892 4650 20913 4653
rect 20856 4631 20913 4650
rect 10144 4517 10300 4521
rect 10144 4499 10164 4517
rect 10182 4499 10300 4517
rect 10144 4478 10300 4499
rect 10200 4477 10300 4478
rect 10257 4441 10299 4477
rect 20852 4515 20913 4531
rect 20852 4511 21008 4515
rect 20852 4493 20872 4511
rect 20890 4493 21008 4511
rect 20852 4472 21008 4493
rect 20908 4471 21008 4472
rect 10148 4418 10299 4441
rect 20965 4435 21007 4471
rect 10148 4400 10166 4418
rect 10184 4403 10299 4418
rect 20856 4412 21007 4435
rect 10184 4400 10205 4403
rect 10148 4381 10205 4400
rect 20856 4394 20874 4412
rect 20892 4397 21007 4412
rect 20892 4394 20913 4397
rect 20856 4375 20913 4394
rect 479 4094 536 4113
rect 479 4091 500 4094
rect 385 4076 500 4091
rect 518 4076 536 4094
rect 11187 4088 11244 4107
rect 11187 4085 11208 4088
rect 385 4053 536 4076
rect 11093 4070 11208 4085
rect 11226 4070 11244 4088
rect 385 4017 427 4053
rect 384 4016 484 4017
rect 384 3995 540 4016
rect 384 3977 502 3995
rect 520 3977 540 3995
rect 11093 4047 11244 4070
rect 384 3973 540 3977
rect 479 3957 540 3973
rect 479 3838 536 3857
rect 479 3835 500 3838
rect 385 3820 500 3835
rect 518 3820 536 3838
rect 385 3797 536 3820
rect 385 3761 427 3797
rect 11093 4011 11135 4047
rect 11092 4010 11192 4011
rect 11092 3989 11248 4010
rect 11092 3971 11210 3989
rect 11228 3971 11248 3989
rect 11092 3967 11248 3971
rect 11187 3951 11248 3967
rect 384 3760 484 3761
rect 384 3739 540 3760
rect 10145 3907 10206 3923
rect 10145 3903 10301 3907
rect 10145 3885 10165 3903
rect 10183 3885 10301 3903
rect 384 3721 502 3739
rect 520 3721 540 3739
rect 384 3717 540 3721
rect 479 3701 540 3717
rect 10145 3864 10301 3885
rect 10201 3863 10301 3864
rect 10258 3827 10300 3863
rect 11187 3832 11244 3851
rect 11187 3829 11208 3832
rect 10149 3804 10300 3827
rect 10149 3786 10167 3804
rect 10185 3789 10300 3804
rect 11093 3814 11208 3829
rect 11226 3814 11244 3832
rect 11093 3791 11244 3814
rect 10185 3786 10206 3789
rect 10149 3767 10206 3786
rect 11093 3755 11135 3791
rect 11092 3754 11192 3755
rect 11092 3733 11248 3754
rect 20853 3901 20914 3917
rect 20853 3897 21009 3901
rect 20853 3879 20873 3897
rect 20891 3879 21009 3897
rect 11092 3715 11210 3733
rect 11228 3715 11248 3733
rect 11092 3711 11248 3715
rect 11187 3695 11248 3711
rect 10145 3652 10206 3668
rect 10145 3648 10301 3652
rect 10145 3630 10165 3648
rect 10183 3630 10301 3648
rect 20853 3858 21009 3879
rect 20909 3857 21009 3858
rect 20966 3821 21008 3857
rect 20857 3798 21008 3821
rect 20857 3780 20875 3798
rect 20893 3783 21008 3798
rect 20893 3780 20914 3783
rect 20857 3761 20914 3780
rect 10145 3609 10301 3630
rect 10201 3608 10301 3609
rect 10258 3572 10300 3608
rect 20853 3646 20914 3662
rect 20853 3642 21009 3646
rect 20853 3624 20873 3642
rect 20891 3624 21009 3642
rect 20853 3603 21009 3624
rect 20909 3602 21009 3603
rect 10149 3549 10300 3572
rect 20966 3566 21008 3602
rect 10149 3531 10167 3549
rect 10185 3534 10300 3549
rect 20857 3543 21008 3566
rect 10185 3531 10206 3534
rect 10149 3512 10206 3531
rect 20857 3525 20875 3543
rect 20893 3528 21008 3543
rect 20893 3525 20914 3528
rect 20857 3506 20914 3525
rect 479 3443 536 3462
rect 479 3440 500 3443
rect 385 3425 500 3440
rect 518 3425 536 3443
rect 11187 3437 11244 3456
rect 11187 3434 11208 3437
rect 385 3402 536 3425
rect 11093 3419 11208 3434
rect 11226 3419 11244 3437
rect 385 3366 427 3402
rect 11093 3396 11244 3419
rect 384 3365 484 3366
rect 384 3344 540 3365
rect 384 3326 502 3344
rect 520 3326 540 3344
rect 384 3322 540 3326
rect 479 3306 540 3322
rect 11093 3360 11135 3396
rect 11092 3359 11192 3360
rect 11092 3338 11248 3359
rect 479 3188 536 3207
rect 479 3185 500 3188
rect 385 3170 500 3185
rect 518 3170 536 3188
rect 11092 3320 11210 3338
rect 11228 3320 11248 3338
rect 11092 3316 11248 3320
rect 11187 3300 11248 3316
rect 385 3147 536 3170
rect 385 3111 427 3147
rect 384 3110 484 3111
rect 384 3089 540 3110
rect 10145 3257 10206 3273
rect 10145 3253 10301 3257
rect 10145 3235 10165 3253
rect 10183 3235 10301 3253
rect 384 3071 502 3089
rect 520 3071 540 3089
rect 384 3067 540 3071
rect 479 3051 540 3067
rect 10145 3214 10301 3235
rect 10201 3213 10301 3214
rect 10258 3177 10300 3213
rect 11187 3182 11244 3201
rect 11187 3179 11208 3182
rect 10149 3154 10300 3177
rect 10149 3136 10167 3154
rect 10185 3139 10300 3154
rect 11093 3164 11208 3179
rect 11226 3164 11244 3182
rect 11093 3141 11244 3164
rect 10185 3136 10206 3139
rect 10149 3117 10206 3136
rect 11093 3105 11135 3141
rect 11092 3104 11192 3105
rect 11092 3083 11248 3104
rect 20853 3251 20914 3267
rect 20853 3247 21009 3251
rect 20853 3229 20873 3247
rect 20891 3229 21009 3247
rect 11092 3065 11210 3083
rect 11228 3065 11248 3083
rect 11092 3061 11248 3065
rect 11187 3045 11248 3061
rect 20853 3208 21009 3229
rect 20909 3207 21009 3208
rect 10145 3001 10206 3017
rect 20966 3171 21008 3207
rect 20857 3148 21008 3171
rect 20857 3130 20875 3148
rect 20893 3133 21008 3148
rect 20893 3130 20914 3133
rect 20857 3111 20914 3130
rect 10145 2997 10301 3001
rect 10145 2979 10165 2997
rect 10183 2979 10301 2997
rect 10145 2958 10301 2979
rect 20853 2995 20914 3011
rect 20853 2991 21009 2995
rect 10201 2957 10301 2958
rect 10258 2921 10300 2957
rect 20853 2973 20873 2991
rect 20891 2973 21009 2991
rect 20853 2952 21009 2973
rect 20909 2951 21009 2952
rect 10149 2898 10300 2921
rect 20966 2915 21008 2951
rect 10149 2880 10167 2898
rect 10185 2883 10300 2898
rect 20857 2892 21008 2915
rect 10185 2880 10206 2883
rect 10149 2861 10206 2880
rect 20857 2874 20875 2892
rect 20893 2877 21008 2892
rect 20893 2874 20914 2877
rect 20857 2855 20914 2874
rect 479 2647 536 2666
rect 479 2644 500 2647
rect 385 2629 500 2644
rect 518 2629 536 2647
rect 11187 2641 11244 2660
rect 11187 2638 11208 2641
rect 385 2606 536 2629
rect 11093 2623 11208 2638
rect 11226 2623 11244 2641
rect 385 2570 427 2606
rect 11093 2600 11244 2623
rect 384 2569 484 2570
rect 384 2548 540 2569
rect 384 2530 502 2548
rect 520 2530 540 2548
rect 11093 2564 11135 2600
rect 11092 2563 11192 2564
rect 384 2526 540 2530
rect 479 2510 540 2526
rect 11092 2542 11248 2563
rect 11092 2524 11210 2542
rect 11228 2524 11248 2542
rect 11092 2520 11248 2524
rect 479 2391 536 2410
rect 479 2388 500 2391
rect 385 2373 500 2388
rect 518 2373 536 2391
rect 385 2350 536 2373
rect 385 2314 427 2350
rect 11187 2504 11248 2520
rect 384 2313 484 2314
rect 384 2292 540 2313
rect 10145 2460 10206 2476
rect 10145 2456 10301 2460
rect 10145 2438 10165 2456
rect 10183 2438 10301 2456
rect 384 2274 502 2292
rect 520 2274 540 2292
rect 384 2270 540 2274
rect 479 2254 540 2270
rect 10145 2417 10301 2438
rect 10201 2416 10301 2417
rect 10258 2380 10300 2416
rect 11187 2385 11244 2404
rect 11187 2382 11208 2385
rect 10149 2357 10300 2380
rect 10149 2339 10167 2357
rect 10185 2342 10300 2357
rect 11093 2367 11208 2382
rect 11226 2367 11244 2385
rect 11093 2344 11244 2367
rect 10185 2339 10206 2342
rect 10149 2320 10206 2339
rect 11093 2308 11135 2344
rect 11092 2307 11192 2308
rect 11092 2286 11248 2307
rect 20853 2454 20914 2470
rect 20853 2450 21009 2454
rect 20853 2432 20873 2450
rect 20891 2432 21009 2450
rect 11092 2268 11210 2286
rect 11228 2268 11248 2286
rect 11092 2264 11248 2268
rect 11187 2248 11248 2264
rect 20853 2411 21009 2432
rect 20909 2410 21009 2411
rect 20966 2374 21008 2410
rect 20857 2351 21008 2374
rect 10145 2205 10206 2221
rect 10145 2201 10301 2205
rect 10145 2183 10165 2201
rect 10183 2183 10301 2201
rect 20857 2333 20875 2351
rect 20893 2336 21008 2351
rect 20893 2333 20914 2336
rect 20857 2314 20914 2333
rect 10145 2162 10301 2183
rect 10201 2161 10301 2162
rect 10258 2125 10300 2161
rect 20853 2199 20914 2215
rect 20853 2195 21009 2199
rect 20853 2177 20873 2195
rect 20891 2177 21009 2195
rect 20853 2156 21009 2177
rect 20909 2155 21009 2156
rect 10149 2102 10300 2125
rect 20966 2119 21008 2155
rect 10149 2084 10167 2102
rect 10185 2087 10300 2102
rect 20857 2096 21008 2119
rect 10185 2084 10206 2087
rect 10149 2065 10206 2084
rect 20857 2078 20875 2096
rect 20893 2081 21008 2096
rect 20893 2078 20914 2081
rect 20857 2059 20914 2078
rect 479 1996 536 2015
rect 479 1993 500 1996
rect 385 1978 500 1993
rect 518 1978 536 1996
rect 11187 1990 11244 2009
rect 11187 1987 11208 1990
rect 385 1955 536 1978
rect 11093 1972 11208 1987
rect 11226 1972 11244 1990
rect 385 1919 427 1955
rect 11093 1949 11244 1972
rect 384 1918 484 1919
rect 384 1897 540 1918
rect 384 1879 502 1897
rect 520 1879 540 1897
rect 384 1875 540 1879
rect 479 1859 540 1875
rect 11093 1913 11135 1949
rect 11092 1912 11192 1913
rect 11092 1891 11248 1912
rect 479 1741 536 1760
rect 479 1738 500 1741
rect 385 1723 500 1738
rect 518 1723 536 1741
rect 11092 1873 11210 1891
rect 11228 1873 11248 1891
rect 11092 1869 11248 1873
rect 11187 1853 11248 1869
rect 10145 1810 10206 1826
rect 10145 1806 10301 1810
rect 10145 1788 10165 1806
rect 10183 1788 10301 1806
rect 385 1700 536 1723
rect 385 1664 427 1700
rect 384 1663 484 1664
rect 384 1642 540 1663
rect 10145 1767 10301 1788
rect 10201 1766 10301 1767
rect 384 1624 502 1642
rect 520 1624 540 1642
rect 384 1620 540 1624
rect 479 1604 540 1620
rect 10258 1730 10300 1766
rect 11187 1735 11244 1754
rect 11187 1732 11208 1735
rect 10149 1707 10300 1730
rect 10149 1689 10167 1707
rect 10185 1692 10300 1707
rect 11093 1717 11208 1732
rect 11226 1717 11244 1735
rect 20853 1804 20914 1820
rect 20853 1800 21009 1804
rect 20853 1782 20873 1800
rect 20891 1782 21009 1800
rect 11093 1694 11244 1717
rect 10185 1689 10206 1692
rect 10149 1670 10206 1689
rect 11093 1658 11135 1694
rect 11092 1657 11192 1658
rect 11092 1636 11248 1657
rect 20853 1761 21009 1782
rect 20909 1760 21009 1761
rect 11092 1618 11210 1636
rect 11228 1618 11248 1636
rect 11092 1614 11248 1618
rect 11187 1598 11248 1614
rect 10145 1554 10206 1570
rect 20966 1724 21008 1760
rect 20857 1701 21008 1724
rect 20857 1683 20875 1701
rect 20893 1686 21008 1701
rect 20893 1683 20914 1686
rect 20857 1664 20914 1683
rect 10145 1550 10301 1554
rect 10145 1532 10165 1550
rect 10183 1532 10301 1550
rect 10145 1511 10301 1532
rect 10201 1510 10301 1511
rect 20853 1548 20914 1564
rect 20853 1544 21009 1548
rect 10258 1474 10300 1510
rect 20853 1526 20873 1544
rect 20891 1526 21009 1544
rect 20853 1505 21009 1526
rect 20909 1504 21009 1505
rect 10149 1451 10300 1474
rect 20966 1468 21008 1504
rect 10149 1433 10167 1451
rect 10185 1436 10300 1451
rect 20857 1445 21008 1468
rect 10185 1433 10206 1436
rect 10149 1414 10206 1433
rect 20857 1427 20875 1445
rect 20893 1430 21008 1445
rect 20893 1427 20914 1430
rect 20857 1408 20914 1427
<< locali >>
rect 2856 13693 2921 13704
rect 2856 13645 2869 13693
rect 2906 13645 2921 13693
rect 2856 13632 2921 13645
rect 479 13069 538 13452
rect 11187 13203 11246 13208
rect 3069 13152 3780 13154
rect 2442 13151 3780 13152
rect 1392 13150 1464 13151
rect 1391 13142 1490 13150
rect 1391 13139 1443 13142
rect 1391 13104 1399 13139
rect 1424 13104 1443 13139
rect 1468 13131 1490 13142
rect 2441 13143 3780 13151
rect 2441 13140 2493 13143
rect 1468 13130 2335 13131
rect 1468 13104 2336 13130
rect 1391 13094 2336 13104
rect 1391 13092 1490 13094
rect 479 13051 501 13069
rect 519 13051 538 13069
rect 479 13029 538 13051
rect 746 13065 1278 13070
rect 746 13045 1632 13065
rect 1652 13045 1655 13065
rect 2291 13061 2336 13094
rect 2441 13105 2449 13140
rect 2474 13105 2493 13140
rect 2518 13105 3780 13143
rect 2441 13096 3780 13105
rect 2441 13093 2530 13096
rect 3069 13094 3780 13096
rect 746 13041 1655 13045
rect 746 12994 789 13041
rect 1239 13040 1655 13041
rect 2287 13041 2680 13061
rect 2700 13041 2703 13061
rect 1239 13039 1580 13040
rect 896 13008 1006 13022
rect 896 13005 939 13008
rect 896 13000 900 13005
rect 734 12993 789 12994
rect 478 12970 789 12993
rect 478 12952 503 12970
rect 521 12958 789 12970
rect 818 12978 900 13000
rect 929 12978 939 13005
rect 967 12981 974 13008
rect 1003 13000 1006 13008
rect 1003 12981 1068 13000
rect 967 12978 1068 12981
rect 818 12976 1068 12978
rect 521 12952 543 12958
rect 478 12813 543 12952
rect 818 12897 855 12976
rect 896 12963 1006 12976
rect 970 12907 1001 12908
rect 818 12877 827 12897
rect 847 12877 855 12897
rect 478 12795 501 12813
rect 519 12795 543 12813
rect 478 12778 543 12795
rect 698 12859 766 12872
rect 818 12867 855 12877
rect 914 12897 1001 12907
rect 914 12877 923 12897
rect 943 12877 1001 12897
rect 914 12868 1001 12877
rect 914 12867 951 12868
rect 698 12817 705 12859
rect 754 12817 766 12859
rect 698 12814 766 12817
rect 970 12815 1001 12868
rect 1031 12897 1068 12976
rect 1183 12907 1214 12908
rect 1031 12877 1040 12897
rect 1060 12877 1068 12897
rect 1031 12867 1068 12877
rect 1127 12900 1214 12907
rect 1127 12897 1188 12900
rect 1127 12877 1136 12897
rect 1156 12880 1188 12897
rect 1209 12880 1214 12900
rect 1156 12877 1214 12880
rect 1127 12870 1214 12877
rect 1239 12897 1276 13039
rect 1542 13038 1579 13039
rect 2287 13036 2703 13041
rect 2287 13035 2628 13036
rect 1944 13004 2054 13018
rect 1944 13001 1987 13004
rect 1944 12996 1948 13001
rect 1866 12974 1948 12996
rect 1977 12974 1987 13001
rect 2015 12977 2022 13004
rect 2051 12996 2054 13004
rect 2051 12977 2116 12996
rect 2015 12974 2116 12977
rect 1866 12972 2116 12974
rect 1391 12907 1427 12908
rect 1239 12877 1248 12897
rect 1268 12877 1276 12897
rect 1127 12868 1183 12870
rect 1127 12867 1164 12868
rect 1239 12867 1276 12877
rect 1335 12897 1483 12907
rect 1583 12904 1679 12906
rect 1335 12877 1344 12897
rect 1364 12877 1454 12897
rect 1474 12877 1483 12897
rect 1335 12871 1483 12877
rect 1335 12868 1399 12871
rect 1335 12867 1372 12868
rect 1391 12841 1399 12868
rect 1420 12868 1483 12871
rect 1541 12897 1679 12904
rect 1541 12877 1550 12897
rect 1570 12877 1679 12897
rect 1541 12868 1679 12877
rect 1866 12893 1903 12972
rect 1944 12959 2054 12972
rect 2018 12903 2049 12904
rect 1866 12873 1875 12893
rect 1895 12873 1903 12893
rect 1420 12841 1427 12868
rect 1446 12867 1483 12868
rect 1542 12867 1579 12868
rect 1391 12816 1427 12841
rect 862 12814 903 12815
rect 698 12807 903 12814
rect 698 12796 872 12807
rect 698 12763 706 12796
rect 699 12754 706 12763
rect 755 12787 872 12796
rect 892 12787 903 12807
rect 755 12779 903 12787
rect 970 12811 1329 12815
rect 970 12806 1292 12811
rect 970 12782 1083 12806
rect 1107 12787 1292 12806
rect 1316 12787 1329 12811
rect 1107 12782 1329 12787
rect 970 12779 1329 12782
rect 1391 12779 1426 12816
rect 1494 12813 1594 12816
rect 1494 12809 1561 12813
rect 1494 12783 1506 12809
rect 1532 12787 1561 12809
rect 1587 12787 1594 12813
rect 1532 12783 1594 12787
rect 1494 12779 1594 12783
rect 755 12763 766 12779
rect 755 12754 763 12763
rect 970 12758 1001 12779
rect 1391 12758 1427 12779
rect 813 12757 850 12758
rect 478 12714 543 12733
rect 478 12696 503 12714
rect 521 12696 543 12714
rect 478 12495 543 12696
rect 699 12570 763 12754
rect 812 12748 850 12757
rect 812 12728 821 12748
rect 841 12728 850 12748
rect 812 12720 850 12728
rect 916 12752 1001 12758
rect 1026 12757 1063 12758
rect 916 12732 924 12752
rect 944 12732 1001 12752
rect 916 12724 1001 12732
rect 1025 12748 1063 12757
rect 1025 12728 1034 12748
rect 1054 12728 1063 12748
rect 916 12723 952 12724
rect 1025 12720 1063 12728
rect 1129 12752 1214 12758
rect 1234 12757 1271 12758
rect 1129 12732 1137 12752
rect 1157 12751 1214 12752
rect 1157 12732 1186 12751
rect 1129 12731 1186 12732
rect 1207 12731 1214 12751
rect 1129 12724 1214 12731
rect 1233 12748 1271 12757
rect 1233 12728 1242 12748
rect 1262 12728 1271 12748
rect 1129 12723 1165 12724
rect 1233 12720 1271 12728
rect 1337 12752 1481 12758
rect 1337 12732 1345 12752
rect 1365 12732 1453 12752
rect 1473 12732 1481 12752
rect 1337 12724 1481 12732
rect 1337 12723 1373 12724
rect 1445 12723 1481 12724
rect 1547 12757 1584 12758
rect 1547 12756 1585 12757
rect 1547 12748 1611 12756
rect 1547 12728 1556 12748
rect 1576 12734 1611 12748
rect 1631 12734 1634 12754
rect 1576 12729 1634 12734
rect 1576 12728 1611 12729
rect 813 12691 850 12720
rect 814 12689 850 12691
rect 1026 12689 1063 12720
rect 814 12667 1063 12689
rect 895 12661 1006 12667
rect 895 12653 936 12661
rect 895 12633 903 12653
rect 922 12633 936 12653
rect 895 12631 936 12633
rect 964 12653 1006 12661
rect 964 12633 980 12653
rect 999 12633 1006 12653
rect 964 12631 1006 12633
rect 895 12616 1006 12631
rect 699 12560 767 12570
rect 699 12527 716 12560
rect 756 12527 767 12560
rect 699 12515 767 12527
rect 699 12513 763 12515
rect 1234 12496 1271 12720
rect 1547 12716 1611 12728
rect 1651 12498 1678 12868
rect 1866 12863 1903 12873
rect 1962 12893 2049 12903
rect 1962 12873 1971 12893
rect 1991 12873 2049 12893
rect 1962 12864 2049 12873
rect 1962 12863 1999 12864
rect 1742 12850 1812 12855
rect 1737 12844 1812 12850
rect 1737 12811 1745 12844
rect 1798 12811 1812 12844
rect 2018 12811 2049 12864
rect 2079 12893 2116 12972
rect 2231 12903 2262 12904
rect 2079 12873 2088 12893
rect 2108 12873 2116 12893
rect 2079 12863 2116 12873
rect 2175 12896 2262 12903
rect 2175 12893 2236 12896
rect 2175 12873 2184 12893
rect 2204 12876 2236 12893
rect 2257 12876 2262 12896
rect 2204 12873 2262 12876
rect 2175 12866 2262 12873
rect 2287 12893 2324 13035
rect 2590 13034 2627 13035
rect 2439 12903 2475 12904
rect 2287 12873 2296 12893
rect 2316 12873 2324 12893
rect 2175 12864 2231 12866
rect 2175 12863 2212 12864
rect 2287 12863 2324 12873
rect 2383 12893 2531 12903
rect 2631 12900 2727 12902
rect 2383 12873 2392 12893
rect 2412 12873 2502 12893
rect 2522 12873 2531 12893
rect 2383 12867 2531 12873
rect 2383 12864 2447 12867
rect 2383 12863 2420 12864
rect 2439 12837 2447 12864
rect 2468 12864 2531 12867
rect 2589 12893 2727 12900
rect 2589 12873 2598 12893
rect 2618 12873 2727 12893
rect 2589 12864 2727 12873
rect 2468 12837 2475 12864
rect 2494 12863 2531 12864
rect 2590 12863 2627 12864
rect 2439 12812 2475 12837
rect 1737 12810 1820 12811
rect 1910 12810 1951 12811
rect 1737 12803 1951 12810
rect 1737 12786 1920 12803
rect 1737 12753 1750 12786
rect 1803 12783 1920 12786
rect 1940 12783 1951 12803
rect 1803 12775 1951 12783
rect 2018 12807 2377 12811
rect 2018 12802 2340 12807
rect 2018 12778 2131 12802
rect 2155 12783 2340 12802
rect 2364 12783 2377 12807
rect 2155 12778 2377 12783
rect 2018 12775 2377 12778
rect 2439 12775 2474 12812
rect 2542 12809 2642 12812
rect 2542 12805 2609 12809
rect 2542 12779 2554 12805
rect 2580 12783 2609 12805
rect 2635 12783 2642 12809
rect 2580 12779 2642 12783
rect 2542 12775 2642 12779
rect 1803 12753 1820 12775
rect 2018 12754 2049 12775
rect 2439 12754 2475 12775
rect 1861 12753 1898 12754
rect 1737 12739 1820 12753
rect 1510 12496 1678 12498
rect 1234 12495 1678 12496
rect 478 12465 1678 12495
rect 1748 12529 1820 12739
rect 1860 12744 1898 12753
rect 1860 12724 1869 12744
rect 1889 12724 1898 12744
rect 1860 12716 1898 12724
rect 1964 12748 2049 12754
rect 2074 12753 2111 12754
rect 1964 12728 1972 12748
rect 1992 12728 2049 12748
rect 1964 12720 2049 12728
rect 2073 12744 2111 12753
rect 2073 12724 2082 12744
rect 2102 12724 2111 12744
rect 1964 12719 2000 12720
rect 2073 12716 2111 12724
rect 2177 12748 2262 12754
rect 2282 12753 2319 12754
rect 2177 12728 2185 12748
rect 2205 12747 2262 12748
rect 2205 12728 2234 12747
rect 2177 12727 2234 12728
rect 2255 12727 2262 12747
rect 2177 12720 2262 12727
rect 2281 12744 2319 12753
rect 2281 12724 2290 12744
rect 2310 12724 2319 12744
rect 2177 12719 2213 12720
rect 2281 12716 2319 12724
rect 2385 12748 2529 12754
rect 2385 12728 2393 12748
rect 2413 12728 2501 12748
rect 2521 12728 2529 12748
rect 2385 12720 2529 12728
rect 2385 12719 2421 12720
rect 2493 12719 2529 12720
rect 2595 12753 2632 12754
rect 2595 12752 2633 12753
rect 2595 12744 2659 12752
rect 2595 12724 2604 12744
rect 2624 12730 2659 12744
rect 2679 12730 2682 12750
rect 2624 12725 2682 12730
rect 2624 12724 2659 12725
rect 1861 12687 1898 12716
rect 1862 12685 1898 12687
rect 2074 12685 2111 12716
rect 1862 12663 2111 12685
rect 1943 12657 2054 12663
rect 1943 12649 1984 12657
rect 1943 12629 1951 12649
rect 1970 12629 1984 12649
rect 1943 12627 1984 12629
rect 2012 12649 2054 12657
rect 2012 12629 2028 12649
rect 2047 12629 2054 12649
rect 2012 12627 2054 12629
rect 1943 12612 2054 12627
rect 1748 12490 1767 12529
rect 1812 12490 1820 12529
rect 1748 12473 1820 12490
rect 2282 12517 2319 12716
rect 2595 12712 2659 12724
rect 2282 12511 2323 12517
rect 2699 12513 2726 12864
rect 3021 12851 3116 12877
rect 2857 12829 2921 12848
rect 2857 12790 2870 12829
rect 2904 12790 2921 12829
rect 2857 12771 2921 12790
rect 2558 12511 2726 12513
rect 2282 12485 2726 12511
rect 478 12418 543 12465
rect 478 12400 501 12418
rect 519 12400 543 12418
rect 1391 12445 1426 12447
rect 1391 12443 1495 12445
rect 2284 12443 2323 12485
rect 2558 12484 2726 12485
rect 1391 12436 2325 12443
rect 1391 12435 1442 12436
rect 1391 12415 1394 12435
rect 1419 12416 1442 12435
rect 1474 12416 2325 12436
rect 1419 12415 2325 12416
rect 1391 12408 2325 12415
rect 1664 12407 2325 12408
rect 478 12379 543 12400
rect 755 12390 795 12393
rect 755 12386 1658 12390
rect 755 12366 1632 12386
rect 1652 12366 1658 12386
rect 755 12363 1658 12366
rect 479 12319 544 12339
rect 479 12301 503 12319
rect 521 12301 544 12319
rect 479 12274 544 12301
rect 755 12274 795 12363
rect 1239 12361 1655 12363
rect 1239 12360 1580 12361
rect 896 12329 1006 12343
rect 896 12326 939 12329
rect 896 12321 900 12326
rect 478 12239 795 12274
rect 818 12299 900 12321
rect 929 12299 939 12326
rect 967 12302 974 12329
rect 1003 12321 1006 12329
rect 1003 12302 1068 12321
rect 967 12299 1068 12302
rect 818 12297 1068 12299
rect 479 12163 544 12239
rect 818 12218 855 12297
rect 896 12284 1006 12297
rect 970 12228 1001 12229
rect 818 12198 827 12218
rect 847 12198 855 12218
rect 818 12188 855 12198
rect 914 12218 1001 12228
rect 914 12198 923 12218
rect 943 12198 1001 12218
rect 914 12189 1001 12198
rect 914 12188 951 12189
rect 479 12145 501 12163
rect 519 12145 544 12163
rect 479 12124 544 12145
rect 692 12143 757 12152
rect 692 12106 702 12143
rect 742 12135 757 12143
rect 970 12136 1001 12189
rect 1031 12218 1068 12297
rect 1183 12228 1214 12229
rect 1031 12198 1040 12218
rect 1060 12198 1068 12218
rect 1031 12188 1068 12198
rect 1127 12221 1214 12228
rect 1127 12218 1188 12221
rect 1127 12198 1136 12218
rect 1156 12201 1188 12218
rect 1209 12201 1214 12221
rect 1156 12198 1214 12201
rect 1127 12191 1214 12198
rect 1239 12218 1276 12360
rect 1542 12359 1579 12360
rect 2859 12300 2921 12771
rect 3021 12810 3047 12851
rect 3083 12810 3116 12851
rect 3021 12514 3116 12810
rect 3021 12470 3036 12514
rect 3096 12470 3116 12514
rect 3021 12450 3116 12470
rect 3733 12381 3776 13094
rect 4809 12984 5702 13024
rect 4809 12917 4842 12984
rect 4928 12917 5710 12984
rect 8875 12920 8945 13173
rect 9414 13170 9455 13172
rect 9686 13170 9790 13172
rect 10126 13170 11249 13203
rect 9007 13135 11249 13170
rect 13777 13146 14488 13148
rect 12100 13144 12172 13145
rect 13658 13144 14488 13146
rect 9007 13121 9035 13135
rect 9009 12990 9035 13121
rect 9414 13133 11249 13135
rect 9414 13132 9557 13133
rect 9815 13132 11249 13133
rect 4809 12849 5710 12917
rect 4818 12848 4924 12849
rect 5593 12755 5710 12849
rect 8867 12869 8947 12920
rect 8867 12843 8883 12869
rect 8923 12843 8947 12869
rect 8867 12824 8947 12843
rect 8867 12798 8886 12824
rect 8926 12798 8947 12824
rect 8867 12771 8947 12798
rect 3733 12361 4127 12381
rect 4147 12361 4150 12381
rect 3734 12356 4150 12361
rect 3734 12355 4075 12356
rect 3391 12324 3501 12338
rect 3391 12321 3434 12324
rect 3391 12316 3395 12321
rect 2854 12248 2929 12300
rect 3313 12294 3395 12316
rect 3424 12294 3434 12321
rect 3462 12297 3469 12324
rect 3498 12316 3501 12324
rect 3498 12297 3563 12316
rect 3462 12294 3563 12297
rect 3313 12292 3563 12294
rect 3223 12248 3269 12249
rect 1391 12228 1427 12229
rect 1239 12198 1248 12218
rect 1268 12198 1276 12218
rect 1127 12189 1183 12191
rect 1127 12188 1164 12189
rect 1239 12188 1276 12198
rect 1335 12218 1483 12228
rect 1583 12225 1679 12227
rect 1335 12198 1344 12218
rect 1364 12198 1454 12218
rect 1474 12198 1483 12218
rect 1335 12192 1483 12198
rect 1335 12189 1399 12192
rect 1335 12188 1372 12189
rect 1391 12162 1399 12189
rect 1420 12189 1483 12192
rect 1541 12218 1679 12225
rect 1541 12198 1550 12218
rect 1570 12198 1679 12218
rect 1541 12189 1679 12198
rect 2854 12213 3269 12248
rect 1420 12162 1427 12189
rect 1446 12188 1483 12189
rect 1542 12188 1579 12189
rect 1391 12137 1427 12162
rect 862 12135 903 12136
rect 742 12128 903 12135
rect 742 12108 872 12128
rect 892 12108 903 12128
rect 742 12106 903 12108
rect 692 12100 903 12106
rect 970 12132 1329 12136
rect 970 12127 1292 12132
rect 970 12103 1083 12127
rect 1107 12108 1292 12127
rect 1316 12108 1329 12132
rect 1107 12103 1329 12108
rect 970 12100 1329 12103
rect 1391 12100 1426 12137
rect 1494 12134 1594 12137
rect 1494 12130 1561 12134
rect 1494 12104 1506 12130
rect 1532 12108 1561 12130
rect 1587 12108 1594 12134
rect 1532 12104 1594 12108
rect 1494 12100 1594 12104
rect 692 12087 759 12100
rect 484 12064 540 12084
rect 484 12046 503 12064
rect 521 12046 540 12064
rect 484 11933 540 12046
rect 692 12066 706 12087
rect 742 12066 759 12087
rect 970 12079 1001 12100
rect 1391 12079 1427 12100
rect 813 12078 850 12079
rect 692 12059 759 12066
rect 812 12069 850 12078
rect 484 11795 539 11933
rect 692 11907 757 12059
rect 812 12049 821 12069
rect 841 12049 850 12069
rect 812 12041 850 12049
rect 916 12073 1001 12079
rect 1026 12078 1063 12079
rect 916 12053 924 12073
rect 944 12053 1001 12073
rect 916 12045 1001 12053
rect 1025 12069 1063 12078
rect 1025 12049 1034 12069
rect 1054 12049 1063 12069
rect 916 12044 952 12045
rect 1025 12041 1063 12049
rect 1129 12073 1214 12079
rect 1234 12078 1271 12079
rect 1129 12053 1137 12073
rect 1157 12072 1214 12073
rect 1157 12053 1186 12072
rect 1129 12052 1186 12053
rect 1207 12052 1214 12072
rect 1129 12045 1214 12052
rect 1233 12069 1271 12078
rect 1233 12049 1242 12069
rect 1262 12049 1271 12069
rect 1129 12044 1165 12045
rect 1233 12041 1271 12049
rect 1337 12073 1481 12079
rect 1337 12053 1345 12073
rect 1365 12053 1453 12073
rect 1473 12053 1481 12073
rect 1337 12045 1481 12053
rect 1337 12044 1373 12045
rect 1445 12044 1481 12045
rect 1547 12078 1584 12079
rect 1547 12077 1585 12078
rect 1547 12069 1611 12077
rect 1547 12049 1556 12069
rect 1576 12055 1611 12069
rect 1631 12055 1634 12075
rect 1576 12050 1634 12055
rect 1576 12049 1611 12050
rect 813 12012 850 12041
rect 814 12010 850 12012
rect 1026 12010 1063 12041
rect 814 11988 1063 12010
rect 895 11982 1006 11988
rect 895 11974 936 11982
rect 895 11954 903 11974
rect 922 11954 936 11974
rect 895 11952 936 11954
rect 964 11974 1006 11982
rect 964 11954 980 11974
rect 999 11954 1006 11974
rect 964 11952 1006 11954
rect 895 11939 1006 11952
rect 1234 11942 1271 12041
rect 1547 12037 1611 12049
rect 685 11897 806 11907
rect 685 11895 754 11897
rect 685 11854 698 11895
rect 735 11856 754 11895
rect 791 11856 806 11897
rect 735 11854 806 11856
rect 685 11836 806 11854
rect 477 11792 541 11795
rect 897 11792 1001 11798
rect 1232 11792 1273 11942
rect 1651 11934 1678 12189
rect 1740 12179 1820 12190
rect 1740 12153 1757 12179
rect 1797 12153 1820 12179
rect 1740 12126 1820 12153
rect 1740 12100 1761 12126
rect 1801 12100 1820 12126
rect 1740 12081 1820 12100
rect 1740 12055 1764 12081
rect 1804 12055 1820 12081
rect 1740 12004 1820 12055
rect 477 11789 1273 11792
rect 1652 11803 1678 11934
rect 1652 11789 1680 11803
rect 477 11754 1680 11789
rect 1742 11796 1812 12004
rect 2854 11929 2929 12213
rect 3223 12130 3269 12213
rect 3313 12213 3350 12292
rect 3391 12279 3501 12292
rect 3465 12223 3496 12224
rect 3313 12193 3322 12213
rect 3342 12193 3350 12213
rect 3313 12183 3350 12193
rect 3409 12213 3496 12223
rect 3409 12193 3418 12213
rect 3438 12193 3496 12213
rect 3409 12184 3496 12193
rect 3409 12183 3446 12184
rect 3465 12131 3496 12184
rect 3526 12213 3563 12292
rect 3678 12223 3709 12224
rect 3526 12193 3535 12213
rect 3555 12193 3563 12213
rect 3526 12183 3563 12193
rect 3622 12216 3709 12223
rect 3622 12213 3683 12216
rect 3622 12193 3631 12213
rect 3651 12196 3683 12213
rect 3704 12196 3709 12216
rect 3651 12193 3709 12196
rect 3622 12186 3709 12193
rect 3734 12213 3771 12355
rect 4037 12354 4074 12355
rect 3886 12223 3922 12224
rect 3734 12193 3743 12213
rect 3763 12193 3771 12213
rect 3622 12184 3678 12186
rect 3622 12183 3659 12184
rect 3734 12183 3771 12193
rect 3830 12213 3978 12223
rect 4078 12220 4174 12222
rect 3830 12193 3839 12213
rect 3859 12193 3949 12213
rect 3969 12193 3978 12213
rect 3830 12187 3978 12193
rect 3830 12184 3894 12187
rect 3830 12183 3867 12184
rect 3886 12157 3894 12184
rect 3915 12184 3978 12187
rect 4036 12213 4174 12220
rect 4036 12193 4045 12213
rect 4065 12193 4174 12213
rect 4036 12184 4174 12193
rect 3915 12157 3922 12184
rect 3941 12183 3978 12184
rect 4037 12183 4074 12184
rect 3886 12132 3922 12157
rect 3357 12130 3398 12131
rect 3223 12123 3398 12130
rect 3021 12097 3107 12116
rect 3021 12056 3036 12097
rect 3090 12056 3107 12097
rect 3223 12103 3367 12123
rect 3387 12103 3398 12123
rect 3223 12095 3398 12103
rect 3465 12127 3824 12131
rect 3465 12122 3787 12127
rect 3465 12098 3578 12122
rect 3602 12103 3787 12122
rect 3811 12103 3824 12127
rect 3602 12098 3824 12103
rect 3465 12095 3824 12098
rect 3886 12095 3921 12132
rect 3989 12129 4089 12132
rect 3989 12125 4056 12129
rect 3989 12099 4001 12125
rect 4027 12103 4056 12125
rect 4082 12103 4089 12129
rect 4027 12099 4089 12103
rect 3989 12095 4089 12099
rect 3223 12091 3269 12095
rect 3465 12074 3496 12095
rect 3886 12074 3922 12095
rect 3308 12073 3345 12074
rect 3021 12020 3107 12056
rect 3307 12064 3345 12073
rect 3307 12044 3316 12064
rect 3336 12044 3345 12064
rect 3307 12036 3345 12044
rect 3411 12068 3496 12074
rect 3521 12073 3558 12074
rect 3411 12048 3419 12068
rect 3439 12048 3496 12068
rect 3411 12040 3496 12048
rect 3520 12064 3558 12073
rect 3520 12044 3529 12064
rect 3549 12044 3558 12064
rect 3411 12039 3447 12040
rect 3520 12036 3558 12044
rect 3624 12068 3709 12074
rect 3729 12073 3766 12074
rect 3624 12048 3632 12068
rect 3652 12067 3709 12068
rect 3652 12048 3681 12067
rect 3624 12047 3681 12048
rect 3702 12047 3709 12067
rect 3624 12040 3709 12047
rect 3728 12064 3766 12073
rect 3728 12044 3737 12064
rect 3757 12044 3766 12064
rect 3624 12039 3660 12040
rect 3728 12036 3766 12044
rect 3832 12068 3976 12074
rect 3832 12048 3840 12068
rect 3860 12048 3948 12068
rect 3968 12048 3976 12068
rect 3832 12040 3976 12048
rect 3832 12039 3868 12040
rect 477 11693 541 11754
rect 897 11752 1001 11754
rect 1232 11752 1273 11754
rect 1742 11751 1763 11796
rect 1743 11730 1763 11751
rect 1793 11751 1812 11796
rect 2849 11887 2929 11929
rect 1793 11730 1810 11751
rect 1743 11711 1810 11730
rect 1392 11703 1464 11704
rect 1391 11695 1490 11703
rect 479 11622 538 11693
rect 1391 11692 1443 11695
rect 1391 11657 1399 11692
rect 1424 11657 1443 11692
rect 1468 11684 1490 11695
rect 1468 11683 2335 11684
rect 1468 11657 2336 11683
rect 1391 11647 2336 11657
rect 1391 11645 1490 11647
rect 479 11604 501 11622
rect 519 11604 538 11622
rect 479 11582 538 11604
rect 746 11618 1278 11623
rect 746 11598 1632 11618
rect 1652 11598 1655 11618
rect 2291 11614 2336 11647
rect 746 11594 1655 11598
rect 746 11547 789 11594
rect 1239 11593 1655 11594
rect 2287 11594 2680 11614
rect 2700 11594 2703 11614
rect 1239 11592 1580 11593
rect 896 11561 1006 11575
rect 896 11558 939 11561
rect 896 11553 900 11558
rect 734 11546 789 11547
rect 478 11523 789 11546
rect 478 11505 503 11523
rect 521 11511 789 11523
rect 818 11531 900 11553
rect 929 11531 939 11558
rect 967 11534 974 11561
rect 1003 11553 1006 11561
rect 1003 11534 1068 11553
rect 967 11531 1068 11534
rect 818 11529 1068 11531
rect 521 11505 543 11511
rect 478 11366 543 11505
rect 818 11450 855 11529
rect 896 11516 1006 11529
rect 970 11460 1001 11461
rect 818 11430 827 11450
rect 847 11430 855 11450
rect 478 11348 501 11366
rect 519 11348 543 11366
rect 478 11331 543 11348
rect 698 11412 766 11425
rect 818 11420 855 11430
rect 914 11450 1001 11460
rect 914 11430 923 11450
rect 943 11430 1001 11450
rect 914 11421 1001 11430
rect 914 11420 951 11421
rect 698 11370 705 11412
rect 754 11370 766 11412
rect 698 11367 766 11370
rect 970 11368 1001 11421
rect 1031 11450 1068 11529
rect 1183 11460 1214 11461
rect 1031 11430 1040 11450
rect 1060 11430 1068 11450
rect 1031 11420 1068 11430
rect 1127 11453 1214 11460
rect 1127 11450 1188 11453
rect 1127 11430 1136 11450
rect 1156 11433 1188 11450
rect 1209 11433 1214 11453
rect 1156 11430 1214 11433
rect 1127 11423 1214 11430
rect 1239 11450 1276 11592
rect 1542 11591 1579 11592
rect 2287 11589 2703 11594
rect 2287 11588 2628 11589
rect 1944 11557 2054 11571
rect 1944 11554 1987 11557
rect 1944 11549 1948 11554
rect 1866 11527 1948 11549
rect 1977 11527 1987 11554
rect 2015 11530 2022 11557
rect 2051 11549 2054 11557
rect 2051 11530 2116 11549
rect 2015 11527 2116 11530
rect 1866 11525 2116 11527
rect 1391 11460 1427 11461
rect 1239 11430 1248 11450
rect 1268 11430 1276 11450
rect 1127 11421 1183 11423
rect 1127 11420 1164 11421
rect 1239 11420 1276 11430
rect 1335 11450 1483 11460
rect 1583 11457 1679 11459
rect 1335 11430 1344 11450
rect 1364 11430 1454 11450
rect 1474 11430 1483 11450
rect 1335 11424 1483 11430
rect 1335 11421 1399 11424
rect 1335 11420 1372 11421
rect 1391 11394 1399 11421
rect 1420 11421 1483 11424
rect 1541 11450 1679 11457
rect 1541 11430 1550 11450
rect 1570 11430 1679 11450
rect 1541 11421 1679 11430
rect 1866 11446 1903 11525
rect 1944 11512 2054 11525
rect 2018 11456 2049 11457
rect 1866 11426 1875 11446
rect 1895 11426 1903 11446
rect 1420 11394 1427 11421
rect 1446 11420 1483 11421
rect 1542 11420 1579 11421
rect 1391 11369 1427 11394
rect 862 11367 903 11368
rect 698 11360 903 11367
rect 698 11349 872 11360
rect 698 11316 706 11349
rect 699 11307 706 11316
rect 755 11340 872 11349
rect 892 11340 903 11360
rect 755 11332 903 11340
rect 970 11364 1329 11368
rect 970 11359 1292 11364
rect 970 11335 1083 11359
rect 1107 11340 1292 11359
rect 1316 11340 1329 11364
rect 1107 11335 1329 11340
rect 970 11332 1329 11335
rect 1391 11332 1426 11369
rect 1494 11366 1594 11369
rect 1494 11362 1561 11366
rect 1494 11336 1506 11362
rect 1532 11340 1561 11362
rect 1587 11340 1594 11366
rect 1532 11336 1594 11340
rect 1494 11332 1594 11336
rect 755 11316 766 11332
rect 755 11307 763 11316
rect 970 11311 1001 11332
rect 1391 11311 1427 11332
rect 813 11310 850 11311
rect 478 11267 543 11286
rect 478 11249 503 11267
rect 521 11249 543 11267
rect 478 11048 543 11249
rect 699 11123 763 11307
rect 812 11301 850 11310
rect 812 11281 821 11301
rect 841 11281 850 11301
rect 812 11273 850 11281
rect 916 11305 1001 11311
rect 1026 11310 1063 11311
rect 916 11285 924 11305
rect 944 11285 1001 11305
rect 916 11277 1001 11285
rect 1025 11301 1063 11310
rect 1025 11281 1034 11301
rect 1054 11281 1063 11301
rect 916 11276 952 11277
rect 1025 11273 1063 11281
rect 1129 11305 1214 11311
rect 1234 11310 1271 11311
rect 1129 11285 1137 11305
rect 1157 11304 1214 11305
rect 1157 11285 1186 11304
rect 1129 11284 1186 11285
rect 1207 11284 1214 11304
rect 1129 11277 1214 11284
rect 1233 11301 1271 11310
rect 1233 11281 1242 11301
rect 1262 11281 1271 11301
rect 1129 11276 1165 11277
rect 1233 11273 1271 11281
rect 1337 11305 1481 11311
rect 1337 11285 1345 11305
rect 1365 11285 1453 11305
rect 1473 11285 1481 11305
rect 1337 11277 1481 11285
rect 1337 11276 1373 11277
rect 1445 11276 1481 11277
rect 1547 11310 1584 11311
rect 1547 11309 1585 11310
rect 1547 11301 1611 11309
rect 1547 11281 1556 11301
rect 1576 11287 1611 11301
rect 1631 11287 1634 11307
rect 1576 11282 1634 11287
rect 1576 11281 1611 11282
rect 813 11244 850 11273
rect 814 11242 850 11244
rect 1026 11242 1063 11273
rect 814 11220 1063 11242
rect 895 11214 1006 11220
rect 895 11206 936 11214
rect 895 11186 903 11206
rect 922 11186 936 11206
rect 895 11184 936 11186
rect 964 11206 1006 11214
rect 964 11186 980 11206
rect 999 11186 1006 11206
rect 964 11184 1006 11186
rect 895 11169 1006 11184
rect 699 11113 767 11123
rect 699 11080 716 11113
rect 756 11080 767 11113
rect 699 11068 767 11080
rect 699 11066 763 11068
rect 1234 11049 1271 11273
rect 1547 11269 1611 11281
rect 1651 11051 1678 11421
rect 1866 11416 1903 11426
rect 1962 11446 2049 11456
rect 1962 11426 1971 11446
rect 1991 11426 2049 11446
rect 1962 11417 2049 11426
rect 1962 11416 1999 11417
rect 1742 11403 1812 11408
rect 1737 11397 1812 11403
rect 1737 11364 1745 11397
rect 1798 11364 1812 11397
rect 2018 11364 2049 11417
rect 2079 11446 2116 11525
rect 2231 11456 2262 11457
rect 2079 11426 2088 11446
rect 2108 11426 2116 11446
rect 2079 11416 2116 11426
rect 2175 11449 2262 11456
rect 2175 11446 2236 11449
rect 2175 11426 2184 11446
rect 2204 11429 2236 11446
rect 2257 11429 2262 11449
rect 2204 11426 2262 11429
rect 2175 11419 2262 11426
rect 2287 11446 2324 11588
rect 2590 11587 2627 11588
rect 2439 11456 2475 11457
rect 2287 11426 2296 11446
rect 2316 11426 2324 11446
rect 2175 11417 2231 11419
rect 2175 11416 2212 11417
rect 2287 11416 2324 11426
rect 2383 11446 2531 11456
rect 2631 11453 2727 11455
rect 2383 11426 2392 11446
rect 2412 11426 2502 11446
rect 2522 11426 2531 11446
rect 2383 11420 2531 11426
rect 2383 11417 2447 11420
rect 2383 11416 2420 11417
rect 2439 11390 2447 11417
rect 2468 11417 2531 11420
rect 2589 11446 2727 11453
rect 2589 11426 2598 11446
rect 2618 11426 2727 11446
rect 2589 11417 2727 11426
rect 2468 11390 2475 11417
rect 2494 11416 2531 11417
rect 2590 11416 2627 11417
rect 2439 11365 2475 11390
rect 1737 11363 1820 11364
rect 1910 11363 1951 11364
rect 1737 11356 1951 11363
rect 1737 11339 1920 11356
rect 1737 11306 1750 11339
rect 1803 11336 1920 11339
rect 1940 11336 1951 11356
rect 1803 11328 1951 11336
rect 2018 11360 2377 11364
rect 2018 11355 2340 11360
rect 2018 11331 2131 11355
rect 2155 11336 2340 11355
rect 2364 11336 2377 11360
rect 2155 11331 2377 11336
rect 2018 11328 2377 11331
rect 2439 11328 2474 11365
rect 2542 11362 2642 11365
rect 2542 11358 2609 11362
rect 2542 11332 2554 11358
rect 2580 11336 2609 11358
rect 2635 11336 2642 11362
rect 2580 11332 2642 11336
rect 2542 11328 2642 11332
rect 1803 11306 1820 11328
rect 2018 11307 2049 11328
rect 2439 11307 2475 11328
rect 1861 11306 1898 11307
rect 1737 11292 1820 11306
rect 1510 11049 1678 11051
rect 1234 11048 1678 11049
rect 478 11018 1678 11048
rect 1748 11082 1820 11292
rect 1860 11297 1898 11306
rect 1860 11277 1869 11297
rect 1889 11277 1898 11297
rect 1860 11269 1898 11277
rect 1964 11301 2049 11307
rect 2074 11306 2111 11307
rect 1964 11281 1972 11301
rect 1992 11281 2049 11301
rect 1964 11273 2049 11281
rect 2073 11297 2111 11306
rect 2073 11277 2082 11297
rect 2102 11277 2111 11297
rect 1964 11272 2000 11273
rect 2073 11269 2111 11277
rect 2177 11301 2262 11307
rect 2282 11306 2319 11307
rect 2177 11281 2185 11301
rect 2205 11300 2262 11301
rect 2205 11281 2234 11300
rect 2177 11280 2234 11281
rect 2255 11280 2262 11300
rect 2177 11273 2262 11280
rect 2281 11297 2319 11306
rect 2281 11277 2290 11297
rect 2310 11277 2319 11297
rect 2177 11272 2213 11273
rect 2281 11269 2319 11277
rect 2385 11301 2529 11307
rect 2385 11281 2393 11301
rect 2413 11281 2501 11301
rect 2521 11281 2529 11301
rect 2385 11273 2529 11281
rect 2385 11272 2421 11273
rect 2493 11272 2529 11273
rect 2595 11306 2632 11307
rect 2595 11305 2633 11306
rect 2595 11297 2659 11305
rect 2595 11277 2604 11297
rect 2624 11283 2659 11297
rect 2679 11283 2682 11303
rect 2624 11278 2682 11283
rect 2624 11277 2659 11278
rect 1861 11240 1898 11269
rect 1862 11238 1898 11240
rect 2074 11238 2111 11269
rect 1862 11216 2111 11238
rect 1943 11210 2054 11216
rect 1943 11202 1984 11210
rect 1943 11182 1951 11202
rect 1970 11182 1984 11202
rect 1943 11180 1984 11182
rect 2012 11202 2054 11210
rect 2012 11182 2028 11202
rect 2047 11182 2054 11202
rect 2012 11180 2054 11182
rect 1943 11165 2054 11180
rect 1748 11043 1767 11082
rect 1812 11043 1820 11082
rect 1748 11026 1820 11043
rect 2282 11070 2319 11269
rect 2595 11265 2659 11277
rect 2282 11064 2323 11070
rect 2699 11066 2726 11417
rect 2849 11287 2928 11887
rect 3025 11435 3104 12020
rect 3308 12007 3345 12036
rect 3309 12005 3345 12007
rect 3521 12005 3558 12036
rect 3309 11983 3558 12005
rect 3390 11977 3501 11983
rect 3390 11969 3431 11977
rect 3390 11949 3398 11969
rect 3417 11949 3431 11969
rect 3390 11947 3431 11949
rect 3459 11969 3501 11977
rect 3459 11949 3475 11969
rect 3494 11949 3501 11969
rect 3459 11947 3501 11949
rect 3390 11932 3501 11947
rect 3729 11921 3766 12036
rect 3722 11809 3769 11921
rect 3890 11881 3920 12040
rect 3940 12039 3976 12040
rect 4042 12073 4079 12074
rect 4042 12072 4080 12073
rect 4042 12064 4106 12072
rect 4042 12044 4051 12064
rect 4071 12050 4106 12064
rect 4126 12050 4129 12070
rect 4071 12045 4129 12050
rect 4071 12044 4106 12045
rect 4042 12032 4106 12044
rect 3890 11877 3976 11881
rect 3890 11859 3905 11877
rect 3957 11859 3976 11877
rect 3890 11850 3976 11859
rect 4146 11811 4173 12184
rect 4005 11809 4173 11811
rect 3722 11783 4173 11809
rect 3722 11705 3769 11783
rect 4005 11782 4173 11783
rect 3667 11704 3769 11705
rect 3666 11696 3769 11704
rect 3666 11693 3718 11696
rect 3666 11658 3674 11693
rect 3699 11658 3718 11693
rect 3743 11658 3769 11696
rect 3666 11652 3769 11658
rect 3929 11697 3965 11701
rect 3929 11674 3937 11697
rect 3961 11674 3965 11697
rect 3929 11653 3965 11674
rect 3666 11648 3765 11652
rect 3929 11630 3937 11653
rect 3961 11630 3965 11653
rect 2558 11064 2726 11066
rect 2282 11038 2726 11064
rect 478 10971 543 11018
rect 478 10953 501 10971
rect 519 10953 543 10971
rect 1391 10998 1426 11000
rect 1391 10996 1495 10998
rect 2284 10996 2323 11038
rect 2558 11037 2726 11038
rect 1391 10989 2325 10996
rect 1391 10988 1442 10989
rect 1391 10968 1394 10988
rect 1419 10969 1442 10988
rect 1474 10969 2325 10989
rect 1419 10968 2325 10969
rect 1391 10961 2325 10968
rect 1664 10960 2325 10961
rect 478 10932 543 10953
rect 755 10943 795 10946
rect 755 10939 1658 10943
rect 755 10919 1632 10939
rect 1652 10919 1658 10939
rect 755 10916 1658 10919
rect 479 10872 544 10892
rect 479 10854 503 10872
rect 521 10854 544 10872
rect 479 10827 544 10854
rect 755 10827 795 10916
rect 1239 10914 1655 10916
rect 1239 10913 1580 10914
rect 896 10882 1006 10896
rect 896 10879 939 10882
rect 896 10874 900 10879
rect 478 10792 795 10827
rect 818 10852 900 10874
rect 929 10852 939 10879
rect 967 10855 974 10882
rect 1003 10874 1006 10882
rect 1003 10855 1068 10874
rect 967 10852 1068 10855
rect 818 10850 1068 10852
rect 479 10716 544 10792
rect 818 10771 855 10850
rect 896 10837 1006 10850
rect 970 10781 1001 10782
rect 818 10751 827 10771
rect 847 10751 855 10771
rect 818 10741 855 10751
rect 914 10771 1001 10781
rect 914 10751 923 10771
rect 943 10751 1001 10771
rect 914 10742 1001 10751
rect 914 10741 951 10742
rect 479 10698 501 10716
rect 519 10698 544 10716
rect 479 10677 544 10698
rect 692 10696 757 10705
rect 692 10659 702 10696
rect 742 10688 757 10696
rect 970 10689 1001 10742
rect 1031 10771 1068 10850
rect 1183 10781 1214 10782
rect 1031 10751 1040 10771
rect 1060 10751 1068 10771
rect 1031 10741 1068 10751
rect 1127 10774 1214 10781
rect 1127 10771 1188 10774
rect 1127 10751 1136 10771
rect 1156 10754 1188 10771
rect 1209 10754 1214 10774
rect 1156 10751 1214 10754
rect 1127 10744 1214 10751
rect 1239 10771 1276 10913
rect 1542 10912 1579 10913
rect 1391 10781 1427 10782
rect 1239 10751 1248 10771
rect 1268 10751 1276 10771
rect 1127 10742 1183 10744
rect 1127 10741 1164 10742
rect 1239 10741 1276 10751
rect 1335 10771 1483 10781
rect 1583 10778 1679 10780
rect 1335 10751 1344 10771
rect 1364 10751 1454 10771
rect 1474 10751 1483 10771
rect 1335 10745 1483 10751
rect 1335 10742 1399 10745
rect 1335 10741 1372 10742
rect 1391 10715 1399 10742
rect 1420 10742 1483 10745
rect 1541 10771 1679 10778
rect 1541 10751 1550 10771
rect 1570 10751 1679 10771
rect 1541 10742 1679 10751
rect 1420 10715 1427 10742
rect 1446 10741 1483 10742
rect 1542 10741 1579 10742
rect 1391 10690 1427 10715
rect 862 10688 903 10689
rect 742 10681 903 10688
rect 742 10661 872 10681
rect 892 10661 903 10681
rect 742 10659 903 10661
rect 692 10653 903 10659
rect 970 10685 1329 10689
rect 970 10680 1292 10685
rect 970 10656 1083 10680
rect 1107 10661 1292 10680
rect 1316 10661 1329 10685
rect 1107 10656 1329 10661
rect 970 10653 1329 10656
rect 1391 10653 1426 10690
rect 1494 10687 1594 10690
rect 1494 10683 1561 10687
rect 1494 10657 1506 10683
rect 1532 10661 1561 10683
rect 1587 10661 1594 10687
rect 1532 10657 1594 10661
rect 1494 10653 1594 10657
rect 692 10640 759 10653
rect 484 10617 540 10637
rect 484 10599 503 10617
rect 521 10599 540 10617
rect 484 10486 540 10599
rect 692 10619 706 10640
rect 742 10619 759 10640
rect 970 10632 1001 10653
rect 1391 10632 1427 10653
rect 813 10631 850 10632
rect 692 10612 759 10619
rect 812 10622 850 10631
rect 484 10357 539 10486
rect 692 10460 757 10612
rect 812 10602 821 10622
rect 841 10602 850 10622
rect 812 10594 850 10602
rect 916 10626 1001 10632
rect 1026 10631 1063 10632
rect 916 10606 924 10626
rect 944 10606 1001 10626
rect 916 10598 1001 10606
rect 1025 10622 1063 10631
rect 1025 10602 1034 10622
rect 1054 10602 1063 10622
rect 916 10597 952 10598
rect 1025 10594 1063 10602
rect 1129 10626 1214 10632
rect 1234 10631 1271 10632
rect 1129 10606 1137 10626
rect 1157 10625 1214 10626
rect 1157 10606 1186 10625
rect 1129 10605 1186 10606
rect 1207 10605 1214 10625
rect 1129 10598 1214 10605
rect 1233 10622 1271 10631
rect 1233 10602 1242 10622
rect 1262 10602 1271 10622
rect 1129 10597 1165 10598
rect 1233 10594 1271 10602
rect 1337 10626 1481 10632
rect 1337 10606 1345 10626
rect 1365 10606 1453 10626
rect 1473 10606 1481 10626
rect 1337 10598 1481 10606
rect 1337 10597 1373 10598
rect 1445 10597 1481 10598
rect 1547 10631 1584 10632
rect 1547 10630 1585 10631
rect 1547 10622 1611 10630
rect 1547 10602 1556 10622
rect 1576 10608 1611 10622
rect 1631 10608 1634 10628
rect 1576 10603 1634 10608
rect 1576 10602 1611 10603
rect 813 10565 850 10594
rect 814 10563 850 10565
rect 1026 10563 1063 10594
rect 814 10541 1063 10563
rect 895 10535 1006 10541
rect 895 10527 936 10535
rect 895 10507 903 10527
rect 922 10507 936 10527
rect 895 10505 936 10507
rect 964 10527 1006 10535
rect 964 10507 980 10527
rect 999 10507 1006 10527
rect 964 10505 1006 10507
rect 895 10490 1006 10505
rect 1234 10495 1271 10594
rect 1547 10590 1611 10602
rect 897 10481 1001 10490
rect 685 10450 806 10460
rect 685 10448 754 10450
rect 685 10407 698 10448
rect 735 10409 754 10448
rect 791 10409 806 10450
rect 735 10407 806 10409
rect 685 10389 806 10407
rect 478 10345 539 10357
rect 1232 10345 1273 10495
rect 1651 10487 1678 10742
rect 1740 10732 1820 10743
rect 1740 10706 1757 10732
rect 1797 10706 1820 10732
rect 1740 10679 1820 10706
rect 1740 10653 1761 10679
rect 1801 10653 1820 10679
rect 1740 10634 1820 10653
rect 1740 10608 1764 10634
rect 1804 10608 1820 10634
rect 1740 10557 1820 10608
rect 478 10342 1273 10345
rect 1652 10356 1678 10487
rect 1742 10401 1812 10557
rect 1741 10385 1817 10401
rect 1652 10342 1680 10356
rect 478 10307 1680 10342
rect 1741 10348 1756 10385
rect 1800 10348 1817 10385
rect 1741 10328 1817 10348
rect 2855 10378 2925 11287
rect 3024 10722 3105 11435
rect 3929 11321 3965 11630
rect 3853 11292 3966 11321
rect 3853 10936 3884 11292
rect 3923 11037 4914 11062
rect 3923 11032 3983 11037
rect 3923 11011 3942 11032
rect 3962 11016 3983 11032
rect 4003 11016 4914 11037
rect 3962 11011 4914 11016
rect 3923 11003 4914 11011
rect 3928 10980 4034 11003
rect 3928 10977 4033 10980
rect 3777 10916 4170 10936
rect 4190 10916 4193 10936
rect 3777 10911 4193 10916
rect 3777 10910 4118 10911
rect 3434 10879 3544 10893
rect 3434 10876 3477 10879
rect 3434 10871 3438 10876
rect 3356 10849 3438 10871
rect 3467 10849 3477 10876
rect 3505 10852 3512 10879
rect 3541 10871 3544 10879
rect 3541 10852 3606 10871
rect 3505 10849 3606 10852
rect 3356 10847 3606 10849
rect 3356 10768 3393 10847
rect 3434 10834 3544 10847
rect 3508 10778 3539 10779
rect 3356 10748 3365 10768
rect 3385 10748 3393 10768
rect 3356 10738 3393 10748
rect 3452 10768 3539 10778
rect 3452 10748 3461 10768
rect 3481 10748 3539 10768
rect 3452 10739 3539 10748
rect 3452 10738 3489 10739
rect 3022 10686 3114 10722
rect 3508 10686 3539 10739
rect 3569 10768 3606 10847
rect 3721 10778 3752 10779
rect 3569 10748 3578 10768
rect 3598 10748 3606 10768
rect 3569 10738 3606 10748
rect 3665 10771 3752 10778
rect 3665 10768 3726 10771
rect 3665 10748 3674 10768
rect 3694 10751 3726 10768
rect 3747 10751 3752 10771
rect 3694 10748 3752 10751
rect 3665 10741 3752 10748
rect 3777 10768 3814 10910
rect 4080 10909 4117 10910
rect 3929 10778 3965 10779
rect 3777 10748 3786 10768
rect 3806 10748 3814 10768
rect 3665 10739 3721 10741
rect 3665 10738 3702 10739
rect 3777 10738 3814 10748
rect 3873 10768 4021 10778
rect 4121 10775 4217 10777
rect 3873 10748 3882 10768
rect 3902 10748 3992 10768
rect 4012 10748 4021 10768
rect 3873 10742 4021 10748
rect 3873 10739 3937 10742
rect 3873 10738 3910 10739
rect 3929 10712 3937 10739
rect 3958 10739 4021 10742
rect 4079 10768 4217 10775
rect 4079 10748 4088 10768
rect 4108 10748 4217 10768
rect 4079 10739 4217 10748
rect 3958 10712 3965 10739
rect 3984 10738 4021 10739
rect 4080 10738 4117 10739
rect 3929 10687 3965 10712
rect 3022 10685 3358 10686
rect 3400 10685 3441 10686
rect 3022 10678 3441 10685
rect 3022 10658 3410 10678
rect 3430 10658 3441 10678
rect 3022 10650 3441 10658
rect 3508 10682 3867 10686
rect 3508 10677 3830 10682
rect 3508 10653 3621 10677
rect 3645 10658 3830 10677
rect 3854 10658 3867 10682
rect 3645 10653 3867 10658
rect 3508 10650 3867 10653
rect 3929 10650 3964 10687
rect 4032 10684 4132 10687
rect 4032 10680 4099 10684
rect 4032 10654 4044 10680
rect 4070 10658 4099 10680
rect 4125 10658 4132 10684
rect 4070 10654 4132 10658
rect 4032 10650 4132 10654
rect 3022 10646 3358 10650
rect 2855 10328 2927 10378
rect 478 10232 539 10307
rect 897 10305 1001 10307
rect 1232 10305 1273 10307
rect 1741 10262 1751 10328
rect 1805 10262 1817 10328
rect 1741 10238 1817 10262
rect 480 10102 539 10232
rect 1393 10183 1465 10184
rect 1392 10175 1491 10183
rect 1392 10172 1444 10175
rect 1392 10137 1400 10172
rect 1425 10137 1444 10172
rect 1469 10164 1491 10175
rect 1469 10163 2336 10164
rect 1469 10137 2337 10163
rect 1392 10127 2337 10137
rect 1392 10125 1491 10127
rect 480 10084 502 10102
rect 520 10084 539 10102
rect 480 10062 539 10084
rect 747 10098 1279 10103
rect 747 10078 1633 10098
rect 1653 10078 1656 10098
rect 2292 10094 2337 10127
rect 747 10074 1656 10078
rect 747 10027 790 10074
rect 1240 10073 1656 10074
rect 2288 10074 2681 10094
rect 2701 10074 2704 10094
rect 1240 10072 1581 10073
rect 897 10041 1007 10055
rect 897 10038 940 10041
rect 897 10033 901 10038
rect 735 10026 790 10027
rect 479 10003 790 10026
rect 479 9985 504 10003
rect 522 9991 790 10003
rect 819 10011 901 10033
rect 930 10011 940 10038
rect 968 10014 975 10041
rect 1004 10033 1007 10041
rect 1004 10014 1069 10033
rect 968 10011 1069 10014
rect 819 10009 1069 10011
rect 522 9985 544 9991
rect 479 9846 544 9985
rect 819 9930 856 10009
rect 897 9996 1007 10009
rect 971 9940 1002 9941
rect 819 9910 828 9930
rect 848 9910 856 9930
rect 479 9828 502 9846
rect 520 9828 544 9846
rect 479 9811 544 9828
rect 699 9892 767 9905
rect 819 9900 856 9910
rect 915 9930 1002 9940
rect 915 9910 924 9930
rect 944 9910 1002 9930
rect 915 9901 1002 9910
rect 915 9900 952 9901
rect 699 9850 706 9892
rect 755 9850 767 9892
rect 699 9847 767 9850
rect 971 9848 1002 9901
rect 1032 9930 1069 10009
rect 1184 9940 1215 9941
rect 1032 9910 1041 9930
rect 1061 9910 1069 9930
rect 1032 9900 1069 9910
rect 1128 9933 1215 9940
rect 1128 9930 1189 9933
rect 1128 9910 1137 9930
rect 1157 9913 1189 9930
rect 1210 9913 1215 9933
rect 1157 9910 1215 9913
rect 1128 9903 1215 9910
rect 1240 9930 1277 10072
rect 1543 10071 1580 10072
rect 2288 10069 2704 10074
rect 2288 10068 2629 10069
rect 1945 10037 2055 10051
rect 1945 10034 1988 10037
rect 1945 10029 1949 10034
rect 1867 10007 1949 10029
rect 1978 10007 1988 10034
rect 2016 10010 2023 10037
rect 2052 10029 2055 10037
rect 2052 10010 2117 10029
rect 2016 10007 2117 10010
rect 1867 10005 2117 10007
rect 1392 9940 1428 9941
rect 1240 9910 1249 9930
rect 1269 9910 1277 9930
rect 1128 9901 1184 9903
rect 1128 9900 1165 9901
rect 1240 9900 1277 9910
rect 1336 9930 1484 9940
rect 1584 9937 1680 9939
rect 1336 9910 1345 9930
rect 1365 9910 1455 9930
rect 1475 9910 1484 9930
rect 1336 9904 1484 9910
rect 1336 9901 1400 9904
rect 1336 9900 1373 9901
rect 1392 9874 1400 9901
rect 1421 9901 1484 9904
rect 1542 9930 1680 9937
rect 1542 9910 1551 9930
rect 1571 9910 1680 9930
rect 1542 9901 1680 9910
rect 1867 9926 1904 10005
rect 1945 9992 2055 10005
rect 2019 9936 2050 9937
rect 1867 9906 1876 9926
rect 1896 9906 1904 9926
rect 1421 9874 1428 9901
rect 1447 9900 1484 9901
rect 1543 9900 1580 9901
rect 1392 9849 1428 9874
rect 863 9847 904 9848
rect 699 9840 904 9847
rect 699 9829 873 9840
rect 699 9796 707 9829
rect 700 9787 707 9796
rect 756 9820 873 9829
rect 893 9820 904 9840
rect 756 9812 904 9820
rect 971 9844 1330 9848
rect 971 9839 1293 9844
rect 971 9815 1084 9839
rect 1108 9820 1293 9839
rect 1317 9820 1330 9844
rect 1108 9815 1330 9820
rect 971 9812 1330 9815
rect 1392 9812 1427 9849
rect 1495 9846 1595 9849
rect 1495 9842 1562 9846
rect 1495 9816 1507 9842
rect 1533 9820 1562 9842
rect 1588 9820 1595 9846
rect 1533 9816 1595 9820
rect 1495 9812 1595 9816
rect 756 9796 767 9812
rect 756 9787 764 9796
rect 971 9791 1002 9812
rect 1392 9791 1428 9812
rect 814 9790 851 9791
rect 479 9747 544 9766
rect 479 9729 504 9747
rect 522 9729 544 9747
rect 479 9528 544 9729
rect 700 9603 764 9787
rect 813 9781 851 9790
rect 813 9761 822 9781
rect 842 9761 851 9781
rect 813 9753 851 9761
rect 917 9785 1002 9791
rect 1027 9790 1064 9791
rect 917 9765 925 9785
rect 945 9765 1002 9785
rect 917 9757 1002 9765
rect 1026 9781 1064 9790
rect 1026 9761 1035 9781
rect 1055 9761 1064 9781
rect 917 9756 953 9757
rect 1026 9753 1064 9761
rect 1130 9785 1215 9791
rect 1235 9790 1272 9791
rect 1130 9765 1138 9785
rect 1158 9784 1215 9785
rect 1158 9765 1187 9784
rect 1130 9764 1187 9765
rect 1208 9764 1215 9784
rect 1130 9757 1215 9764
rect 1234 9781 1272 9790
rect 1234 9761 1243 9781
rect 1263 9761 1272 9781
rect 1130 9756 1166 9757
rect 1234 9753 1272 9761
rect 1338 9785 1482 9791
rect 1338 9765 1346 9785
rect 1366 9765 1454 9785
rect 1474 9765 1482 9785
rect 1338 9757 1482 9765
rect 1338 9756 1374 9757
rect 1446 9756 1482 9757
rect 1548 9790 1585 9791
rect 1548 9789 1586 9790
rect 1548 9781 1612 9789
rect 1548 9761 1557 9781
rect 1577 9767 1612 9781
rect 1632 9767 1635 9787
rect 1577 9762 1635 9767
rect 1577 9761 1612 9762
rect 814 9724 851 9753
rect 815 9722 851 9724
rect 1027 9722 1064 9753
rect 815 9700 1064 9722
rect 896 9694 1007 9700
rect 896 9686 937 9694
rect 896 9666 904 9686
rect 923 9666 937 9686
rect 896 9664 937 9666
rect 965 9686 1007 9694
rect 965 9666 981 9686
rect 1000 9666 1007 9686
rect 965 9664 1007 9666
rect 896 9649 1007 9664
rect 700 9593 768 9603
rect 700 9560 717 9593
rect 757 9560 768 9593
rect 700 9548 768 9560
rect 700 9546 764 9548
rect 1235 9529 1272 9753
rect 1548 9749 1612 9761
rect 1652 9531 1679 9901
rect 1867 9896 1904 9906
rect 1963 9926 2050 9936
rect 1963 9906 1972 9926
rect 1992 9906 2050 9926
rect 1963 9897 2050 9906
rect 1963 9896 2000 9897
rect 1743 9883 1813 9888
rect 1738 9877 1813 9883
rect 1738 9844 1746 9877
rect 1799 9844 1813 9877
rect 2019 9844 2050 9897
rect 2080 9926 2117 10005
rect 2232 9936 2263 9937
rect 2080 9906 2089 9926
rect 2109 9906 2117 9926
rect 2080 9896 2117 9906
rect 2176 9929 2263 9936
rect 2176 9926 2237 9929
rect 2176 9906 2185 9926
rect 2205 9909 2237 9926
rect 2258 9909 2263 9929
rect 2205 9906 2263 9909
rect 2176 9899 2263 9906
rect 2288 9926 2325 10068
rect 2591 10067 2628 10068
rect 2440 9936 2476 9937
rect 2288 9906 2297 9926
rect 2317 9906 2325 9926
rect 2176 9897 2232 9899
rect 2176 9896 2213 9897
rect 2288 9896 2325 9906
rect 2384 9926 2532 9936
rect 2632 9933 2728 9935
rect 2384 9906 2393 9926
rect 2413 9906 2503 9926
rect 2523 9906 2532 9926
rect 2384 9900 2532 9906
rect 2384 9897 2448 9900
rect 2384 9896 2421 9897
rect 2440 9870 2448 9897
rect 2469 9897 2532 9900
rect 2590 9926 2728 9933
rect 2590 9906 2599 9926
rect 2619 9906 2728 9926
rect 2590 9897 2728 9906
rect 2469 9870 2476 9897
rect 2495 9896 2532 9897
rect 2591 9896 2628 9897
rect 2440 9845 2476 9870
rect 1738 9843 1821 9844
rect 1911 9843 1952 9844
rect 1738 9836 1952 9843
rect 1738 9819 1921 9836
rect 1738 9786 1751 9819
rect 1804 9816 1921 9819
rect 1941 9816 1952 9836
rect 1804 9808 1952 9816
rect 2019 9840 2378 9844
rect 2019 9835 2341 9840
rect 2019 9811 2132 9835
rect 2156 9816 2341 9835
rect 2365 9816 2378 9840
rect 2156 9811 2378 9816
rect 2019 9808 2378 9811
rect 2440 9808 2475 9845
rect 2543 9842 2643 9845
rect 2543 9838 2610 9842
rect 2543 9812 2555 9838
rect 2581 9816 2610 9838
rect 2636 9816 2643 9842
rect 2581 9812 2643 9816
rect 2543 9808 2643 9812
rect 1804 9786 1821 9808
rect 2019 9787 2050 9808
rect 2440 9787 2476 9808
rect 1862 9786 1899 9787
rect 1738 9772 1821 9786
rect 1511 9529 1679 9531
rect 1235 9528 1679 9529
rect 479 9498 1679 9528
rect 1749 9562 1821 9772
rect 1861 9777 1899 9786
rect 1861 9757 1870 9777
rect 1890 9757 1899 9777
rect 1861 9749 1899 9757
rect 1965 9781 2050 9787
rect 2075 9786 2112 9787
rect 1965 9761 1973 9781
rect 1993 9761 2050 9781
rect 1965 9753 2050 9761
rect 2074 9777 2112 9786
rect 2074 9757 2083 9777
rect 2103 9757 2112 9777
rect 1965 9752 2001 9753
rect 2074 9749 2112 9757
rect 2178 9781 2263 9787
rect 2283 9786 2320 9787
rect 2178 9761 2186 9781
rect 2206 9780 2263 9781
rect 2206 9761 2235 9780
rect 2178 9760 2235 9761
rect 2256 9760 2263 9780
rect 2178 9753 2263 9760
rect 2282 9777 2320 9786
rect 2282 9757 2291 9777
rect 2311 9757 2320 9777
rect 2178 9752 2214 9753
rect 2282 9749 2320 9757
rect 2386 9781 2530 9787
rect 2386 9761 2394 9781
rect 2414 9761 2502 9781
rect 2522 9761 2530 9781
rect 2386 9753 2530 9761
rect 2386 9752 2422 9753
rect 2494 9752 2530 9753
rect 2596 9786 2633 9787
rect 2596 9785 2634 9786
rect 2596 9777 2660 9785
rect 2596 9757 2605 9777
rect 2625 9763 2660 9777
rect 2680 9763 2683 9783
rect 2625 9758 2683 9763
rect 2625 9757 2660 9758
rect 1862 9720 1899 9749
rect 1863 9718 1899 9720
rect 2075 9718 2112 9749
rect 1863 9696 2112 9718
rect 1944 9690 2055 9696
rect 1944 9682 1985 9690
rect 1944 9662 1952 9682
rect 1971 9662 1985 9682
rect 1944 9660 1985 9662
rect 2013 9682 2055 9690
rect 2013 9662 2029 9682
rect 2048 9662 2055 9682
rect 2013 9660 2055 9662
rect 1944 9645 2055 9660
rect 1749 9523 1768 9562
rect 1813 9523 1821 9562
rect 1749 9506 1821 9523
rect 2283 9550 2320 9749
rect 2596 9745 2660 9757
rect 2283 9544 2324 9550
rect 2700 9546 2727 9897
rect 2856 9849 2927 10328
rect 2856 9765 2925 9849
rect 2559 9544 2727 9546
rect 2283 9518 2727 9544
rect 479 9451 544 9498
rect 479 9433 502 9451
rect 520 9433 544 9451
rect 1392 9478 1427 9480
rect 1392 9476 1496 9478
rect 2285 9476 2324 9518
rect 2559 9517 2727 9518
rect 1392 9469 2326 9476
rect 1392 9468 1443 9469
rect 1392 9448 1395 9468
rect 1420 9449 1443 9468
rect 1475 9449 2326 9469
rect 1420 9448 2326 9449
rect 1392 9441 2326 9448
rect 1665 9440 2326 9441
rect 479 9412 544 9433
rect 756 9423 796 9426
rect 756 9419 1659 9423
rect 756 9399 1633 9419
rect 1653 9399 1659 9419
rect 756 9396 1659 9399
rect 480 9352 545 9372
rect 480 9334 504 9352
rect 522 9334 545 9352
rect 480 9307 545 9334
rect 756 9307 796 9396
rect 1240 9394 1656 9396
rect 1240 9393 1581 9394
rect 897 9362 1007 9376
rect 897 9359 940 9362
rect 897 9354 901 9359
rect 479 9272 796 9307
rect 819 9332 901 9354
rect 930 9332 940 9359
rect 968 9335 975 9362
rect 1004 9354 1007 9362
rect 1004 9335 1069 9354
rect 968 9332 1069 9335
rect 819 9330 1069 9332
rect 480 9196 545 9272
rect 819 9251 856 9330
rect 897 9317 1007 9330
rect 971 9261 1002 9262
rect 819 9231 828 9251
rect 848 9231 856 9251
rect 819 9221 856 9231
rect 915 9251 1002 9261
rect 915 9231 924 9251
rect 944 9231 1002 9251
rect 915 9222 1002 9231
rect 915 9221 952 9222
rect 480 9178 502 9196
rect 520 9178 545 9196
rect 480 9157 545 9178
rect 693 9176 758 9185
rect 693 9139 703 9176
rect 743 9168 758 9176
rect 971 9169 1002 9222
rect 1032 9251 1069 9330
rect 1184 9261 1215 9262
rect 1032 9231 1041 9251
rect 1061 9231 1069 9251
rect 1032 9221 1069 9231
rect 1128 9254 1215 9261
rect 1128 9251 1189 9254
rect 1128 9231 1137 9251
rect 1157 9234 1189 9251
rect 1210 9234 1215 9254
rect 1157 9231 1215 9234
rect 1128 9224 1215 9231
rect 1240 9251 1277 9393
rect 1543 9392 1580 9393
rect 1392 9261 1428 9262
rect 1240 9231 1249 9251
rect 1269 9231 1277 9251
rect 1128 9222 1184 9224
rect 1128 9221 1165 9222
rect 1240 9221 1277 9231
rect 1336 9251 1484 9261
rect 1584 9258 1680 9260
rect 1336 9231 1345 9251
rect 1365 9231 1455 9251
rect 1475 9231 1484 9251
rect 1336 9225 1484 9231
rect 1336 9222 1400 9225
rect 1336 9221 1373 9222
rect 1392 9195 1400 9222
rect 1421 9222 1484 9225
rect 1542 9251 1680 9258
rect 1542 9231 1551 9251
rect 1571 9231 1680 9251
rect 2860 9249 2922 9765
rect 1542 9222 1680 9231
rect 1421 9195 1428 9222
rect 1447 9221 1484 9222
rect 1543 9221 1580 9222
rect 1392 9170 1428 9195
rect 863 9168 904 9169
rect 743 9161 904 9168
rect 743 9141 873 9161
rect 893 9141 904 9161
rect 743 9139 904 9141
rect 693 9133 904 9139
rect 971 9165 1330 9169
rect 971 9160 1293 9165
rect 971 9136 1084 9160
rect 1108 9141 1293 9160
rect 1317 9141 1330 9165
rect 1108 9136 1330 9141
rect 971 9133 1330 9136
rect 1392 9133 1427 9170
rect 1495 9167 1595 9170
rect 1495 9163 1562 9167
rect 1495 9137 1507 9163
rect 1533 9141 1562 9163
rect 1588 9141 1595 9167
rect 1533 9137 1595 9141
rect 1495 9133 1595 9137
rect 693 9120 760 9133
rect 485 9097 541 9117
rect 485 9079 504 9097
rect 522 9079 541 9097
rect 485 8966 541 9079
rect 693 9099 707 9120
rect 743 9099 760 9120
rect 971 9112 1002 9133
rect 1392 9112 1428 9133
rect 814 9111 851 9112
rect 693 9092 760 9099
rect 813 9102 851 9111
rect 485 8828 540 8966
rect 693 8940 758 9092
rect 813 9082 822 9102
rect 842 9082 851 9102
rect 813 9074 851 9082
rect 917 9106 1002 9112
rect 1027 9111 1064 9112
rect 917 9086 925 9106
rect 945 9086 1002 9106
rect 917 9078 1002 9086
rect 1026 9102 1064 9111
rect 1026 9082 1035 9102
rect 1055 9082 1064 9102
rect 917 9077 953 9078
rect 1026 9074 1064 9082
rect 1130 9106 1215 9112
rect 1235 9111 1272 9112
rect 1130 9086 1138 9106
rect 1158 9105 1215 9106
rect 1158 9086 1187 9105
rect 1130 9085 1187 9086
rect 1208 9085 1215 9105
rect 1130 9078 1215 9085
rect 1234 9102 1272 9111
rect 1234 9082 1243 9102
rect 1263 9082 1272 9102
rect 1130 9077 1166 9078
rect 1234 9074 1272 9082
rect 1338 9106 1482 9112
rect 1338 9086 1346 9106
rect 1366 9086 1454 9106
rect 1474 9086 1482 9106
rect 1338 9078 1482 9086
rect 1338 9077 1374 9078
rect 1446 9077 1482 9078
rect 1548 9111 1585 9112
rect 1548 9110 1586 9111
rect 1548 9102 1612 9110
rect 1548 9082 1557 9102
rect 1577 9088 1612 9102
rect 1632 9088 1635 9108
rect 1577 9083 1635 9088
rect 1577 9082 1612 9083
rect 814 9045 851 9074
rect 815 9043 851 9045
rect 1027 9043 1064 9074
rect 815 9021 1064 9043
rect 896 9015 1007 9021
rect 896 9007 937 9015
rect 896 8987 904 9007
rect 923 8987 937 9007
rect 896 8985 937 8987
rect 965 9007 1007 9015
rect 965 8987 981 9007
rect 1000 8987 1007 9007
rect 965 8985 1007 8987
rect 896 8972 1007 8985
rect 1235 8975 1272 9074
rect 1548 9070 1612 9082
rect 686 8930 807 8940
rect 686 8928 755 8930
rect 686 8887 699 8928
rect 736 8889 755 8928
rect 792 8889 807 8930
rect 736 8887 807 8889
rect 686 8869 807 8887
rect 478 8825 542 8828
rect 898 8825 1002 8831
rect 1233 8825 1274 8975
rect 1652 8967 1679 9222
rect 1741 9212 1821 9223
rect 1741 9186 1758 9212
rect 1798 9186 1821 9212
rect 1741 9159 1821 9186
rect 1741 9133 1762 9159
rect 1802 9133 1821 9159
rect 1741 9114 1821 9133
rect 1741 9088 1765 9114
rect 1805 9088 1821 9114
rect 1741 9037 1821 9088
rect 2844 9214 2922 9249
rect 2844 9152 2926 9214
rect 2844 9129 2872 9152
rect 2898 9129 2926 9152
rect 2844 9109 2926 9129
rect 478 8822 1274 8825
rect 1653 8836 1679 8967
rect 1653 8822 1681 8836
rect 478 8787 1681 8822
rect 1743 8829 1813 9037
rect 478 8726 542 8787
rect 898 8785 1002 8787
rect 1233 8785 1274 8787
rect 1743 8784 1764 8829
rect 1744 8763 1764 8784
rect 1794 8784 1813 8829
rect 1794 8763 1811 8784
rect 1744 8744 1811 8763
rect 1393 8736 1465 8737
rect 1392 8728 1491 8736
rect 480 8655 539 8726
rect 1392 8725 1444 8728
rect 1392 8690 1400 8725
rect 1425 8690 1444 8725
rect 1469 8717 1491 8728
rect 1469 8716 2336 8717
rect 1469 8690 2337 8716
rect 1392 8680 2337 8690
rect 1392 8678 1491 8680
rect 480 8637 502 8655
rect 520 8637 539 8655
rect 480 8615 539 8637
rect 747 8651 1279 8656
rect 747 8631 1633 8651
rect 1653 8631 1656 8651
rect 2292 8647 2337 8680
rect 747 8627 1656 8631
rect 747 8580 790 8627
rect 1240 8626 1656 8627
rect 2288 8627 2681 8647
rect 2701 8627 2704 8647
rect 1240 8625 1581 8626
rect 897 8594 1007 8608
rect 897 8591 940 8594
rect 897 8586 901 8591
rect 735 8579 790 8580
rect 479 8556 790 8579
rect 479 8538 504 8556
rect 522 8544 790 8556
rect 819 8564 901 8586
rect 930 8564 940 8591
rect 968 8567 975 8594
rect 1004 8586 1007 8594
rect 1004 8567 1069 8586
rect 968 8564 1069 8567
rect 819 8562 1069 8564
rect 522 8538 544 8544
rect 479 8399 544 8538
rect 819 8483 856 8562
rect 897 8549 1007 8562
rect 971 8493 1002 8494
rect 819 8463 828 8483
rect 848 8463 856 8483
rect 479 8381 502 8399
rect 520 8381 544 8399
rect 479 8364 544 8381
rect 699 8445 767 8458
rect 819 8453 856 8463
rect 915 8483 1002 8493
rect 915 8463 924 8483
rect 944 8463 1002 8483
rect 915 8454 1002 8463
rect 915 8453 952 8454
rect 699 8403 706 8445
rect 755 8403 767 8445
rect 699 8400 767 8403
rect 971 8401 1002 8454
rect 1032 8483 1069 8562
rect 1184 8493 1215 8494
rect 1032 8463 1041 8483
rect 1061 8463 1069 8483
rect 1032 8453 1069 8463
rect 1128 8486 1215 8493
rect 1128 8483 1189 8486
rect 1128 8463 1137 8483
rect 1157 8466 1189 8483
rect 1210 8466 1215 8486
rect 1157 8463 1215 8466
rect 1128 8456 1215 8463
rect 1240 8483 1277 8625
rect 1543 8624 1580 8625
rect 2288 8622 2704 8627
rect 2288 8621 2629 8622
rect 1945 8590 2055 8604
rect 1945 8587 1988 8590
rect 1945 8582 1949 8587
rect 1867 8560 1949 8582
rect 1978 8560 1988 8587
rect 2016 8563 2023 8590
rect 2052 8582 2055 8590
rect 2052 8563 2117 8582
rect 2016 8560 2117 8563
rect 1867 8558 2117 8560
rect 1392 8493 1428 8494
rect 1240 8463 1249 8483
rect 1269 8463 1277 8483
rect 1128 8454 1184 8456
rect 1128 8453 1165 8454
rect 1240 8453 1277 8463
rect 1336 8483 1484 8493
rect 1584 8490 1680 8492
rect 1336 8463 1345 8483
rect 1365 8463 1455 8483
rect 1475 8463 1484 8483
rect 1336 8457 1484 8463
rect 1336 8454 1400 8457
rect 1336 8453 1373 8454
rect 1392 8427 1400 8454
rect 1421 8454 1484 8457
rect 1542 8483 1680 8490
rect 1542 8463 1551 8483
rect 1571 8463 1680 8483
rect 1542 8454 1680 8463
rect 1867 8479 1904 8558
rect 1945 8545 2055 8558
rect 2019 8489 2050 8490
rect 1867 8459 1876 8479
rect 1896 8459 1904 8479
rect 1421 8427 1428 8454
rect 1447 8453 1484 8454
rect 1543 8453 1580 8454
rect 1392 8402 1428 8427
rect 863 8400 904 8401
rect 699 8393 904 8400
rect 699 8382 873 8393
rect 699 8349 707 8382
rect 700 8340 707 8349
rect 756 8373 873 8382
rect 893 8373 904 8393
rect 756 8365 904 8373
rect 971 8397 1330 8401
rect 971 8392 1293 8397
rect 971 8368 1084 8392
rect 1108 8373 1293 8392
rect 1317 8373 1330 8397
rect 1108 8368 1330 8373
rect 971 8365 1330 8368
rect 1392 8365 1427 8402
rect 1495 8399 1595 8402
rect 1495 8395 1562 8399
rect 1495 8369 1507 8395
rect 1533 8373 1562 8395
rect 1588 8373 1595 8399
rect 1533 8369 1595 8373
rect 1495 8365 1595 8369
rect 756 8349 767 8365
rect 756 8340 764 8349
rect 971 8344 1002 8365
rect 1392 8344 1428 8365
rect 814 8343 851 8344
rect 479 8300 544 8319
rect 479 8282 504 8300
rect 522 8282 544 8300
rect 479 8081 544 8282
rect 700 8156 764 8340
rect 813 8334 851 8343
rect 813 8314 822 8334
rect 842 8314 851 8334
rect 813 8306 851 8314
rect 917 8338 1002 8344
rect 1027 8343 1064 8344
rect 917 8318 925 8338
rect 945 8318 1002 8338
rect 917 8310 1002 8318
rect 1026 8334 1064 8343
rect 1026 8314 1035 8334
rect 1055 8314 1064 8334
rect 917 8309 953 8310
rect 1026 8306 1064 8314
rect 1130 8338 1215 8344
rect 1235 8343 1272 8344
rect 1130 8318 1138 8338
rect 1158 8337 1215 8338
rect 1158 8318 1187 8337
rect 1130 8317 1187 8318
rect 1208 8317 1215 8337
rect 1130 8310 1215 8317
rect 1234 8334 1272 8343
rect 1234 8314 1243 8334
rect 1263 8314 1272 8334
rect 1130 8309 1166 8310
rect 1234 8306 1272 8314
rect 1338 8338 1482 8344
rect 1338 8318 1346 8338
rect 1366 8318 1454 8338
rect 1474 8318 1482 8338
rect 1338 8310 1482 8318
rect 1338 8309 1374 8310
rect 1446 8309 1482 8310
rect 1548 8343 1585 8344
rect 1548 8342 1586 8343
rect 1548 8334 1612 8342
rect 1548 8314 1557 8334
rect 1577 8320 1612 8334
rect 1632 8320 1635 8340
rect 1577 8315 1635 8320
rect 1577 8314 1612 8315
rect 814 8277 851 8306
rect 815 8275 851 8277
rect 1027 8275 1064 8306
rect 815 8253 1064 8275
rect 896 8247 1007 8253
rect 896 8239 937 8247
rect 896 8219 904 8239
rect 923 8219 937 8239
rect 896 8217 937 8219
rect 965 8239 1007 8247
rect 965 8219 981 8239
rect 1000 8219 1007 8239
rect 965 8217 1007 8219
rect 896 8202 1007 8217
rect 700 8146 768 8156
rect 700 8113 717 8146
rect 757 8113 768 8146
rect 700 8101 768 8113
rect 700 8099 764 8101
rect 1235 8082 1272 8306
rect 1548 8302 1612 8314
rect 1652 8084 1679 8454
rect 1867 8449 1904 8459
rect 1963 8479 2050 8489
rect 1963 8459 1972 8479
rect 1992 8459 2050 8479
rect 1963 8450 2050 8459
rect 1963 8449 2000 8450
rect 1743 8436 1813 8441
rect 1738 8430 1813 8436
rect 1738 8397 1746 8430
rect 1799 8397 1813 8430
rect 2019 8397 2050 8450
rect 2080 8479 2117 8558
rect 2232 8489 2263 8490
rect 2080 8459 2089 8479
rect 2109 8459 2117 8479
rect 2080 8449 2117 8459
rect 2176 8482 2263 8489
rect 2176 8479 2237 8482
rect 2176 8459 2185 8479
rect 2205 8462 2237 8479
rect 2258 8462 2263 8482
rect 2205 8459 2263 8462
rect 2176 8452 2263 8459
rect 2288 8479 2325 8621
rect 2591 8620 2628 8621
rect 2440 8489 2476 8490
rect 2288 8459 2297 8479
rect 2317 8459 2325 8479
rect 2176 8450 2232 8452
rect 2176 8449 2213 8450
rect 2288 8449 2325 8459
rect 2384 8479 2532 8489
rect 2632 8486 2728 8488
rect 2384 8459 2393 8479
rect 2413 8459 2503 8479
rect 2523 8459 2532 8479
rect 2384 8453 2532 8459
rect 2384 8450 2448 8453
rect 2384 8449 2421 8450
rect 2440 8423 2448 8450
rect 2469 8450 2532 8453
rect 2590 8479 2728 8486
rect 2590 8459 2599 8479
rect 2619 8459 2728 8479
rect 2590 8450 2728 8459
rect 2469 8423 2476 8450
rect 2495 8449 2532 8450
rect 2591 8449 2628 8450
rect 2440 8398 2476 8423
rect 1738 8396 1821 8397
rect 1911 8396 1952 8397
rect 1738 8389 1952 8396
rect 1738 8372 1921 8389
rect 1738 8339 1751 8372
rect 1804 8369 1921 8372
rect 1941 8369 1952 8389
rect 1804 8361 1952 8369
rect 2019 8393 2378 8397
rect 2019 8388 2341 8393
rect 2019 8364 2132 8388
rect 2156 8369 2341 8388
rect 2365 8369 2378 8393
rect 2156 8364 2378 8369
rect 2019 8361 2378 8364
rect 2440 8361 2475 8398
rect 2543 8395 2643 8398
rect 2543 8391 2610 8395
rect 2543 8365 2555 8391
rect 2581 8369 2610 8391
rect 2636 8369 2643 8395
rect 2581 8365 2643 8369
rect 2543 8361 2643 8365
rect 1804 8339 1821 8361
rect 2019 8340 2050 8361
rect 2440 8340 2476 8361
rect 1862 8339 1899 8340
rect 1738 8325 1821 8339
rect 1511 8082 1679 8084
rect 1235 8081 1679 8082
rect 479 8051 1679 8081
rect 1749 8115 1821 8325
rect 1861 8330 1899 8339
rect 1861 8310 1870 8330
rect 1890 8310 1899 8330
rect 1861 8302 1899 8310
rect 1965 8334 2050 8340
rect 2075 8339 2112 8340
rect 1965 8314 1973 8334
rect 1993 8314 2050 8334
rect 1965 8306 2050 8314
rect 2074 8330 2112 8339
rect 2074 8310 2083 8330
rect 2103 8310 2112 8330
rect 1965 8305 2001 8306
rect 2074 8302 2112 8310
rect 2178 8334 2263 8340
rect 2283 8339 2320 8340
rect 2178 8314 2186 8334
rect 2206 8333 2263 8334
rect 2206 8314 2235 8333
rect 2178 8313 2235 8314
rect 2256 8313 2263 8333
rect 2178 8306 2263 8313
rect 2282 8330 2320 8339
rect 2282 8310 2291 8330
rect 2311 8310 2320 8330
rect 2178 8305 2214 8306
rect 2282 8302 2320 8310
rect 2386 8334 2530 8340
rect 2386 8314 2394 8334
rect 2414 8314 2502 8334
rect 2522 8314 2530 8334
rect 2386 8306 2530 8314
rect 2386 8305 2422 8306
rect 2494 8305 2530 8306
rect 2596 8339 2633 8340
rect 2596 8338 2634 8339
rect 2596 8330 2660 8338
rect 2596 8310 2605 8330
rect 2625 8316 2660 8330
rect 2680 8316 2683 8336
rect 2625 8311 2683 8316
rect 2625 8310 2660 8311
rect 1862 8273 1899 8302
rect 1863 8271 1899 8273
rect 2075 8271 2112 8302
rect 1863 8249 2112 8271
rect 1944 8243 2055 8249
rect 1944 8235 1985 8243
rect 1944 8215 1952 8235
rect 1971 8215 1985 8235
rect 1944 8213 1985 8215
rect 2013 8235 2055 8243
rect 2013 8215 2029 8235
rect 2048 8215 2055 8235
rect 2013 8213 2055 8215
rect 1944 8198 2055 8213
rect 1749 8076 1768 8115
rect 1813 8076 1821 8115
rect 1749 8059 1821 8076
rect 2283 8103 2320 8302
rect 2596 8298 2660 8310
rect 2283 8097 2324 8103
rect 2700 8099 2727 8450
rect 2559 8097 2727 8099
rect 2283 8071 2727 8097
rect 479 8004 544 8051
rect 479 7986 502 8004
rect 520 7986 544 8004
rect 1392 8031 1427 8033
rect 1392 8029 1496 8031
rect 2285 8029 2324 8071
rect 2559 8070 2727 8071
rect 1392 8022 2326 8029
rect 1392 8021 1443 8022
rect 1392 8001 1395 8021
rect 1420 8002 1443 8021
rect 1475 8002 2326 8022
rect 1420 8001 2326 8002
rect 1392 7994 2326 8001
rect 1665 7993 2326 7994
rect 479 7965 544 7986
rect 756 7976 796 7979
rect 756 7972 1659 7976
rect 756 7952 1633 7972
rect 1653 7952 1659 7972
rect 756 7949 1659 7952
rect 480 7905 545 7925
rect 480 7887 504 7905
rect 522 7887 545 7905
rect 480 7860 545 7887
rect 756 7860 796 7949
rect 1240 7947 1656 7949
rect 1240 7946 1581 7947
rect 897 7915 1007 7929
rect 897 7912 940 7915
rect 897 7907 901 7912
rect 479 7825 796 7860
rect 819 7885 901 7907
rect 930 7885 940 7912
rect 968 7888 975 7915
rect 1004 7907 1007 7915
rect 1004 7888 1069 7907
rect 968 7885 1069 7888
rect 819 7883 1069 7885
rect 480 7749 545 7825
rect 819 7804 856 7883
rect 897 7870 1007 7883
rect 971 7814 1002 7815
rect 819 7784 828 7804
rect 848 7784 856 7804
rect 819 7774 856 7784
rect 915 7804 1002 7814
rect 915 7784 924 7804
rect 944 7784 1002 7804
rect 915 7775 1002 7784
rect 915 7774 952 7775
rect 480 7731 502 7749
rect 520 7731 545 7749
rect 480 7710 545 7731
rect 693 7729 758 7738
rect 693 7692 703 7729
rect 743 7721 758 7729
rect 971 7722 1002 7775
rect 1032 7804 1069 7883
rect 1184 7814 1215 7815
rect 1032 7784 1041 7804
rect 1061 7784 1069 7804
rect 1032 7774 1069 7784
rect 1128 7807 1215 7814
rect 1128 7804 1189 7807
rect 1128 7784 1137 7804
rect 1157 7787 1189 7804
rect 1210 7787 1215 7807
rect 1157 7784 1215 7787
rect 1128 7777 1215 7784
rect 1240 7804 1277 7946
rect 1543 7945 1580 7946
rect 1392 7814 1428 7815
rect 1240 7784 1249 7804
rect 1269 7784 1277 7804
rect 1128 7775 1184 7777
rect 1128 7774 1165 7775
rect 1240 7774 1277 7784
rect 1336 7804 1484 7814
rect 1584 7811 1680 7813
rect 1336 7784 1345 7804
rect 1365 7784 1455 7804
rect 1475 7784 1484 7804
rect 1336 7778 1484 7784
rect 1336 7775 1400 7778
rect 1336 7774 1373 7775
rect 1392 7748 1400 7775
rect 1421 7775 1484 7778
rect 1542 7804 1680 7811
rect 1542 7784 1551 7804
rect 1571 7784 1680 7804
rect 1542 7775 1680 7784
rect 1421 7748 1428 7775
rect 1447 7774 1484 7775
rect 1543 7774 1580 7775
rect 1392 7723 1428 7748
rect 863 7721 904 7722
rect 743 7714 904 7721
rect 743 7694 873 7714
rect 893 7694 904 7714
rect 743 7692 904 7694
rect 693 7686 904 7692
rect 971 7718 1330 7722
rect 971 7713 1293 7718
rect 971 7689 1084 7713
rect 1108 7694 1293 7713
rect 1317 7694 1330 7718
rect 1108 7689 1330 7694
rect 971 7686 1330 7689
rect 1392 7686 1427 7723
rect 1495 7720 1595 7723
rect 1495 7716 1562 7720
rect 1495 7690 1507 7716
rect 1533 7694 1562 7716
rect 1588 7694 1595 7720
rect 1533 7690 1595 7694
rect 1495 7686 1595 7690
rect 693 7673 760 7686
rect 485 7650 541 7670
rect 485 7632 504 7650
rect 522 7632 541 7650
rect 485 7519 541 7632
rect 693 7652 707 7673
rect 743 7652 760 7673
rect 971 7665 1002 7686
rect 1392 7665 1428 7686
rect 814 7664 851 7665
rect 693 7645 760 7652
rect 813 7655 851 7664
rect 485 7412 540 7519
rect 693 7493 758 7645
rect 813 7635 822 7655
rect 842 7635 851 7655
rect 813 7627 851 7635
rect 917 7659 1002 7665
rect 1027 7664 1064 7665
rect 917 7639 925 7659
rect 945 7639 1002 7659
rect 917 7631 1002 7639
rect 1026 7655 1064 7664
rect 1026 7635 1035 7655
rect 1055 7635 1064 7655
rect 917 7630 953 7631
rect 1026 7627 1064 7635
rect 1130 7659 1215 7665
rect 1235 7664 1272 7665
rect 1130 7639 1138 7659
rect 1158 7658 1215 7659
rect 1158 7639 1187 7658
rect 1130 7638 1187 7639
rect 1208 7638 1215 7658
rect 1130 7631 1215 7638
rect 1234 7655 1272 7664
rect 1234 7635 1243 7655
rect 1263 7635 1272 7655
rect 1130 7630 1166 7631
rect 1234 7627 1272 7635
rect 1338 7659 1482 7665
rect 1338 7639 1346 7659
rect 1366 7639 1454 7659
rect 1474 7639 1482 7659
rect 1338 7631 1482 7639
rect 1338 7630 1374 7631
rect 1446 7630 1482 7631
rect 1548 7664 1585 7665
rect 1548 7663 1586 7664
rect 1548 7655 1612 7663
rect 1548 7635 1557 7655
rect 1577 7641 1612 7655
rect 1632 7641 1635 7661
rect 1577 7636 1635 7641
rect 1577 7635 1612 7636
rect 814 7598 851 7627
rect 815 7596 851 7598
rect 1027 7596 1064 7627
rect 815 7574 1064 7596
rect 896 7568 1007 7574
rect 896 7560 937 7568
rect 896 7540 904 7560
rect 923 7540 937 7560
rect 896 7538 937 7540
rect 965 7560 1007 7568
rect 965 7540 981 7560
rect 1000 7540 1007 7560
rect 965 7538 1007 7540
rect 896 7523 1007 7538
rect 1235 7528 1272 7627
rect 1548 7623 1612 7635
rect 898 7520 1002 7523
rect 686 7483 807 7493
rect 686 7481 755 7483
rect 686 7440 699 7481
rect 736 7442 755 7481
rect 792 7442 807 7483
rect 736 7440 807 7442
rect 686 7422 807 7440
rect 478 7378 543 7412
rect 898 7378 1002 7380
rect 1233 7378 1274 7528
rect 1652 7520 1679 7775
rect 1741 7765 1821 7776
rect 1741 7739 1758 7765
rect 1798 7739 1821 7765
rect 1741 7712 1821 7739
rect 1741 7686 1762 7712
rect 1802 7686 1821 7712
rect 1741 7667 1821 7686
rect 1741 7641 1765 7667
rect 1805 7641 1821 7667
rect 1741 7590 1821 7641
rect 478 7375 1274 7378
rect 1653 7389 1679 7520
rect 1743 7390 1813 7590
rect 1653 7375 1681 7389
rect 478 7340 1681 7375
rect 1742 7368 1814 7390
rect 478 7183 543 7340
rect 898 7338 1002 7340
rect 1233 7338 1274 7340
rect 1742 7320 1756 7368
rect 1802 7320 1814 7368
rect 1742 7303 1814 7320
rect 2844 7270 2916 9109
rect 3022 7342 3114 10646
rect 3508 10629 3539 10650
rect 3929 10629 3965 10650
rect 3351 10628 3388 10629
rect 3350 10619 3388 10628
rect 3350 10599 3359 10619
rect 3379 10599 3388 10619
rect 3350 10591 3388 10599
rect 3454 10623 3539 10629
rect 3564 10628 3601 10629
rect 3454 10603 3462 10623
rect 3482 10603 3539 10623
rect 3454 10595 3539 10603
rect 3563 10619 3601 10628
rect 3563 10599 3572 10619
rect 3592 10599 3601 10619
rect 3454 10594 3490 10595
rect 3563 10591 3601 10599
rect 3667 10623 3752 10629
rect 3772 10628 3809 10629
rect 3667 10603 3675 10623
rect 3695 10622 3752 10623
rect 3695 10603 3724 10622
rect 3667 10602 3724 10603
rect 3745 10602 3752 10622
rect 3667 10595 3752 10602
rect 3771 10619 3809 10628
rect 3771 10599 3780 10619
rect 3800 10599 3809 10619
rect 3667 10594 3703 10595
rect 3771 10591 3809 10599
rect 3875 10623 4019 10629
rect 3875 10603 3883 10623
rect 3903 10603 3991 10623
rect 4011 10603 4019 10623
rect 3875 10595 4019 10603
rect 3875 10594 3911 10595
rect 3983 10594 4019 10595
rect 4085 10628 4122 10629
rect 4085 10627 4123 10628
rect 4085 10619 4149 10627
rect 4085 10599 4094 10619
rect 4114 10605 4149 10619
rect 4169 10605 4172 10625
rect 4114 10600 4172 10605
rect 4114 10599 4149 10600
rect 3351 10562 3388 10591
rect 3352 10560 3388 10562
rect 3564 10560 3601 10591
rect 3352 10538 3601 10560
rect 3433 10532 3544 10538
rect 3433 10524 3474 10532
rect 3433 10504 3441 10524
rect 3460 10504 3474 10524
rect 3433 10502 3474 10504
rect 3502 10524 3544 10532
rect 3502 10504 3518 10524
rect 3537 10504 3544 10524
rect 3502 10502 3544 10504
rect 3433 10487 3544 10502
rect 3772 10470 3809 10591
rect 4085 10587 4149 10599
rect 3890 10470 3919 10474
rect 4189 10472 4216 10739
rect 4048 10470 4216 10472
rect 3772 10444 4216 10470
rect 3731 10176 3776 10185
rect 3731 10138 3741 10176
rect 3766 10138 3776 10176
rect 3731 10127 3776 10138
rect 3734 10119 3776 10127
rect 3734 9414 3777 10119
rect 3890 9505 3919 10444
rect 4048 10443 4216 10444
rect 3888 9484 3925 9505
rect 3888 9447 3899 9484
rect 3916 9447 3925 9484
rect 3888 9437 3925 9447
rect 3734 9394 4128 9414
rect 4148 9394 4151 9414
rect 3735 9389 4151 9394
rect 3735 9388 4076 9389
rect 3392 9357 3502 9371
rect 3392 9354 3435 9357
rect 3392 9349 3396 9354
rect 3314 9327 3396 9349
rect 3425 9327 3435 9354
rect 3463 9330 3470 9357
rect 3499 9349 3502 9357
rect 3499 9330 3564 9349
rect 3463 9327 3564 9330
rect 3314 9325 3564 9327
rect 3314 9246 3351 9325
rect 3392 9312 3502 9325
rect 3466 9256 3497 9257
rect 3314 9226 3323 9246
rect 3343 9226 3351 9246
rect 3314 9216 3351 9226
rect 3410 9246 3497 9256
rect 3410 9226 3419 9246
rect 3439 9226 3497 9246
rect 3410 9217 3497 9226
rect 3410 9216 3447 9217
rect 3466 9164 3497 9217
rect 3527 9246 3564 9325
rect 3679 9256 3710 9257
rect 3527 9226 3536 9246
rect 3556 9226 3564 9246
rect 3527 9216 3564 9226
rect 3623 9249 3710 9256
rect 3623 9246 3684 9249
rect 3623 9226 3632 9246
rect 3652 9229 3684 9246
rect 3705 9229 3710 9249
rect 3652 9226 3710 9229
rect 3623 9219 3710 9226
rect 3735 9246 3772 9388
rect 4038 9387 4075 9388
rect 3887 9256 3923 9257
rect 3735 9226 3744 9246
rect 3764 9226 3772 9246
rect 3623 9217 3679 9219
rect 3623 9216 3660 9217
rect 3735 9216 3772 9226
rect 3831 9246 3979 9256
rect 4079 9253 4175 9255
rect 3831 9226 3840 9246
rect 3860 9226 3950 9246
rect 3970 9226 3979 9246
rect 3831 9220 3979 9226
rect 3831 9217 3895 9220
rect 3831 9216 3868 9217
rect 3887 9190 3895 9217
rect 3916 9217 3979 9220
rect 4037 9246 4175 9253
rect 4037 9226 4046 9246
rect 4066 9226 4175 9246
rect 4037 9217 4175 9226
rect 3916 9190 3923 9217
rect 3942 9216 3979 9217
rect 4038 9216 4075 9217
rect 3887 9165 3923 9190
rect 3358 9163 3399 9164
rect 3278 9158 3399 9163
rect 3229 9156 3399 9158
rect 3229 9145 3368 9156
rect 3229 9122 3252 9145
rect 3278 9136 3368 9145
rect 3388 9136 3399 9156
rect 3278 9128 3399 9136
rect 3466 9160 3825 9164
rect 3466 9155 3788 9160
rect 3466 9131 3579 9155
rect 3603 9136 3788 9155
rect 3812 9136 3825 9160
rect 3603 9131 3825 9136
rect 3466 9128 3825 9131
rect 3887 9128 3922 9165
rect 3990 9162 4090 9165
rect 3990 9158 4057 9162
rect 3990 9132 4002 9158
rect 4028 9136 4057 9158
rect 4083 9136 4090 9162
rect 4028 9132 4090 9136
rect 3990 9128 4090 9132
rect 3278 9122 3286 9128
rect 3229 9114 3286 9122
rect 3466 9107 3497 9128
rect 3887 9107 3923 9128
rect 3309 9106 3346 9107
rect 3308 9097 3346 9106
rect 3308 9077 3317 9097
rect 3337 9077 3346 9097
rect 3308 9069 3346 9077
rect 3412 9101 3497 9107
rect 3522 9106 3559 9107
rect 3412 9081 3420 9101
rect 3440 9081 3497 9101
rect 3412 9073 3497 9081
rect 3521 9097 3559 9106
rect 3521 9077 3530 9097
rect 3550 9077 3559 9097
rect 3412 9072 3448 9073
rect 3521 9069 3559 9077
rect 3625 9101 3710 9107
rect 3730 9106 3767 9107
rect 3625 9081 3633 9101
rect 3653 9100 3710 9101
rect 3653 9081 3682 9100
rect 3625 9080 3682 9081
rect 3703 9080 3710 9100
rect 3625 9073 3710 9080
rect 3729 9097 3767 9106
rect 3729 9077 3738 9097
rect 3758 9077 3767 9097
rect 3625 9072 3661 9073
rect 3729 9069 3767 9077
rect 3833 9101 3977 9107
rect 3833 9081 3841 9101
rect 3861 9081 3949 9101
rect 3969 9081 3977 9101
rect 3833 9073 3977 9081
rect 3833 9072 3869 9073
rect 3941 9072 3977 9073
rect 4043 9106 4080 9107
rect 4043 9105 4081 9106
rect 4043 9097 4107 9105
rect 4043 9077 4052 9097
rect 4072 9083 4107 9097
rect 4127 9083 4130 9103
rect 4072 9078 4130 9083
rect 4072 9077 4107 9078
rect 3309 9040 3346 9069
rect 3310 9038 3346 9040
rect 3522 9038 3559 9069
rect 3310 9016 3559 9038
rect 3391 9010 3502 9016
rect 3391 9002 3432 9010
rect 3391 8982 3399 9002
rect 3418 8982 3432 9002
rect 3391 8980 3432 8982
rect 3460 9002 3502 9010
rect 3460 8982 3476 9002
rect 3495 8982 3502 9002
rect 3460 8980 3502 8982
rect 3391 8965 3502 8980
rect 3730 8954 3767 9069
rect 4043 9065 4107 9077
rect 3723 8948 3770 8954
rect 4147 8950 4174 9217
rect 4006 8948 4174 8950
rect 3723 8922 4174 8948
rect 3723 8787 3770 8922
rect 4006 8921 4174 8922
rect 3721 8738 3780 8787
rect 3721 8710 3739 8738
rect 3767 8710 3780 8738
rect 3721 8700 3780 8710
rect 4836 7963 4914 11003
rect 4836 7943 5236 7963
rect 5256 7943 5259 7963
rect 4836 7941 5259 7943
rect 4843 7938 5259 7941
rect 4843 7937 5184 7938
rect 4500 7906 4610 7920
rect 4500 7903 4543 7906
rect 4500 7898 4504 7903
rect 4422 7876 4504 7898
rect 4533 7876 4543 7903
rect 4571 7879 4578 7906
rect 4607 7898 4610 7906
rect 4607 7879 4672 7898
rect 4571 7876 4672 7879
rect 4422 7874 4672 7876
rect 4422 7795 4459 7874
rect 4500 7861 4610 7874
rect 4574 7805 4605 7806
rect 4422 7775 4431 7795
rect 4451 7775 4459 7795
rect 4422 7765 4459 7775
rect 4518 7795 4605 7805
rect 4518 7775 4527 7795
rect 4547 7775 4605 7795
rect 4518 7766 4605 7775
rect 4518 7765 4555 7766
rect 4292 7712 4403 7715
rect 4574 7713 4605 7766
rect 4635 7795 4672 7874
rect 4787 7805 4818 7806
rect 4635 7775 4644 7795
rect 4664 7775 4672 7795
rect 4635 7765 4672 7775
rect 4731 7798 4818 7805
rect 4731 7795 4792 7798
rect 4731 7775 4740 7795
rect 4760 7778 4792 7795
rect 4813 7778 4818 7798
rect 4760 7775 4818 7778
rect 4731 7768 4818 7775
rect 4843 7795 4880 7937
rect 5146 7936 5183 7937
rect 4995 7805 5031 7806
rect 4843 7775 4852 7795
rect 4872 7775 4880 7795
rect 4731 7766 4787 7768
rect 4731 7765 4768 7766
rect 4843 7765 4880 7775
rect 4939 7795 5087 7805
rect 5187 7802 5283 7804
rect 4939 7775 4948 7795
rect 4968 7775 5058 7795
rect 5078 7775 5087 7795
rect 4939 7769 5087 7775
rect 4939 7766 5003 7769
rect 4939 7765 4976 7766
rect 4995 7739 5003 7766
rect 5024 7766 5087 7769
rect 5145 7795 5283 7802
rect 5145 7775 5154 7795
rect 5174 7775 5283 7795
rect 5145 7766 5283 7775
rect 5024 7739 5031 7766
rect 5050 7765 5087 7766
rect 5146 7765 5183 7766
rect 4995 7714 5031 7739
rect 4466 7712 4507 7713
rect 4292 7705 4507 7712
rect 4292 7704 4357 7705
rect 4292 7680 4300 7704
rect 4324 7681 4357 7704
rect 4381 7685 4476 7705
rect 4496 7685 4507 7705
rect 4381 7681 4507 7685
rect 4324 7680 4507 7681
rect 4292 7677 4507 7680
rect 4574 7709 4933 7713
rect 4574 7704 4896 7709
rect 4574 7680 4687 7704
rect 4711 7685 4896 7704
rect 4920 7685 4933 7709
rect 4711 7680 4933 7685
rect 4574 7677 4933 7680
rect 4995 7677 5030 7714
rect 5098 7711 5198 7714
rect 5098 7707 5165 7711
rect 5098 7681 5110 7707
rect 5136 7685 5165 7707
rect 5191 7685 5198 7711
rect 5136 7681 5198 7685
rect 5098 7677 5198 7681
rect 4292 7673 4403 7677
rect 4574 7656 4605 7677
rect 4995 7656 5031 7677
rect 4417 7655 4454 7656
rect 4416 7646 4454 7655
rect 4416 7626 4425 7646
rect 4445 7626 4454 7646
rect 4416 7618 4454 7626
rect 4520 7650 4605 7656
rect 4630 7655 4667 7656
rect 4520 7630 4528 7650
rect 4548 7630 4605 7650
rect 4520 7622 4605 7630
rect 4629 7646 4667 7655
rect 4629 7626 4638 7646
rect 4658 7626 4667 7646
rect 4520 7621 4556 7622
rect 4629 7618 4667 7626
rect 4733 7650 4818 7656
rect 4838 7655 4875 7656
rect 4733 7630 4741 7650
rect 4761 7649 4818 7650
rect 4761 7630 4790 7649
rect 4733 7629 4790 7630
rect 4811 7629 4818 7649
rect 4733 7622 4818 7629
rect 4837 7646 4875 7655
rect 4837 7626 4846 7646
rect 4866 7626 4875 7646
rect 4733 7621 4769 7622
rect 4837 7618 4875 7626
rect 4941 7650 5085 7656
rect 4941 7630 4949 7650
rect 4969 7649 5057 7650
rect 4969 7630 5003 7649
rect 4941 7627 5003 7630
rect 5027 7630 5057 7649
rect 5077 7630 5085 7650
rect 5027 7627 5085 7630
rect 4941 7622 5085 7627
rect 4941 7621 4977 7622
rect 5049 7621 5085 7622
rect 5151 7655 5188 7656
rect 5151 7654 5189 7655
rect 5151 7646 5215 7654
rect 5151 7626 5160 7646
rect 5180 7632 5215 7646
rect 5235 7632 5238 7652
rect 5180 7627 5238 7632
rect 5180 7626 5215 7627
rect 4417 7589 4454 7618
rect 4418 7587 4454 7589
rect 4630 7587 4667 7618
rect 4418 7565 4667 7587
rect 4499 7559 4610 7565
rect 4499 7551 4540 7559
rect 4499 7531 4507 7551
rect 4526 7531 4540 7551
rect 4499 7529 4540 7531
rect 4568 7551 4610 7559
rect 4568 7531 4584 7551
rect 4603 7531 4610 7551
rect 4568 7529 4610 7531
rect 4499 7514 4610 7529
rect 4838 7503 4875 7618
rect 5151 7614 5215 7626
rect 4834 7497 4889 7503
rect 5255 7499 5282 7766
rect 5114 7497 5282 7499
rect 4834 7472 5282 7497
rect 5595 7557 5701 12755
rect 8867 12745 8890 12771
rect 8930 12745 8947 12771
rect 8867 12734 8947 12745
rect 9009 12735 9036 12990
rect 9414 12982 9455 13132
rect 10126 13101 11249 13132
rect 12099 13136 12198 13144
rect 12099 13133 12151 13136
rect 9881 13070 10002 13088
rect 9881 13068 9952 13070
rect 9881 13027 9896 13068
rect 9933 13029 9952 13068
rect 9989 13029 10002 13070
rect 9933 13027 10002 13029
rect 9881 13017 10002 13027
rect 9076 12875 9140 12887
rect 9416 12883 9453 12982
rect 9681 12972 9792 12983
rect 9681 12970 9723 12972
rect 9681 12950 9688 12970
rect 9707 12950 9723 12970
rect 9681 12942 9723 12950
rect 9751 12970 9792 12972
rect 9751 12950 9765 12970
rect 9784 12950 9792 12970
rect 9751 12942 9792 12950
rect 9681 12936 9792 12942
rect 9624 12914 9873 12936
rect 9624 12883 9661 12914
rect 9837 12912 9873 12914
rect 9837 12883 9874 12912
rect 9076 12874 9111 12875
rect 9053 12869 9111 12874
rect 9053 12849 9056 12869
rect 9076 12855 9111 12869
rect 9131 12855 9140 12875
rect 9076 12847 9140 12855
rect 9102 12846 9140 12847
rect 9103 12845 9140 12846
rect 9206 12879 9242 12880
rect 9314 12879 9350 12880
rect 9206 12871 9350 12879
rect 9206 12851 9214 12871
rect 9234 12851 9322 12871
rect 9342 12851 9350 12871
rect 9206 12845 9350 12851
rect 9416 12875 9454 12883
rect 9522 12879 9558 12880
rect 9416 12855 9425 12875
rect 9445 12855 9454 12875
rect 9416 12846 9454 12855
rect 9473 12872 9558 12879
rect 9473 12852 9480 12872
rect 9501 12871 9558 12872
rect 9501 12852 9530 12871
rect 9473 12851 9530 12852
rect 9550 12851 9558 12871
rect 9416 12845 9453 12846
rect 9473 12845 9558 12851
rect 9624 12875 9662 12883
rect 9735 12879 9771 12880
rect 9624 12855 9633 12875
rect 9653 12855 9662 12875
rect 9624 12846 9662 12855
rect 9686 12871 9771 12879
rect 9686 12851 9743 12871
rect 9763 12851 9771 12871
rect 9624 12845 9661 12846
rect 9686 12845 9771 12851
rect 9837 12875 9875 12883
rect 9837 12855 9846 12875
rect 9866 12855 9875 12875
rect 9930 12865 9995 13017
rect 10148 12991 10203 13101
rect 11187 13063 11246 13101
rect 12099 13098 12107 13133
rect 12132 13098 12151 13133
rect 12176 13125 12198 13136
rect 13149 13137 14488 13144
rect 13149 13134 13201 13137
rect 12176 13124 13043 13125
rect 12176 13098 13044 13124
rect 12099 13088 13044 13098
rect 12099 13086 12198 13088
rect 11187 13045 11209 13063
rect 11227 13045 11246 13063
rect 11187 13023 11246 13045
rect 11454 13059 11986 13064
rect 11454 13039 12340 13059
rect 12360 13039 12363 13059
rect 12999 13055 13044 13088
rect 13149 13099 13157 13134
rect 13182 13099 13201 13134
rect 13226 13099 14488 13137
rect 13149 13090 14488 13099
rect 13149 13087 13238 13090
rect 13777 13088 14488 13090
rect 11454 13035 12363 13039
rect 9837 12846 9875 12855
rect 9928 12858 9995 12865
rect 9837 12845 9874 12846
rect 9260 12824 9296 12845
rect 9686 12824 9717 12845
rect 9928 12837 9945 12858
rect 9981 12837 9995 12858
rect 10147 12878 10203 12991
rect 11454 12988 11497 13035
rect 11947 13034 12363 13035
rect 12995 13035 13388 13055
rect 13408 13035 13411 13055
rect 11947 13033 12288 13034
rect 11604 13002 11714 13016
rect 11604 12999 11647 13002
rect 11604 12994 11608 12999
rect 11442 12987 11497 12988
rect 10147 12860 10166 12878
rect 10184 12860 10203 12878
rect 10147 12840 10203 12860
rect 11186 12964 11497 12987
rect 11186 12946 11211 12964
rect 11229 12952 11497 12964
rect 11526 12972 11608 12994
rect 11637 12972 11647 12999
rect 11675 12975 11682 13002
rect 11711 12994 11714 13002
rect 11711 12975 11776 12994
rect 11675 12972 11776 12975
rect 11526 12970 11776 12972
rect 11229 12946 11251 12952
rect 9928 12824 9995 12837
rect 9093 12820 9193 12824
rect 9093 12816 9155 12820
rect 9093 12790 9100 12816
rect 9126 12794 9155 12816
rect 9181 12794 9193 12820
rect 9126 12790 9193 12794
rect 9093 12787 9193 12790
rect 9261 12787 9296 12824
rect 9358 12821 9717 12824
rect 9358 12816 9580 12821
rect 9358 12792 9371 12816
rect 9395 12797 9580 12816
rect 9604 12797 9717 12821
rect 9395 12792 9717 12797
rect 9358 12788 9717 12792
rect 9784 12818 9995 12824
rect 9784 12816 9945 12818
rect 9784 12796 9795 12816
rect 9815 12796 9945 12816
rect 9784 12789 9945 12796
rect 9784 12788 9825 12789
rect 9260 12762 9296 12787
rect 9108 12735 9145 12736
rect 9204 12735 9241 12736
rect 9260 12735 9267 12762
rect 9008 12726 9146 12735
rect 9008 12706 9117 12726
rect 9137 12706 9146 12726
rect 9008 12699 9146 12706
rect 9204 12732 9267 12735
rect 9288 12735 9296 12762
rect 9315 12735 9352 12736
rect 9288 12732 9352 12735
rect 9204 12726 9352 12732
rect 9204 12706 9213 12726
rect 9233 12706 9323 12726
rect 9343 12706 9352 12726
rect 9008 12697 9104 12699
rect 9204 12696 9352 12706
rect 9411 12726 9448 12736
rect 9523 12735 9560 12736
rect 9504 12733 9560 12735
rect 9411 12706 9419 12726
rect 9439 12706 9448 12726
rect 9260 12695 9296 12696
rect 9108 12564 9145 12565
rect 9411 12564 9448 12706
rect 9473 12726 9560 12733
rect 9473 12723 9531 12726
rect 9473 12703 9478 12723
rect 9499 12706 9531 12723
rect 9551 12706 9560 12726
rect 9499 12703 9560 12706
rect 9473 12696 9560 12703
rect 9619 12726 9656 12736
rect 9619 12706 9627 12726
rect 9647 12706 9656 12726
rect 9473 12695 9504 12696
rect 9619 12627 9656 12706
rect 9686 12735 9717 12788
rect 9930 12781 9945 12789
rect 9985 12781 9995 12818
rect 11186 12807 11251 12946
rect 11526 12891 11563 12970
rect 11604 12957 11714 12970
rect 11678 12901 11709 12902
rect 11526 12871 11535 12891
rect 11555 12871 11563 12891
rect 9930 12772 9995 12781
rect 10143 12779 10208 12800
rect 10143 12761 10168 12779
rect 10186 12761 10208 12779
rect 11186 12789 11209 12807
rect 11227 12789 11251 12807
rect 11186 12772 11251 12789
rect 11406 12853 11474 12866
rect 11526 12861 11563 12871
rect 11622 12891 11709 12901
rect 11622 12871 11631 12891
rect 11651 12871 11709 12891
rect 11622 12862 11709 12871
rect 11622 12861 11659 12862
rect 11406 12811 11413 12853
rect 11462 12811 11474 12853
rect 11406 12808 11474 12811
rect 11678 12809 11709 12862
rect 11739 12891 11776 12970
rect 11891 12901 11922 12902
rect 11739 12871 11748 12891
rect 11768 12871 11776 12891
rect 11739 12861 11776 12871
rect 11835 12894 11922 12901
rect 11835 12891 11896 12894
rect 11835 12871 11844 12891
rect 11864 12874 11896 12891
rect 11917 12874 11922 12894
rect 11864 12871 11922 12874
rect 11835 12864 11922 12871
rect 11947 12891 11984 13033
rect 12250 13032 12287 13033
rect 12995 13030 13411 13035
rect 12995 13029 13336 13030
rect 12652 12998 12762 13012
rect 12652 12995 12695 12998
rect 12652 12990 12656 12995
rect 12574 12968 12656 12990
rect 12685 12968 12695 12995
rect 12723 12971 12730 12998
rect 12759 12990 12762 12998
rect 12759 12971 12824 12990
rect 12723 12968 12824 12971
rect 12574 12966 12824 12968
rect 12099 12901 12135 12902
rect 11947 12871 11956 12891
rect 11976 12871 11984 12891
rect 11835 12862 11891 12864
rect 11835 12861 11872 12862
rect 11947 12861 11984 12871
rect 12043 12891 12191 12901
rect 12291 12898 12387 12900
rect 12043 12871 12052 12891
rect 12072 12871 12162 12891
rect 12182 12871 12191 12891
rect 12043 12865 12191 12871
rect 12043 12862 12107 12865
rect 12043 12861 12080 12862
rect 12099 12835 12107 12862
rect 12128 12862 12191 12865
rect 12249 12891 12387 12898
rect 12249 12871 12258 12891
rect 12278 12871 12387 12891
rect 12249 12862 12387 12871
rect 12574 12887 12611 12966
rect 12652 12953 12762 12966
rect 12726 12897 12757 12898
rect 12574 12867 12583 12887
rect 12603 12867 12611 12887
rect 12128 12835 12135 12862
rect 12154 12861 12191 12862
rect 12250 12861 12287 12862
rect 12099 12810 12135 12835
rect 11570 12808 11611 12809
rect 11406 12801 11611 12808
rect 11406 12790 11580 12801
rect 9736 12735 9773 12736
rect 9686 12726 9773 12735
rect 9686 12706 9744 12726
rect 9764 12706 9773 12726
rect 9686 12696 9773 12706
rect 9832 12726 9869 12736
rect 9832 12706 9840 12726
rect 9860 12706 9869 12726
rect 9686 12695 9717 12696
rect 9681 12627 9791 12640
rect 9832 12627 9869 12706
rect 10143 12685 10208 12761
rect 11406 12757 11414 12790
rect 11407 12748 11414 12757
rect 11463 12781 11580 12790
rect 11600 12781 11611 12801
rect 11463 12773 11611 12781
rect 11678 12805 12037 12809
rect 11678 12800 12000 12805
rect 11678 12776 11791 12800
rect 11815 12781 12000 12800
rect 12024 12781 12037 12805
rect 11815 12776 12037 12781
rect 11678 12773 12037 12776
rect 12099 12773 12134 12810
rect 12202 12807 12302 12810
rect 12202 12803 12269 12807
rect 12202 12777 12214 12803
rect 12240 12781 12269 12803
rect 12295 12781 12302 12807
rect 12240 12777 12302 12781
rect 12202 12773 12302 12777
rect 11463 12757 11474 12773
rect 11463 12748 11471 12757
rect 11678 12752 11709 12773
rect 12099 12752 12135 12773
rect 11521 12751 11558 12752
rect 11186 12708 11251 12727
rect 11186 12690 11211 12708
rect 11229 12690 11251 12708
rect 9619 12625 9869 12627
rect 9619 12622 9720 12625
rect 9619 12603 9684 12622
rect 9681 12595 9684 12603
rect 9713 12595 9720 12622
rect 9748 12598 9758 12625
rect 9787 12603 9869 12625
rect 9892 12650 10209 12685
rect 9787 12598 9791 12603
rect 9748 12595 9791 12598
rect 9681 12581 9791 12595
rect 9107 12563 9448 12564
rect 9032 12561 9448 12563
rect 9892 12561 9932 12650
rect 10143 12623 10208 12650
rect 10143 12605 10166 12623
rect 10184 12605 10208 12623
rect 10143 12585 10208 12605
rect 9029 12558 9932 12561
rect 9029 12538 9035 12558
rect 9055 12538 9932 12558
rect 9029 12534 9932 12538
rect 9892 12531 9932 12534
rect 10144 12524 10209 12545
rect 8362 12516 9023 12517
rect 8362 12509 9296 12516
rect 8362 12508 9268 12509
rect 8362 12488 9213 12508
rect 9245 12489 9268 12508
rect 9293 12489 9296 12509
rect 9245 12488 9296 12489
rect 8362 12481 9296 12488
rect 7961 12439 8129 12440
rect 8364 12439 8403 12481
rect 9192 12479 9296 12481
rect 9261 12477 9296 12479
rect 10144 12506 10168 12524
rect 10186 12506 10209 12524
rect 10144 12459 10209 12506
rect 7961 12413 8405 12439
rect 7961 12411 8129 12413
rect 7961 12060 7988 12411
rect 8364 12407 8405 12413
rect 8028 12200 8092 12212
rect 8368 12208 8405 12407
rect 8867 12434 8939 12451
rect 8867 12395 8875 12434
rect 8920 12395 8939 12434
rect 8633 12297 8744 12312
rect 8633 12295 8675 12297
rect 8633 12275 8640 12295
rect 8659 12275 8675 12295
rect 8633 12267 8675 12275
rect 8703 12295 8744 12297
rect 8703 12275 8717 12295
rect 8736 12275 8744 12295
rect 8703 12267 8744 12275
rect 8633 12261 8744 12267
rect 8576 12239 8825 12261
rect 8576 12208 8613 12239
rect 8789 12237 8825 12239
rect 8789 12208 8826 12237
rect 8028 12199 8063 12200
rect 8005 12194 8063 12199
rect 8005 12174 8008 12194
rect 8028 12180 8063 12194
rect 8083 12180 8092 12200
rect 8028 12172 8092 12180
rect 8054 12171 8092 12172
rect 8055 12170 8092 12171
rect 8158 12204 8194 12205
rect 8266 12204 8302 12205
rect 8158 12196 8302 12204
rect 8158 12176 8166 12196
rect 8186 12176 8274 12196
rect 8294 12176 8302 12196
rect 8158 12170 8302 12176
rect 8368 12200 8406 12208
rect 8474 12204 8510 12205
rect 8368 12180 8377 12200
rect 8397 12180 8406 12200
rect 8368 12171 8406 12180
rect 8425 12197 8510 12204
rect 8425 12177 8432 12197
rect 8453 12196 8510 12197
rect 8453 12177 8482 12196
rect 8425 12176 8482 12177
rect 8502 12176 8510 12196
rect 8368 12170 8405 12171
rect 8425 12170 8510 12176
rect 8576 12200 8614 12208
rect 8687 12204 8723 12205
rect 8576 12180 8585 12200
rect 8605 12180 8614 12200
rect 8576 12171 8614 12180
rect 8638 12196 8723 12204
rect 8638 12176 8695 12196
rect 8715 12176 8723 12196
rect 8576 12170 8613 12171
rect 8638 12170 8723 12176
rect 8789 12200 8827 12208
rect 8789 12180 8798 12200
rect 8818 12180 8827 12200
rect 8789 12171 8827 12180
rect 8867 12185 8939 12395
rect 9009 12429 10209 12459
rect 9009 12428 9453 12429
rect 9009 12426 9177 12428
rect 8867 12171 8950 12185
rect 8789 12170 8826 12171
rect 8212 12149 8248 12170
rect 8638 12149 8669 12170
rect 8867 12149 8884 12171
rect 8045 12145 8145 12149
rect 8045 12141 8107 12145
rect 8045 12115 8052 12141
rect 8078 12119 8107 12141
rect 8133 12119 8145 12145
rect 8078 12115 8145 12119
rect 8045 12112 8145 12115
rect 8213 12112 8248 12149
rect 8310 12146 8669 12149
rect 8310 12141 8532 12146
rect 8310 12117 8323 12141
rect 8347 12122 8532 12141
rect 8556 12122 8669 12146
rect 8347 12117 8669 12122
rect 8310 12113 8669 12117
rect 8736 12141 8884 12149
rect 8736 12121 8747 12141
rect 8767 12138 8884 12141
rect 8937 12138 8950 12171
rect 8767 12121 8950 12138
rect 8736 12114 8950 12121
rect 8736 12113 8777 12114
rect 8867 12113 8950 12114
rect 8212 12087 8248 12112
rect 8060 12060 8097 12061
rect 8156 12060 8193 12061
rect 8212 12060 8219 12087
rect 7960 12051 8098 12060
rect 7960 12031 8069 12051
rect 8089 12031 8098 12051
rect 7960 12024 8098 12031
rect 8156 12057 8219 12060
rect 8240 12060 8248 12087
rect 8267 12060 8304 12061
rect 8240 12057 8304 12060
rect 8156 12051 8304 12057
rect 8156 12031 8165 12051
rect 8185 12031 8275 12051
rect 8295 12031 8304 12051
rect 7960 12022 8056 12024
rect 8156 12021 8304 12031
rect 8363 12051 8400 12061
rect 8475 12060 8512 12061
rect 8456 12058 8512 12060
rect 8363 12031 8371 12051
rect 8391 12031 8400 12051
rect 8212 12020 8248 12021
rect 8060 11889 8097 11890
rect 8363 11889 8400 12031
rect 8425 12051 8512 12058
rect 8425 12048 8483 12051
rect 8425 12028 8430 12048
rect 8451 12031 8483 12048
rect 8503 12031 8512 12051
rect 8451 12028 8512 12031
rect 8425 12021 8512 12028
rect 8571 12051 8608 12061
rect 8571 12031 8579 12051
rect 8599 12031 8608 12051
rect 8425 12020 8456 12021
rect 8571 11952 8608 12031
rect 8638 12060 8669 12113
rect 8875 12080 8889 12113
rect 8942 12080 8950 12113
rect 8875 12074 8950 12080
rect 8875 12069 8945 12074
rect 8688 12060 8725 12061
rect 8638 12051 8725 12060
rect 8638 12031 8696 12051
rect 8716 12031 8725 12051
rect 8638 12021 8725 12031
rect 8784 12051 8821 12061
rect 9009 12056 9036 12426
rect 9076 12196 9140 12208
rect 9416 12204 9453 12428
rect 9924 12409 9988 12411
rect 9920 12397 9988 12409
rect 9920 12364 9931 12397
rect 9971 12364 9988 12397
rect 9920 12354 9988 12364
rect 9681 12293 9792 12308
rect 9681 12291 9723 12293
rect 9681 12271 9688 12291
rect 9707 12271 9723 12291
rect 9681 12263 9723 12271
rect 9751 12291 9792 12293
rect 9751 12271 9765 12291
rect 9784 12271 9792 12291
rect 9751 12263 9792 12271
rect 9681 12257 9792 12263
rect 9624 12235 9873 12257
rect 9624 12204 9661 12235
rect 9837 12233 9873 12235
rect 9837 12204 9874 12233
rect 9076 12195 9111 12196
rect 9053 12190 9111 12195
rect 9053 12170 9056 12190
rect 9076 12176 9111 12190
rect 9131 12176 9140 12196
rect 9076 12168 9140 12176
rect 9102 12167 9140 12168
rect 9103 12166 9140 12167
rect 9206 12200 9242 12201
rect 9314 12200 9350 12201
rect 9206 12192 9350 12200
rect 9206 12172 9214 12192
rect 9234 12172 9322 12192
rect 9342 12172 9350 12192
rect 9206 12166 9350 12172
rect 9416 12196 9454 12204
rect 9522 12200 9558 12201
rect 9416 12176 9425 12196
rect 9445 12176 9454 12196
rect 9416 12167 9454 12176
rect 9473 12193 9558 12200
rect 9473 12173 9480 12193
rect 9501 12192 9558 12193
rect 9501 12173 9530 12192
rect 9473 12172 9530 12173
rect 9550 12172 9558 12192
rect 9416 12166 9453 12167
rect 9473 12166 9558 12172
rect 9624 12196 9662 12204
rect 9735 12200 9771 12201
rect 9624 12176 9633 12196
rect 9653 12176 9662 12196
rect 9624 12167 9662 12176
rect 9686 12192 9771 12200
rect 9686 12172 9743 12192
rect 9763 12172 9771 12192
rect 9624 12166 9661 12167
rect 9686 12166 9771 12172
rect 9837 12196 9875 12204
rect 9837 12176 9846 12196
rect 9866 12176 9875 12196
rect 9837 12167 9875 12176
rect 9924 12170 9988 12354
rect 10144 12228 10209 12429
rect 11186 12489 11251 12690
rect 11407 12564 11471 12748
rect 11520 12742 11558 12751
rect 11520 12722 11529 12742
rect 11549 12722 11558 12742
rect 11520 12714 11558 12722
rect 11624 12746 11709 12752
rect 11734 12751 11771 12752
rect 11624 12726 11632 12746
rect 11652 12726 11709 12746
rect 11624 12718 11709 12726
rect 11733 12742 11771 12751
rect 11733 12722 11742 12742
rect 11762 12722 11771 12742
rect 11624 12717 11660 12718
rect 11733 12714 11771 12722
rect 11837 12746 11922 12752
rect 11942 12751 11979 12752
rect 11837 12726 11845 12746
rect 11865 12745 11922 12746
rect 11865 12726 11894 12745
rect 11837 12725 11894 12726
rect 11915 12725 11922 12745
rect 11837 12718 11922 12725
rect 11941 12742 11979 12751
rect 11941 12722 11950 12742
rect 11970 12722 11979 12742
rect 11837 12717 11873 12718
rect 11941 12714 11979 12722
rect 12045 12746 12189 12752
rect 12045 12726 12053 12746
rect 12073 12726 12161 12746
rect 12181 12726 12189 12746
rect 12045 12718 12189 12726
rect 12045 12717 12081 12718
rect 12153 12717 12189 12718
rect 12255 12751 12292 12752
rect 12255 12750 12293 12751
rect 12255 12742 12319 12750
rect 12255 12722 12264 12742
rect 12284 12728 12319 12742
rect 12339 12728 12342 12748
rect 12284 12723 12342 12728
rect 12284 12722 12319 12723
rect 11521 12685 11558 12714
rect 11522 12683 11558 12685
rect 11734 12683 11771 12714
rect 11522 12661 11771 12683
rect 11603 12655 11714 12661
rect 11603 12647 11644 12655
rect 11603 12627 11611 12647
rect 11630 12627 11644 12647
rect 11603 12625 11644 12627
rect 11672 12647 11714 12655
rect 11672 12627 11688 12647
rect 11707 12627 11714 12647
rect 11672 12625 11714 12627
rect 11603 12610 11714 12625
rect 11407 12554 11475 12564
rect 11407 12521 11424 12554
rect 11464 12521 11475 12554
rect 11407 12509 11475 12521
rect 11407 12507 11471 12509
rect 11942 12490 11979 12714
rect 12255 12710 12319 12722
rect 12359 12492 12386 12862
rect 12574 12857 12611 12867
rect 12670 12887 12757 12897
rect 12670 12867 12679 12887
rect 12699 12867 12757 12887
rect 12670 12858 12757 12867
rect 12670 12857 12707 12858
rect 12450 12844 12520 12849
rect 12445 12838 12520 12844
rect 12445 12805 12453 12838
rect 12506 12805 12520 12838
rect 12726 12805 12757 12858
rect 12787 12887 12824 12966
rect 12939 12897 12970 12898
rect 12787 12867 12796 12887
rect 12816 12867 12824 12887
rect 12787 12857 12824 12867
rect 12883 12890 12970 12897
rect 12883 12887 12944 12890
rect 12883 12867 12892 12887
rect 12912 12870 12944 12887
rect 12965 12870 12970 12890
rect 12912 12867 12970 12870
rect 12883 12860 12970 12867
rect 12995 12887 13032 13029
rect 13298 13028 13335 13029
rect 13147 12897 13183 12898
rect 12995 12867 13004 12887
rect 13024 12867 13032 12887
rect 12883 12858 12939 12860
rect 12883 12857 12920 12858
rect 12995 12857 13032 12867
rect 13091 12887 13239 12897
rect 13339 12894 13435 12896
rect 13091 12867 13100 12887
rect 13120 12867 13210 12887
rect 13230 12867 13239 12887
rect 13091 12861 13239 12867
rect 13091 12858 13155 12861
rect 13091 12857 13128 12858
rect 13147 12831 13155 12858
rect 13176 12858 13239 12861
rect 13297 12887 13435 12894
rect 13297 12867 13306 12887
rect 13326 12867 13435 12887
rect 13297 12858 13435 12867
rect 13176 12831 13183 12858
rect 13202 12857 13239 12858
rect 13298 12857 13335 12858
rect 13147 12806 13183 12831
rect 12445 12804 12528 12805
rect 12618 12804 12659 12805
rect 12445 12797 12659 12804
rect 12445 12780 12628 12797
rect 12445 12747 12458 12780
rect 12511 12777 12628 12780
rect 12648 12777 12659 12797
rect 12511 12769 12659 12777
rect 12726 12801 13085 12805
rect 12726 12796 13048 12801
rect 12726 12772 12839 12796
rect 12863 12777 13048 12796
rect 13072 12777 13085 12801
rect 12863 12772 13085 12777
rect 12726 12769 13085 12772
rect 13147 12769 13182 12806
rect 13250 12803 13350 12806
rect 13250 12799 13317 12803
rect 13250 12773 13262 12799
rect 13288 12777 13317 12799
rect 13343 12777 13350 12803
rect 13288 12773 13350 12777
rect 13250 12769 13350 12773
rect 12511 12747 12528 12769
rect 12726 12748 12757 12769
rect 13147 12748 13183 12769
rect 12569 12747 12606 12748
rect 12445 12733 12528 12747
rect 12218 12490 12386 12492
rect 11942 12489 12386 12490
rect 11186 12459 12386 12489
rect 12456 12523 12528 12733
rect 12568 12738 12606 12747
rect 12568 12718 12577 12738
rect 12597 12718 12606 12738
rect 12568 12710 12606 12718
rect 12672 12742 12757 12748
rect 12782 12747 12819 12748
rect 12672 12722 12680 12742
rect 12700 12722 12757 12742
rect 12672 12714 12757 12722
rect 12781 12738 12819 12747
rect 12781 12718 12790 12738
rect 12810 12718 12819 12738
rect 12672 12713 12708 12714
rect 12781 12710 12819 12718
rect 12885 12742 12970 12748
rect 12990 12747 13027 12748
rect 12885 12722 12893 12742
rect 12913 12741 12970 12742
rect 12913 12722 12942 12741
rect 12885 12721 12942 12722
rect 12963 12721 12970 12741
rect 12885 12714 12970 12721
rect 12989 12738 13027 12747
rect 12989 12718 12998 12738
rect 13018 12718 13027 12738
rect 12885 12713 12921 12714
rect 12989 12710 13027 12718
rect 13093 12742 13237 12748
rect 13093 12722 13101 12742
rect 13121 12722 13209 12742
rect 13229 12722 13237 12742
rect 13093 12714 13237 12722
rect 13093 12713 13129 12714
rect 13201 12713 13237 12714
rect 13303 12747 13340 12748
rect 13303 12746 13341 12747
rect 13303 12738 13367 12746
rect 13303 12718 13312 12738
rect 13332 12724 13367 12738
rect 13387 12724 13390 12744
rect 13332 12719 13390 12724
rect 13332 12718 13367 12719
rect 12569 12681 12606 12710
rect 12570 12679 12606 12681
rect 12782 12679 12819 12710
rect 12570 12657 12819 12679
rect 12651 12651 12762 12657
rect 12651 12643 12692 12651
rect 12651 12623 12659 12643
rect 12678 12623 12692 12643
rect 12651 12621 12692 12623
rect 12720 12643 12762 12651
rect 12720 12623 12736 12643
rect 12755 12623 12762 12643
rect 12720 12621 12762 12623
rect 12651 12606 12762 12621
rect 12456 12484 12475 12523
rect 12520 12484 12528 12523
rect 12456 12467 12528 12484
rect 12990 12511 13027 12710
rect 13303 12706 13367 12718
rect 12990 12505 13031 12511
rect 13407 12507 13434 12858
rect 13729 12845 13824 12871
rect 13565 12823 13629 12842
rect 13565 12784 13578 12823
rect 13612 12784 13629 12823
rect 13565 12765 13629 12784
rect 13266 12505 13434 12507
rect 12990 12479 13434 12505
rect 11186 12412 11251 12459
rect 11186 12394 11209 12412
rect 11227 12394 11251 12412
rect 12099 12439 12134 12441
rect 12099 12437 12203 12439
rect 12992 12437 13031 12479
rect 13266 12478 13434 12479
rect 12099 12430 13033 12437
rect 12099 12429 12150 12430
rect 12099 12409 12102 12429
rect 12127 12410 12150 12429
rect 12182 12410 13033 12430
rect 12127 12409 13033 12410
rect 12099 12402 13033 12409
rect 12372 12401 13033 12402
rect 11186 12373 11251 12394
rect 11463 12384 11503 12387
rect 11463 12380 12366 12384
rect 11463 12360 12340 12380
rect 12360 12360 12366 12380
rect 11463 12357 12366 12360
rect 11187 12313 11252 12333
rect 11187 12295 11211 12313
rect 11229 12295 11252 12313
rect 11187 12268 11252 12295
rect 11463 12268 11503 12357
rect 11947 12355 12363 12357
rect 11947 12354 12288 12355
rect 11604 12323 11714 12337
rect 11604 12320 11647 12323
rect 11604 12315 11608 12320
rect 11186 12233 11503 12268
rect 11526 12293 11608 12315
rect 11637 12293 11647 12320
rect 11675 12296 11682 12323
rect 11711 12315 11714 12323
rect 11711 12296 11776 12315
rect 11675 12293 11776 12296
rect 11526 12291 11776 12293
rect 10144 12210 10166 12228
rect 10184 12210 10209 12228
rect 10144 12191 10209 12210
rect 9837 12166 9874 12167
rect 9260 12145 9296 12166
rect 9686 12145 9717 12166
rect 9924 12161 9932 12170
rect 9921 12145 9932 12161
rect 9093 12141 9193 12145
rect 9093 12137 9155 12141
rect 9093 12111 9100 12137
rect 9126 12115 9155 12137
rect 9181 12115 9193 12141
rect 9126 12111 9193 12115
rect 9093 12108 9193 12111
rect 9261 12108 9296 12145
rect 9358 12142 9717 12145
rect 9358 12137 9580 12142
rect 9358 12113 9371 12137
rect 9395 12118 9580 12137
rect 9604 12118 9717 12142
rect 9395 12113 9717 12118
rect 9358 12109 9717 12113
rect 9784 12137 9932 12145
rect 9784 12117 9795 12137
rect 9815 12128 9932 12137
rect 9981 12161 9988 12170
rect 9981 12128 9989 12161
rect 11187 12157 11252 12233
rect 11526 12212 11563 12291
rect 11604 12278 11714 12291
rect 11678 12222 11709 12223
rect 11526 12192 11535 12212
rect 11555 12192 11563 12212
rect 11526 12182 11563 12192
rect 11622 12212 11709 12222
rect 11622 12192 11631 12212
rect 11651 12192 11709 12212
rect 11622 12183 11709 12192
rect 11622 12182 11659 12183
rect 9815 12117 9989 12128
rect 9784 12110 9989 12117
rect 9784 12109 9825 12110
rect 9260 12083 9296 12108
rect 9108 12056 9145 12057
rect 9204 12056 9241 12057
rect 9260 12056 9267 12083
rect 8784 12031 8792 12051
rect 8812 12031 8821 12051
rect 8638 12020 8669 12021
rect 8633 11952 8743 11965
rect 8784 11952 8821 12031
rect 9008 12047 9146 12056
rect 9008 12027 9117 12047
rect 9137 12027 9146 12047
rect 9008 12020 9146 12027
rect 9204 12053 9267 12056
rect 9288 12056 9296 12083
rect 9315 12056 9352 12057
rect 9288 12053 9352 12056
rect 9204 12047 9352 12053
rect 9204 12027 9213 12047
rect 9233 12027 9323 12047
rect 9343 12027 9352 12047
rect 9008 12018 9104 12020
rect 9204 12017 9352 12027
rect 9411 12047 9448 12057
rect 9523 12056 9560 12057
rect 9504 12054 9560 12056
rect 9411 12027 9419 12047
rect 9439 12027 9448 12047
rect 9260 12016 9296 12017
rect 8571 11950 8821 11952
rect 8571 11947 8672 11950
rect 8571 11928 8636 11947
rect 8633 11920 8636 11928
rect 8665 11920 8672 11947
rect 8700 11923 8710 11950
rect 8739 11928 8821 11950
rect 8739 11923 8743 11928
rect 8700 11920 8743 11923
rect 8633 11906 8743 11920
rect 8059 11888 8400 11889
rect 7984 11883 8400 11888
rect 9108 11885 9145 11886
rect 9411 11885 9448 12027
rect 9473 12047 9560 12054
rect 9473 12044 9531 12047
rect 9473 12024 9478 12044
rect 9499 12027 9531 12044
rect 9551 12027 9560 12047
rect 9499 12024 9560 12027
rect 9473 12017 9560 12024
rect 9619 12047 9656 12057
rect 9619 12027 9627 12047
rect 9647 12027 9656 12047
rect 9473 12016 9504 12017
rect 9619 11948 9656 12027
rect 9686 12056 9717 12109
rect 9921 12107 9989 12110
rect 9921 12065 9933 12107
rect 9982 12065 9989 12107
rect 9736 12056 9773 12057
rect 9686 12047 9773 12056
rect 9686 12027 9744 12047
rect 9764 12027 9773 12047
rect 9686 12017 9773 12027
rect 9832 12047 9869 12057
rect 9921 12052 9989 12065
rect 10144 12129 10209 12146
rect 10144 12111 10168 12129
rect 10186 12111 10209 12129
rect 11187 12139 11209 12157
rect 11227 12139 11252 12157
rect 11187 12118 11252 12139
rect 11400 12137 11465 12146
rect 9832 12027 9840 12047
rect 9860 12027 9869 12047
rect 9686 12016 9717 12017
rect 9681 11948 9791 11961
rect 9832 11948 9869 12027
rect 10144 11972 10209 12111
rect 11400 12100 11410 12137
rect 11450 12129 11465 12137
rect 11678 12130 11709 12183
rect 11739 12212 11776 12291
rect 11891 12222 11922 12223
rect 11739 12192 11748 12212
rect 11768 12192 11776 12212
rect 11739 12182 11776 12192
rect 11835 12215 11922 12222
rect 11835 12212 11896 12215
rect 11835 12192 11844 12212
rect 11864 12195 11896 12212
rect 11917 12195 11922 12215
rect 11864 12192 11922 12195
rect 11835 12185 11922 12192
rect 11947 12212 11984 12354
rect 12250 12353 12287 12354
rect 13567 12294 13629 12765
rect 13729 12804 13755 12845
rect 13791 12804 13824 12845
rect 13729 12508 13824 12804
rect 13729 12464 13744 12508
rect 13804 12464 13824 12508
rect 13729 12444 13824 12464
rect 14441 12375 14484 13088
rect 15024 13030 15170 13041
rect 15024 13014 16406 13030
rect 15024 13009 16433 13014
rect 15024 13003 15116 13009
rect 15024 12906 15056 13003
rect 15094 12912 15116 13003
rect 15154 12912 16433 13009
rect 19583 12914 19653 13167
rect 20122 13164 20163 13166
rect 20394 13164 20498 13166
rect 19715 13162 20909 13164
rect 19715 13129 20911 13162
rect 19715 13115 19743 13129
rect 19717 12984 19743 13115
rect 20122 13126 20911 13129
rect 15094 12906 16433 12912
rect 15024 12879 16433 12906
rect 16303 12804 16433 12879
rect 19575 12863 19655 12914
rect 19575 12837 19591 12863
rect 19631 12837 19655 12863
rect 19575 12818 19655 12837
rect 14441 12355 14835 12375
rect 14855 12355 14858 12375
rect 14442 12350 14858 12355
rect 14442 12349 14783 12350
rect 14099 12318 14209 12332
rect 14099 12315 14142 12318
rect 14099 12310 14103 12315
rect 13562 12242 13637 12294
rect 14021 12288 14103 12310
rect 14132 12288 14142 12315
rect 14170 12291 14177 12318
rect 14206 12310 14209 12318
rect 14206 12291 14271 12310
rect 14170 12288 14271 12291
rect 14021 12286 14271 12288
rect 13931 12242 13977 12243
rect 12099 12222 12135 12223
rect 11947 12192 11956 12212
rect 11976 12192 11984 12212
rect 11835 12183 11891 12185
rect 11835 12182 11872 12183
rect 11947 12182 11984 12192
rect 12043 12212 12191 12222
rect 12291 12219 12387 12221
rect 12043 12192 12052 12212
rect 12072 12192 12162 12212
rect 12182 12192 12191 12212
rect 12043 12186 12191 12192
rect 12043 12183 12107 12186
rect 12043 12182 12080 12183
rect 12099 12156 12107 12183
rect 12128 12183 12191 12186
rect 12249 12212 12387 12219
rect 12249 12192 12258 12212
rect 12278 12192 12387 12212
rect 12249 12183 12387 12192
rect 13562 12207 13977 12242
rect 12128 12156 12135 12183
rect 12154 12182 12191 12183
rect 12250 12182 12287 12183
rect 12099 12131 12135 12156
rect 11570 12129 11611 12130
rect 11450 12122 11611 12129
rect 11450 12102 11580 12122
rect 11600 12102 11611 12122
rect 11450 12100 11611 12102
rect 11400 12094 11611 12100
rect 11678 12126 12037 12130
rect 11678 12121 12000 12126
rect 11678 12097 11791 12121
rect 11815 12102 12000 12121
rect 12024 12102 12037 12126
rect 11815 12097 12037 12102
rect 11678 12094 12037 12097
rect 12099 12094 12134 12131
rect 12202 12128 12302 12131
rect 12202 12124 12269 12128
rect 12202 12098 12214 12124
rect 12240 12102 12269 12124
rect 12295 12102 12302 12128
rect 12240 12098 12302 12102
rect 12202 12094 12302 12098
rect 11400 12081 11467 12094
rect 10144 11966 10166 11972
rect 9619 11946 9869 11948
rect 9619 11943 9720 11946
rect 9619 11924 9684 11943
rect 9681 11916 9684 11924
rect 9713 11916 9720 11943
rect 9748 11919 9758 11946
rect 9787 11924 9869 11946
rect 9898 11954 10166 11966
rect 10184 11954 10209 11972
rect 9898 11931 10209 11954
rect 11192 12058 11248 12078
rect 11192 12040 11211 12058
rect 11229 12040 11248 12058
rect 9898 11930 9953 11931
rect 9787 11919 9791 11924
rect 9748 11916 9791 11919
rect 9681 11902 9791 11916
rect 9107 11884 9448 11885
rect 7984 11863 7987 11883
rect 8007 11863 8400 11883
rect 9032 11883 9448 11884
rect 9898 11883 9941 11930
rect 11192 11927 11248 12040
rect 11400 12060 11414 12081
rect 11450 12060 11467 12081
rect 11678 12073 11709 12094
rect 12099 12073 12135 12094
rect 11521 12072 11558 12073
rect 11400 12053 11467 12060
rect 11520 12063 11558 12072
rect 9032 11879 9941 11883
rect 8351 11830 8396 11863
rect 9032 11859 9035 11879
rect 9055 11859 9941 11879
rect 9409 11854 9941 11859
rect 10149 11873 10208 11895
rect 10149 11855 10168 11873
rect 10186 11855 10208 11873
rect 9197 11830 9296 11832
rect 8351 11820 9296 11830
rect 6908 11800 6967 11810
rect 6908 11772 6921 11800
rect 6949 11772 6967 11800
rect 8351 11794 9219 11820
rect 8352 11793 9219 11794
rect 9197 11782 9219 11793
rect 9244 11785 9263 11820
rect 9288 11785 9296 11820
rect 9244 11782 9296 11785
rect 10149 11784 10208 11855
rect 11192 11789 11247 11927
rect 11400 11901 11465 12053
rect 11520 12043 11529 12063
rect 11549 12043 11558 12063
rect 11520 12035 11558 12043
rect 11624 12067 11709 12073
rect 11734 12072 11771 12073
rect 11624 12047 11632 12067
rect 11652 12047 11709 12067
rect 11624 12039 11709 12047
rect 11733 12063 11771 12072
rect 11733 12043 11742 12063
rect 11762 12043 11771 12063
rect 11624 12038 11660 12039
rect 11733 12035 11771 12043
rect 11837 12067 11922 12073
rect 11942 12072 11979 12073
rect 11837 12047 11845 12067
rect 11865 12066 11922 12067
rect 11865 12047 11894 12066
rect 11837 12046 11894 12047
rect 11915 12046 11922 12066
rect 11837 12039 11922 12046
rect 11941 12063 11979 12072
rect 11941 12043 11950 12063
rect 11970 12043 11979 12063
rect 11837 12038 11873 12039
rect 11941 12035 11979 12043
rect 12045 12067 12189 12073
rect 12045 12047 12053 12067
rect 12073 12047 12161 12067
rect 12181 12047 12189 12067
rect 12045 12039 12189 12047
rect 12045 12038 12081 12039
rect 12153 12038 12189 12039
rect 12255 12072 12292 12073
rect 12255 12071 12293 12072
rect 12255 12063 12319 12071
rect 12255 12043 12264 12063
rect 12284 12049 12319 12063
rect 12339 12049 12342 12069
rect 12284 12044 12342 12049
rect 12284 12043 12319 12044
rect 11521 12006 11558 12035
rect 11522 12004 11558 12006
rect 11734 12004 11771 12035
rect 11522 11982 11771 12004
rect 11603 11976 11714 11982
rect 11603 11968 11644 11976
rect 11603 11948 11611 11968
rect 11630 11948 11644 11968
rect 11603 11946 11644 11948
rect 11672 11968 11714 11976
rect 11672 11948 11688 11968
rect 11707 11948 11714 11968
rect 11672 11946 11714 11948
rect 11603 11933 11714 11946
rect 11942 11936 11979 12035
rect 12255 12031 12319 12043
rect 11393 11891 11514 11901
rect 11393 11889 11462 11891
rect 11393 11848 11406 11889
rect 11443 11850 11462 11889
rect 11499 11850 11514 11891
rect 11443 11848 11514 11850
rect 11393 11830 11514 11848
rect 11185 11786 11249 11789
rect 11605 11786 11709 11792
rect 11940 11786 11981 11936
rect 12359 11928 12386 12183
rect 12448 12173 12528 12184
rect 12448 12147 12465 12173
rect 12505 12147 12528 12173
rect 12448 12120 12528 12147
rect 12448 12094 12469 12120
rect 12509 12094 12528 12120
rect 12448 12075 12528 12094
rect 12448 12049 12472 12075
rect 12512 12049 12528 12075
rect 12448 11998 12528 12049
rect 9197 11774 9296 11782
rect 9223 11773 9295 11774
rect 6908 11723 6967 11772
rect 8877 11747 8944 11766
rect 8877 11726 8894 11747
rect 6514 11588 6682 11589
rect 6918 11588 6965 11723
rect 6514 11562 6965 11588
rect 6514 11560 6682 11562
rect 6514 11293 6541 11560
rect 6918 11556 6965 11562
rect 8875 11681 8894 11726
rect 8924 11726 8944 11747
rect 8924 11681 8945 11726
rect 9414 11723 9455 11725
rect 9686 11723 9790 11725
rect 10146 11723 10210 11784
rect 6581 11433 6645 11445
rect 6921 11441 6958 11556
rect 7186 11530 7297 11545
rect 7186 11528 7228 11530
rect 7186 11508 7193 11528
rect 7212 11508 7228 11528
rect 7186 11500 7228 11508
rect 7256 11528 7297 11530
rect 7256 11508 7270 11528
rect 7289 11508 7297 11528
rect 7256 11500 7297 11508
rect 7186 11494 7297 11500
rect 7129 11472 7378 11494
rect 8875 11473 8945 11681
rect 9007 11688 10210 11723
rect 9007 11674 9035 11688
rect 9009 11543 9035 11674
rect 9414 11685 10210 11688
rect 11185 11783 11981 11786
rect 12360 11797 12386 11928
rect 12360 11783 12388 11797
rect 11185 11748 12388 11783
rect 12450 11790 12520 11998
rect 13562 11923 13637 12207
rect 13931 12124 13977 12207
rect 14021 12207 14058 12286
rect 14099 12273 14209 12286
rect 14173 12217 14204 12218
rect 14021 12187 14030 12207
rect 14050 12187 14058 12207
rect 14021 12177 14058 12187
rect 14117 12207 14204 12217
rect 14117 12187 14126 12207
rect 14146 12187 14204 12207
rect 14117 12178 14204 12187
rect 14117 12177 14154 12178
rect 14173 12125 14204 12178
rect 14234 12207 14271 12286
rect 14386 12217 14417 12218
rect 14234 12187 14243 12207
rect 14263 12187 14271 12207
rect 14234 12177 14271 12187
rect 14330 12210 14417 12217
rect 14330 12207 14391 12210
rect 14330 12187 14339 12207
rect 14359 12190 14391 12207
rect 14412 12190 14417 12210
rect 14359 12187 14417 12190
rect 14330 12180 14417 12187
rect 14442 12207 14479 12349
rect 14745 12348 14782 12349
rect 14594 12217 14630 12218
rect 14442 12187 14451 12207
rect 14471 12187 14479 12207
rect 14330 12178 14386 12180
rect 14330 12177 14367 12178
rect 14442 12177 14479 12187
rect 14538 12207 14686 12217
rect 14786 12214 14882 12216
rect 14538 12187 14547 12207
rect 14567 12187 14657 12207
rect 14677 12187 14686 12207
rect 14538 12181 14686 12187
rect 14538 12178 14602 12181
rect 14538 12177 14575 12178
rect 14594 12151 14602 12178
rect 14623 12178 14686 12181
rect 14744 12207 14882 12214
rect 14744 12187 14753 12207
rect 14773 12187 14882 12207
rect 14744 12178 14882 12187
rect 14623 12151 14630 12178
rect 14649 12177 14686 12178
rect 14745 12177 14782 12178
rect 14594 12126 14630 12151
rect 14065 12124 14106 12125
rect 13931 12117 14106 12124
rect 13729 12091 13815 12110
rect 13729 12050 13744 12091
rect 13798 12050 13815 12091
rect 13931 12097 14075 12117
rect 14095 12097 14106 12117
rect 13931 12089 14106 12097
rect 14173 12121 14532 12125
rect 14173 12116 14495 12121
rect 14173 12092 14286 12116
rect 14310 12097 14495 12116
rect 14519 12097 14532 12121
rect 14310 12092 14532 12097
rect 14173 12089 14532 12092
rect 14594 12089 14629 12126
rect 14697 12123 14797 12126
rect 14697 12119 14764 12123
rect 14697 12093 14709 12119
rect 14735 12097 14764 12119
rect 14790 12097 14797 12123
rect 14735 12093 14797 12097
rect 14697 12089 14797 12093
rect 13931 12085 13977 12089
rect 14173 12068 14204 12089
rect 14594 12068 14630 12089
rect 14016 12067 14053 12068
rect 13729 12014 13815 12050
rect 14015 12058 14053 12067
rect 14015 12038 14024 12058
rect 14044 12038 14053 12058
rect 14015 12030 14053 12038
rect 14119 12062 14204 12068
rect 14229 12067 14266 12068
rect 14119 12042 14127 12062
rect 14147 12042 14204 12062
rect 14119 12034 14204 12042
rect 14228 12058 14266 12067
rect 14228 12038 14237 12058
rect 14257 12038 14266 12058
rect 14119 12033 14155 12034
rect 14228 12030 14266 12038
rect 14332 12062 14417 12068
rect 14437 12067 14474 12068
rect 14332 12042 14340 12062
rect 14360 12061 14417 12062
rect 14360 12042 14389 12061
rect 14332 12041 14389 12042
rect 14410 12041 14417 12061
rect 14332 12034 14417 12041
rect 14436 12058 14474 12067
rect 14436 12038 14445 12058
rect 14465 12038 14474 12058
rect 14332 12033 14368 12034
rect 14436 12030 14474 12038
rect 14540 12062 14684 12068
rect 14540 12042 14548 12062
rect 14568 12042 14656 12062
rect 14676 12042 14684 12062
rect 14540 12034 14684 12042
rect 14540 12033 14576 12034
rect 11185 11687 11249 11748
rect 11605 11746 11709 11748
rect 11940 11746 11981 11748
rect 12450 11745 12471 11790
rect 12451 11724 12471 11745
rect 12501 11745 12520 11790
rect 13557 11881 13637 11923
rect 12501 11724 12518 11745
rect 12451 11705 12518 11724
rect 12100 11697 12172 11698
rect 12099 11689 12198 11697
rect 7129 11441 7166 11472
rect 7342 11470 7378 11472
rect 7342 11441 7379 11470
rect 6581 11432 6616 11433
rect 6558 11427 6616 11432
rect 6558 11407 6561 11427
rect 6581 11413 6616 11427
rect 6636 11413 6645 11433
rect 6581 11405 6645 11413
rect 6607 11404 6645 11405
rect 6608 11403 6645 11404
rect 6711 11437 6747 11438
rect 6819 11437 6855 11438
rect 6711 11429 6855 11437
rect 6711 11409 6719 11429
rect 6739 11409 6827 11429
rect 6847 11409 6855 11429
rect 6711 11403 6855 11409
rect 6921 11433 6959 11441
rect 7027 11437 7063 11438
rect 6921 11413 6930 11433
rect 6950 11413 6959 11433
rect 6921 11404 6959 11413
rect 6978 11430 7063 11437
rect 6978 11410 6985 11430
rect 7006 11429 7063 11430
rect 7006 11410 7035 11429
rect 6978 11409 7035 11410
rect 7055 11409 7063 11429
rect 6921 11403 6958 11404
rect 6978 11403 7063 11409
rect 7129 11433 7167 11441
rect 7240 11437 7276 11438
rect 7129 11413 7138 11433
rect 7158 11413 7167 11433
rect 7129 11404 7167 11413
rect 7191 11429 7276 11437
rect 7191 11409 7248 11429
rect 7268 11409 7276 11429
rect 7129 11403 7166 11404
rect 7191 11403 7276 11409
rect 7342 11433 7380 11441
rect 7342 11413 7351 11433
rect 7371 11413 7380 11433
rect 7342 11404 7380 11413
rect 8867 11422 8947 11473
rect 7342 11403 7379 11404
rect 6765 11382 6801 11403
rect 7191 11382 7222 11403
rect 7402 11388 7459 11396
rect 7402 11382 7410 11388
rect 6598 11378 6698 11382
rect 6598 11374 6660 11378
rect 6598 11348 6605 11374
rect 6631 11352 6660 11374
rect 6686 11352 6698 11378
rect 6631 11348 6698 11352
rect 6598 11345 6698 11348
rect 6766 11345 6801 11382
rect 6863 11379 7222 11382
rect 6863 11374 7085 11379
rect 6863 11350 6876 11374
rect 6900 11355 7085 11374
rect 7109 11355 7222 11379
rect 6900 11350 7222 11355
rect 6863 11346 7222 11350
rect 7289 11374 7410 11382
rect 7289 11354 7300 11374
rect 7320 11365 7410 11374
rect 7436 11365 7459 11388
rect 7320 11354 7459 11365
rect 7289 11352 7459 11354
rect 7762 11381 7834 11401
rect 7762 11358 7790 11381
rect 7816 11358 7834 11381
rect 7289 11347 7410 11352
rect 7289 11346 7330 11347
rect 6765 11320 6801 11345
rect 6613 11293 6650 11294
rect 6709 11293 6746 11294
rect 6765 11293 6772 11320
rect 6513 11284 6651 11293
rect 6513 11264 6622 11284
rect 6642 11264 6651 11284
rect 6513 11257 6651 11264
rect 6709 11290 6772 11293
rect 6793 11293 6801 11320
rect 6820 11293 6857 11294
rect 6793 11290 6857 11293
rect 6709 11284 6857 11290
rect 6709 11264 6718 11284
rect 6738 11264 6828 11284
rect 6848 11264 6857 11284
rect 6513 11255 6609 11257
rect 6709 11254 6857 11264
rect 6916 11284 6953 11294
rect 7028 11293 7065 11294
rect 7009 11291 7065 11293
rect 6916 11264 6924 11284
rect 6944 11264 6953 11284
rect 6765 11253 6801 11254
rect 6613 11122 6650 11123
rect 6916 11122 6953 11264
rect 6978 11284 7065 11291
rect 6978 11281 7036 11284
rect 6978 11261 6983 11281
rect 7004 11264 7036 11281
rect 7056 11264 7065 11284
rect 7004 11261 7065 11264
rect 6978 11254 7065 11261
rect 7124 11284 7161 11294
rect 7124 11264 7132 11284
rect 7152 11264 7161 11284
rect 6978 11253 7009 11254
rect 7124 11185 7161 11264
rect 7191 11293 7222 11346
rect 7762 11296 7834 11358
rect 8867 11396 8883 11422
rect 8923 11396 8947 11422
rect 8867 11377 8947 11396
rect 8867 11351 8886 11377
rect 8926 11351 8947 11377
rect 8867 11324 8947 11351
rect 8867 11298 8890 11324
rect 8930 11298 8947 11324
rect 7241 11293 7278 11294
rect 7191 11284 7278 11293
rect 7191 11264 7249 11284
rect 7269 11264 7278 11284
rect 7191 11254 7278 11264
rect 7337 11284 7374 11294
rect 7337 11264 7345 11284
rect 7365 11264 7374 11284
rect 7191 11253 7222 11254
rect 7186 11185 7296 11198
rect 7337 11185 7374 11264
rect 7124 11183 7374 11185
rect 7124 11180 7225 11183
rect 7124 11161 7189 11180
rect 7186 11153 7189 11161
rect 7218 11153 7225 11180
rect 7253 11156 7263 11183
rect 7292 11161 7374 11183
rect 7292 11156 7296 11161
rect 7253 11153 7296 11156
rect 7186 11139 7296 11153
rect 6612 11121 6953 11122
rect 6537 11116 6953 11121
rect 6537 11096 6540 11116
rect 6560 11096 6954 11116
rect 6763 11063 6800 11073
rect 6763 11026 6772 11063
rect 6789 11026 6800 11063
rect 6763 11005 6800 11026
rect 6472 10066 6640 10067
rect 6769 10066 6798 11005
rect 6911 10391 6954 11096
rect 7766 10745 7828 11296
rect 8867 11287 8947 11298
rect 9009 11288 9036 11543
rect 9414 11535 9455 11685
rect 9686 11679 9790 11685
rect 10146 11682 10210 11685
rect 9881 11623 10002 11641
rect 9881 11621 9952 11623
rect 9881 11580 9896 11621
rect 9933 11582 9952 11621
rect 9989 11582 10002 11623
rect 9933 11580 10002 11582
rect 9881 11570 10002 11580
rect 9076 11428 9140 11440
rect 9416 11436 9453 11535
rect 9681 11525 9792 11538
rect 9681 11523 9723 11525
rect 9681 11503 9688 11523
rect 9707 11503 9723 11523
rect 9681 11495 9723 11503
rect 9751 11523 9792 11525
rect 9751 11503 9765 11523
rect 9784 11503 9792 11523
rect 9751 11495 9792 11503
rect 9681 11489 9792 11495
rect 9624 11467 9873 11489
rect 9624 11436 9661 11467
rect 9837 11465 9873 11467
rect 9837 11436 9874 11465
rect 9076 11427 9111 11428
rect 9053 11422 9111 11427
rect 9053 11402 9056 11422
rect 9076 11408 9111 11422
rect 9131 11408 9140 11428
rect 9076 11400 9140 11408
rect 9102 11399 9140 11400
rect 9103 11398 9140 11399
rect 9206 11432 9242 11433
rect 9314 11432 9350 11433
rect 9206 11424 9350 11432
rect 9206 11404 9214 11424
rect 9234 11404 9322 11424
rect 9342 11404 9350 11424
rect 9206 11398 9350 11404
rect 9416 11428 9454 11436
rect 9522 11432 9558 11433
rect 9416 11408 9425 11428
rect 9445 11408 9454 11428
rect 9416 11399 9454 11408
rect 9473 11425 9558 11432
rect 9473 11405 9480 11425
rect 9501 11424 9558 11425
rect 9501 11405 9530 11424
rect 9473 11404 9530 11405
rect 9550 11404 9558 11424
rect 9416 11398 9453 11399
rect 9473 11398 9558 11404
rect 9624 11428 9662 11436
rect 9735 11432 9771 11433
rect 9624 11408 9633 11428
rect 9653 11408 9662 11428
rect 9624 11399 9662 11408
rect 9686 11424 9771 11432
rect 9686 11404 9743 11424
rect 9763 11404 9771 11424
rect 9624 11398 9661 11399
rect 9686 11398 9771 11404
rect 9837 11428 9875 11436
rect 9837 11408 9846 11428
rect 9866 11408 9875 11428
rect 9930 11418 9995 11570
rect 10148 11544 10203 11682
rect 11187 11616 11246 11687
rect 12099 11686 12151 11689
rect 12099 11651 12107 11686
rect 12132 11651 12151 11686
rect 12176 11678 12198 11689
rect 12176 11677 13043 11678
rect 12176 11651 13044 11677
rect 12099 11641 13044 11651
rect 12099 11639 12198 11641
rect 11187 11598 11209 11616
rect 11227 11598 11246 11616
rect 11187 11576 11246 11598
rect 11454 11612 11986 11617
rect 11454 11592 12340 11612
rect 12360 11592 12363 11612
rect 12999 11608 13044 11641
rect 11454 11588 12363 11592
rect 9837 11399 9875 11408
rect 9928 11411 9995 11418
rect 9837 11398 9874 11399
rect 9260 11377 9296 11398
rect 9686 11377 9717 11398
rect 9928 11390 9945 11411
rect 9981 11390 9995 11411
rect 10147 11431 10203 11544
rect 11454 11541 11497 11588
rect 11947 11587 12363 11588
rect 12995 11588 13388 11608
rect 13408 11588 13411 11608
rect 11947 11586 12288 11587
rect 11604 11555 11714 11569
rect 11604 11552 11647 11555
rect 11604 11547 11608 11552
rect 11442 11540 11497 11541
rect 10147 11413 10166 11431
rect 10184 11413 10203 11431
rect 10147 11393 10203 11413
rect 11186 11517 11497 11540
rect 11186 11499 11211 11517
rect 11229 11505 11497 11517
rect 11526 11525 11608 11547
rect 11637 11525 11647 11552
rect 11675 11528 11682 11555
rect 11711 11547 11714 11555
rect 11711 11528 11776 11547
rect 11675 11525 11776 11528
rect 11526 11523 11776 11525
rect 11229 11499 11251 11505
rect 9928 11377 9995 11390
rect 9093 11373 9193 11377
rect 9093 11369 9155 11373
rect 9093 11343 9100 11369
rect 9126 11347 9155 11369
rect 9181 11347 9193 11373
rect 9126 11343 9193 11347
rect 9093 11340 9193 11343
rect 9261 11340 9296 11377
rect 9358 11374 9717 11377
rect 9358 11369 9580 11374
rect 9358 11345 9371 11369
rect 9395 11350 9580 11369
rect 9604 11350 9717 11374
rect 9395 11345 9717 11350
rect 9358 11341 9717 11345
rect 9784 11371 9995 11377
rect 9784 11369 9945 11371
rect 9784 11349 9795 11369
rect 9815 11349 9945 11369
rect 9784 11342 9945 11349
rect 9784 11341 9825 11342
rect 9260 11315 9296 11340
rect 9108 11288 9145 11289
rect 9204 11288 9241 11289
rect 9260 11288 9267 11315
rect 9008 11279 9146 11288
rect 9008 11259 9117 11279
rect 9137 11259 9146 11279
rect 9008 11252 9146 11259
rect 9204 11285 9267 11288
rect 9288 11288 9296 11315
rect 9315 11288 9352 11289
rect 9288 11285 9352 11288
rect 9204 11279 9352 11285
rect 9204 11259 9213 11279
rect 9233 11259 9323 11279
rect 9343 11259 9352 11279
rect 9008 11250 9104 11252
rect 9204 11249 9352 11259
rect 9411 11279 9448 11289
rect 9523 11288 9560 11289
rect 9504 11286 9560 11288
rect 9411 11259 9419 11279
rect 9439 11259 9448 11279
rect 9260 11248 9296 11249
rect 9108 11117 9145 11118
rect 9411 11117 9448 11259
rect 9473 11279 9560 11286
rect 9473 11276 9531 11279
rect 9473 11256 9478 11276
rect 9499 11259 9531 11276
rect 9551 11259 9560 11279
rect 9499 11256 9560 11259
rect 9473 11249 9560 11256
rect 9619 11279 9656 11289
rect 9619 11259 9627 11279
rect 9647 11259 9656 11279
rect 9473 11248 9504 11249
rect 9619 11180 9656 11259
rect 9686 11288 9717 11341
rect 9930 11334 9945 11342
rect 9985 11334 9995 11371
rect 11186 11360 11251 11499
rect 11526 11444 11563 11523
rect 11604 11510 11714 11523
rect 11678 11454 11709 11455
rect 11526 11424 11535 11444
rect 11555 11424 11563 11444
rect 9930 11325 9995 11334
rect 10143 11332 10208 11353
rect 10143 11314 10168 11332
rect 10186 11314 10208 11332
rect 11186 11342 11209 11360
rect 11227 11342 11251 11360
rect 11186 11325 11251 11342
rect 11406 11406 11474 11419
rect 11526 11414 11563 11424
rect 11622 11444 11709 11454
rect 11622 11424 11631 11444
rect 11651 11424 11709 11444
rect 11622 11415 11709 11424
rect 11622 11414 11659 11415
rect 11406 11364 11413 11406
rect 11462 11364 11474 11406
rect 11406 11361 11474 11364
rect 11678 11362 11709 11415
rect 11739 11444 11776 11523
rect 11891 11454 11922 11455
rect 11739 11424 11748 11444
rect 11768 11424 11776 11444
rect 11739 11414 11776 11424
rect 11835 11447 11922 11454
rect 11835 11444 11896 11447
rect 11835 11424 11844 11444
rect 11864 11427 11896 11444
rect 11917 11427 11922 11447
rect 11864 11424 11922 11427
rect 11835 11417 11922 11424
rect 11947 11444 11984 11586
rect 12250 11585 12287 11586
rect 12995 11583 13411 11588
rect 12995 11582 13336 11583
rect 12652 11551 12762 11565
rect 12652 11548 12695 11551
rect 12652 11543 12656 11548
rect 12574 11521 12656 11543
rect 12685 11521 12695 11548
rect 12723 11524 12730 11551
rect 12759 11543 12762 11551
rect 12759 11524 12824 11543
rect 12723 11521 12824 11524
rect 12574 11519 12824 11521
rect 12099 11454 12135 11455
rect 11947 11424 11956 11444
rect 11976 11424 11984 11444
rect 11835 11415 11891 11417
rect 11835 11414 11872 11415
rect 11947 11414 11984 11424
rect 12043 11444 12191 11454
rect 12291 11451 12387 11453
rect 12043 11424 12052 11444
rect 12072 11424 12162 11444
rect 12182 11424 12191 11444
rect 12043 11418 12191 11424
rect 12043 11415 12107 11418
rect 12043 11414 12080 11415
rect 12099 11388 12107 11415
rect 12128 11415 12191 11418
rect 12249 11444 12387 11451
rect 12249 11424 12258 11444
rect 12278 11424 12387 11444
rect 12249 11415 12387 11424
rect 12574 11440 12611 11519
rect 12652 11506 12762 11519
rect 12726 11450 12757 11451
rect 12574 11420 12583 11440
rect 12603 11420 12611 11440
rect 12128 11388 12135 11415
rect 12154 11414 12191 11415
rect 12250 11414 12287 11415
rect 12099 11363 12135 11388
rect 11570 11361 11611 11362
rect 11406 11354 11611 11361
rect 11406 11343 11580 11354
rect 9736 11288 9773 11289
rect 9686 11279 9773 11288
rect 9686 11259 9744 11279
rect 9764 11259 9773 11279
rect 9686 11249 9773 11259
rect 9832 11279 9869 11289
rect 9832 11259 9840 11279
rect 9860 11259 9869 11279
rect 9686 11248 9717 11249
rect 9681 11180 9791 11193
rect 9832 11180 9869 11259
rect 10143 11238 10208 11314
rect 11406 11310 11414 11343
rect 11407 11301 11414 11310
rect 11463 11334 11580 11343
rect 11600 11334 11611 11354
rect 11463 11326 11611 11334
rect 11678 11358 12037 11362
rect 11678 11353 12000 11358
rect 11678 11329 11791 11353
rect 11815 11334 12000 11353
rect 12024 11334 12037 11358
rect 11815 11329 12037 11334
rect 11678 11326 12037 11329
rect 12099 11326 12134 11363
rect 12202 11360 12302 11363
rect 12202 11356 12269 11360
rect 12202 11330 12214 11356
rect 12240 11334 12269 11356
rect 12295 11334 12302 11360
rect 12240 11330 12302 11334
rect 12202 11326 12302 11330
rect 11463 11310 11474 11326
rect 11463 11301 11471 11310
rect 11678 11305 11709 11326
rect 12099 11305 12135 11326
rect 11521 11304 11558 11305
rect 11186 11261 11251 11280
rect 11186 11243 11211 11261
rect 11229 11243 11251 11261
rect 9619 11178 9869 11180
rect 9619 11175 9720 11178
rect 9619 11156 9684 11175
rect 9681 11148 9684 11156
rect 9713 11148 9720 11175
rect 9748 11151 9758 11178
rect 9787 11156 9869 11178
rect 9892 11203 10209 11238
rect 9787 11151 9791 11156
rect 9748 11148 9791 11151
rect 9681 11134 9791 11148
rect 9107 11116 9448 11117
rect 9032 11114 9448 11116
rect 9892 11114 9932 11203
rect 10143 11176 10208 11203
rect 10143 11158 10166 11176
rect 10184 11158 10208 11176
rect 10143 11138 10208 11158
rect 9029 11111 9932 11114
rect 9029 11091 9035 11111
rect 9055 11091 9932 11111
rect 9029 11087 9932 11091
rect 9892 11084 9932 11087
rect 10144 11077 10209 11098
rect 8362 11069 9023 11070
rect 8362 11062 9296 11069
rect 8362 11061 9268 11062
rect 8362 11041 9213 11061
rect 9245 11042 9268 11061
rect 9293 11042 9296 11062
rect 9245 11041 9296 11042
rect 8362 11034 9296 11041
rect 7961 10992 8129 10993
rect 8364 10992 8403 11034
rect 9192 11032 9296 11034
rect 9261 11030 9296 11032
rect 10144 11059 10168 11077
rect 10186 11059 10209 11077
rect 10144 11012 10209 11059
rect 7961 10966 8405 10992
rect 7961 10964 8129 10966
rect 7763 10661 7832 10745
rect 6912 10383 6954 10391
rect 6912 10372 6957 10383
rect 6912 10334 6922 10372
rect 6947 10334 6957 10372
rect 6912 10325 6957 10334
rect 7761 10182 7832 10661
rect 7961 10613 7988 10964
rect 8364 10960 8405 10966
rect 8028 10753 8092 10765
rect 8368 10761 8405 10960
rect 8867 10987 8939 11004
rect 8867 10948 8875 10987
rect 8920 10948 8939 10987
rect 8633 10850 8744 10865
rect 8633 10848 8675 10850
rect 8633 10828 8640 10848
rect 8659 10828 8675 10848
rect 8633 10820 8675 10828
rect 8703 10848 8744 10850
rect 8703 10828 8717 10848
rect 8736 10828 8744 10848
rect 8703 10820 8744 10828
rect 8633 10814 8744 10820
rect 8576 10792 8825 10814
rect 8576 10761 8613 10792
rect 8789 10790 8825 10792
rect 8789 10761 8826 10790
rect 8028 10752 8063 10753
rect 8005 10747 8063 10752
rect 8005 10727 8008 10747
rect 8028 10733 8063 10747
rect 8083 10733 8092 10753
rect 8028 10725 8092 10733
rect 8054 10724 8092 10725
rect 8055 10723 8092 10724
rect 8158 10757 8194 10758
rect 8266 10757 8302 10758
rect 8158 10749 8302 10757
rect 8158 10729 8166 10749
rect 8186 10729 8274 10749
rect 8294 10729 8302 10749
rect 8158 10723 8302 10729
rect 8368 10753 8406 10761
rect 8474 10757 8510 10758
rect 8368 10733 8377 10753
rect 8397 10733 8406 10753
rect 8368 10724 8406 10733
rect 8425 10750 8510 10757
rect 8425 10730 8432 10750
rect 8453 10749 8510 10750
rect 8453 10730 8482 10749
rect 8425 10729 8482 10730
rect 8502 10729 8510 10749
rect 8368 10723 8405 10724
rect 8425 10723 8510 10729
rect 8576 10753 8614 10761
rect 8687 10757 8723 10758
rect 8576 10733 8585 10753
rect 8605 10733 8614 10753
rect 8576 10724 8614 10733
rect 8638 10749 8723 10757
rect 8638 10729 8695 10749
rect 8715 10729 8723 10749
rect 8576 10723 8613 10724
rect 8638 10723 8723 10729
rect 8789 10753 8827 10761
rect 8789 10733 8798 10753
rect 8818 10733 8827 10753
rect 8789 10724 8827 10733
rect 8867 10738 8939 10948
rect 9009 10982 10209 11012
rect 9009 10981 9453 10982
rect 9009 10979 9177 10981
rect 8867 10724 8950 10738
rect 8789 10723 8826 10724
rect 8212 10702 8248 10723
rect 8638 10702 8669 10723
rect 8867 10702 8884 10724
rect 8045 10698 8145 10702
rect 8045 10694 8107 10698
rect 8045 10668 8052 10694
rect 8078 10672 8107 10694
rect 8133 10672 8145 10698
rect 8078 10668 8145 10672
rect 8045 10665 8145 10668
rect 8213 10665 8248 10702
rect 8310 10699 8669 10702
rect 8310 10694 8532 10699
rect 8310 10670 8323 10694
rect 8347 10675 8532 10694
rect 8556 10675 8669 10699
rect 8347 10670 8669 10675
rect 8310 10666 8669 10670
rect 8736 10694 8884 10702
rect 8736 10674 8747 10694
rect 8767 10691 8884 10694
rect 8937 10691 8950 10724
rect 8767 10674 8950 10691
rect 8736 10667 8950 10674
rect 8736 10666 8777 10667
rect 8867 10666 8950 10667
rect 8212 10640 8248 10665
rect 8060 10613 8097 10614
rect 8156 10613 8193 10614
rect 8212 10613 8219 10640
rect 7960 10604 8098 10613
rect 7960 10584 8069 10604
rect 8089 10584 8098 10604
rect 7960 10577 8098 10584
rect 8156 10610 8219 10613
rect 8240 10613 8248 10640
rect 8267 10613 8304 10614
rect 8240 10610 8304 10613
rect 8156 10604 8304 10610
rect 8156 10584 8165 10604
rect 8185 10584 8275 10604
rect 8295 10584 8304 10604
rect 7960 10575 8056 10577
rect 8156 10574 8304 10584
rect 8363 10604 8400 10614
rect 8475 10613 8512 10614
rect 8456 10611 8512 10613
rect 8363 10584 8371 10604
rect 8391 10584 8400 10604
rect 8212 10573 8248 10574
rect 8060 10442 8097 10443
rect 8363 10442 8400 10584
rect 8425 10604 8512 10611
rect 8425 10601 8483 10604
rect 8425 10581 8430 10601
rect 8451 10584 8483 10601
rect 8503 10584 8512 10604
rect 8451 10581 8512 10584
rect 8425 10574 8512 10581
rect 8571 10604 8608 10614
rect 8571 10584 8579 10604
rect 8599 10584 8608 10604
rect 8425 10573 8456 10574
rect 8571 10505 8608 10584
rect 8638 10613 8669 10666
rect 8875 10633 8889 10666
rect 8942 10633 8950 10666
rect 8875 10627 8950 10633
rect 8875 10622 8945 10627
rect 8688 10613 8725 10614
rect 8638 10604 8725 10613
rect 8638 10584 8696 10604
rect 8716 10584 8725 10604
rect 8638 10574 8725 10584
rect 8784 10604 8821 10614
rect 9009 10609 9036 10979
rect 9076 10749 9140 10761
rect 9416 10757 9453 10981
rect 9924 10962 9988 10964
rect 9920 10950 9988 10962
rect 9920 10917 9931 10950
rect 9971 10917 9988 10950
rect 9920 10907 9988 10917
rect 9681 10846 9792 10861
rect 9681 10844 9723 10846
rect 9681 10824 9688 10844
rect 9707 10824 9723 10844
rect 9681 10816 9723 10824
rect 9751 10844 9792 10846
rect 9751 10824 9765 10844
rect 9784 10824 9792 10844
rect 9751 10816 9792 10824
rect 9681 10810 9792 10816
rect 9624 10788 9873 10810
rect 9624 10757 9661 10788
rect 9837 10786 9873 10788
rect 9837 10757 9874 10786
rect 9076 10748 9111 10749
rect 9053 10743 9111 10748
rect 9053 10723 9056 10743
rect 9076 10729 9111 10743
rect 9131 10729 9140 10749
rect 9076 10721 9140 10729
rect 9102 10720 9140 10721
rect 9103 10719 9140 10720
rect 9206 10753 9242 10754
rect 9314 10753 9350 10754
rect 9206 10745 9350 10753
rect 9206 10725 9214 10745
rect 9234 10725 9322 10745
rect 9342 10725 9350 10745
rect 9206 10719 9350 10725
rect 9416 10749 9454 10757
rect 9522 10753 9558 10754
rect 9416 10729 9425 10749
rect 9445 10729 9454 10749
rect 9416 10720 9454 10729
rect 9473 10746 9558 10753
rect 9473 10726 9480 10746
rect 9501 10745 9558 10746
rect 9501 10726 9530 10745
rect 9473 10725 9530 10726
rect 9550 10725 9558 10745
rect 9416 10719 9453 10720
rect 9473 10719 9558 10725
rect 9624 10749 9662 10757
rect 9735 10753 9771 10754
rect 9624 10729 9633 10749
rect 9653 10729 9662 10749
rect 9624 10720 9662 10729
rect 9686 10745 9771 10753
rect 9686 10725 9743 10745
rect 9763 10725 9771 10745
rect 9624 10719 9661 10720
rect 9686 10719 9771 10725
rect 9837 10749 9875 10757
rect 9837 10729 9846 10749
rect 9866 10729 9875 10749
rect 9837 10720 9875 10729
rect 9924 10723 9988 10907
rect 10144 10781 10209 10982
rect 11186 11042 11251 11243
rect 11407 11117 11471 11301
rect 11520 11295 11558 11304
rect 11520 11275 11529 11295
rect 11549 11275 11558 11295
rect 11520 11267 11558 11275
rect 11624 11299 11709 11305
rect 11734 11304 11771 11305
rect 11624 11279 11632 11299
rect 11652 11279 11709 11299
rect 11624 11271 11709 11279
rect 11733 11295 11771 11304
rect 11733 11275 11742 11295
rect 11762 11275 11771 11295
rect 11624 11270 11660 11271
rect 11733 11267 11771 11275
rect 11837 11299 11922 11305
rect 11942 11304 11979 11305
rect 11837 11279 11845 11299
rect 11865 11298 11922 11299
rect 11865 11279 11894 11298
rect 11837 11278 11894 11279
rect 11915 11278 11922 11298
rect 11837 11271 11922 11278
rect 11941 11295 11979 11304
rect 11941 11275 11950 11295
rect 11970 11275 11979 11295
rect 11837 11270 11873 11271
rect 11941 11267 11979 11275
rect 12045 11299 12189 11305
rect 12045 11279 12053 11299
rect 12073 11279 12161 11299
rect 12181 11279 12189 11299
rect 12045 11271 12189 11279
rect 12045 11270 12081 11271
rect 12153 11270 12189 11271
rect 12255 11304 12292 11305
rect 12255 11303 12293 11304
rect 12255 11295 12319 11303
rect 12255 11275 12264 11295
rect 12284 11281 12319 11295
rect 12339 11281 12342 11301
rect 12284 11276 12342 11281
rect 12284 11275 12319 11276
rect 11521 11238 11558 11267
rect 11522 11236 11558 11238
rect 11734 11236 11771 11267
rect 11522 11214 11771 11236
rect 11603 11208 11714 11214
rect 11603 11200 11644 11208
rect 11603 11180 11611 11200
rect 11630 11180 11644 11200
rect 11603 11178 11644 11180
rect 11672 11200 11714 11208
rect 11672 11180 11688 11200
rect 11707 11180 11714 11200
rect 11672 11178 11714 11180
rect 11603 11163 11714 11178
rect 11407 11107 11475 11117
rect 11407 11074 11424 11107
rect 11464 11074 11475 11107
rect 11407 11062 11475 11074
rect 11407 11060 11471 11062
rect 11942 11043 11979 11267
rect 12255 11263 12319 11275
rect 12359 11045 12386 11415
rect 12574 11410 12611 11420
rect 12670 11440 12757 11450
rect 12670 11420 12679 11440
rect 12699 11420 12757 11440
rect 12670 11411 12757 11420
rect 12670 11410 12707 11411
rect 12450 11397 12520 11402
rect 12445 11391 12520 11397
rect 12445 11358 12453 11391
rect 12506 11358 12520 11391
rect 12726 11358 12757 11411
rect 12787 11440 12824 11519
rect 12939 11450 12970 11451
rect 12787 11420 12796 11440
rect 12816 11420 12824 11440
rect 12787 11410 12824 11420
rect 12883 11443 12970 11450
rect 12883 11440 12944 11443
rect 12883 11420 12892 11440
rect 12912 11423 12944 11440
rect 12965 11423 12970 11443
rect 12912 11420 12970 11423
rect 12883 11413 12970 11420
rect 12995 11440 13032 11582
rect 13298 11581 13335 11582
rect 13147 11450 13183 11451
rect 12995 11420 13004 11440
rect 13024 11420 13032 11440
rect 12883 11411 12939 11413
rect 12883 11410 12920 11411
rect 12995 11410 13032 11420
rect 13091 11440 13239 11450
rect 13339 11447 13435 11449
rect 13091 11420 13100 11440
rect 13120 11420 13210 11440
rect 13230 11420 13239 11440
rect 13091 11414 13239 11420
rect 13091 11411 13155 11414
rect 13091 11410 13128 11411
rect 13147 11384 13155 11411
rect 13176 11411 13239 11414
rect 13297 11440 13435 11447
rect 13297 11420 13306 11440
rect 13326 11420 13435 11440
rect 13297 11411 13435 11420
rect 13176 11384 13183 11411
rect 13202 11410 13239 11411
rect 13298 11410 13335 11411
rect 13147 11359 13183 11384
rect 12445 11357 12528 11358
rect 12618 11357 12659 11358
rect 12445 11350 12659 11357
rect 12445 11333 12628 11350
rect 12445 11300 12458 11333
rect 12511 11330 12628 11333
rect 12648 11330 12659 11350
rect 12511 11322 12659 11330
rect 12726 11354 13085 11358
rect 12726 11349 13048 11354
rect 12726 11325 12839 11349
rect 12863 11330 13048 11349
rect 13072 11330 13085 11354
rect 12863 11325 13085 11330
rect 12726 11322 13085 11325
rect 13147 11322 13182 11359
rect 13250 11356 13350 11359
rect 13250 11352 13317 11356
rect 13250 11326 13262 11352
rect 13288 11330 13317 11352
rect 13343 11330 13350 11356
rect 13288 11326 13350 11330
rect 13250 11322 13350 11326
rect 12511 11300 12528 11322
rect 12726 11301 12757 11322
rect 13147 11301 13183 11322
rect 12569 11300 12606 11301
rect 12445 11286 12528 11300
rect 12218 11043 12386 11045
rect 11942 11042 12386 11043
rect 11186 11012 12386 11042
rect 12456 11076 12528 11286
rect 12568 11291 12606 11300
rect 12568 11271 12577 11291
rect 12597 11271 12606 11291
rect 12568 11263 12606 11271
rect 12672 11295 12757 11301
rect 12782 11300 12819 11301
rect 12672 11275 12680 11295
rect 12700 11275 12757 11295
rect 12672 11267 12757 11275
rect 12781 11291 12819 11300
rect 12781 11271 12790 11291
rect 12810 11271 12819 11291
rect 12672 11266 12708 11267
rect 12781 11263 12819 11271
rect 12885 11295 12970 11301
rect 12990 11300 13027 11301
rect 12885 11275 12893 11295
rect 12913 11294 12970 11295
rect 12913 11275 12942 11294
rect 12885 11274 12942 11275
rect 12963 11274 12970 11294
rect 12885 11267 12970 11274
rect 12989 11291 13027 11300
rect 12989 11271 12998 11291
rect 13018 11271 13027 11291
rect 12885 11266 12921 11267
rect 12989 11263 13027 11271
rect 13093 11295 13237 11301
rect 13093 11275 13101 11295
rect 13121 11275 13209 11295
rect 13229 11275 13237 11295
rect 13093 11267 13237 11275
rect 13093 11266 13129 11267
rect 13201 11266 13237 11267
rect 13303 11300 13340 11301
rect 13303 11299 13341 11300
rect 13303 11291 13367 11299
rect 13303 11271 13312 11291
rect 13332 11277 13367 11291
rect 13387 11277 13390 11297
rect 13332 11272 13390 11277
rect 13332 11271 13367 11272
rect 12569 11234 12606 11263
rect 12570 11232 12606 11234
rect 12782 11232 12819 11263
rect 12570 11210 12819 11232
rect 12651 11204 12762 11210
rect 12651 11196 12692 11204
rect 12651 11176 12659 11196
rect 12678 11176 12692 11196
rect 12651 11174 12692 11176
rect 12720 11196 12762 11204
rect 12720 11176 12736 11196
rect 12755 11176 12762 11196
rect 12720 11174 12762 11176
rect 12651 11159 12762 11174
rect 12456 11037 12475 11076
rect 12520 11037 12528 11076
rect 12456 11020 12528 11037
rect 12990 11064 13027 11263
rect 13303 11259 13367 11271
rect 12990 11058 13031 11064
rect 13407 11060 13434 11411
rect 13557 11281 13636 11881
rect 13733 11429 13812 12014
rect 14016 12001 14053 12030
rect 14017 11999 14053 12001
rect 14229 11999 14266 12030
rect 14017 11977 14266 11999
rect 14098 11971 14209 11977
rect 14098 11963 14139 11971
rect 14098 11943 14106 11963
rect 14125 11943 14139 11963
rect 14098 11941 14139 11943
rect 14167 11963 14209 11971
rect 14167 11943 14183 11963
rect 14202 11943 14209 11963
rect 14167 11941 14209 11943
rect 14098 11926 14209 11941
rect 14437 11915 14474 12030
rect 14430 11803 14477 11915
rect 14598 11875 14628 12034
rect 14648 12033 14684 12034
rect 14750 12067 14787 12068
rect 14750 12066 14788 12067
rect 14750 12058 14814 12066
rect 14750 12038 14759 12058
rect 14779 12044 14814 12058
rect 14834 12044 14837 12064
rect 14779 12039 14837 12044
rect 14779 12038 14814 12039
rect 14750 12026 14814 12038
rect 14598 11871 14684 11875
rect 14598 11853 14613 11871
rect 14665 11853 14684 11871
rect 14598 11844 14684 11853
rect 14854 11805 14881 12178
rect 14713 11803 14881 11805
rect 14430 11777 14881 11803
rect 14430 11699 14477 11777
rect 14713 11776 14881 11777
rect 14375 11698 14477 11699
rect 14374 11690 14477 11698
rect 14374 11687 14426 11690
rect 14374 11652 14382 11687
rect 14407 11652 14426 11687
rect 14451 11652 14477 11690
rect 14374 11646 14477 11652
rect 14637 11691 14673 11695
rect 14637 11668 14645 11691
rect 14669 11668 14673 11691
rect 14637 11647 14673 11668
rect 14374 11642 14473 11646
rect 14637 11624 14645 11647
rect 14669 11624 14673 11647
rect 13266 11058 13434 11060
rect 12990 11032 13434 11058
rect 11186 10965 11251 11012
rect 11186 10947 11209 10965
rect 11227 10947 11251 10965
rect 12099 10992 12134 10994
rect 12099 10990 12203 10992
rect 12992 10990 13031 11032
rect 13266 11031 13434 11032
rect 12099 10983 13033 10990
rect 12099 10982 12150 10983
rect 12099 10962 12102 10982
rect 12127 10963 12150 10982
rect 12182 10963 13033 10983
rect 12127 10962 13033 10963
rect 12099 10955 13033 10962
rect 12372 10954 13033 10955
rect 11186 10926 11251 10947
rect 11463 10937 11503 10940
rect 11463 10933 12366 10937
rect 11463 10913 12340 10933
rect 12360 10913 12366 10933
rect 11463 10910 12366 10913
rect 11187 10866 11252 10886
rect 11187 10848 11211 10866
rect 11229 10848 11252 10866
rect 11187 10821 11252 10848
rect 11463 10821 11503 10910
rect 11947 10908 12363 10910
rect 11947 10907 12288 10908
rect 11604 10876 11714 10890
rect 11604 10873 11647 10876
rect 11604 10868 11608 10873
rect 11186 10786 11503 10821
rect 11526 10846 11608 10868
rect 11637 10846 11647 10873
rect 11675 10849 11682 10876
rect 11711 10868 11714 10876
rect 11711 10849 11776 10868
rect 11675 10846 11776 10849
rect 11526 10844 11776 10846
rect 10144 10763 10166 10781
rect 10184 10763 10209 10781
rect 10144 10744 10209 10763
rect 9837 10719 9874 10720
rect 9260 10698 9296 10719
rect 9686 10698 9717 10719
rect 9924 10714 9932 10723
rect 9921 10698 9932 10714
rect 9093 10694 9193 10698
rect 9093 10690 9155 10694
rect 9093 10664 9100 10690
rect 9126 10668 9155 10690
rect 9181 10668 9193 10694
rect 9126 10664 9193 10668
rect 9093 10661 9193 10664
rect 9261 10661 9296 10698
rect 9358 10695 9717 10698
rect 9358 10690 9580 10695
rect 9358 10666 9371 10690
rect 9395 10671 9580 10690
rect 9604 10671 9717 10695
rect 9395 10666 9717 10671
rect 9358 10662 9717 10666
rect 9784 10690 9932 10698
rect 9784 10670 9795 10690
rect 9815 10681 9932 10690
rect 9981 10714 9988 10723
rect 9981 10681 9989 10714
rect 11187 10710 11252 10786
rect 11526 10765 11563 10844
rect 11604 10831 11714 10844
rect 11678 10775 11709 10776
rect 11526 10745 11535 10765
rect 11555 10745 11563 10765
rect 11526 10735 11563 10745
rect 11622 10765 11709 10775
rect 11622 10745 11631 10765
rect 11651 10745 11709 10765
rect 11622 10736 11709 10745
rect 11622 10735 11659 10736
rect 9815 10670 9989 10681
rect 9784 10663 9989 10670
rect 9784 10662 9825 10663
rect 9260 10636 9296 10661
rect 9108 10609 9145 10610
rect 9204 10609 9241 10610
rect 9260 10609 9267 10636
rect 8784 10584 8792 10604
rect 8812 10584 8821 10604
rect 8638 10573 8669 10574
rect 8633 10505 8743 10518
rect 8784 10505 8821 10584
rect 9008 10600 9146 10609
rect 9008 10580 9117 10600
rect 9137 10580 9146 10600
rect 9008 10573 9146 10580
rect 9204 10606 9267 10609
rect 9288 10609 9296 10636
rect 9315 10609 9352 10610
rect 9288 10606 9352 10609
rect 9204 10600 9352 10606
rect 9204 10580 9213 10600
rect 9233 10580 9323 10600
rect 9343 10580 9352 10600
rect 9008 10571 9104 10573
rect 9204 10570 9352 10580
rect 9411 10600 9448 10610
rect 9523 10609 9560 10610
rect 9504 10607 9560 10609
rect 9411 10580 9419 10600
rect 9439 10580 9448 10600
rect 9260 10569 9296 10570
rect 8571 10503 8821 10505
rect 8571 10500 8672 10503
rect 8571 10481 8636 10500
rect 8633 10473 8636 10481
rect 8665 10473 8672 10500
rect 8700 10476 8710 10503
rect 8739 10481 8821 10503
rect 8739 10476 8743 10481
rect 8700 10473 8743 10476
rect 8633 10459 8743 10473
rect 8059 10441 8400 10442
rect 7984 10436 8400 10441
rect 9108 10438 9145 10439
rect 9411 10438 9448 10580
rect 9473 10600 9560 10607
rect 9473 10597 9531 10600
rect 9473 10577 9478 10597
rect 9499 10580 9531 10597
rect 9551 10580 9560 10600
rect 9499 10577 9560 10580
rect 9473 10570 9560 10577
rect 9619 10600 9656 10610
rect 9619 10580 9627 10600
rect 9647 10580 9656 10600
rect 9473 10569 9504 10570
rect 9619 10501 9656 10580
rect 9686 10609 9717 10662
rect 9921 10660 9989 10663
rect 9921 10618 9933 10660
rect 9982 10618 9989 10660
rect 9736 10609 9773 10610
rect 9686 10600 9773 10609
rect 9686 10580 9744 10600
rect 9764 10580 9773 10600
rect 9686 10570 9773 10580
rect 9832 10600 9869 10610
rect 9921 10605 9989 10618
rect 10144 10682 10209 10699
rect 10144 10664 10168 10682
rect 10186 10664 10209 10682
rect 11187 10692 11209 10710
rect 11227 10692 11252 10710
rect 11187 10671 11252 10692
rect 11400 10690 11465 10699
rect 9832 10580 9840 10600
rect 9860 10580 9869 10600
rect 9686 10569 9717 10570
rect 9681 10501 9791 10514
rect 9832 10501 9869 10580
rect 10144 10525 10209 10664
rect 11400 10653 11410 10690
rect 11450 10682 11465 10690
rect 11678 10683 11709 10736
rect 11739 10765 11776 10844
rect 11891 10775 11922 10776
rect 11739 10745 11748 10765
rect 11768 10745 11776 10765
rect 11739 10735 11776 10745
rect 11835 10768 11922 10775
rect 11835 10765 11896 10768
rect 11835 10745 11844 10765
rect 11864 10748 11896 10765
rect 11917 10748 11922 10768
rect 11864 10745 11922 10748
rect 11835 10738 11922 10745
rect 11947 10765 11984 10907
rect 12250 10906 12287 10907
rect 12099 10775 12135 10776
rect 11947 10745 11956 10765
rect 11976 10745 11984 10765
rect 11835 10736 11891 10738
rect 11835 10735 11872 10736
rect 11947 10735 11984 10745
rect 12043 10765 12191 10775
rect 12291 10772 12387 10774
rect 12043 10745 12052 10765
rect 12072 10745 12162 10765
rect 12182 10745 12191 10765
rect 12043 10739 12191 10745
rect 12043 10736 12107 10739
rect 12043 10735 12080 10736
rect 12099 10709 12107 10736
rect 12128 10736 12191 10739
rect 12249 10765 12387 10772
rect 12249 10745 12258 10765
rect 12278 10745 12387 10765
rect 12249 10736 12387 10745
rect 12128 10709 12135 10736
rect 12154 10735 12191 10736
rect 12250 10735 12287 10736
rect 12099 10684 12135 10709
rect 11570 10682 11611 10683
rect 11450 10675 11611 10682
rect 11450 10655 11580 10675
rect 11600 10655 11611 10675
rect 11450 10653 11611 10655
rect 11400 10647 11611 10653
rect 11678 10679 12037 10683
rect 11678 10674 12000 10679
rect 11678 10650 11791 10674
rect 11815 10655 12000 10674
rect 12024 10655 12037 10679
rect 11815 10650 12037 10655
rect 11678 10647 12037 10650
rect 12099 10647 12134 10684
rect 12202 10681 12302 10684
rect 12202 10677 12269 10681
rect 12202 10651 12214 10677
rect 12240 10655 12269 10677
rect 12295 10655 12302 10681
rect 12240 10651 12302 10655
rect 12202 10647 12302 10651
rect 11400 10634 11467 10647
rect 10144 10519 10166 10525
rect 9619 10499 9869 10501
rect 9619 10496 9720 10499
rect 9619 10477 9684 10496
rect 9681 10469 9684 10477
rect 9713 10469 9720 10496
rect 9748 10472 9758 10499
rect 9787 10477 9869 10499
rect 9898 10507 10166 10519
rect 10184 10507 10209 10525
rect 9898 10484 10209 10507
rect 11192 10611 11248 10631
rect 11192 10593 11211 10611
rect 11229 10593 11248 10611
rect 9898 10483 9953 10484
rect 9787 10472 9791 10477
rect 9748 10469 9791 10472
rect 9681 10455 9791 10469
rect 9107 10437 9448 10438
rect 7984 10416 7987 10436
rect 8007 10416 8400 10436
rect 9032 10436 9448 10437
rect 9898 10436 9941 10483
rect 11192 10480 11248 10593
rect 11400 10613 11414 10634
rect 11450 10613 11467 10634
rect 11678 10626 11709 10647
rect 12099 10626 12135 10647
rect 11521 10625 11558 10626
rect 11400 10606 11467 10613
rect 11520 10616 11558 10625
rect 9032 10432 9941 10436
rect 8351 10383 8396 10416
rect 9032 10412 9035 10432
rect 9055 10412 9941 10432
rect 9409 10407 9941 10412
rect 10149 10426 10208 10448
rect 10149 10408 10168 10426
rect 10186 10408 10208 10426
rect 9197 10383 9296 10385
rect 8351 10373 9296 10383
rect 8351 10347 9219 10373
rect 8352 10346 9219 10347
rect 9197 10335 9219 10346
rect 9244 10338 9263 10373
rect 9288 10338 9296 10373
rect 9244 10335 9296 10338
rect 9197 10327 9296 10335
rect 9223 10326 9295 10327
rect 10149 10278 10208 10408
rect 11192 10351 11247 10480
rect 11400 10454 11465 10606
rect 11520 10596 11529 10616
rect 11549 10596 11558 10616
rect 11520 10588 11558 10596
rect 11624 10620 11709 10626
rect 11734 10625 11771 10626
rect 11624 10600 11632 10620
rect 11652 10600 11709 10620
rect 11624 10592 11709 10600
rect 11733 10616 11771 10625
rect 11733 10596 11742 10616
rect 11762 10596 11771 10616
rect 11624 10591 11660 10592
rect 11733 10588 11771 10596
rect 11837 10620 11922 10626
rect 11942 10625 11979 10626
rect 11837 10600 11845 10620
rect 11865 10619 11922 10620
rect 11865 10600 11894 10619
rect 11837 10599 11894 10600
rect 11915 10599 11922 10619
rect 11837 10592 11922 10599
rect 11941 10616 11979 10625
rect 11941 10596 11950 10616
rect 11970 10596 11979 10616
rect 11837 10591 11873 10592
rect 11941 10588 11979 10596
rect 12045 10620 12189 10626
rect 12045 10600 12053 10620
rect 12073 10600 12161 10620
rect 12181 10600 12189 10620
rect 12045 10592 12189 10600
rect 12045 10591 12081 10592
rect 12153 10591 12189 10592
rect 12255 10625 12292 10626
rect 12255 10624 12293 10625
rect 12255 10616 12319 10624
rect 12255 10596 12264 10616
rect 12284 10602 12319 10616
rect 12339 10602 12342 10622
rect 12284 10597 12342 10602
rect 12284 10596 12319 10597
rect 11521 10559 11558 10588
rect 11522 10557 11558 10559
rect 11734 10557 11771 10588
rect 11522 10535 11771 10557
rect 11603 10529 11714 10535
rect 11603 10521 11644 10529
rect 11603 10501 11611 10521
rect 11630 10501 11644 10521
rect 11603 10499 11644 10501
rect 11672 10521 11714 10529
rect 11672 10501 11688 10521
rect 11707 10501 11714 10521
rect 11672 10499 11714 10501
rect 11603 10484 11714 10499
rect 11942 10489 11979 10588
rect 12255 10584 12319 10596
rect 11605 10475 11709 10484
rect 11393 10444 11514 10454
rect 11393 10442 11462 10444
rect 11393 10401 11406 10442
rect 11443 10403 11462 10442
rect 11499 10403 11514 10444
rect 11443 10401 11514 10403
rect 11393 10383 11514 10401
rect 11186 10339 11247 10351
rect 11940 10339 11981 10489
rect 12359 10481 12386 10736
rect 12448 10726 12528 10737
rect 12448 10700 12465 10726
rect 12505 10700 12528 10726
rect 12448 10673 12528 10700
rect 12448 10647 12469 10673
rect 12509 10647 12528 10673
rect 12448 10628 12528 10647
rect 12448 10602 12472 10628
rect 12512 10602 12528 10628
rect 12448 10551 12528 10602
rect 11186 10336 11981 10339
rect 12360 10350 12386 10481
rect 12450 10395 12520 10551
rect 12449 10379 12525 10395
rect 12360 10336 12388 10350
rect 11186 10301 12388 10336
rect 12449 10342 12464 10379
rect 12508 10342 12525 10379
rect 12449 10322 12525 10342
rect 13563 10372 13633 11281
rect 13732 10716 13813 11429
rect 14637 11315 14673 11624
rect 14561 11286 14674 11315
rect 14561 10930 14592 11286
rect 14631 11031 15622 11056
rect 14631 11026 14691 11031
rect 14631 11005 14650 11026
rect 14670 11010 14691 11026
rect 14711 11010 15622 11031
rect 14670 11005 15622 11010
rect 14631 10997 15622 11005
rect 14636 10974 14742 10997
rect 14636 10971 14741 10974
rect 14485 10910 14878 10930
rect 14898 10910 14901 10930
rect 14485 10905 14901 10910
rect 14485 10904 14826 10905
rect 14142 10873 14252 10887
rect 14142 10870 14185 10873
rect 14142 10865 14146 10870
rect 14064 10843 14146 10865
rect 14175 10843 14185 10870
rect 14213 10846 14220 10873
rect 14249 10865 14252 10873
rect 14249 10846 14314 10865
rect 14213 10843 14314 10846
rect 14064 10841 14314 10843
rect 14064 10762 14101 10841
rect 14142 10828 14252 10841
rect 14216 10772 14247 10773
rect 14064 10742 14073 10762
rect 14093 10742 14101 10762
rect 14064 10732 14101 10742
rect 14160 10762 14247 10772
rect 14160 10742 14169 10762
rect 14189 10742 14247 10762
rect 14160 10733 14247 10742
rect 14160 10732 14197 10733
rect 13730 10680 13822 10716
rect 14216 10680 14247 10733
rect 14277 10762 14314 10841
rect 14429 10772 14460 10773
rect 14277 10742 14286 10762
rect 14306 10742 14314 10762
rect 14277 10732 14314 10742
rect 14373 10765 14460 10772
rect 14373 10762 14434 10765
rect 14373 10742 14382 10762
rect 14402 10745 14434 10762
rect 14455 10745 14460 10765
rect 14402 10742 14460 10745
rect 14373 10735 14460 10742
rect 14485 10762 14522 10904
rect 14788 10903 14825 10904
rect 14637 10772 14673 10773
rect 14485 10742 14494 10762
rect 14514 10742 14522 10762
rect 14373 10733 14429 10735
rect 14373 10732 14410 10733
rect 14485 10732 14522 10742
rect 14581 10762 14729 10772
rect 14829 10769 14925 10771
rect 14581 10742 14590 10762
rect 14610 10742 14700 10762
rect 14720 10742 14729 10762
rect 14581 10736 14729 10742
rect 14581 10733 14645 10736
rect 14581 10732 14618 10733
rect 14637 10706 14645 10733
rect 14666 10733 14729 10736
rect 14787 10762 14925 10769
rect 14787 10742 14796 10762
rect 14816 10742 14925 10762
rect 14787 10733 14925 10742
rect 14666 10706 14673 10733
rect 14692 10732 14729 10733
rect 14788 10732 14825 10733
rect 14637 10681 14673 10706
rect 13730 10679 14066 10680
rect 14108 10679 14149 10680
rect 13730 10672 14149 10679
rect 13730 10652 14118 10672
rect 14138 10652 14149 10672
rect 13730 10644 14149 10652
rect 14216 10676 14575 10680
rect 14216 10671 14538 10676
rect 14216 10647 14329 10671
rect 14353 10652 14538 10671
rect 14562 10652 14575 10676
rect 14353 10647 14575 10652
rect 14216 10644 14575 10647
rect 14637 10644 14672 10681
rect 14740 10678 14840 10681
rect 14740 10674 14807 10678
rect 14740 10648 14752 10674
rect 14778 10652 14807 10674
rect 14833 10652 14840 10678
rect 14778 10648 14840 10652
rect 14740 10644 14840 10648
rect 13730 10640 14066 10644
rect 13563 10322 13635 10372
rect 8871 10248 8947 10272
rect 8871 10182 8883 10248
rect 8937 10182 8947 10248
rect 9415 10203 9456 10205
rect 9687 10203 9791 10205
rect 10149 10203 10210 10278
rect 11186 10226 11247 10301
rect 11605 10299 11709 10301
rect 11940 10299 11981 10301
rect 12449 10256 12459 10322
rect 12513 10256 12525 10322
rect 12449 10232 12525 10256
rect 7761 10132 7833 10182
rect 6472 10040 6916 10066
rect 6472 10038 6640 10040
rect 6472 9771 6499 10038
rect 6769 10036 6798 10040
rect 6539 9911 6603 9923
rect 6879 9919 6916 10040
rect 7144 10008 7255 10023
rect 7144 10006 7186 10008
rect 7144 9986 7151 10006
rect 7170 9986 7186 10006
rect 7144 9978 7186 9986
rect 7214 10006 7255 10008
rect 7214 9986 7228 10006
rect 7247 9986 7255 10006
rect 7214 9978 7255 9986
rect 7144 9972 7255 9978
rect 7087 9950 7336 9972
rect 7087 9919 7124 9950
rect 7300 9948 7336 9950
rect 7300 9919 7337 9948
rect 6539 9910 6574 9911
rect 6516 9905 6574 9910
rect 6516 9885 6519 9905
rect 6539 9891 6574 9905
rect 6594 9891 6603 9911
rect 6539 9883 6603 9891
rect 6565 9882 6603 9883
rect 6566 9881 6603 9882
rect 6669 9915 6705 9916
rect 6777 9915 6813 9916
rect 6669 9907 6813 9915
rect 6669 9887 6677 9907
rect 6697 9887 6785 9907
rect 6805 9887 6813 9907
rect 6669 9881 6813 9887
rect 6879 9911 6917 9919
rect 6985 9915 7021 9916
rect 6879 9891 6888 9911
rect 6908 9891 6917 9911
rect 6879 9882 6917 9891
rect 6936 9908 7021 9915
rect 6936 9888 6943 9908
rect 6964 9907 7021 9908
rect 6964 9888 6993 9907
rect 6936 9887 6993 9888
rect 7013 9887 7021 9907
rect 6879 9881 6916 9882
rect 6936 9881 7021 9887
rect 7087 9911 7125 9919
rect 7198 9915 7234 9916
rect 7087 9891 7096 9911
rect 7116 9891 7125 9911
rect 7087 9882 7125 9891
rect 7149 9907 7234 9915
rect 7149 9887 7206 9907
rect 7226 9887 7234 9907
rect 7087 9881 7124 9882
rect 7149 9881 7234 9887
rect 7300 9911 7338 9919
rect 7300 9891 7309 9911
rect 7329 9891 7338 9911
rect 7300 9882 7338 9891
rect 7300 9881 7337 9882
rect 6723 9860 6759 9881
rect 7149 9860 7180 9881
rect 7330 9860 7664 9864
rect 6556 9856 6656 9860
rect 6556 9852 6618 9856
rect 6556 9826 6563 9852
rect 6589 9830 6618 9852
rect 6644 9830 6656 9856
rect 6589 9826 6656 9830
rect 6556 9823 6656 9826
rect 6724 9823 6759 9860
rect 6821 9857 7180 9860
rect 6821 9852 7043 9857
rect 6821 9828 6834 9852
rect 6858 9833 7043 9852
rect 7067 9833 7180 9857
rect 6858 9828 7180 9833
rect 6821 9824 7180 9828
rect 7247 9852 7664 9860
rect 7247 9832 7258 9852
rect 7278 9832 7664 9852
rect 7247 9825 7664 9832
rect 7247 9824 7288 9825
rect 7330 9824 7664 9825
rect 6723 9798 6759 9823
rect 6571 9771 6608 9772
rect 6667 9771 6704 9772
rect 6723 9771 6730 9798
rect 6471 9762 6609 9771
rect 6471 9742 6580 9762
rect 6600 9742 6609 9762
rect 6471 9735 6609 9742
rect 6667 9768 6730 9771
rect 6751 9771 6759 9798
rect 6778 9771 6815 9772
rect 6751 9768 6815 9771
rect 6667 9762 6815 9768
rect 6667 9742 6676 9762
rect 6696 9742 6786 9762
rect 6806 9742 6815 9762
rect 6471 9733 6567 9735
rect 6667 9732 6815 9742
rect 6874 9762 6911 9772
rect 6986 9771 7023 9772
rect 6967 9769 7023 9771
rect 6874 9742 6882 9762
rect 6902 9742 6911 9762
rect 6723 9731 6759 9732
rect 6571 9600 6608 9601
rect 6874 9600 6911 9742
rect 6936 9762 7023 9769
rect 6936 9759 6994 9762
rect 6936 9739 6941 9759
rect 6962 9742 6994 9759
rect 7014 9742 7023 9762
rect 6962 9739 7023 9742
rect 6936 9732 7023 9739
rect 7082 9762 7119 9772
rect 7082 9742 7090 9762
rect 7110 9742 7119 9762
rect 6936 9731 6967 9732
rect 7082 9663 7119 9742
rect 7149 9771 7180 9824
rect 7199 9771 7236 9772
rect 7149 9762 7236 9771
rect 7149 9742 7207 9762
rect 7227 9742 7236 9762
rect 7149 9732 7236 9742
rect 7295 9762 7332 9772
rect 7295 9742 7303 9762
rect 7323 9742 7332 9762
rect 7149 9731 7180 9732
rect 7144 9663 7254 9676
rect 7295 9663 7332 9742
rect 7082 9661 7332 9663
rect 7082 9658 7183 9661
rect 7082 9639 7147 9658
rect 7144 9631 7147 9639
rect 7176 9631 7183 9658
rect 7211 9634 7221 9661
rect 7250 9639 7332 9661
rect 7250 9634 7254 9639
rect 7211 9631 7254 9634
rect 7144 9617 7254 9631
rect 6570 9599 6911 9600
rect 6495 9594 6911 9599
rect 6495 9574 6498 9594
rect 6518 9574 6911 9594
rect 6804 9209 6835 9574
rect 6722 9180 6835 9209
rect 6723 8880 6759 9180
rect 7583 9075 7664 9824
rect 7763 9223 7833 10132
rect 8871 10162 8947 10182
rect 8871 10125 8888 10162
rect 8932 10125 8947 10162
rect 9008 10168 10210 10203
rect 9008 10154 9036 10168
rect 8871 10109 8947 10125
rect 8876 9953 8946 10109
rect 9010 10023 9036 10154
rect 9415 10165 10210 10168
rect 8868 9902 8948 9953
rect 8868 9876 8884 9902
rect 8924 9876 8948 9902
rect 8868 9857 8948 9876
rect 8868 9831 8887 9857
rect 8927 9831 8948 9857
rect 8868 9804 8948 9831
rect 8868 9778 8891 9804
rect 8931 9778 8948 9804
rect 8868 9767 8948 9778
rect 9010 9768 9037 10023
rect 9415 10015 9456 10165
rect 10149 10153 10210 10165
rect 9882 10103 10003 10121
rect 9882 10101 9953 10103
rect 9882 10060 9897 10101
rect 9934 10062 9953 10101
rect 9990 10062 10003 10103
rect 9934 10060 10003 10062
rect 9882 10050 10003 10060
rect 9687 10020 9791 10029
rect 9077 9908 9141 9920
rect 9417 9916 9454 10015
rect 9682 10005 9793 10020
rect 9682 10003 9724 10005
rect 9682 9983 9689 10003
rect 9708 9983 9724 10003
rect 9682 9975 9724 9983
rect 9752 10003 9793 10005
rect 9752 9983 9766 10003
rect 9785 9983 9793 10003
rect 9752 9975 9793 9983
rect 9682 9969 9793 9975
rect 9625 9947 9874 9969
rect 9625 9916 9662 9947
rect 9838 9945 9874 9947
rect 9838 9916 9875 9945
rect 9077 9907 9112 9908
rect 9054 9902 9112 9907
rect 9054 9882 9057 9902
rect 9077 9888 9112 9902
rect 9132 9888 9141 9908
rect 9077 9880 9141 9888
rect 9103 9879 9141 9880
rect 9104 9878 9141 9879
rect 9207 9912 9243 9913
rect 9315 9912 9351 9913
rect 9207 9904 9351 9912
rect 9207 9884 9215 9904
rect 9235 9884 9323 9904
rect 9343 9884 9351 9904
rect 9207 9878 9351 9884
rect 9417 9908 9455 9916
rect 9523 9912 9559 9913
rect 9417 9888 9426 9908
rect 9446 9888 9455 9908
rect 9417 9879 9455 9888
rect 9474 9905 9559 9912
rect 9474 9885 9481 9905
rect 9502 9904 9559 9905
rect 9502 9885 9531 9904
rect 9474 9884 9531 9885
rect 9551 9884 9559 9904
rect 9417 9878 9454 9879
rect 9474 9878 9559 9884
rect 9625 9908 9663 9916
rect 9736 9912 9772 9913
rect 9625 9888 9634 9908
rect 9654 9888 9663 9908
rect 9625 9879 9663 9888
rect 9687 9904 9772 9912
rect 9687 9884 9744 9904
rect 9764 9884 9772 9904
rect 9625 9878 9662 9879
rect 9687 9878 9772 9884
rect 9838 9908 9876 9916
rect 9838 9888 9847 9908
rect 9867 9888 9876 9908
rect 9931 9898 9996 10050
rect 10149 10024 10204 10153
rect 11188 10096 11247 10226
rect 12101 10177 12173 10178
rect 12100 10169 12199 10177
rect 12100 10166 12152 10169
rect 12100 10131 12108 10166
rect 12133 10131 12152 10166
rect 12177 10158 12199 10169
rect 12177 10157 13044 10158
rect 12177 10131 13045 10157
rect 12100 10121 13045 10131
rect 12100 10119 12199 10121
rect 11188 10078 11210 10096
rect 11228 10078 11247 10096
rect 11188 10056 11247 10078
rect 11455 10092 11987 10097
rect 11455 10072 12341 10092
rect 12361 10072 12364 10092
rect 13000 10088 13045 10121
rect 11455 10068 12364 10072
rect 9838 9879 9876 9888
rect 9929 9891 9996 9898
rect 9838 9878 9875 9879
rect 9261 9857 9297 9878
rect 9687 9857 9718 9878
rect 9929 9870 9946 9891
rect 9982 9870 9996 9891
rect 10148 9911 10204 10024
rect 11455 10021 11498 10068
rect 11948 10067 12364 10068
rect 12996 10068 13389 10088
rect 13409 10068 13412 10088
rect 11948 10066 12289 10067
rect 11605 10035 11715 10049
rect 11605 10032 11648 10035
rect 11605 10027 11609 10032
rect 11443 10020 11498 10021
rect 10148 9893 10167 9911
rect 10185 9893 10204 9911
rect 10148 9873 10204 9893
rect 11187 9997 11498 10020
rect 11187 9979 11212 9997
rect 11230 9985 11498 9997
rect 11527 10005 11609 10027
rect 11638 10005 11648 10032
rect 11676 10008 11683 10035
rect 11712 10027 11715 10035
rect 11712 10008 11777 10027
rect 11676 10005 11777 10008
rect 11527 10003 11777 10005
rect 11230 9979 11252 9985
rect 9929 9857 9996 9870
rect 9094 9853 9194 9857
rect 9094 9849 9156 9853
rect 9094 9823 9101 9849
rect 9127 9827 9156 9849
rect 9182 9827 9194 9853
rect 9127 9823 9194 9827
rect 9094 9820 9194 9823
rect 9262 9820 9297 9857
rect 9359 9854 9718 9857
rect 9359 9849 9581 9854
rect 9359 9825 9372 9849
rect 9396 9830 9581 9849
rect 9605 9830 9718 9854
rect 9396 9825 9718 9830
rect 9359 9821 9718 9825
rect 9785 9851 9996 9857
rect 9785 9849 9946 9851
rect 9785 9829 9796 9849
rect 9816 9829 9946 9849
rect 9785 9822 9946 9829
rect 9785 9821 9826 9822
rect 9261 9795 9297 9820
rect 9109 9768 9146 9769
rect 9205 9768 9242 9769
rect 9261 9768 9268 9795
rect 9009 9759 9147 9768
rect 9009 9739 9118 9759
rect 9138 9739 9147 9759
rect 9009 9732 9147 9739
rect 9205 9765 9268 9768
rect 9289 9768 9297 9795
rect 9316 9768 9353 9769
rect 9289 9765 9353 9768
rect 9205 9759 9353 9765
rect 9205 9739 9214 9759
rect 9234 9739 9324 9759
rect 9344 9739 9353 9759
rect 9009 9730 9105 9732
rect 9205 9729 9353 9739
rect 9412 9759 9449 9769
rect 9524 9768 9561 9769
rect 9505 9766 9561 9768
rect 9412 9739 9420 9759
rect 9440 9739 9449 9759
rect 9261 9728 9297 9729
rect 9109 9597 9146 9598
rect 9412 9597 9449 9739
rect 9474 9759 9561 9766
rect 9474 9756 9532 9759
rect 9474 9736 9479 9756
rect 9500 9739 9532 9756
rect 9552 9739 9561 9759
rect 9500 9736 9561 9739
rect 9474 9729 9561 9736
rect 9620 9759 9657 9769
rect 9620 9739 9628 9759
rect 9648 9739 9657 9759
rect 9474 9728 9505 9729
rect 9620 9660 9657 9739
rect 9687 9768 9718 9821
rect 9931 9814 9946 9822
rect 9986 9814 9996 9851
rect 11187 9840 11252 9979
rect 11527 9924 11564 10003
rect 11605 9990 11715 10003
rect 11679 9934 11710 9935
rect 11527 9904 11536 9924
rect 11556 9904 11564 9924
rect 9931 9805 9996 9814
rect 10144 9812 10209 9833
rect 10144 9794 10169 9812
rect 10187 9794 10209 9812
rect 11187 9822 11210 9840
rect 11228 9822 11252 9840
rect 11187 9805 11252 9822
rect 11407 9886 11475 9899
rect 11527 9894 11564 9904
rect 11623 9924 11710 9934
rect 11623 9904 11632 9924
rect 11652 9904 11710 9924
rect 11623 9895 11710 9904
rect 11623 9894 11660 9895
rect 11407 9844 11414 9886
rect 11463 9844 11475 9886
rect 11407 9841 11475 9844
rect 11679 9842 11710 9895
rect 11740 9924 11777 10003
rect 11892 9934 11923 9935
rect 11740 9904 11749 9924
rect 11769 9904 11777 9924
rect 11740 9894 11777 9904
rect 11836 9927 11923 9934
rect 11836 9924 11897 9927
rect 11836 9904 11845 9924
rect 11865 9907 11897 9924
rect 11918 9907 11923 9927
rect 11865 9904 11923 9907
rect 11836 9897 11923 9904
rect 11948 9924 11985 10066
rect 12251 10065 12288 10066
rect 12996 10063 13412 10068
rect 12996 10062 13337 10063
rect 12653 10031 12763 10045
rect 12653 10028 12696 10031
rect 12653 10023 12657 10028
rect 12575 10001 12657 10023
rect 12686 10001 12696 10028
rect 12724 10004 12731 10031
rect 12760 10023 12763 10031
rect 12760 10004 12825 10023
rect 12724 10001 12825 10004
rect 12575 9999 12825 10001
rect 12100 9934 12136 9935
rect 11948 9904 11957 9924
rect 11977 9904 11985 9924
rect 11836 9895 11892 9897
rect 11836 9894 11873 9895
rect 11948 9894 11985 9904
rect 12044 9924 12192 9934
rect 12292 9931 12388 9933
rect 12044 9904 12053 9924
rect 12073 9904 12163 9924
rect 12183 9904 12192 9924
rect 12044 9898 12192 9904
rect 12044 9895 12108 9898
rect 12044 9894 12081 9895
rect 12100 9868 12108 9895
rect 12129 9895 12192 9898
rect 12250 9924 12388 9931
rect 12250 9904 12259 9924
rect 12279 9904 12388 9924
rect 12250 9895 12388 9904
rect 12575 9920 12612 9999
rect 12653 9986 12763 9999
rect 12727 9930 12758 9931
rect 12575 9900 12584 9920
rect 12604 9900 12612 9920
rect 12129 9868 12136 9895
rect 12155 9894 12192 9895
rect 12251 9894 12288 9895
rect 12100 9843 12136 9868
rect 11571 9841 11612 9842
rect 11407 9834 11612 9841
rect 11407 9823 11581 9834
rect 9737 9768 9774 9769
rect 9687 9759 9774 9768
rect 9687 9739 9745 9759
rect 9765 9739 9774 9759
rect 9687 9729 9774 9739
rect 9833 9759 9870 9769
rect 9833 9739 9841 9759
rect 9861 9739 9870 9759
rect 9687 9728 9718 9729
rect 9682 9660 9792 9673
rect 9833 9660 9870 9739
rect 10144 9718 10209 9794
rect 11407 9790 11415 9823
rect 11408 9781 11415 9790
rect 11464 9814 11581 9823
rect 11601 9814 11612 9834
rect 11464 9806 11612 9814
rect 11679 9838 12038 9842
rect 11679 9833 12001 9838
rect 11679 9809 11792 9833
rect 11816 9814 12001 9833
rect 12025 9814 12038 9838
rect 11816 9809 12038 9814
rect 11679 9806 12038 9809
rect 12100 9806 12135 9843
rect 12203 9840 12303 9843
rect 12203 9836 12270 9840
rect 12203 9810 12215 9836
rect 12241 9814 12270 9836
rect 12296 9814 12303 9840
rect 12241 9810 12303 9814
rect 12203 9806 12303 9810
rect 11464 9790 11475 9806
rect 11464 9781 11472 9790
rect 11679 9785 11710 9806
rect 12100 9785 12136 9806
rect 11522 9784 11559 9785
rect 11187 9741 11252 9760
rect 11187 9723 11212 9741
rect 11230 9723 11252 9741
rect 9620 9658 9870 9660
rect 9620 9655 9721 9658
rect 9620 9636 9685 9655
rect 9682 9628 9685 9636
rect 9714 9628 9721 9655
rect 9749 9631 9759 9658
rect 9788 9636 9870 9658
rect 9893 9683 10210 9718
rect 9788 9631 9792 9636
rect 9749 9628 9792 9631
rect 9682 9614 9792 9628
rect 9108 9596 9449 9597
rect 9033 9594 9449 9596
rect 9893 9594 9933 9683
rect 10144 9656 10209 9683
rect 10144 9638 10167 9656
rect 10185 9638 10209 9656
rect 10144 9618 10209 9638
rect 9030 9591 9933 9594
rect 9030 9571 9036 9591
rect 9056 9571 9933 9591
rect 9030 9567 9933 9571
rect 9893 9564 9933 9567
rect 10145 9557 10210 9578
rect 8363 9549 9024 9550
rect 8363 9542 9297 9549
rect 8363 9541 9269 9542
rect 8363 9521 9214 9541
rect 9246 9522 9269 9541
rect 9294 9522 9297 9542
rect 9246 9521 9297 9522
rect 8363 9514 9297 9521
rect 7962 9472 8130 9473
rect 8365 9472 8404 9514
rect 9193 9512 9297 9514
rect 9262 9510 9297 9512
rect 10145 9539 10169 9557
rect 10187 9539 10210 9557
rect 10145 9492 10210 9539
rect 7962 9446 8406 9472
rect 7962 9444 8130 9446
rect 6723 8857 6727 8880
rect 6751 8857 6759 8880
rect 6923 8858 7022 8862
rect 6723 8836 6759 8857
rect 6723 8813 6727 8836
rect 6751 8813 6759 8836
rect 6723 8809 6759 8813
rect 6919 8852 7022 8858
rect 6919 8814 6945 8852
rect 6970 8817 6989 8852
rect 7014 8817 7022 8852
rect 6970 8814 7022 8817
rect 6919 8806 7022 8814
rect 6919 8805 7021 8806
rect 6515 8727 6683 8728
rect 6919 8727 6966 8805
rect 6515 8701 6966 8727
rect 6515 8699 6683 8701
rect 6515 8326 6542 8699
rect 6712 8651 6798 8660
rect 6712 8633 6731 8651
rect 6783 8633 6798 8651
rect 6712 8629 6798 8633
rect 6582 8466 6646 8478
rect 6582 8465 6617 8466
rect 6559 8460 6617 8465
rect 6559 8440 6562 8460
rect 6582 8446 6617 8460
rect 6637 8446 6646 8466
rect 6582 8438 6646 8446
rect 6608 8437 6646 8438
rect 6609 8436 6646 8437
rect 6712 8470 6748 8471
rect 6768 8470 6798 8629
rect 6919 8589 6966 8701
rect 6922 8474 6959 8589
rect 7187 8563 7298 8578
rect 7187 8561 7229 8563
rect 7187 8541 7194 8561
rect 7213 8541 7229 8561
rect 7187 8533 7229 8541
rect 7257 8561 7298 8563
rect 7257 8541 7271 8561
rect 7290 8541 7298 8561
rect 7257 8533 7298 8541
rect 7187 8527 7298 8533
rect 7130 8505 7379 8527
rect 7130 8474 7167 8505
rect 7343 8503 7379 8505
rect 7343 8474 7380 8503
rect 7584 8490 7663 9075
rect 7760 8623 7839 9223
rect 7962 9093 7989 9444
rect 8365 9440 8406 9446
rect 8029 9233 8093 9245
rect 8369 9241 8406 9440
rect 8868 9467 8940 9484
rect 8868 9428 8876 9467
rect 8921 9428 8940 9467
rect 8634 9330 8745 9345
rect 8634 9328 8676 9330
rect 8634 9308 8641 9328
rect 8660 9308 8676 9328
rect 8634 9300 8676 9308
rect 8704 9328 8745 9330
rect 8704 9308 8718 9328
rect 8737 9308 8745 9328
rect 8704 9300 8745 9308
rect 8634 9294 8745 9300
rect 8577 9272 8826 9294
rect 8577 9241 8614 9272
rect 8790 9270 8826 9272
rect 8790 9241 8827 9270
rect 8029 9232 8064 9233
rect 8006 9227 8064 9232
rect 8006 9207 8009 9227
rect 8029 9213 8064 9227
rect 8084 9213 8093 9233
rect 8029 9205 8093 9213
rect 8055 9204 8093 9205
rect 8056 9203 8093 9204
rect 8159 9237 8195 9238
rect 8267 9237 8303 9238
rect 8159 9229 8303 9237
rect 8159 9209 8167 9229
rect 8187 9209 8275 9229
rect 8295 9209 8303 9229
rect 8159 9203 8303 9209
rect 8369 9233 8407 9241
rect 8475 9237 8511 9238
rect 8369 9213 8378 9233
rect 8398 9213 8407 9233
rect 8369 9204 8407 9213
rect 8426 9230 8511 9237
rect 8426 9210 8433 9230
rect 8454 9229 8511 9230
rect 8454 9210 8483 9229
rect 8426 9209 8483 9210
rect 8503 9209 8511 9229
rect 8369 9203 8406 9204
rect 8426 9203 8511 9209
rect 8577 9233 8615 9241
rect 8688 9237 8724 9238
rect 8577 9213 8586 9233
rect 8606 9213 8615 9233
rect 8577 9204 8615 9213
rect 8639 9229 8724 9237
rect 8639 9209 8696 9229
rect 8716 9209 8724 9229
rect 8577 9203 8614 9204
rect 8639 9203 8724 9209
rect 8790 9233 8828 9241
rect 8790 9213 8799 9233
rect 8819 9213 8828 9233
rect 8790 9204 8828 9213
rect 8868 9218 8940 9428
rect 9010 9462 10210 9492
rect 9010 9461 9454 9462
rect 9010 9459 9178 9461
rect 8868 9204 8951 9218
rect 8790 9203 8827 9204
rect 8213 9182 8249 9203
rect 8639 9182 8670 9203
rect 8868 9182 8885 9204
rect 8046 9178 8146 9182
rect 8046 9174 8108 9178
rect 8046 9148 8053 9174
rect 8079 9152 8108 9174
rect 8134 9152 8146 9178
rect 8079 9148 8146 9152
rect 8046 9145 8146 9148
rect 8214 9145 8249 9182
rect 8311 9179 8670 9182
rect 8311 9174 8533 9179
rect 8311 9150 8324 9174
rect 8348 9155 8533 9174
rect 8557 9155 8670 9179
rect 8348 9150 8670 9155
rect 8311 9146 8670 9150
rect 8737 9174 8885 9182
rect 8737 9154 8748 9174
rect 8768 9171 8885 9174
rect 8938 9171 8951 9204
rect 8768 9154 8951 9171
rect 8737 9147 8951 9154
rect 8737 9146 8778 9147
rect 8868 9146 8951 9147
rect 8213 9120 8249 9145
rect 8061 9093 8098 9094
rect 8157 9093 8194 9094
rect 8213 9093 8220 9120
rect 7961 9084 8099 9093
rect 7961 9064 8070 9084
rect 8090 9064 8099 9084
rect 7961 9057 8099 9064
rect 8157 9090 8220 9093
rect 8241 9093 8249 9120
rect 8268 9093 8305 9094
rect 8241 9090 8305 9093
rect 8157 9084 8305 9090
rect 8157 9064 8166 9084
rect 8186 9064 8276 9084
rect 8296 9064 8305 9084
rect 7961 9055 8057 9057
rect 8157 9054 8305 9064
rect 8364 9084 8401 9094
rect 8476 9093 8513 9094
rect 8457 9091 8513 9093
rect 8364 9064 8372 9084
rect 8392 9064 8401 9084
rect 8213 9053 8249 9054
rect 8061 8922 8098 8923
rect 8364 8922 8401 9064
rect 8426 9084 8513 9091
rect 8426 9081 8484 9084
rect 8426 9061 8431 9081
rect 8452 9064 8484 9081
rect 8504 9064 8513 9084
rect 8452 9061 8513 9064
rect 8426 9054 8513 9061
rect 8572 9084 8609 9094
rect 8572 9064 8580 9084
rect 8600 9064 8609 9084
rect 8426 9053 8457 9054
rect 8572 8985 8609 9064
rect 8639 9093 8670 9146
rect 8876 9113 8890 9146
rect 8943 9113 8951 9146
rect 8876 9107 8951 9113
rect 8876 9102 8946 9107
rect 8689 9093 8726 9094
rect 8639 9084 8726 9093
rect 8639 9064 8697 9084
rect 8717 9064 8726 9084
rect 8639 9054 8726 9064
rect 8785 9084 8822 9094
rect 9010 9089 9037 9459
rect 9077 9229 9141 9241
rect 9417 9237 9454 9461
rect 9925 9442 9989 9444
rect 9921 9430 9989 9442
rect 9921 9397 9932 9430
rect 9972 9397 9989 9430
rect 9921 9387 9989 9397
rect 9682 9326 9793 9341
rect 9682 9324 9724 9326
rect 9682 9304 9689 9324
rect 9708 9304 9724 9324
rect 9682 9296 9724 9304
rect 9752 9324 9793 9326
rect 9752 9304 9766 9324
rect 9785 9304 9793 9324
rect 9752 9296 9793 9304
rect 9682 9290 9793 9296
rect 9625 9268 9874 9290
rect 9625 9237 9662 9268
rect 9838 9266 9874 9268
rect 9838 9237 9875 9266
rect 9077 9228 9112 9229
rect 9054 9223 9112 9228
rect 9054 9203 9057 9223
rect 9077 9209 9112 9223
rect 9132 9209 9141 9229
rect 9077 9201 9141 9209
rect 9103 9200 9141 9201
rect 9104 9199 9141 9200
rect 9207 9233 9243 9234
rect 9315 9233 9351 9234
rect 9207 9225 9351 9233
rect 9207 9205 9215 9225
rect 9235 9205 9323 9225
rect 9343 9205 9351 9225
rect 9207 9199 9351 9205
rect 9417 9229 9455 9237
rect 9523 9233 9559 9234
rect 9417 9209 9426 9229
rect 9446 9209 9455 9229
rect 9417 9200 9455 9209
rect 9474 9226 9559 9233
rect 9474 9206 9481 9226
rect 9502 9225 9559 9226
rect 9502 9206 9531 9225
rect 9474 9205 9531 9206
rect 9551 9205 9559 9225
rect 9417 9199 9454 9200
rect 9474 9199 9559 9205
rect 9625 9229 9663 9237
rect 9736 9233 9772 9234
rect 9625 9209 9634 9229
rect 9654 9209 9663 9229
rect 9625 9200 9663 9209
rect 9687 9225 9772 9233
rect 9687 9205 9744 9225
rect 9764 9205 9772 9225
rect 9625 9199 9662 9200
rect 9687 9199 9772 9205
rect 9838 9229 9876 9237
rect 9838 9209 9847 9229
rect 9867 9209 9876 9229
rect 9838 9200 9876 9209
rect 9925 9203 9989 9387
rect 10145 9261 10210 9462
rect 11187 9522 11252 9723
rect 11408 9597 11472 9781
rect 11521 9775 11559 9784
rect 11521 9755 11530 9775
rect 11550 9755 11559 9775
rect 11521 9747 11559 9755
rect 11625 9779 11710 9785
rect 11735 9784 11772 9785
rect 11625 9759 11633 9779
rect 11653 9759 11710 9779
rect 11625 9751 11710 9759
rect 11734 9775 11772 9784
rect 11734 9755 11743 9775
rect 11763 9755 11772 9775
rect 11625 9750 11661 9751
rect 11734 9747 11772 9755
rect 11838 9779 11923 9785
rect 11943 9784 11980 9785
rect 11838 9759 11846 9779
rect 11866 9778 11923 9779
rect 11866 9759 11895 9778
rect 11838 9758 11895 9759
rect 11916 9758 11923 9778
rect 11838 9751 11923 9758
rect 11942 9775 11980 9784
rect 11942 9755 11951 9775
rect 11971 9755 11980 9775
rect 11838 9750 11874 9751
rect 11942 9747 11980 9755
rect 12046 9779 12190 9785
rect 12046 9759 12054 9779
rect 12074 9759 12162 9779
rect 12182 9759 12190 9779
rect 12046 9751 12190 9759
rect 12046 9750 12082 9751
rect 12154 9750 12190 9751
rect 12256 9784 12293 9785
rect 12256 9783 12294 9784
rect 12256 9775 12320 9783
rect 12256 9755 12265 9775
rect 12285 9761 12320 9775
rect 12340 9761 12343 9781
rect 12285 9756 12343 9761
rect 12285 9755 12320 9756
rect 11522 9718 11559 9747
rect 11523 9716 11559 9718
rect 11735 9716 11772 9747
rect 11523 9694 11772 9716
rect 11604 9688 11715 9694
rect 11604 9680 11645 9688
rect 11604 9660 11612 9680
rect 11631 9660 11645 9680
rect 11604 9658 11645 9660
rect 11673 9680 11715 9688
rect 11673 9660 11689 9680
rect 11708 9660 11715 9680
rect 11673 9658 11715 9660
rect 11604 9643 11715 9658
rect 11408 9587 11476 9597
rect 11408 9554 11425 9587
rect 11465 9554 11476 9587
rect 11408 9542 11476 9554
rect 11408 9540 11472 9542
rect 11943 9523 11980 9747
rect 12256 9743 12320 9755
rect 12360 9525 12387 9895
rect 12575 9890 12612 9900
rect 12671 9920 12758 9930
rect 12671 9900 12680 9920
rect 12700 9900 12758 9920
rect 12671 9891 12758 9900
rect 12671 9890 12708 9891
rect 12451 9877 12521 9882
rect 12446 9871 12521 9877
rect 12446 9838 12454 9871
rect 12507 9838 12521 9871
rect 12727 9838 12758 9891
rect 12788 9920 12825 9999
rect 12940 9930 12971 9931
rect 12788 9900 12797 9920
rect 12817 9900 12825 9920
rect 12788 9890 12825 9900
rect 12884 9923 12971 9930
rect 12884 9920 12945 9923
rect 12884 9900 12893 9920
rect 12913 9903 12945 9920
rect 12966 9903 12971 9923
rect 12913 9900 12971 9903
rect 12884 9893 12971 9900
rect 12996 9920 13033 10062
rect 13299 10061 13336 10062
rect 13148 9930 13184 9931
rect 12996 9900 13005 9920
rect 13025 9900 13033 9920
rect 12884 9891 12940 9893
rect 12884 9890 12921 9891
rect 12996 9890 13033 9900
rect 13092 9920 13240 9930
rect 13340 9927 13436 9929
rect 13092 9900 13101 9920
rect 13121 9900 13211 9920
rect 13231 9900 13240 9920
rect 13092 9894 13240 9900
rect 13092 9891 13156 9894
rect 13092 9890 13129 9891
rect 13148 9864 13156 9891
rect 13177 9891 13240 9894
rect 13298 9920 13436 9927
rect 13298 9900 13307 9920
rect 13327 9900 13436 9920
rect 13298 9891 13436 9900
rect 13177 9864 13184 9891
rect 13203 9890 13240 9891
rect 13299 9890 13336 9891
rect 13148 9839 13184 9864
rect 12446 9837 12529 9838
rect 12619 9837 12660 9838
rect 12446 9830 12660 9837
rect 12446 9813 12629 9830
rect 12446 9780 12459 9813
rect 12512 9810 12629 9813
rect 12649 9810 12660 9830
rect 12512 9802 12660 9810
rect 12727 9834 13086 9838
rect 12727 9829 13049 9834
rect 12727 9805 12840 9829
rect 12864 9810 13049 9829
rect 13073 9810 13086 9834
rect 12864 9805 13086 9810
rect 12727 9802 13086 9805
rect 13148 9802 13183 9839
rect 13251 9836 13351 9839
rect 13251 9832 13318 9836
rect 13251 9806 13263 9832
rect 13289 9810 13318 9832
rect 13344 9810 13351 9836
rect 13289 9806 13351 9810
rect 13251 9802 13351 9806
rect 12512 9780 12529 9802
rect 12727 9781 12758 9802
rect 13148 9781 13184 9802
rect 12570 9780 12607 9781
rect 12446 9766 12529 9780
rect 12219 9523 12387 9525
rect 11943 9522 12387 9523
rect 11187 9492 12387 9522
rect 12457 9556 12529 9766
rect 12569 9771 12607 9780
rect 12569 9751 12578 9771
rect 12598 9751 12607 9771
rect 12569 9743 12607 9751
rect 12673 9775 12758 9781
rect 12783 9780 12820 9781
rect 12673 9755 12681 9775
rect 12701 9755 12758 9775
rect 12673 9747 12758 9755
rect 12782 9771 12820 9780
rect 12782 9751 12791 9771
rect 12811 9751 12820 9771
rect 12673 9746 12709 9747
rect 12782 9743 12820 9751
rect 12886 9775 12971 9781
rect 12991 9780 13028 9781
rect 12886 9755 12894 9775
rect 12914 9774 12971 9775
rect 12914 9755 12943 9774
rect 12886 9754 12943 9755
rect 12964 9754 12971 9774
rect 12886 9747 12971 9754
rect 12990 9771 13028 9780
rect 12990 9751 12999 9771
rect 13019 9751 13028 9771
rect 12886 9746 12922 9747
rect 12990 9743 13028 9751
rect 13094 9775 13238 9781
rect 13094 9755 13102 9775
rect 13122 9755 13210 9775
rect 13230 9755 13238 9775
rect 13094 9747 13238 9755
rect 13094 9746 13130 9747
rect 13202 9746 13238 9747
rect 13304 9780 13341 9781
rect 13304 9779 13342 9780
rect 13304 9771 13368 9779
rect 13304 9751 13313 9771
rect 13333 9757 13368 9771
rect 13388 9757 13391 9777
rect 13333 9752 13391 9757
rect 13333 9751 13368 9752
rect 12570 9714 12607 9743
rect 12571 9712 12607 9714
rect 12783 9712 12820 9743
rect 12571 9690 12820 9712
rect 12652 9684 12763 9690
rect 12652 9676 12693 9684
rect 12652 9656 12660 9676
rect 12679 9656 12693 9676
rect 12652 9654 12693 9656
rect 12721 9676 12763 9684
rect 12721 9656 12737 9676
rect 12756 9656 12763 9676
rect 12721 9654 12763 9656
rect 12652 9639 12763 9654
rect 12457 9517 12476 9556
rect 12521 9517 12529 9556
rect 12457 9500 12529 9517
rect 12991 9544 13028 9743
rect 13304 9739 13368 9751
rect 12991 9538 13032 9544
rect 13408 9540 13435 9891
rect 13564 9843 13635 10322
rect 13564 9759 13633 9843
rect 13267 9538 13435 9540
rect 12991 9512 13435 9538
rect 11187 9445 11252 9492
rect 11187 9427 11210 9445
rect 11228 9427 11252 9445
rect 12100 9472 12135 9474
rect 12100 9470 12204 9472
rect 12993 9470 13032 9512
rect 13267 9511 13435 9512
rect 12100 9463 13034 9470
rect 12100 9462 12151 9463
rect 12100 9442 12103 9462
rect 12128 9443 12151 9462
rect 12183 9443 13034 9463
rect 12128 9442 13034 9443
rect 12100 9435 13034 9442
rect 12373 9434 13034 9435
rect 11187 9406 11252 9427
rect 11464 9417 11504 9420
rect 11464 9413 12367 9417
rect 11464 9393 12341 9413
rect 12361 9393 12367 9413
rect 11464 9390 12367 9393
rect 11188 9346 11253 9366
rect 11188 9328 11212 9346
rect 11230 9328 11253 9346
rect 11188 9301 11253 9328
rect 11464 9301 11504 9390
rect 11948 9388 12364 9390
rect 11948 9387 12289 9388
rect 11605 9356 11715 9370
rect 11605 9353 11648 9356
rect 11605 9348 11609 9353
rect 11187 9266 11504 9301
rect 11527 9326 11609 9348
rect 11638 9326 11648 9353
rect 11676 9329 11683 9356
rect 11712 9348 11715 9356
rect 11712 9329 11777 9348
rect 11676 9326 11777 9329
rect 11527 9324 11777 9326
rect 10145 9243 10167 9261
rect 10185 9243 10210 9261
rect 10145 9224 10210 9243
rect 9838 9199 9875 9200
rect 9261 9178 9297 9199
rect 9687 9178 9718 9199
rect 9925 9194 9933 9203
rect 9922 9178 9933 9194
rect 9094 9174 9194 9178
rect 9094 9170 9156 9174
rect 9094 9144 9101 9170
rect 9127 9148 9156 9170
rect 9182 9148 9194 9174
rect 9127 9144 9194 9148
rect 9094 9141 9194 9144
rect 9262 9141 9297 9178
rect 9359 9175 9718 9178
rect 9359 9170 9581 9175
rect 9359 9146 9372 9170
rect 9396 9151 9581 9170
rect 9605 9151 9718 9175
rect 9396 9146 9718 9151
rect 9359 9142 9718 9146
rect 9785 9170 9933 9178
rect 9785 9150 9796 9170
rect 9816 9161 9933 9170
rect 9982 9194 9989 9203
rect 9982 9161 9990 9194
rect 11188 9190 11253 9266
rect 11527 9245 11564 9324
rect 11605 9311 11715 9324
rect 11679 9255 11710 9256
rect 11527 9225 11536 9245
rect 11556 9225 11564 9245
rect 11527 9215 11564 9225
rect 11623 9245 11710 9255
rect 11623 9225 11632 9245
rect 11652 9225 11710 9245
rect 11623 9216 11710 9225
rect 11623 9215 11660 9216
rect 9816 9150 9990 9161
rect 9785 9143 9990 9150
rect 9785 9142 9826 9143
rect 9261 9116 9297 9141
rect 9109 9089 9146 9090
rect 9205 9089 9242 9090
rect 9261 9089 9268 9116
rect 8785 9064 8793 9084
rect 8813 9064 8822 9084
rect 8639 9053 8670 9054
rect 8634 8985 8744 8998
rect 8785 8985 8822 9064
rect 9009 9080 9147 9089
rect 9009 9060 9118 9080
rect 9138 9060 9147 9080
rect 9009 9053 9147 9060
rect 9205 9086 9268 9089
rect 9289 9089 9297 9116
rect 9316 9089 9353 9090
rect 9289 9086 9353 9089
rect 9205 9080 9353 9086
rect 9205 9060 9214 9080
rect 9234 9060 9324 9080
rect 9344 9060 9353 9080
rect 9009 9051 9105 9053
rect 9205 9050 9353 9060
rect 9412 9080 9449 9090
rect 9524 9089 9561 9090
rect 9505 9087 9561 9089
rect 9412 9060 9420 9080
rect 9440 9060 9449 9080
rect 9261 9049 9297 9050
rect 8572 8983 8822 8985
rect 8572 8980 8673 8983
rect 8572 8961 8637 8980
rect 8634 8953 8637 8961
rect 8666 8953 8673 8980
rect 8701 8956 8711 8983
rect 8740 8961 8822 8983
rect 8740 8956 8744 8961
rect 8701 8953 8744 8956
rect 8634 8939 8744 8953
rect 8060 8921 8401 8922
rect 7985 8916 8401 8921
rect 9109 8918 9146 8919
rect 9412 8918 9449 9060
rect 9474 9080 9561 9087
rect 9474 9077 9532 9080
rect 9474 9057 9479 9077
rect 9500 9060 9532 9077
rect 9552 9060 9561 9080
rect 9500 9057 9561 9060
rect 9474 9050 9561 9057
rect 9620 9080 9657 9090
rect 9620 9060 9628 9080
rect 9648 9060 9657 9080
rect 9474 9049 9505 9050
rect 9620 8981 9657 9060
rect 9687 9089 9718 9142
rect 9922 9140 9990 9143
rect 9922 9098 9934 9140
rect 9983 9098 9990 9140
rect 9737 9089 9774 9090
rect 9687 9080 9774 9089
rect 9687 9060 9745 9080
rect 9765 9060 9774 9080
rect 9687 9050 9774 9060
rect 9833 9080 9870 9090
rect 9922 9085 9990 9098
rect 10145 9162 10210 9179
rect 10145 9144 10169 9162
rect 10187 9144 10210 9162
rect 11188 9172 11210 9190
rect 11228 9172 11253 9190
rect 11188 9151 11253 9172
rect 11401 9170 11466 9179
rect 9833 9060 9841 9080
rect 9861 9060 9870 9080
rect 9687 9049 9718 9050
rect 9682 8981 9792 8994
rect 9833 8981 9870 9060
rect 10145 9005 10210 9144
rect 11401 9133 11411 9170
rect 11451 9162 11466 9170
rect 11679 9163 11710 9216
rect 11740 9245 11777 9324
rect 11892 9255 11923 9256
rect 11740 9225 11749 9245
rect 11769 9225 11777 9245
rect 11740 9215 11777 9225
rect 11836 9248 11923 9255
rect 11836 9245 11897 9248
rect 11836 9225 11845 9245
rect 11865 9228 11897 9245
rect 11918 9228 11923 9248
rect 11865 9225 11923 9228
rect 11836 9218 11923 9225
rect 11948 9245 11985 9387
rect 12251 9386 12288 9387
rect 12100 9255 12136 9256
rect 11948 9225 11957 9245
rect 11977 9225 11985 9245
rect 11836 9216 11892 9218
rect 11836 9215 11873 9216
rect 11948 9215 11985 9225
rect 12044 9245 12192 9255
rect 12292 9252 12388 9254
rect 12044 9225 12053 9245
rect 12073 9225 12163 9245
rect 12183 9225 12192 9245
rect 12044 9219 12192 9225
rect 12044 9216 12108 9219
rect 12044 9215 12081 9216
rect 12100 9189 12108 9216
rect 12129 9216 12192 9219
rect 12250 9245 12388 9252
rect 12250 9225 12259 9245
rect 12279 9225 12388 9245
rect 13568 9243 13630 9759
rect 12250 9216 12388 9225
rect 12129 9189 12136 9216
rect 12155 9215 12192 9216
rect 12251 9215 12288 9216
rect 12100 9164 12136 9189
rect 11571 9162 11612 9163
rect 11451 9155 11612 9162
rect 11451 9135 11581 9155
rect 11601 9135 11612 9155
rect 11451 9133 11612 9135
rect 11401 9127 11612 9133
rect 11679 9159 12038 9163
rect 11679 9154 12001 9159
rect 11679 9130 11792 9154
rect 11816 9135 12001 9154
rect 12025 9135 12038 9159
rect 11816 9130 12038 9135
rect 11679 9127 12038 9130
rect 12100 9127 12135 9164
rect 12203 9161 12303 9164
rect 12203 9157 12270 9161
rect 12203 9131 12215 9157
rect 12241 9135 12270 9157
rect 12296 9135 12303 9161
rect 12241 9131 12303 9135
rect 12203 9127 12303 9131
rect 11401 9114 11468 9127
rect 10145 8999 10167 9005
rect 9620 8979 9870 8981
rect 9620 8976 9721 8979
rect 9620 8957 9685 8976
rect 9682 8949 9685 8957
rect 9714 8949 9721 8976
rect 9749 8952 9759 8979
rect 9788 8957 9870 8979
rect 9899 8987 10167 8999
rect 10185 8987 10210 9005
rect 9899 8964 10210 8987
rect 11193 9091 11249 9111
rect 11193 9073 11212 9091
rect 11230 9073 11249 9091
rect 9899 8963 9954 8964
rect 9788 8952 9792 8957
rect 9749 8949 9792 8952
rect 9682 8935 9792 8949
rect 9108 8917 9449 8918
rect 7985 8896 7988 8916
rect 8008 8896 8401 8916
rect 9033 8916 9449 8917
rect 9899 8916 9942 8963
rect 11193 8960 11249 9073
rect 11401 9093 11415 9114
rect 11451 9093 11468 9114
rect 11679 9106 11710 9127
rect 12100 9106 12136 9127
rect 11522 9105 11559 9106
rect 11401 9086 11468 9093
rect 11521 9096 11559 9105
rect 9033 8912 9942 8916
rect 8352 8863 8397 8896
rect 9033 8892 9036 8912
rect 9056 8892 9942 8912
rect 9410 8887 9942 8892
rect 10150 8906 10209 8928
rect 10150 8888 10169 8906
rect 10187 8888 10209 8906
rect 9198 8863 9297 8865
rect 8352 8853 9297 8863
rect 8352 8827 9220 8853
rect 8353 8826 9220 8827
rect 9198 8815 9220 8826
rect 9245 8818 9264 8853
rect 9289 8818 9297 8853
rect 9245 8815 9297 8818
rect 10150 8817 10209 8888
rect 11193 8822 11248 8960
rect 11401 8934 11466 9086
rect 11521 9076 11530 9096
rect 11550 9076 11559 9096
rect 11521 9068 11559 9076
rect 11625 9100 11710 9106
rect 11735 9105 11772 9106
rect 11625 9080 11633 9100
rect 11653 9080 11710 9100
rect 11625 9072 11710 9080
rect 11734 9096 11772 9105
rect 11734 9076 11743 9096
rect 11763 9076 11772 9096
rect 11625 9071 11661 9072
rect 11734 9068 11772 9076
rect 11838 9100 11923 9106
rect 11943 9105 11980 9106
rect 11838 9080 11846 9100
rect 11866 9099 11923 9100
rect 11866 9080 11895 9099
rect 11838 9079 11895 9080
rect 11916 9079 11923 9099
rect 11838 9072 11923 9079
rect 11942 9096 11980 9105
rect 11942 9076 11951 9096
rect 11971 9076 11980 9096
rect 11838 9071 11874 9072
rect 11942 9068 11980 9076
rect 12046 9100 12190 9106
rect 12046 9080 12054 9100
rect 12074 9080 12162 9100
rect 12182 9080 12190 9100
rect 12046 9072 12190 9080
rect 12046 9071 12082 9072
rect 12154 9071 12190 9072
rect 12256 9105 12293 9106
rect 12256 9104 12294 9105
rect 12256 9096 12320 9104
rect 12256 9076 12265 9096
rect 12285 9082 12320 9096
rect 12340 9082 12343 9102
rect 12285 9077 12343 9082
rect 12285 9076 12320 9077
rect 11522 9039 11559 9068
rect 11523 9037 11559 9039
rect 11735 9037 11772 9068
rect 11523 9015 11772 9037
rect 11604 9009 11715 9015
rect 11604 9001 11645 9009
rect 11604 8981 11612 9001
rect 11631 8981 11645 9001
rect 11604 8979 11645 8981
rect 11673 9001 11715 9009
rect 11673 8981 11689 9001
rect 11708 8981 11715 9001
rect 11673 8979 11715 8981
rect 11604 8966 11715 8979
rect 11943 8969 11980 9068
rect 12256 9064 12320 9076
rect 11394 8924 11515 8934
rect 11394 8922 11463 8924
rect 11394 8881 11407 8922
rect 11444 8883 11463 8922
rect 11500 8883 11515 8924
rect 11444 8881 11515 8883
rect 11394 8863 11515 8881
rect 11186 8819 11250 8822
rect 11606 8819 11710 8825
rect 11941 8819 11982 8969
rect 12360 8961 12387 9216
rect 12449 9206 12529 9217
rect 12449 9180 12466 9206
rect 12506 9180 12529 9206
rect 12449 9153 12529 9180
rect 12449 9127 12470 9153
rect 12510 9127 12529 9153
rect 12449 9108 12529 9127
rect 12449 9082 12473 9108
rect 12513 9082 12529 9108
rect 12449 9031 12529 9082
rect 13552 9208 13630 9243
rect 13552 9146 13634 9208
rect 13552 9123 13580 9146
rect 13606 9123 13634 9146
rect 13552 9103 13634 9123
rect 9198 8807 9297 8815
rect 9224 8806 9296 8807
rect 8878 8780 8945 8799
rect 8878 8759 8895 8780
rect 7759 8581 7839 8623
rect 8876 8714 8895 8759
rect 8925 8759 8945 8780
rect 8925 8714 8946 8759
rect 9415 8756 9456 8758
rect 9687 8756 9791 8758
rect 10147 8756 10211 8817
rect 6820 8470 6856 8471
rect 6712 8462 6856 8470
rect 6712 8442 6720 8462
rect 6740 8442 6828 8462
rect 6848 8442 6856 8462
rect 6712 8436 6856 8442
rect 6922 8466 6960 8474
rect 7028 8470 7064 8471
rect 6922 8446 6931 8466
rect 6951 8446 6960 8466
rect 6922 8437 6960 8446
rect 6979 8463 7064 8470
rect 6979 8443 6986 8463
rect 7007 8462 7064 8463
rect 7007 8443 7036 8462
rect 6979 8442 7036 8443
rect 7056 8442 7064 8462
rect 6922 8436 6959 8437
rect 6979 8436 7064 8442
rect 7130 8466 7168 8474
rect 7241 8470 7277 8471
rect 7130 8446 7139 8466
rect 7159 8446 7168 8466
rect 7130 8437 7168 8446
rect 7192 8462 7277 8470
rect 7192 8442 7249 8462
rect 7269 8442 7277 8462
rect 7130 8436 7167 8437
rect 7192 8436 7277 8442
rect 7343 8466 7381 8474
rect 7343 8446 7352 8466
rect 7372 8446 7381 8466
rect 7343 8437 7381 8446
rect 7581 8454 7667 8490
rect 7343 8436 7380 8437
rect 6766 8415 6802 8436
rect 7192 8415 7223 8436
rect 7419 8415 7465 8419
rect 6599 8411 6699 8415
rect 6599 8407 6661 8411
rect 6599 8381 6606 8407
rect 6632 8385 6661 8407
rect 6687 8385 6699 8411
rect 6632 8381 6699 8385
rect 6599 8378 6699 8381
rect 6767 8378 6802 8415
rect 6864 8412 7223 8415
rect 6864 8407 7086 8412
rect 6864 8383 6877 8407
rect 6901 8388 7086 8407
rect 7110 8388 7223 8412
rect 6901 8383 7223 8388
rect 6864 8379 7223 8383
rect 7290 8407 7465 8415
rect 7290 8387 7301 8407
rect 7321 8387 7465 8407
rect 7581 8413 7598 8454
rect 7652 8413 7667 8454
rect 7581 8394 7667 8413
rect 7290 8380 7465 8387
rect 7290 8379 7331 8380
rect 6766 8353 6802 8378
rect 6614 8326 6651 8327
rect 6710 8326 6747 8327
rect 6766 8326 6773 8353
rect 6514 8317 6652 8326
rect 6514 8297 6623 8317
rect 6643 8297 6652 8317
rect 6514 8290 6652 8297
rect 6710 8323 6773 8326
rect 6794 8326 6802 8353
rect 6821 8326 6858 8327
rect 6794 8323 6858 8326
rect 6710 8317 6858 8323
rect 6710 8297 6719 8317
rect 6739 8297 6829 8317
rect 6849 8297 6858 8317
rect 6514 8288 6610 8290
rect 6710 8287 6858 8297
rect 6917 8317 6954 8327
rect 7029 8326 7066 8327
rect 7010 8324 7066 8326
rect 6917 8297 6925 8317
rect 6945 8297 6954 8317
rect 6766 8286 6802 8287
rect 6614 8155 6651 8156
rect 6917 8155 6954 8297
rect 6979 8317 7066 8324
rect 6979 8314 7037 8317
rect 6979 8294 6984 8314
rect 7005 8297 7037 8314
rect 7057 8297 7066 8317
rect 7005 8294 7066 8297
rect 6979 8287 7066 8294
rect 7125 8317 7162 8327
rect 7125 8297 7133 8317
rect 7153 8297 7162 8317
rect 6979 8286 7010 8287
rect 7125 8218 7162 8297
rect 7192 8326 7223 8379
rect 7242 8326 7279 8327
rect 7192 8317 7279 8326
rect 7192 8297 7250 8317
rect 7270 8297 7279 8317
rect 7192 8287 7279 8297
rect 7338 8317 7375 8327
rect 7338 8297 7346 8317
rect 7366 8297 7375 8317
rect 7192 8286 7223 8287
rect 7187 8218 7297 8231
rect 7338 8218 7375 8297
rect 7419 8297 7465 8380
rect 7759 8297 7834 8581
rect 8876 8506 8946 8714
rect 9008 8721 10211 8756
rect 9008 8707 9036 8721
rect 9010 8576 9036 8707
rect 9415 8718 10211 8721
rect 11186 8816 11982 8819
rect 12361 8830 12387 8961
rect 12361 8816 12389 8830
rect 11186 8781 12389 8816
rect 12451 8823 12521 9031
rect 11186 8720 11250 8781
rect 11606 8779 11710 8781
rect 11941 8779 11982 8781
rect 12451 8778 12472 8823
rect 12452 8757 12472 8778
rect 12502 8778 12521 8823
rect 12502 8757 12519 8778
rect 12452 8738 12519 8757
rect 12101 8730 12173 8731
rect 12100 8722 12199 8730
rect 8868 8455 8948 8506
rect 8868 8429 8884 8455
rect 8924 8429 8948 8455
rect 8868 8410 8948 8429
rect 8868 8384 8887 8410
rect 8927 8384 8948 8410
rect 8868 8357 8948 8384
rect 8868 8331 8891 8357
rect 8931 8331 8948 8357
rect 8868 8320 8948 8331
rect 9010 8321 9037 8576
rect 9415 8568 9456 8718
rect 9687 8712 9791 8718
rect 10147 8715 10211 8718
rect 9882 8656 10003 8674
rect 9882 8654 9953 8656
rect 9882 8613 9897 8654
rect 9934 8615 9953 8654
rect 9990 8615 10003 8656
rect 9934 8613 10003 8615
rect 9882 8603 10003 8613
rect 9077 8461 9141 8473
rect 9417 8469 9454 8568
rect 9682 8558 9793 8571
rect 9682 8556 9724 8558
rect 9682 8536 9689 8556
rect 9708 8536 9724 8556
rect 9682 8528 9724 8536
rect 9752 8556 9793 8558
rect 9752 8536 9766 8556
rect 9785 8536 9793 8556
rect 9752 8528 9793 8536
rect 9682 8522 9793 8528
rect 9625 8500 9874 8522
rect 9625 8469 9662 8500
rect 9838 8498 9874 8500
rect 9838 8469 9875 8498
rect 9077 8460 9112 8461
rect 9054 8455 9112 8460
rect 9054 8435 9057 8455
rect 9077 8441 9112 8455
rect 9132 8441 9141 8461
rect 9077 8433 9141 8441
rect 9103 8432 9141 8433
rect 9104 8431 9141 8432
rect 9207 8465 9243 8466
rect 9315 8465 9351 8466
rect 9207 8457 9351 8465
rect 9207 8437 9215 8457
rect 9235 8437 9323 8457
rect 9343 8437 9351 8457
rect 9207 8431 9351 8437
rect 9417 8461 9455 8469
rect 9523 8465 9559 8466
rect 9417 8441 9426 8461
rect 9446 8441 9455 8461
rect 9417 8432 9455 8441
rect 9474 8458 9559 8465
rect 9474 8438 9481 8458
rect 9502 8457 9559 8458
rect 9502 8438 9531 8457
rect 9474 8437 9531 8438
rect 9551 8437 9559 8457
rect 9417 8431 9454 8432
rect 9474 8431 9559 8437
rect 9625 8461 9663 8469
rect 9736 8465 9772 8466
rect 9625 8441 9634 8461
rect 9654 8441 9663 8461
rect 9625 8432 9663 8441
rect 9687 8457 9772 8465
rect 9687 8437 9744 8457
rect 9764 8437 9772 8457
rect 9625 8431 9662 8432
rect 9687 8431 9772 8437
rect 9838 8461 9876 8469
rect 9838 8441 9847 8461
rect 9867 8441 9876 8461
rect 9931 8451 9996 8603
rect 10149 8577 10204 8715
rect 11188 8649 11247 8720
rect 12100 8719 12152 8722
rect 12100 8684 12108 8719
rect 12133 8684 12152 8719
rect 12177 8711 12199 8722
rect 12177 8710 13044 8711
rect 12177 8684 13045 8710
rect 12100 8674 13045 8684
rect 12100 8672 12199 8674
rect 11188 8631 11210 8649
rect 11228 8631 11247 8649
rect 11188 8609 11247 8631
rect 11455 8645 11987 8650
rect 11455 8625 12341 8645
rect 12361 8625 12364 8645
rect 13000 8641 13045 8674
rect 11455 8621 12364 8625
rect 9838 8432 9876 8441
rect 9929 8444 9996 8451
rect 9838 8431 9875 8432
rect 9261 8410 9297 8431
rect 9687 8410 9718 8431
rect 9929 8423 9946 8444
rect 9982 8423 9996 8444
rect 10148 8464 10204 8577
rect 11455 8574 11498 8621
rect 11948 8620 12364 8621
rect 12996 8621 13389 8641
rect 13409 8621 13412 8641
rect 11948 8619 12289 8620
rect 11605 8588 11715 8602
rect 11605 8585 11648 8588
rect 11605 8580 11609 8585
rect 11443 8573 11498 8574
rect 10148 8446 10167 8464
rect 10185 8446 10204 8464
rect 10148 8426 10204 8446
rect 11187 8550 11498 8573
rect 11187 8532 11212 8550
rect 11230 8538 11498 8550
rect 11527 8558 11609 8580
rect 11638 8558 11648 8585
rect 11676 8561 11683 8588
rect 11712 8580 11715 8588
rect 11712 8561 11777 8580
rect 11676 8558 11777 8561
rect 11527 8556 11777 8558
rect 11230 8532 11252 8538
rect 9929 8410 9996 8423
rect 9094 8406 9194 8410
rect 9094 8402 9156 8406
rect 9094 8376 9101 8402
rect 9127 8380 9156 8402
rect 9182 8380 9194 8406
rect 9127 8376 9194 8380
rect 9094 8373 9194 8376
rect 9262 8373 9297 8410
rect 9359 8407 9718 8410
rect 9359 8402 9581 8407
rect 9359 8378 9372 8402
rect 9396 8383 9581 8402
rect 9605 8383 9718 8407
rect 9396 8378 9718 8383
rect 9359 8374 9718 8378
rect 9785 8404 9996 8410
rect 9785 8402 9946 8404
rect 9785 8382 9796 8402
rect 9816 8382 9946 8402
rect 9785 8375 9946 8382
rect 9785 8374 9826 8375
rect 9261 8348 9297 8373
rect 9109 8321 9146 8322
rect 9205 8321 9242 8322
rect 9261 8321 9268 8348
rect 7419 8262 7834 8297
rect 9009 8312 9147 8321
rect 9009 8292 9118 8312
rect 9138 8292 9147 8312
rect 9009 8285 9147 8292
rect 9205 8318 9268 8321
rect 9289 8321 9297 8348
rect 9316 8321 9353 8322
rect 9289 8318 9353 8321
rect 9205 8312 9353 8318
rect 9205 8292 9214 8312
rect 9234 8292 9324 8312
rect 9344 8292 9353 8312
rect 9009 8283 9105 8285
rect 9205 8282 9353 8292
rect 9412 8312 9449 8322
rect 9524 8321 9561 8322
rect 9505 8319 9561 8321
rect 9412 8292 9420 8312
rect 9440 8292 9449 8312
rect 9261 8281 9297 8282
rect 7419 8261 7465 8262
rect 7125 8216 7375 8218
rect 7125 8213 7226 8216
rect 7125 8194 7190 8213
rect 7187 8186 7190 8194
rect 7219 8186 7226 8213
rect 7254 8189 7264 8216
rect 7293 8194 7375 8216
rect 7759 8210 7834 8262
rect 7293 8189 7297 8194
rect 7254 8186 7297 8189
rect 7187 8172 7297 8186
rect 6613 8154 6954 8155
rect 6538 8149 6954 8154
rect 6538 8129 6541 8149
rect 6561 8129 6955 8149
rect 5595 7482 6401 7557
rect 4834 7438 4843 7472
rect 4872 7471 5282 7472
rect 4872 7438 4889 7471
rect 5114 7470 5282 7471
rect 4834 7412 4889 7438
rect 4834 7378 4842 7412
rect 4871 7378 4889 7412
rect 4834 7366 4889 7378
rect 3030 7321 3114 7342
rect 3030 7293 3058 7321
rect 3102 7293 3114 7321
rect 2844 7242 2918 7270
rect 2844 7194 2867 7242
rect 2904 7194 2918 7242
rect 3030 7264 3114 7293
rect 3030 7236 3055 7264
rect 3099 7236 3114 7264
rect 3030 7211 3114 7236
rect 5170 7225 5258 7229
rect 2844 7185 2918 7194
rect 477 7135 543 7183
rect 2854 7181 2918 7185
rect 5170 7208 5434 7225
rect 5170 7154 5350 7208
rect 5413 7154 5434 7208
rect 3067 7144 3778 7146
rect 2440 7143 3778 7144
rect 1390 7142 1462 7143
rect 477 7061 536 7135
rect 1389 7134 1488 7142
rect 1389 7131 1441 7134
rect 1389 7096 1397 7131
rect 1422 7096 1441 7131
rect 1466 7123 1488 7134
rect 2439 7135 3778 7143
rect 2439 7132 2491 7135
rect 1466 7122 2333 7123
rect 1466 7096 2334 7122
rect 1389 7086 2334 7096
rect 1389 7084 1488 7086
rect 477 7043 499 7061
rect 517 7043 536 7061
rect 477 7021 536 7043
rect 744 7057 1276 7062
rect 744 7037 1630 7057
rect 1650 7037 1653 7057
rect 2289 7053 2334 7086
rect 2439 7097 2447 7132
rect 2472 7097 2491 7132
rect 2516 7097 3778 7135
rect 2439 7088 3778 7097
rect 2439 7085 2528 7088
rect 3067 7086 3778 7088
rect 5170 7137 5434 7154
rect 744 7033 1653 7037
rect 744 6986 787 7033
rect 1237 7032 1653 7033
rect 2285 7033 2678 7053
rect 2698 7033 2701 7053
rect 1237 7031 1578 7032
rect 894 7000 1004 7014
rect 894 6997 937 7000
rect 894 6992 898 6997
rect 732 6985 787 6986
rect 476 6962 787 6985
rect 476 6944 501 6962
rect 519 6950 787 6962
rect 816 6970 898 6992
rect 927 6970 937 6997
rect 965 6973 972 7000
rect 1001 6992 1004 7000
rect 1001 6973 1066 6992
rect 965 6970 1066 6973
rect 816 6968 1066 6970
rect 519 6944 541 6950
rect 476 6805 541 6944
rect 816 6889 853 6968
rect 894 6955 1004 6968
rect 968 6899 999 6900
rect 816 6869 825 6889
rect 845 6869 853 6889
rect 476 6787 499 6805
rect 517 6787 541 6805
rect 476 6770 541 6787
rect 696 6851 764 6864
rect 816 6859 853 6869
rect 912 6889 999 6899
rect 912 6869 921 6889
rect 941 6869 999 6889
rect 912 6860 999 6869
rect 912 6859 949 6860
rect 696 6809 703 6851
rect 752 6809 764 6851
rect 696 6806 764 6809
rect 968 6807 999 6860
rect 1029 6889 1066 6968
rect 1181 6899 1212 6900
rect 1029 6869 1038 6889
rect 1058 6869 1066 6889
rect 1029 6859 1066 6869
rect 1125 6892 1212 6899
rect 1125 6889 1186 6892
rect 1125 6869 1134 6889
rect 1154 6872 1186 6889
rect 1207 6872 1212 6892
rect 1154 6869 1212 6872
rect 1125 6862 1212 6869
rect 1237 6889 1274 7031
rect 1540 7030 1577 7031
rect 2285 7028 2701 7033
rect 2285 7027 2626 7028
rect 1942 6996 2052 7010
rect 1942 6993 1985 6996
rect 1942 6988 1946 6993
rect 1864 6966 1946 6988
rect 1975 6966 1985 6993
rect 2013 6969 2020 6996
rect 2049 6988 2052 6996
rect 2049 6969 2114 6988
rect 2013 6966 2114 6969
rect 1864 6964 2114 6966
rect 1389 6899 1425 6900
rect 1237 6869 1246 6889
rect 1266 6869 1274 6889
rect 1125 6860 1181 6862
rect 1125 6859 1162 6860
rect 1237 6859 1274 6869
rect 1333 6889 1481 6899
rect 1581 6896 1677 6898
rect 1333 6869 1342 6889
rect 1362 6869 1452 6889
rect 1472 6869 1481 6889
rect 1333 6863 1481 6869
rect 1333 6860 1397 6863
rect 1333 6859 1370 6860
rect 1389 6833 1397 6860
rect 1418 6860 1481 6863
rect 1539 6889 1677 6896
rect 1539 6869 1548 6889
rect 1568 6869 1677 6889
rect 1539 6860 1677 6869
rect 1864 6885 1901 6964
rect 1942 6951 2052 6964
rect 2016 6895 2047 6896
rect 1864 6865 1873 6885
rect 1893 6865 1901 6885
rect 1418 6833 1425 6860
rect 1444 6859 1481 6860
rect 1540 6859 1577 6860
rect 1389 6808 1425 6833
rect 860 6806 901 6807
rect 696 6799 901 6806
rect 696 6788 870 6799
rect 696 6755 704 6788
rect 697 6746 704 6755
rect 753 6779 870 6788
rect 890 6779 901 6799
rect 753 6771 901 6779
rect 968 6803 1327 6807
rect 968 6798 1290 6803
rect 968 6774 1081 6798
rect 1105 6779 1290 6798
rect 1314 6779 1327 6803
rect 1105 6774 1327 6779
rect 968 6771 1327 6774
rect 1389 6771 1424 6808
rect 1492 6805 1592 6808
rect 1492 6801 1559 6805
rect 1492 6775 1504 6801
rect 1530 6779 1559 6801
rect 1585 6779 1592 6805
rect 1530 6775 1592 6779
rect 1492 6771 1592 6775
rect 753 6755 764 6771
rect 753 6746 761 6755
rect 968 6750 999 6771
rect 1389 6750 1425 6771
rect 811 6749 848 6750
rect 476 6706 541 6725
rect 476 6688 501 6706
rect 519 6688 541 6706
rect 476 6487 541 6688
rect 697 6562 761 6746
rect 810 6740 848 6749
rect 810 6720 819 6740
rect 839 6720 848 6740
rect 810 6712 848 6720
rect 914 6744 999 6750
rect 1024 6749 1061 6750
rect 914 6724 922 6744
rect 942 6724 999 6744
rect 914 6716 999 6724
rect 1023 6740 1061 6749
rect 1023 6720 1032 6740
rect 1052 6720 1061 6740
rect 914 6715 950 6716
rect 1023 6712 1061 6720
rect 1127 6744 1212 6750
rect 1232 6749 1269 6750
rect 1127 6724 1135 6744
rect 1155 6743 1212 6744
rect 1155 6724 1184 6743
rect 1127 6723 1184 6724
rect 1205 6723 1212 6743
rect 1127 6716 1212 6723
rect 1231 6740 1269 6749
rect 1231 6720 1240 6740
rect 1260 6720 1269 6740
rect 1127 6715 1163 6716
rect 1231 6712 1269 6720
rect 1335 6744 1479 6750
rect 1335 6724 1343 6744
rect 1363 6724 1451 6744
rect 1471 6724 1479 6744
rect 1335 6716 1479 6724
rect 1335 6715 1371 6716
rect 1443 6715 1479 6716
rect 1545 6749 1582 6750
rect 1545 6748 1583 6749
rect 1545 6740 1609 6748
rect 1545 6720 1554 6740
rect 1574 6726 1609 6740
rect 1629 6726 1632 6746
rect 1574 6721 1632 6726
rect 1574 6720 1609 6721
rect 811 6683 848 6712
rect 812 6681 848 6683
rect 1024 6681 1061 6712
rect 812 6659 1061 6681
rect 893 6653 1004 6659
rect 893 6645 934 6653
rect 893 6625 901 6645
rect 920 6625 934 6645
rect 893 6623 934 6625
rect 962 6645 1004 6653
rect 962 6625 978 6645
rect 997 6625 1004 6645
rect 962 6623 1004 6625
rect 893 6608 1004 6623
rect 697 6552 765 6562
rect 697 6519 714 6552
rect 754 6519 765 6552
rect 697 6507 765 6519
rect 697 6505 761 6507
rect 1232 6488 1269 6712
rect 1545 6708 1609 6720
rect 1649 6490 1676 6860
rect 1864 6855 1901 6865
rect 1960 6885 2047 6895
rect 1960 6865 1969 6885
rect 1989 6865 2047 6885
rect 1960 6856 2047 6865
rect 1960 6855 1997 6856
rect 1740 6842 1810 6847
rect 1735 6836 1810 6842
rect 1735 6803 1743 6836
rect 1796 6803 1810 6836
rect 2016 6803 2047 6856
rect 2077 6885 2114 6964
rect 2229 6895 2260 6896
rect 2077 6865 2086 6885
rect 2106 6865 2114 6885
rect 2077 6855 2114 6865
rect 2173 6888 2260 6895
rect 2173 6885 2234 6888
rect 2173 6865 2182 6885
rect 2202 6868 2234 6885
rect 2255 6868 2260 6888
rect 2202 6865 2260 6868
rect 2173 6858 2260 6865
rect 2285 6885 2322 7027
rect 2588 7026 2625 7027
rect 2437 6895 2473 6896
rect 2285 6865 2294 6885
rect 2314 6865 2322 6885
rect 2173 6856 2229 6858
rect 2173 6855 2210 6856
rect 2285 6855 2322 6865
rect 2381 6885 2529 6895
rect 2629 6892 2725 6894
rect 2381 6865 2390 6885
rect 2410 6865 2500 6885
rect 2520 6865 2529 6885
rect 2381 6859 2529 6865
rect 2381 6856 2445 6859
rect 2381 6855 2418 6856
rect 2437 6829 2445 6856
rect 2466 6856 2529 6859
rect 2587 6885 2725 6892
rect 2587 6865 2596 6885
rect 2616 6865 2725 6885
rect 2587 6856 2725 6865
rect 2466 6829 2473 6856
rect 2492 6855 2529 6856
rect 2588 6855 2625 6856
rect 2437 6804 2473 6829
rect 1735 6802 1818 6803
rect 1908 6802 1949 6803
rect 1735 6795 1949 6802
rect 1735 6778 1918 6795
rect 1735 6745 1748 6778
rect 1801 6775 1918 6778
rect 1938 6775 1949 6795
rect 1801 6767 1949 6775
rect 2016 6799 2375 6803
rect 2016 6794 2338 6799
rect 2016 6770 2129 6794
rect 2153 6775 2338 6794
rect 2362 6775 2375 6799
rect 2153 6770 2375 6775
rect 2016 6767 2375 6770
rect 2437 6767 2472 6804
rect 2540 6801 2640 6804
rect 2540 6797 2607 6801
rect 2540 6771 2552 6797
rect 2578 6775 2607 6797
rect 2633 6775 2640 6801
rect 2578 6771 2640 6775
rect 2540 6767 2640 6771
rect 1801 6745 1818 6767
rect 2016 6746 2047 6767
rect 2437 6746 2473 6767
rect 1859 6745 1896 6746
rect 1735 6731 1818 6745
rect 1508 6488 1676 6490
rect 1232 6487 1676 6488
rect 476 6457 1676 6487
rect 1746 6521 1818 6731
rect 1858 6736 1896 6745
rect 1858 6716 1867 6736
rect 1887 6716 1896 6736
rect 1858 6708 1896 6716
rect 1962 6740 2047 6746
rect 2072 6745 2109 6746
rect 1962 6720 1970 6740
rect 1990 6720 2047 6740
rect 1962 6712 2047 6720
rect 2071 6736 2109 6745
rect 2071 6716 2080 6736
rect 2100 6716 2109 6736
rect 1962 6711 1998 6712
rect 2071 6708 2109 6716
rect 2175 6740 2260 6746
rect 2280 6745 2317 6746
rect 2175 6720 2183 6740
rect 2203 6739 2260 6740
rect 2203 6720 2232 6739
rect 2175 6719 2232 6720
rect 2253 6719 2260 6739
rect 2175 6712 2260 6719
rect 2279 6736 2317 6745
rect 2279 6716 2288 6736
rect 2308 6716 2317 6736
rect 2175 6711 2211 6712
rect 2279 6708 2317 6716
rect 2383 6740 2527 6746
rect 2383 6720 2391 6740
rect 2411 6720 2499 6740
rect 2519 6720 2527 6740
rect 2383 6712 2527 6720
rect 2383 6711 2419 6712
rect 2491 6711 2527 6712
rect 2593 6745 2630 6746
rect 2593 6744 2631 6745
rect 2593 6736 2657 6744
rect 2593 6716 2602 6736
rect 2622 6722 2657 6736
rect 2677 6722 2680 6742
rect 2622 6717 2680 6722
rect 2622 6716 2657 6717
rect 1859 6679 1896 6708
rect 1860 6677 1896 6679
rect 2072 6677 2109 6708
rect 1860 6655 2109 6677
rect 1941 6649 2052 6655
rect 1941 6641 1982 6649
rect 1941 6621 1949 6641
rect 1968 6621 1982 6641
rect 1941 6619 1982 6621
rect 2010 6641 2052 6649
rect 2010 6621 2026 6641
rect 2045 6621 2052 6641
rect 2010 6619 2052 6621
rect 1941 6604 2052 6619
rect 1746 6482 1765 6521
rect 1810 6482 1818 6521
rect 1746 6465 1818 6482
rect 2280 6509 2317 6708
rect 2593 6704 2657 6716
rect 2280 6503 2321 6509
rect 2697 6505 2724 6856
rect 3019 6843 3114 6869
rect 2855 6821 2919 6840
rect 2855 6782 2868 6821
rect 2902 6782 2919 6821
rect 2855 6763 2919 6782
rect 2556 6503 2724 6505
rect 2280 6477 2724 6503
rect 476 6410 541 6457
rect 476 6392 499 6410
rect 517 6392 541 6410
rect 1389 6437 1424 6439
rect 1389 6435 1493 6437
rect 2282 6435 2321 6477
rect 2556 6476 2724 6477
rect 1389 6428 2323 6435
rect 1389 6427 1440 6428
rect 1389 6407 1392 6427
rect 1417 6408 1440 6427
rect 1472 6408 2323 6428
rect 1417 6407 2323 6408
rect 1389 6400 2323 6407
rect 1662 6399 2323 6400
rect 476 6371 541 6392
rect 753 6382 793 6385
rect 753 6378 1656 6382
rect 753 6358 1630 6378
rect 1650 6358 1656 6378
rect 753 6355 1656 6358
rect 477 6311 542 6331
rect 477 6293 501 6311
rect 519 6293 542 6311
rect 477 6266 542 6293
rect 753 6266 793 6355
rect 1237 6353 1653 6355
rect 1237 6352 1578 6353
rect 894 6321 1004 6335
rect 894 6318 937 6321
rect 894 6313 898 6318
rect 476 6231 793 6266
rect 816 6291 898 6313
rect 927 6291 937 6318
rect 965 6294 972 6321
rect 1001 6313 1004 6321
rect 1001 6294 1066 6313
rect 965 6291 1066 6294
rect 816 6289 1066 6291
rect 477 6155 542 6231
rect 816 6210 853 6289
rect 894 6276 1004 6289
rect 968 6220 999 6221
rect 816 6190 825 6210
rect 845 6190 853 6210
rect 816 6180 853 6190
rect 912 6210 999 6220
rect 912 6190 921 6210
rect 941 6190 999 6210
rect 912 6181 999 6190
rect 912 6180 949 6181
rect 477 6137 499 6155
rect 517 6137 542 6155
rect 477 6116 542 6137
rect 690 6135 755 6144
rect 690 6098 700 6135
rect 740 6127 755 6135
rect 968 6128 999 6181
rect 1029 6210 1066 6289
rect 1181 6220 1212 6221
rect 1029 6190 1038 6210
rect 1058 6190 1066 6210
rect 1029 6180 1066 6190
rect 1125 6213 1212 6220
rect 1125 6210 1186 6213
rect 1125 6190 1134 6210
rect 1154 6193 1186 6210
rect 1207 6193 1212 6213
rect 1154 6190 1212 6193
rect 1125 6183 1212 6190
rect 1237 6210 1274 6352
rect 1540 6351 1577 6352
rect 2857 6292 2919 6763
rect 3019 6802 3045 6843
rect 3081 6802 3114 6843
rect 3019 6506 3114 6802
rect 3019 6462 3034 6506
rect 3094 6462 3114 6506
rect 3019 6442 3114 6462
rect 3731 6373 3774 7086
rect 3731 6353 4125 6373
rect 4145 6353 4148 6373
rect 3732 6348 4148 6353
rect 3732 6347 4073 6348
rect 3389 6316 3499 6330
rect 3389 6313 3432 6316
rect 3389 6308 3393 6313
rect 2852 6240 2927 6292
rect 3311 6286 3393 6308
rect 3422 6286 3432 6313
rect 3460 6289 3467 6316
rect 3496 6308 3499 6316
rect 3496 6289 3561 6308
rect 3460 6286 3561 6289
rect 3311 6284 3561 6286
rect 3221 6240 3267 6241
rect 1389 6220 1425 6221
rect 1237 6190 1246 6210
rect 1266 6190 1274 6210
rect 1125 6181 1181 6183
rect 1125 6180 1162 6181
rect 1237 6180 1274 6190
rect 1333 6210 1481 6220
rect 1581 6217 1677 6219
rect 1333 6190 1342 6210
rect 1362 6190 1452 6210
rect 1472 6190 1481 6210
rect 1333 6184 1481 6190
rect 1333 6181 1397 6184
rect 1333 6180 1370 6181
rect 1389 6154 1397 6181
rect 1418 6181 1481 6184
rect 1539 6210 1677 6217
rect 1539 6190 1548 6210
rect 1568 6190 1677 6210
rect 1539 6181 1677 6190
rect 2852 6205 3267 6240
rect 1418 6154 1425 6181
rect 1444 6180 1481 6181
rect 1540 6180 1577 6181
rect 1389 6129 1425 6154
rect 860 6127 901 6128
rect 740 6120 901 6127
rect 740 6100 870 6120
rect 890 6100 901 6120
rect 740 6098 901 6100
rect 690 6092 901 6098
rect 968 6124 1327 6128
rect 968 6119 1290 6124
rect 968 6095 1081 6119
rect 1105 6100 1290 6119
rect 1314 6100 1327 6124
rect 1105 6095 1327 6100
rect 968 6092 1327 6095
rect 1389 6092 1424 6129
rect 1492 6126 1592 6129
rect 1492 6122 1559 6126
rect 1492 6096 1504 6122
rect 1530 6100 1559 6122
rect 1585 6100 1592 6126
rect 1530 6096 1592 6100
rect 1492 6092 1592 6096
rect 690 6079 757 6092
rect 482 6056 538 6076
rect 482 6038 501 6056
rect 519 6038 538 6056
rect 482 5925 538 6038
rect 690 6058 704 6079
rect 740 6058 757 6079
rect 968 6071 999 6092
rect 1389 6071 1425 6092
rect 811 6070 848 6071
rect 690 6051 757 6058
rect 810 6061 848 6070
rect 482 5787 537 5925
rect 690 5899 755 6051
rect 810 6041 819 6061
rect 839 6041 848 6061
rect 810 6033 848 6041
rect 914 6065 999 6071
rect 1024 6070 1061 6071
rect 914 6045 922 6065
rect 942 6045 999 6065
rect 914 6037 999 6045
rect 1023 6061 1061 6070
rect 1023 6041 1032 6061
rect 1052 6041 1061 6061
rect 914 6036 950 6037
rect 1023 6033 1061 6041
rect 1127 6065 1212 6071
rect 1232 6070 1269 6071
rect 1127 6045 1135 6065
rect 1155 6064 1212 6065
rect 1155 6045 1184 6064
rect 1127 6044 1184 6045
rect 1205 6044 1212 6064
rect 1127 6037 1212 6044
rect 1231 6061 1269 6070
rect 1231 6041 1240 6061
rect 1260 6041 1269 6061
rect 1127 6036 1163 6037
rect 1231 6033 1269 6041
rect 1335 6065 1479 6071
rect 1335 6045 1343 6065
rect 1363 6045 1451 6065
rect 1471 6045 1479 6065
rect 1335 6037 1479 6045
rect 1335 6036 1371 6037
rect 1443 6036 1479 6037
rect 1545 6070 1582 6071
rect 1545 6069 1583 6070
rect 1545 6061 1609 6069
rect 1545 6041 1554 6061
rect 1574 6047 1609 6061
rect 1629 6047 1632 6067
rect 1574 6042 1632 6047
rect 1574 6041 1609 6042
rect 811 6004 848 6033
rect 812 6002 848 6004
rect 1024 6002 1061 6033
rect 812 5980 1061 6002
rect 893 5974 1004 5980
rect 893 5966 934 5974
rect 893 5946 901 5966
rect 920 5946 934 5966
rect 893 5944 934 5946
rect 962 5966 1004 5974
rect 962 5946 978 5966
rect 997 5946 1004 5966
rect 962 5944 1004 5946
rect 893 5931 1004 5944
rect 1232 5934 1269 6033
rect 1545 6029 1609 6041
rect 683 5889 804 5899
rect 683 5887 752 5889
rect 683 5846 696 5887
rect 733 5848 752 5887
rect 789 5848 804 5889
rect 733 5846 804 5848
rect 683 5828 804 5846
rect 475 5784 539 5787
rect 895 5784 999 5790
rect 1230 5784 1271 5934
rect 1649 5926 1676 6181
rect 1738 6171 1818 6182
rect 1738 6145 1755 6171
rect 1795 6145 1818 6171
rect 1738 6118 1818 6145
rect 1738 6092 1759 6118
rect 1799 6092 1818 6118
rect 1738 6073 1818 6092
rect 1738 6047 1762 6073
rect 1802 6047 1818 6073
rect 1738 5996 1818 6047
rect 475 5781 1271 5784
rect 1650 5795 1676 5926
rect 1650 5781 1678 5795
rect 475 5746 1678 5781
rect 1740 5788 1810 5996
rect 2852 5921 2927 6205
rect 3221 6122 3267 6205
rect 3311 6205 3348 6284
rect 3389 6271 3499 6284
rect 3463 6215 3494 6216
rect 3311 6185 3320 6205
rect 3340 6185 3348 6205
rect 3311 6175 3348 6185
rect 3407 6205 3494 6215
rect 3407 6185 3416 6205
rect 3436 6185 3494 6205
rect 3407 6176 3494 6185
rect 3407 6175 3444 6176
rect 3463 6123 3494 6176
rect 3524 6205 3561 6284
rect 3676 6215 3707 6216
rect 3524 6185 3533 6205
rect 3553 6185 3561 6205
rect 3524 6175 3561 6185
rect 3620 6208 3707 6215
rect 3620 6205 3681 6208
rect 3620 6185 3629 6205
rect 3649 6188 3681 6205
rect 3702 6188 3707 6208
rect 3649 6185 3707 6188
rect 3620 6178 3707 6185
rect 3732 6205 3769 6347
rect 4035 6346 4072 6347
rect 3884 6215 3920 6216
rect 3732 6185 3741 6205
rect 3761 6185 3769 6205
rect 3620 6176 3676 6178
rect 3620 6175 3657 6176
rect 3732 6175 3769 6185
rect 3828 6205 3976 6215
rect 4076 6212 4172 6214
rect 3828 6185 3837 6205
rect 3857 6185 3947 6205
rect 3967 6185 3976 6205
rect 3828 6179 3976 6185
rect 3828 6176 3892 6179
rect 3828 6175 3865 6176
rect 3884 6149 3892 6176
rect 3913 6176 3976 6179
rect 4034 6205 4172 6212
rect 4034 6185 4043 6205
rect 4063 6185 4172 6205
rect 4034 6176 4172 6185
rect 3913 6149 3920 6176
rect 3939 6175 3976 6176
rect 4035 6175 4072 6176
rect 3884 6124 3920 6149
rect 3355 6122 3396 6123
rect 3221 6115 3396 6122
rect 3019 6089 3105 6108
rect 3019 6048 3034 6089
rect 3088 6048 3105 6089
rect 3221 6095 3365 6115
rect 3385 6095 3396 6115
rect 3221 6087 3396 6095
rect 3463 6119 3822 6123
rect 3463 6114 3785 6119
rect 3463 6090 3576 6114
rect 3600 6095 3785 6114
rect 3809 6095 3822 6119
rect 3600 6090 3822 6095
rect 3463 6087 3822 6090
rect 3884 6087 3919 6124
rect 3987 6121 4087 6124
rect 3987 6117 4054 6121
rect 3987 6091 3999 6117
rect 4025 6095 4054 6117
rect 4080 6095 4087 6121
rect 4025 6091 4087 6095
rect 3987 6087 4087 6091
rect 3221 6083 3267 6087
rect 3463 6066 3494 6087
rect 3884 6066 3920 6087
rect 3306 6065 3343 6066
rect 3019 6012 3105 6048
rect 3305 6056 3343 6065
rect 3305 6036 3314 6056
rect 3334 6036 3343 6056
rect 3305 6028 3343 6036
rect 3409 6060 3494 6066
rect 3519 6065 3556 6066
rect 3409 6040 3417 6060
rect 3437 6040 3494 6060
rect 3409 6032 3494 6040
rect 3518 6056 3556 6065
rect 3518 6036 3527 6056
rect 3547 6036 3556 6056
rect 3409 6031 3445 6032
rect 3518 6028 3556 6036
rect 3622 6060 3707 6066
rect 3727 6065 3764 6066
rect 3622 6040 3630 6060
rect 3650 6059 3707 6060
rect 3650 6040 3679 6059
rect 3622 6039 3679 6040
rect 3700 6039 3707 6059
rect 3622 6032 3707 6039
rect 3726 6056 3764 6065
rect 3726 6036 3735 6056
rect 3755 6036 3764 6056
rect 3622 6031 3658 6032
rect 3726 6028 3764 6036
rect 3830 6060 3974 6066
rect 3830 6040 3838 6060
rect 3858 6040 3946 6060
rect 3966 6040 3974 6060
rect 3830 6032 3974 6040
rect 3830 6031 3866 6032
rect 475 5685 539 5746
rect 895 5744 999 5746
rect 1230 5744 1271 5746
rect 1740 5743 1761 5788
rect 1741 5722 1761 5743
rect 1791 5743 1810 5788
rect 2847 5879 2927 5921
rect 1791 5722 1808 5743
rect 1741 5703 1808 5722
rect 1390 5695 1462 5696
rect 1389 5687 1488 5695
rect 477 5614 536 5685
rect 1389 5684 1441 5687
rect 1389 5649 1397 5684
rect 1422 5649 1441 5684
rect 1466 5676 1488 5687
rect 1466 5675 2333 5676
rect 1466 5649 2334 5675
rect 1389 5639 2334 5649
rect 1389 5637 1488 5639
rect 477 5596 499 5614
rect 517 5596 536 5614
rect 477 5574 536 5596
rect 744 5610 1276 5615
rect 744 5590 1630 5610
rect 1650 5590 1653 5610
rect 2289 5606 2334 5639
rect 744 5586 1653 5590
rect 744 5539 787 5586
rect 1237 5585 1653 5586
rect 2285 5586 2678 5606
rect 2698 5586 2701 5606
rect 1237 5584 1578 5585
rect 894 5553 1004 5567
rect 894 5550 937 5553
rect 894 5545 898 5550
rect 732 5538 787 5539
rect 476 5515 787 5538
rect 476 5497 501 5515
rect 519 5503 787 5515
rect 816 5523 898 5545
rect 927 5523 937 5550
rect 965 5526 972 5553
rect 1001 5545 1004 5553
rect 1001 5526 1066 5545
rect 965 5523 1066 5526
rect 816 5521 1066 5523
rect 519 5497 541 5503
rect 476 5358 541 5497
rect 816 5442 853 5521
rect 894 5508 1004 5521
rect 968 5452 999 5453
rect 816 5422 825 5442
rect 845 5422 853 5442
rect 476 5340 499 5358
rect 517 5340 541 5358
rect 476 5323 541 5340
rect 696 5404 764 5417
rect 816 5412 853 5422
rect 912 5442 999 5452
rect 912 5422 921 5442
rect 941 5422 999 5442
rect 912 5413 999 5422
rect 912 5412 949 5413
rect 696 5362 703 5404
rect 752 5362 764 5404
rect 696 5359 764 5362
rect 968 5360 999 5413
rect 1029 5442 1066 5521
rect 1181 5452 1212 5453
rect 1029 5422 1038 5442
rect 1058 5422 1066 5442
rect 1029 5412 1066 5422
rect 1125 5445 1212 5452
rect 1125 5442 1186 5445
rect 1125 5422 1134 5442
rect 1154 5425 1186 5442
rect 1207 5425 1212 5445
rect 1154 5422 1212 5425
rect 1125 5415 1212 5422
rect 1237 5442 1274 5584
rect 1540 5583 1577 5584
rect 2285 5581 2701 5586
rect 2285 5580 2626 5581
rect 1942 5549 2052 5563
rect 1942 5546 1985 5549
rect 1942 5541 1946 5546
rect 1864 5519 1946 5541
rect 1975 5519 1985 5546
rect 2013 5522 2020 5549
rect 2049 5541 2052 5549
rect 2049 5522 2114 5541
rect 2013 5519 2114 5522
rect 1864 5517 2114 5519
rect 1389 5452 1425 5453
rect 1237 5422 1246 5442
rect 1266 5422 1274 5442
rect 1125 5413 1181 5415
rect 1125 5412 1162 5413
rect 1237 5412 1274 5422
rect 1333 5442 1481 5452
rect 1581 5449 1677 5451
rect 1333 5422 1342 5442
rect 1362 5422 1452 5442
rect 1472 5422 1481 5442
rect 1333 5416 1481 5422
rect 1333 5413 1397 5416
rect 1333 5412 1370 5413
rect 1389 5386 1397 5413
rect 1418 5413 1481 5416
rect 1539 5442 1677 5449
rect 1539 5422 1548 5442
rect 1568 5422 1677 5442
rect 1539 5413 1677 5422
rect 1864 5438 1901 5517
rect 1942 5504 2052 5517
rect 2016 5448 2047 5449
rect 1864 5418 1873 5438
rect 1893 5418 1901 5438
rect 1418 5386 1425 5413
rect 1444 5412 1481 5413
rect 1540 5412 1577 5413
rect 1389 5361 1425 5386
rect 860 5359 901 5360
rect 696 5352 901 5359
rect 696 5341 870 5352
rect 696 5308 704 5341
rect 697 5299 704 5308
rect 753 5332 870 5341
rect 890 5332 901 5352
rect 753 5324 901 5332
rect 968 5356 1327 5360
rect 968 5351 1290 5356
rect 968 5327 1081 5351
rect 1105 5332 1290 5351
rect 1314 5332 1327 5356
rect 1105 5327 1327 5332
rect 968 5324 1327 5327
rect 1389 5324 1424 5361
rect 1492 5358 1592 5361
rect 1492 5354 1559 5358
rect 1492 5328 1504 5354
rect 1530 5332 1559 5354
rect 1585 5332 1592 5358
rect 1530 5328 1592 5332
rect 1492 5324 1592 5328
rect 753 5308 764 5324
rect 753 5299 761 5308
rect 968 5303 999 5324
rect 1389 5303 1425 5324
rect 811 5302 848 5303
rect 476 5259 541 5278
rect 476 5241 501 5259
rect 519 5241 541 5259
rect 476 5040 541 5241
rect 697 5115 761 5299
rect 810 5293 848 5302
rect 810 5273 819 5293
rect 839 5273 848 5293
rect 810 5265 848 5273
rect 914 5297 999 5303
rect 1024 5302 1061 5303
rect 914 5277 922 5297
rect 942 5277 999 5297
rect 914 5269 999 5277
rect 1023 5293 1061 5302
rect 1023 5273 1032 5293
rect 1052 5273 1061 5293
rect 914 5268 950 5269
rect 1023 5265 1061 5273
rect 1127 5297 1212 5303
rect 1232 5302 1269 5303
rect 1127 5277 1135 5297
rect 1155 5296 1212 5297
rect 1155 5277 1184 5296
rect 1127 5276 1184 5277
rect 1205 5276 1212 5296
rect 1127 5269 1212 5276
rect 1231 5293 1269 5302
rect 1231 5273 1240 5293
rect 1260 5273 1269 5293
rect 1127 5268 1163 5269
rect 1231 5265 1269 5273
rect 1335 5297 1479 5303
rect 1335 5277 1343 5297
rect 1363 5277 1451 5297
rect 1471 5277 1479 5297
rect 1335 5269 1479 5277
rect 1335 5268 1371 5269
rect 1443 5268 1479 5269
rect 1545 5302 1582 5303
rect 1545 5301 1583 5302
rect 1545 5293 1609 5301
rect 1545 5273 1554 5293
rect 1574 5279 1609 5293
rect 1629 5279 1632 5299
rect 1574 5274 1632 5279
rect 1574 5273 1609 5274
rect 811 5236 848 5265
rect 812 5234 848 5236
rect 1024 5234 1061 5265
rect 812 5212 1061 5234
rect 893 5206 1004 5212
rect 893 5198 934 5206
rect 893 5178 901 5198
rect 920 5178 934 5198
rect 893 5176 934 5178
rect 962 5198 1004 5206
rect 962 5178 978 5198
rect 997 5178 1004 5198
rect 962 5176 1004 5178
rect 893 5161 1004 5176
rect 697 5105 765 5115
rect 697 5072 714 5105
rect 754 5072 765 5105
rect 697 5060 765 5072
rect 697 5058 761 5060
rect 1232 5041 1269 5265
rect 1545 5261 1609 5273
rect 1649 5043 1676 5413
rect 1864 5408 1901 5418
rect 1960 5438 2047 5448
rect 1960 5418 1969 5438
rect 1989 5418 2047 5438
rect 1960 5409 2047 5418
rect 1960 5408 1997 5409
rect 1740 5395 1810 5400
rect 1735 5389 1810 5395
rect 1735 5356 1743 5389
rect 1796 5356 1810 5389
rect 2016 5356 2047 5409
rect 2077 5438 2114 5517
rect 2229 5448 2260 5449
rect 2077 5418 2086 5438
rect 2106 5418 2114 5438
rect 2077 5408 2114 5418
rect 2173 5441 2260 5448
rect 2173 5438 2234 5441
rect 2173 5418 2182 5438
rect 2202 5421 2234 5438
rect 2255 5421 2260 5441
rect 2202 5418 2260 5421
rect 2173 5411 2260 5418
rect 2285 5438 2322 5580
rect 2588 5579 2625 5580
rect 2437 5448 2473 5449
rect 2285 5418 2294 5438
rect 2314 5418 2322 5438
rect 2173 5409 2229 5411
rect 2173 5408 2210 5409
rect 2285 5408 2322 5418
rect 2381 5438 2529 5448
rect 2629 5445 2725 5447
rect 2381 5418 2390 5438
rect 2410 5418 2500 5438
rect 2520 5418 2529 5438
rect 2381 5412 2529 5418
rect 2381 5409 2445 5412
rect 2381 5408 2418 5409
rect 2437 5382 2445 5409
rect 2466 5409 2529 5412
rect 2587 5438 2725 5445
rect 2587 5418 2596 5438
rect 2616 5418 2725 5438
rect 2587 5409 2725 5418
rect 2466 5382 2473 5409
rect 2492 5408 2529 5409
rect 2588 5408 2625 5409
rect 2437 5357 2473 5382
rect 1735 5355 1818 5356
rect 1908 5355 1949 5356
rect 1735 5348 1949 5355
rect 1735 5331 1918 5348
rect 1735 5298 1748 5331
rect 1801 5328 1918 5331
rect 1938 5328 1949 5348
rect 1801 5320 1949 5328
rect 2016 5352 2375 5356
rect 2016 5347 2338 5352
rect 2016 5323 2129 5347
rect 2153 5328 2338 5347
rect 2362 5328 2375 5352
rect 2153 5323 2375 5328
rect 2016 5320 2375 5323
rect 2437 5320 2472 5357
rect 2540 5354 2640 5357
rect 2540 5350 2607 5354
rect 2540 5324 2552 5350
rect 2578 5328 2607 5350
rect 2633 5328 2640 5354
rect 2578 5324 2640 5328
rect 2540 5320 2640 5324
rect 1801 5298 1818 5320
rect 2016 5299 2047 5320
rect 2437 5299 2473 5320
rect 1859 5298 1896 5299
rect 1735 5284 1818 5298
rect 1508 5041 1676 5043
rect 1232 5040 1676 5041
rect 476 5010 1676 5040
rect 1746 5074 1818 5284
rect 1858 5289 1896 5298
rect 1858 5269 1867 5289
rect 1887 5269 1896 5289
rect 1858 5261 1896 5269
rect 1962 5293 2047 5299
rect 2072 5298 2109 5299
rect 1962 5273 1970 5293
rect 1990 5273 2047 5293
rect 1962 5265 2047 5273
rect 2071 5289 2109 5298
rect 2071 5269 2080 5289
rect 2100 5269 2109 5289
rect 1962 5264 1998 5265
rect 2071 5261 2109 5269
rect 2175 5293 2260 5299
rect 2280 5298 2317 5299
rect 2175 5273 2183 5293
rect 2203 5292 2260 5293
rect 2203 5273 2232 5292
rect 2175 5272 2232 5273
rect 2253 5272 2260 5292
rect 2175 5265 2260 5272
rect 2279 5289 2317 5298
rect 2279 5269 2288 5289
rect 2308 5269 2317 5289
rect 2175 5264 2211 5265
rect 2279 5261 2317 5269
rect 2383 5293 2527 5299
rect 2383 5273 2391 5293
rect 2411 5273 2499 5293
rect 2519 5273 2527 5293
rect 2383 5265 2527 5273
rect 2383 5264 2419 5265
rect 2491 5264 2527 5265
rect 2593 5298 2630 5299
rect 2593 5297 2631 5298
rect 2593 5289 2657 5297
rect 2593 5269 2602 5289
rect 2622 5275 2657 5289
rect 2677 5275 2680 5295
rect 2622 5270 2680 5275
rect 2622 5269 2657 5270
rect 1859 5232 1896 5261
rect 1860 5230 1896 5232
rect 2072 5230 2109 5261
rect 1860 5208 2109 5230
rect 1941 5202 2052 5208
rect 1941 5194 1982 5202
rect 1941 5174 1949 5194
rect 1968 5174 1982 5194
rect 1941 5172 1982 5174
rect 2010 5194 2052 5202
rect 2010 5174 2026 5194
rect 2045 5174 2052 5194
rect 2010 5172 2052 5174
rect 1941 5157 2052 5172
rect 1746 5035 1765 5074
rect 1810 5035 1818 5074
rect 1746 5018 1818 5035
rect 2280 5062 2317 5261
rect 2593 5257 2657 5269
rect 2280 5056 2321 5062
rect 2697 5058 2724 5409
rect 2847 5279 2926 5879
rect 3023 5427 3102 6012
rect 3306 5999 3343 6028
rect 3307 5997 3343 5999
rect 3519 5997 3556 6028
rect 3307 5975 3556 5997
rect 3388 5969 3499 5975
rect 3388 5961 3429 5969
rect 3388 5941 3396 5961
rect 3415 5941 3429 5961
rect 3388 5939 3429 5941
rect 3457 5961 3499 5969
rect 3457 5941 3473 5961
rect 3492 5941 3499 5961
rect 3457 5939 3499 5941
rect 3388 5924 3499 5939
rect 3727 5913 3764 6028
rect 3720 5801 3767 5913
rect 3888 5873 3918 6032
rect 3938 6031 3974 6032
rect 4040 6065 4077 6066
rect 4040 6064 4078 6065
rect 4040 6056 4104 6064
rect 4040 6036 4049 6056
rect 4069 6042 4104 6056
rect 4124 6042 4127 6062
rect 4069 6037 4127 6042
rect 4069 6036 4104 6037
rect 4040 6024 4104 6036
rect 3888 5869 3974 5873
rect 3888 5851 3903 5869
rect 3955 5851 3974 5869
rect 3888 5842 3974 5851
rect 4144 5803 4171 6176
rect 4003 5801 4171 5803
rect 3720 5775 4171 5801
rect 3720 5697 3767 5775
rect 4003 5774 4171 5775
rect 3665 5696 3767 5697
rect 3664 5688 3767 5696
rect 3664 5685 3716 5688
rect 3664 5650 3672 5685
rect 3697 5650 3716 5685
rect 3741 5650 3767 5688
rect 3664 5644 3767 5650
rect 3927 5689 3963 5693
rect 3927 5666 3935 5689
rect 3959 5666 3963 5689
rect 3927 5645 3963 5666
rect 3664 5640 3763 5644
rect 3927 5622 3935 5645
rect 3959 5622 3963 5645
rect 2556 5056 2724 5058
rect 2280 5030 2724 5056
rect 476 4963 541 5010
rect 476 4945 499 4963
rect 517 4945 541 4963
rect 1389 4990 1424 4992
rect 1389 4988 1493 4990
rect 2282 4988 2321 5030
rect 2556 5029 2724 5030
rect 1389 4981 2323 4988
rect 1389 4980 1440 4981
rect 1389 4960 1392 4980
rect 1417 4961 1440 4980
rect 1472 4961 2323 4981
rect 1417 4960 2323 4961
rect 1389 4953 2323 4960
rect 1662 4952 2323 4953
rect 476 4924 541 4945
rect 753 4935 793 4938
rect 753 4931 1656 4935
rect 753 4911 1630 4931
rect 1650 4911 1656 4931
rect 753 4908 1656 4911
rect 477 4864 542 4884
rect 477 4846 501 4864
rect 519 4846 542 4864
rect 477 4819 542 4846
rect 753 4819 793 4908
rect 1237 4906 1653 4908
rect 1237 4905 1578 4906
rect 894 4874 1004 4888
rect 894 4871 937 4874
rect 894 4866 898 4871
rect 476 4784 793 4819
rect 816 4844 898 4866
rect 927 4844 937 4871
rect 965 4847 972 4874
rect 1001 4866 1004 4874
rect 1001 4847 1066 4866
rect 965 4844 1066 4847
rect 816 4842 1066 4844
rect 477 4708 542 4784
rect 816 4763 853 4842
rect 894 4829 1004 4842
rect 968 4773 999 4774
rect 816 4743 825 4763
rect 845 4743 853 4763
rect 816 4733 853 4743
rect 912 4763 999 4773
rect 912 4743 921 4763
rect 941 4743 999 4763
rect 912 4734 999 4743
rect 912 4733 949 4734
rect 477 4690 499 4708
rect 517 4690 542 4708
rect 477 4669 542 4690
rect 690 4688 755 4697
rect 690 4651 700 4688
rect 740 4680 755 4688
rect 968 4681 999 4734
rect 1029 4763 1066 4842
rect 1181 4773 1212 4774
rect 1029 4743 1038 4763
rect 1058 4743 1066 4763
rect 1029 4733 1066 4743
rect 1125 4766 1212 4773
rect 1125 4763 1186 4766
rect 1125 4743 1134 4763
rect 1154 4746 1186 4763
rect 1207 4746 1212 4766
rect 1154 4743 1212 4746
rect 1125 4736 1212 4743
rect 1237 4763 1274 4905
rect 1540 4904 1577 4905
rect 1389 4773 1425 4774
rect 1237 4743 1246 4763
rect 1266 4743 1274 4763
rect 1125 4734 1181 4736
rect 1125 4733 1162 4734
rect 1237 4733 1274 4743
rect 1333 4763 1481 4773
rect 1581 4770 1677 4772
rect 1333 4743 1342 4763
rect 1362 4743 1452 4763
rect 1472 4743 1481 4763
rect 1333 4737 1481 4743
rect 1333 4734 1397 4737
rect 1333 4733 1370 4734
rect 1389 4707 1397 4734
rect 1418 4734 1481 4737
rect 1539 4763 1677 4770
rect 1539 4743 1548 4763
rect 1568 4743 1677 4763
rect 1539 4734 1677 4743
rect 1418 4707 1425 4734
rect 1444 4733 1481 4734
rect 1540 4733 1577 4734
rect 1389 4682 1425 4707
rect 860 4680 901 4681
rect 740 4673 901 4680
rect 740 4653 870 4673
rect 890 4653 901 4673
rect 740 4651 901 4653
rect 690 4645 901 4651
rect 968 4677 1327 4681
rect 968 4672 1290 4677
rect 968 4648 1081 4672
rect 1105 4653 1290 4672
rect 1314 4653 1327 4677
rect 1105 4648 1327 4653
rect 968 4645 1327 4648
rect 1389 4645 1424 4682
rect 1492 4679 1592 4682
rect 1492 4675 1559 4679
rect 1492 4649 1504 4675
rect 1530 4653 1559 4675
rect 1585 4653 1592 4679
rect 1530 4649 1592 4653
rect 1492 4645 1592 4649
rect 690 4632 757 4645
rect 482 4609 538 4629
rect 482 4591 501 4609
rect 519 4591 538 4609
rect 482 4478 538 4591
rect 690 4611 704 4632
rect 740 4611 757 4632
rect 968 4624 999 4645
rect 1389 4624 1425 4645
rect 811 4623 848 4624
rect 690 4604 757 4611
rect 810 4614 848 4623
rect 482 4349 537 4478
rect 690 4452 755 4604
rect 810 4594 819 4614
rect 839 4594 848 4614
rect 810 4586 848 4594
rect 914 4618 999 4624
rect 1024 4623 1061 4624
rect 914 4598 922 4618
rect 942 4598 999 4618
rect 914 4590 999 4598
rect 1023 4614 1061 4623
rect 1023 4594 1032 4614
rect 1052 4594 1061 4614
rect 914 4589 950 4590
rect 1023 4586 1061 4594
rect 1127 4618 1212 4624
rect 1232 4623 1269 4624
rect 1127 4598 1135 4618
rect 1155 4617 1212 4618
rect 1155 4598 1184 4617
rect 1127 4597 1184 4598
rect 1205 4597 1212 4617
rect 1127 4590 1212 4597
rect 1231 4614 1269 4623
rect 1231 4594 1240 4614
rect 1260 4594 1269 4614
rect 1127 4589 1163 4590
rect 1231 4586 1269 4594
rect 1335 4618 1479 4624
rect 1335 4598 1343 4618
rect 1363 4598 1451 4618
rect 1471 4598 1479 4618
rect 1335 4590 1479 4598
rect 1335 4589 1371 4590
rect 1443 4589 1479 4590
rect 1545 4623 1582 4624
rect 1545 4622 1583 4623
rect 1545 4614 1609 4622
rect 1545 4594 1554 4614
rect 1574 4600 1609 4614
rect 1629 4600 1632 4620
rect 1574 4595 1632 4600
rect 1574 4594 1609 4595
rect 811 4557 848 4586
rect 812 4555 848 4557
rect 1024 4555 1061 4586
rect 812 4533 1061 4555
rect 893 4527 1004 4533
rect 893 4519 934 4527
rect 893 4499 901 4519
rect 920 4499 934 4519
rect 893 4497 934 4499
rect 962 4519 1004 4527
rect 962 4499 978 4519
rect 997 4499 1004 4519
rect 962 4497 1004 4499
rect 893 4482 1004 4497
rect 1232 4487 1269 4586
rect 1545 4582 1609 4594
rect 895 4473 999 4482
rect 683 4442 804 4452
rect 683 4440 752 4442
rect 683 4399 696 4440
rect 733 4401 752 4440
rect 789 4401 804 4442
rect 733 4399 804 4401
rect 683 4381 804 4399
rect 476 4337 537 4349
rect 1230 4337 1271 4487
rect 1649 4479 1676 4734
rect 1738 4724 1818 4735
rect 1738 4698 1755 4724
rect 1795 4698 1818 4724
rect 1738 4671 1818 4698
rect 1738 4645 1759 4671
rect 1799 4645 1818 4671
rect 1738 4626 1818 4645
rect 1738 4600 1762 4626
rect 1802 4600 1818 4626
rect 1738 4549 1818 4600
rect 476 4334 1271 4337
rect 1650 4348 1676 4479
rect 1740 4393 1810 4549
rect 1739 4377 1815 4393
rect 1650 4334 1678 4348
rect 476 4299 1678 4334
rect 1739 4340 1754 4377
rect 1798 4340 1815 4377
rect 1739 4320 1815 4340
rect 2853 4370 2923 5279
rect 3022 4758 3103 5427
rect 3927 5322 3963 5622
rect 3851 5293 3964 5322
rect 3851 4928 3882 5293
rect 3775 4908 4168 4928
rect 4188 4908 4191 4928
rect 3775 4903 4191 4908
rect 3775 4902 4116 4903
rect 3432 4871 3542 4885
rect 3432 4868 3475 4871
rect 3432 4863 3436 4868
rect 3354 4841 3436 4863
rect 3465 4841 3475 4868
rect 3503 4844 3510 4871
rect 3539 4863 3542 4871
rect 3539 4844 3604 4863
rect 3503 4841 3604 4844
rect 3354 4839 3604 4841
rect 3354 4760 3391 4839
rect 3432 4826 3542 4839
rect 3506 4770 3537 4771
rect 3016 4678 3115 4758
rect 3354 4740 3363 4760
rect 3383 4740 3391 4760
rect 3354 4730 3391 4740
rect 3450 4760 3537 4770
rect 3450 4740 3459 4760
rect 3479 4740 3537 4760
rect 3450 4731 3537 4740
rect 3450 4730 3487 4731
rect 3506 4678 3537 4731
rect 3567 4760 3604 4839
rect 3719 4770 3750 4771
rect 3567 4740 3576 4760
rect 3596 4740 3604 4760
rect 3567 4730 3604 4740
rect 3663 4763 3750 4770
rect 3663 4760 3724 4763
rect 3663 4740 3672 4760
rect 3692 4743 3724 4760
rect 3745 4743 3750 4763
rect 3692 4740 3750 4743
rect 3663 4733 3750 4740
rect 3775 4760 3812 4902
rect 4078 4901 4115 4902
rect 3927 4770 3963 4771
rect 3775 4740 3784 4760
rect 3804 4740 3812 4760
rect 3663 4731 3719 4733
rect 3663 4730 3700 4731
rect 3775 4730 3812 4740
rect 3871 4760 4019 4770
rect 4119 4767 4215 4769
rect 3871 4740 3880 4760
rect 3900 4740 3990 4760
rect 4010 4740 4019 4760
rect 3871 4734 4019 4740
rect 3871 4731 3935 4734
rect 3871 4730 3908 4731
rect 3927 4704 3935 4731
rect 3956 4731 4019 4734
rect 4077 4760 4215 4767
rect 4077 4740 4086 4760
rect 4106 4740 4215 4760
rect 4077 4731 4215 4740
rect 3956 4704 3963 4731
rect 3982 4730 4019 4731
rect 4078 4730 4115 4731
rect 3927 4679 3963 4704
rect 3016 4677 3356 4678
rect 3398 4677 3439 4678
rect 3016 4670 3439 4677
rect 3016 4650 3408 4670
rect 3428 4650 3439 4670
rect 3016 4642 3439 4650
rect 3506 4674 3865 4678
rect 3506 4669 3828 4674
rect 3506 4645 3619 4669
rect 3643 4650 3828 4669
rect 3852 4650 3865 4674
rect 3643 4645 3865 4650
rect 3506 4642 3865 4645
rect 3927 4642 3962 4679
rect 4030 4676 4130 4679
rect 4030 4672 4097 4676
rect 4030 4646 4042 4672
rect 4068 4650 4097 4672
rect 4123 4650 4130 4676
rect 4068 4646 4130 4650
rect 4030 4642 4130 4646
rect 3016 4638 3356 4642
rect 2853 4320 2925 4370
rect 476 4224 537 4299
rect 895 4297 999 4299
rect 1230 4297 1271 4299
rect 1739 4254 1749 4320
rect 1803 4254 1815 4320
rect 1739 4230 1815 4254
rect 478 4094 537 4224
rect 1391 4175 1463 4176
rect 1390 4167 1489 4175
rect 1390 4164 1442 4167
rect 1390 4129 1398 4164
rect 1423 4129 1442 4164
rect 1467 4156 1489 4167
rect 1467 4155 2334 4156
rect 1467 4129 2335 4155
rect 1390 4119 2335 4129
rect 1390 4117 1489 4119
rect 478 4076 500 4094
rect 518 4076 537 4094
rect 478 4054 537 4076
rect 745 4090 1277 4095
rect 745 4070 1631 4090
rect 1651 4070 1654 4090
rect 2290 4086 2335 4119
rect 745 4066 1654 4070
rect 745 4019 788 4066
rect 1238 4065 1654 4066
rect 2286 4066 2679 4086
rect 2699 4066 2702 4086
rect 1238 4064 1579 4065
rect 895 4033 1005 4047
rect 895 4030 938 4033
rect 895 4025 899 4030
rect 733 4018 788 4019
rect 477 3995 788 4018
rect 477 3977 502 3995
rect 520 3983 788 3995
rect 817 4003 899 4025
rect 928 4003 938 4030
rect 966 4006 973 4033
rect 1002 4025 1005 4033
rect 1002 4006 1067 4025
rect 966 4003 1067 4006
rect 817 4001 1067 4003
rect 520 3977 542 3983
rect 477 3838 542 3977
rect 817 3922 854 4001
rect 895 3988 1005 4001
rect 969 3932 1000 3933
rect 817 3902 826 3922
rect 846 3902 854 3922
rect 477 3820 500 3838
rect 518 3820 542 3838
rect 477 3803 542 3820
rect 697 3884 765 3897
rect 817 3892 854 3902
rect 913 3922 1000 3932
rect 913 3902 922 3922
rect 942 3902 1000 3922
rect 913 3893 1000 3902
rect 913 3892 950 3893
rect 697 3842 704 3884
rect 753 3842 765 3884
rect 697 3839 765 3842
rect 969 3840 1000 3893
rect 1030 3922 1067 4001
rect 1182 3932 1213 3933
rect 1030 3902 1039 3922
rect 1059 3902 1067 3922
rect 1030 3892 1067 3902
rect 1126 3925 1213 3932
rect 1126 3922 1187 3925
rect 1126 3902 1135 3922
rect 1155 3905 1187 3922
rect 1208 3905 1213 3925
rect 1155 3902 1213 3905
rect 1126 3895 1213 3902
rect 1238 3922 1275 4064
rect 1541 4063 1578 4064
rect 2286 4061 2702 4066
rect 2286 4060 2627 4061
rect 1943 4029 2053 4043
rect 1943 4026 1986 4029
rect 1943 4021 1947 4026
rect 1865 3999 1947 4021
rect 1976 3999 1986 4026
rect 2014 4002 2021 4029
rect 2050 4021 2053 4029
rect 2050 4002 2115 4021
rect 2014 3999 2115 4002
rect 1865 3997 2115 3999
rect 1390 3932 1426 3933
rect 1238 3902 1247 3922
rect 1267 3902 1275 3922
rect 1126 3893 1182 3895
rect 1126 3892 1163 3893
rect 1238 3892 1275 3902
rect 1334 3922 1482 3932
rect 1582 3929 1678 3931
rect 1334 3902 1343 3922
rect 1363 3902 1453 3922
rect 1473 3902 1482 3922
rect 1334 3896 1482 3902
rect 1334 3893 1398 3896
rect 1334 3892 1371 3893
rect 1390 3866 1398 3893
rect 1419 3893 1482 3896
rect 1540 3922 1678 3929
rect 1540 3902 1549 3922
rect 1569 3902 1678 3922
rect 1540 3893 1678 3902
rect 1865 3918 1902 3997
rect 1943 3984 2053 3997
rect 2017 3928 2048 3929
rect 1865 3898 1874 3918
rect 1894 3898 1902 3918
rect 1419 3866 1426 3893
rect 1445 3892 1482 3893
rect 1541 3892 1578 3893
rect 1390 3841 1426 3866
rect 861 3839 902 3840
rect 697 3832 902 3839
rect 697 3821 871 3832
rect 697 3788 705 3821
rect 698 3779 705 3788
rect 754 3812 871 3821
rect 891 3812 902 3832
rect 754 3804 902 3812
rect 969 3836 1328 3840
rect 969 3831 1291 3836
rect 969 3807 1082 3831
rect 1106 3812 1291 3831
rect 1315 3812 1328 3836
rect 1106 3807 1328 3812
rect 969 3804 1328 3807
rect 1390 3804 1425 3841
rect 1493 3838 1593 3841
rect 1493 3834 1560 3838
rect 1493 3808 1505 3834
rect 1531 3812 1560 3834
rect 1586 3812 1593 3838
rect 1531 3808 1593 3812
rect 1493 3804 1593 3808
rect 754 3788 765 3804
rect 754 3779 762 3788
rect 969 3783 1000 3804
rect 1390 3783 1426 3804
rect 812 3782 849 3783
rect 477 3739 542 3758
rect 477 3721 502 3739
rect 520 3721 542 3739
rect 477 3520 542 3721
rect 698 3595 762 3779
rect 811 3773 849 3782
rect 811 3753 820 3773
rect 840 3753 849 3773
rect 811 3745 849 3753
rect 915 3777 1000 3783
rect 1025 3782 1062 3783
rect 915 3757 923 3777
rect 943 3757 1000 3777
rect 915 3749 1000 3757
rect 1024 3773 1062 3782
rect 1024 3753 1033 3773
rect 1053 3753 1062 3773
rect 915 3748 951 3749
rect 1024 3745 1062 3753
rect 1128 3777 1213 3783
rect 1233 3782 1270 3783
rect 1128 3757 1136 3777
rect 1156 3776 1213 3777
rect 1156 3757 1185 3776
rect 1128 3756 1185 3757
rect 1206 3756 1213 3776
rect 1128 3749 1213 3756
rect 1232 3773 1270 3782
rect 1232 3753 1241 3773
rect 1261 3753 1270 3773
rect 1128 3748 1164 3749
rect 1232 3745 1270 3753
rect 1336 3777 1480 3783
rect 1336 3757 1344 3777
rect 1364 3757 1452 3777
rect 1472 3757 1480 3777
rect 1336 3749 1480 3757
rect 1336 3748 1372 3749
rect 1444 3748 1480 3749
rect 1546 3782 1583 3783
rect 1546 3781 1584 3782
rect 1546 3773 1610 3781
rect 1546 3753 1555 3773
rect 1575 3759 1610 3773
rect 1630 3759 1633 3779
rect 1575 3754 1633 3759
rect 1575 3753 1610 3754
rect 812 3716 849 3745
rect 813 3714 849 3716
rect 1025 3714 1062 3745
rect 813 3692 1062 3714
rect 894 3686 1005 3692
rect 894 3678 935 3686
rect 894 3658 902 3678
rect 921 3658 935 3678
rect 894 3656 935 3658
rect 963 3678 1005 3686
rect 963 3658 979 3678
rect 998 3658 1005 3678
rect 963 3656 1005 3658
rect 894 3641 1005 3656
rect 698 3585 766 3595
rect 698 3552 715 3585
rect 755 3552 766 3585
rect 698 3540 766 3552
rect 698 3538 762 3540
rect 1233 3521 1270 3745
rect 1546 3741 1610 3753
rect 1650 3523 1677 3893
rect 1865 3888 1902 3898
rect 1961 3918 2048 3928
rect 1961 3898 1970 3918
rect 1990 3898 2048 3918
rect 1961 3889 2048 3898
rect 1961 3888 1998 3889
rect 1741 3875 1811 3880
rect 1736 3869 1811 3875
rect 1736 3836 1744 3869
rect 1797 3836 1811 3869
rect 2017 3836 2048 3889
rect 2078 3918 2115 3997
rect 2230 3928 2261 3929
rect 2078 3898 2087 3918
rect 2107 3898 2115 3918
rect 2078 3888 2115 3898
rect 2174 3921 2261 3928
rect 2174 3918 2235 3921
rect 2174 3898 2183 3918
rect 2203 3901 2235 3918
rect 2256 3901 2261 3921
rect 2203 3898 2261 3901
rect 2174 3891 2261 3898
rect 2286 3918 2323 4060
rect 2589 4059 2626 4060
rect 2438 3928 2474 3929
rect 2286 3898 2295 3918
rect 2315 3898 2323 3918
rect 2174 3889 2230 3891
rect 2174 3888 2211 3889
rect 2286 3888 2323 3898
rect 2382 3918 2530 3928
rect 2630 3925 2726 3927
rect 2382 3898 2391 3918
rect 2411 3898 2501 3918
rect 2521 3898 2530 3918
rect 2382 3892 2530 3898
rect 2382 3889 2446 3892
rect 2382 3888 2419 3889
rect 2438 3862 2446 3889
rect 2467 3889 2530 3892
rect 2588 3918 2726 3925
rect 2588 3898 2597 3918
rect 2617 3898 2726 3918
rect 2588 3889 2726 3898
rect 2467 3862 2474 3889
rect 2493 3888 2530 3889
rect 2589 3888 2626 3889
rect 2438 3837 2474 3862
rect 1736 3835 1819 3836
rect 1909 3835 1950 3836
rect 1736 3828 1950 3835
rect 1736 3811 1919 3828
rect 1736 3778 1749 3811
rect 1802 3808 1919 3811
rect 1939 3808 1950 3828
rect 1802 3800 1950 3808
rect 2017 3832 2376 3836
rect 2017 3827 2339 3832
rect 2017 3803 2130 3827
rect 2154 3808 2339 3827
rect 2363 3808 2376 3832
rect 2154 3803 2376 3808
rect 2017 3800 2376 3803
rect 2438 3800 2473 3837
rect 2541 3834 2641 3837
rect 2541 3830 2608 3834
rect 2541 3804 2553 3830
rect 2579 3808 2608 3830
rect 2634 3808 2641 3834
rect 2579 3804 2641 3808
rect 2541 3800 2641 3804
rect 1802 3778 1819 3800
rect 2017 3779 2048 3800
rect 2438 3779 2474 3800
rect 1860 3778 1897 3779
rect 1736 3764 1819 3778
rect 1509 3521 1677 3523
rect 1233 3520 1677 3521
rect 477 3490 1677 3520
rect 1747 3554 1819 3764
rect 1859 3769 1897 3778
rect 1859 3749 1868 3769
rect 1888 3749 1897 3769
rect 1859 3741 1897 3749
rect 1963 3773 2048 3779
rect 2073 3778 2110 3779
rect 1963 3753 1971 3773
rect 1991 3753 2048 3773
rect 1963 3745 2048 3753
rect 2072 3769 2110 3778
rect 2072 3749 2081 3769
rect 2101 3749 2110 3769
rect 1963 3744 1999 3745
rect 2072 3741 2110 3749
rect 2176 3773 2261 3779
rect 2281 3778 2318 3779
rect 2176 3753 2184 3773
rect 2204 3772 2261 3773
rect 2204 3753 2233 3772
rect 2176 3752 2233 3753
rect 2254 3752 2261 3772
rect 2176 3745 2261 3752
rect 2280 3769 2318 3778
rect 2280 3749 2289 3769
rect 2309 3749 2318 3769
rect 2176 3744 2212 3745
rect 2280 3741 2318 3749
rect 2384 3773 2528 3779
rect 2384 3753 2392 3773
rect 2412 3753 2500 3773
rect 2520 3753 2528 3773
rect 2384 3745 2528 3753
rect 2384 3744 2420 3745
rect 2492 3744 2528 3745
rect 2594 3778 2631 3779
rect 2594 3777 2632 3778
rect 2594 3769 2658 3777
rect 2594 3749 2603 3769
rect 2623 3755 2658 3769
rect 2678 3755 2681 3775
rect 2623 3750 2681 3755
rect 2623 3749 2658 3750
rect 1860 3712 1897 3741
rect 1861 3710 1897 3712
rect 2073 3710 2110 3741
rect 1861 3688 2110 3710
rect 1942 3682 2053 3688
rect 1942 3674 1983 3682
rect 1942 3654 1950 3674
rect 1969 3654 1983 3674
rect 1942 3652 1983 3654
rect 2011 3674 2053 3682
rect 2011 3654 2027 3674
rect 2046 3654 2053 3674
rect 2011 3652 2053 3654
rect 1942 3637 2053 3652
rect 1747 3515 1766 3554
rect 1811 3515 1819 3554
rect 1747 3498 1819 3515
rect 2281 3542 2318 3741
rect 2594 3737 2658 3749
rect 2281 3536 2322 3542
rect 2698 3538 2725 3889
rect 2854 3841 2925 4320
rect 2854 3757 2923 3841
rect 2557 3536 2725 3538
rect 2281 3510 2725 3536
rect 477 3443 542 3490
rect 477 3425 500 3443
rect 518 3425 542 3443
rect 1390 3470 1425 3472
rect 1390 3468 1494 3470
rect 2283 3468 2322 3510
rect 2557 3509 2725 3510
rect 1390 3461 2324 3468
rect 1390 3460 1441 3461
rect 1390 3440 1393 3460
rect 1418 3441 1441 3460
rect 1473 3441 2324 3461
rect 1418 3440 2324 3441
rect 1390 3433 2324 3440
rect 1663 3432 2324 3433
rect 477 3404 542 3425
rect 754 3415 794 3418
rect 754 3411 1657 3415
rect 754 3391 1631 3411
rect 1651 3391 1657 3411
rect 754 3388 1657 3391
rect 478 3344 543 3364
rect 478 3326 502 3344
rect 520 3326 543 3344
rect 478 3299 543 3326
rect 754 3299 794 3388
rect 1238 3386 1654 3388
rect 1238 3385 1579 3386
rect 895 3354 1005 3368
rect 895 3351 938 3354
rect 895 3346 899 3351
rect 477 3264 794 3299
rect 817 3324 899 3346
rect 928 3324 938 3351
rect 966 3327 973 3354
rect 1002 3346 1005 3354
rect 1002 3327 1067 3346
rect 966 3324 1067 3327
rect 817 3322 1067 3324
rect 478 3188 543 3264
rect 817 3243 854 3322
rect 895 3309 1005 3322
rect 969 3253 1000 3254
rect 817 3223 826 3243
rect 846 3223 854 3243
rect 817 3213 854 3223
rect 913 3243 1000 3253
rect 913 3223 922 3243
rect 942 3223 1000 3243
rect 913 3214 1000 3223
rect 913 3213 950 3214
rect 478 3170 500 3188
rect 518 3170 543 3188
rect 478 3149 543 3170
rect 691 3168 756 3177
rect 691 3131 701 3168
rect 741 3160 756 3168
rect 969 3161 1000 3214
rect 1030 3243 1067 3322
rect 1182 3253 1213 3254
rect 1030 3223 1039 3243
rect 1059 3223 1067 3243
rect 1030 3213 1067 3223
rect 1126 3246 1213 3253
rect 1126 3243 1187 3246
rect 1126 3223 1135 3243
rect 1155 3226 1187 3243
rect 1208 3226 1213 3246
rect 1155 3223 1213 3226
rect 1126 3216 1213 3223
rect 1238 3243 1275 3385
rect 1541 3384 1578 3385
rect 1390 3253 1426 3254
rect 1238 3223 1247 3243
rect 1267 3223 1275 3243
rect 1126 3214 1182 3216
rect 1126 3213 1163 3214
rect 1238 3213 1275 3223
rect 1334 3243 1482 3253
rect 1582 3250 1678 3252
rect 1334 3223 1343 3243
rect 1363 3223 1453 3243
rect 1473 3223 1482 3243
rect 1334 3217 1482 3223
rect 1334 3214 1398 3217
rect 1334 3213 1371 3214
rect 1390 3187 1398 3214
rect 1419 3214 1482 3217
rect 1540 3243 1678 3250
rect 2858 3245 2920 3757
rect 1540 3223 1549 3243
rect 1569 3223 1678 3243
rect 1540 3214 1678 3223
rect 1419 3187 1426 3214
rect 1445 3213 1482 3214
rect 1541 3213 1578 3214
rect 1390 3162 1426 3187
rect 861 3160 902 3161
rect 741 3153 902 3160
rect 741 3133 871 3153
rect 891 3133 902 3153
rect 741 3131 902 3133
rect 691 3125 902 3131
rect 969 3157 1328 3161
rect 969 3152 1291 3157
rect 969 3128 1082 3152
rect 1106 3133 1291 3152
rect 1315 3133 1328 3157
rect 1106 3128 1328 3133
rect 969 3125 1328 3128
rect 1390 3125 1425 3162
rect 1493 3159 1593 3162
rect 1493 3155 1560 3159
rect 1493 3129 1505 3155
rect 1531 3133 1560 3155
rect 1586 3133 1593 3159
rect 1531 3129 1593 3133
rect 1493 3125 1593 3129
rect 691 3112 758 3125
rect 483 3089 539 3109
rect 483 3071 502 3089
rect 520 3071 539 3089
rect 483 2958 539 3071
rect 691 3091 705 3112
rect 741 3091 758 3112
rect 969 3104 1000 3125
rect 1390 3104 1426 3125
rect 812 3103 849 3104
rect 691 3084 758 3091
rect 811 3094 849 3103
rect 483 2820 538 2958
rect 691 2932 756 3084
rect 811 3074 820 3094
rect 840 3074 849 3094
rect 811 3066 849 3074
rect 915 3098 1000 3104
rect 1025 3103 1062 3104
rect 915 3078 923 3098
rect 943 3078 1000 3098
rect 915 3070 1000 3078
rect 1024 3094 1062 3103
rect 1024 3074 1033 3094
rect 1053 3074 1062 3094
rect 915 3069 951 3070
rect 1024 3066 1062 3074
rect 1128 3098 1213 3104
rect 1233 3103 1270 3104
rect 1128 3078 1136 3098
rect 1156 3097 1213 3098
rect 1156 3078 1185 3097
rect 1128 3077 1185 3078
rect 1206 3077 1213 3097
rect 1128 3070 1213 3077
rect 1232 3094 1270 3103
rect 1232 3074 1241 3094
rect 1261 3074 1270 3094
rect 1128 3069 1164 3070
rect 1232 3066 1270 3074
rect 1336 3098 1480 3104
rect 1336 3078 1344 3098
rect 1364 3078 1452 3098
rect 1472 3078 1480 3098
rect 1336 3070 1480 3078
rect 1336 3069 1372 3070
rect 1444 3069 1480 3070
rect 1546 3103 1583 3104
rect 1546 3102 1584 3103
rect 1546 3094 1610 3102
rect 1546 3074 1555 3094
rect 1575 3080 1610 3094
rect 1630 3080 1633 3100
rect 1575 3075 1633 3080
rect 1575 3074 1610 3075
rect 812 3037 849 3066
rect 813 3035 849 3037
rect 1025 3035 1062 3066
rect 813 3013 1062 3035
rect 894 3007 1005 3013
rect 894 2999 935 3007
rect 894 2979 902 2999
rect 921 2979 935 2999
rect 894 2977 935 2979
rect 963 2999 1005 3007
rect 963 2979 979 2999
rect 998 2979 1005 2999
rect 963 2977 1005 2979
rect 894 2964 1005 2977
rect 1233 2967 1270 3066
rect 1546 3062 1610 3074
rect 684 2922 805 2932
rect 684 2920 753 2922
rect 684 2879 697 2920
rect 734 2881 753 2920
rect 790 2881 805 2922
rect 734 2879 805 2881
rect 684 2861 805 2879
rect 476 2817 540 2820
rect 896 2817 1000 2823
rect 1231 2817 1272 2967
rect 1650 2959 1677 3214
rect 1739 3204 1819 3215
rect 1739 3178 1756 3204
rect 1796 3178 1819 3204
rect 1739 3151 1819 3178
rect 2862 3206 2920 3245
rect 2862 3171 2924 3206
rect 1739 3125 1760 3151
rect 1800 3125 1819 3151
rect 1739 3106 1819 3125
rect 1739 3080 1763 3106
rect 1803 3080 1819 3106
rect 1739 3029 1819 3080
rect 2811 3144 2924 3171
rect 2811 3142 2870 3144
rect 2811 3111 2825 3142
rect 2850 3121 2870 3142
rect 2896 3121 2924 3144
rect 2850 3111 2924 3121
rect 2811 3101 2924 3111
rect 476 2814 1272 2817
rect 1651 2828 1677 2959
rect 1651 2814 1679 2828
rect 476 2779 1679 2814
rect 1741 2821 1811 3029
rect 476 2718 540 2779
rect 896 2777 1000 2779
rect 1231 2777 1272 2779
rect 1741 2776 1762 2821
rect 1742 2755 1762 2776
rect 1792 2776 1811 2821
rect 1792 2755 1809 2776
rect 1742 2736 1809 2755
rect 1391 2728 1463 2729
rect 1390 2720 1489 2728
rect 478 2647 537 2718
rect 1390 2717 1442 2720
rect 1390 2682 1398 2717
rect 1423 2682 1442 2717
rect 1467 2709 1489 2720
rect 1467 2708 2334 2709
rect 1467 2682 2335 2708
rect 1390 2672 2335 2682
rect 1390 2670 1489 2672
rect 478 2629 500 2647
rect 518 2629 537 2647
rect 478 2607 537 2629
rect 745 2643 1277 2648
rect 745 2623 1631 2643
rect 1651 2623 1654 2643
rect 2290 2639 2335 2672
rect 745 2619 1654 2623
rect 745 2572 788 2619
rect 1238 2618 1654 2619
rect 2286 2619 2679 2639
rect 2699 2619 2702 2639
rect 1238 2617 1579 2618
rect 895 2586 1005 2600
rect 895 2583 938 2586
rect 895 2578 899 2583
rect 733 2571 788 2572
rect 477 2548 788 2571
rect 477 2530 502 2548
rect 520 2536 788 2548
rect 817 2556 899 2578
rect 928 2556 938 2583
rect 966 2559 973 2586
rect 1002 2578 1005 2586
rect 1002 2559 1067 2578
rect 966 2556 1067 2559
rect 817 2554 1067 2556
rect 520 2530 542 2536
rect 477 2391 542 2530
rect 817 2475 854 2554
rect 895 2541 1005 2554
rect 969 2485 1000 2486
rect 817 2455 826 2475
rect 846 2455 854 2475
rect 477 2373 500 2391
rect 518 2373 542 2391
rect 477 2356 542 2373
rect 697 2437 765 2450
rect 817 2445 854 2455
rect 913 2475 1000 2485
rect 913 2455 922 2475
rect 942 2455 1000 2475
rect 913 2446 1000 2455
rect 913 2445 950 2446
rect 697 2395 704 2437
rect 753 2395 765 2437
rect 697 2392 765 2395
rect 969 2393 1000 2446
rect 1030 2475 1067 2554
rect 1182 2485 1213 2486
rect 1030 2455 1039 2475
rect 1059 2455 1067 2475
rect 1030 2445 1067 2455
rect 1126 2478 1213 2485
rect 1126 2475 1187 2478
rect 1126 2455 1135 2475
rect 1155 2458 1187 2475
rect 1208 2458 1213 2478
rect 1155 2455 1213 2458
rect 1126 2448 1213 2455
rect 1238 2475 1275 2617
rect 1541 2616 1578 2617
rect 2286 2614 2702 2619
rect 2286 2613 2627 2614
rect 1943 2582 2053 2596
rect 1943 2579 1986 2582
rect 1943 2574 1947 2579
rect 1865 2552 1947 2574
rect 1976 2552 1986 2579
rect 2014 2555 2021 2582
rect 2050 2574 2053 2582
rect 2050 2555 2115 2574
rect 2014 2552 2115 2555
rect 1865 2550 2115 2552
rect 1390 2485 1426 2486
rect 1238 2455 1247 2475
rect 1267 2455 1275 2475
rect 1126 2446 1182 2448
rect 1126 2445 1163 2446
rect 1238 2445 1275 2455
rect 1334 2475 1482 2485
rect 1582 2482 1678 2484
rect 1334 2455 1343 2475
rect 1363 2455 1453 2475
rect 1473 2455 1482 2475
rect 1334 2449 1482 2455
rect 1334 2446 1398 2449
rect 1334 2445 1371 2446
rect 1390 2419 1398 2446
rect 1419 2446 1482 2449
rect 1540 2475 1678 2482
rect 1540 2455 1549 2475
rect 1569 2455 1678 2475
rect 1540 2446 1678 2455
rect 1865 2471 1902 2550
rect 1943 2537 2053 2550
rect 2017 2481 2048 2482
rect 1865 2451 1874 2471
rect 1894 2451 1902 2471
rect 1419 2419 1426 2446
rect 1445 2445 1482 2446
rect 1541 2445 1578 2446
rect 1390 2394 1426 2419
rect 861 2392 902 2393
rect 697 2385 902 2392
rect 697 2374 871 2385
rect 697 2341 705 2374
rect 698 2332 705 2341
rect 754 2365 871 2374
rect 891 2365 902 2385
rect 754 2357 902 2365
rect 969 2389 1328 2393
rect 969 2384 1291 2389
rect 969 2360 1082 2384
rect 1106 2365 1291 2384
rect 1315 2365 1328 2389
rect 1106 2360 1328 2365
rect 969 2357 1328 2360
rect 1390 2357 1425 2394
rect 1493 2391 1593 2394
rect 1493 2387 1560 2391
rect 1493 2361 1505 2387
rect 1531 2365 1560 2387
rect 1586 2365 1593 2391
rect 1531 2361 1593 2365
rect 1493 2357 1593 2361
rect 754 2341 765 2357
rect 754 2332 762 2341
rect 969 2336 1000 2357
rect 1390 2336 1426 2357
rect 812 2335 849 2336
rect 477 2292 542 2311
rect 477 2274 502 2292
rect 520 2274 542 2292
rect 477 2073 542 2274
rect 698 2148 762 2332
rect 811 2326 849 2335
rect 811 2306 820 2326
rect 840 2306 849 2326
rect 811 2298 849 2306
rect 915 2330 1000 2336
rect 1025 2335 1062 2336
rect 915 2310 923 2330
rect 943 2310 1000 2330
rect 915 2302 1000 2310
rect 1024 2326 1062 2335
rect 1024 2306 1033 2326
rect 1053 2306 1062 2326
rect 915 2301 951 2302
rect 1024 2298 1062 2306
rect 1128 2330 1213 2336
rect 1233 2335 1270 2336
rect 1128 2310 1136 2330
rect 1156 2329 1213 2330
rect 1156 2310 1185 2329
rect 1128 2309 1185 2310
rect 1206 2309 1213 2329
rect 1128 2302 1213 2309
rect 1232 2326 1270 2335
rect 1232 2306 1241 2326
rect 1261 2306 1270 2326
rect 1128 2301 1164 2302
rect 1232 2298 1270 2306
rect 1336 2330 1480 2336
rect 1336 2310 1344 2330
rect 1364 2310 1452 2330
rect 1472 2310 1480 2330
rect 1336 2302 1480 2310
rect 1336 2301 1372 2302
rect 1444 2301 1480 2302
rect 1546 2335 1583 2336
rect 1546 2334 1584 2335
rect 1546 2326 1610 2334
rect 1546 2306 1555 2326
rect 1575 2312 1610 2326
rect 1630 2312 1633 2332
rect 1575 2307 1633 2312
rect 1575 2306 1610 2307
rect 812 2269 849 2298
rect 813 2267 849 2269
rect 1025 2267 1062 2298
rect 813 2245 1062 2267
rect 894 2239 1005 2245
rect 894 2231 935 2239
rect 894 2211 902 2231
rect 921 2211 935 2231
rect 894 2209 935 2211
rect 963 2231 1005 2239
rect 963 2211 979 2231
rect 998 2211 1005 2231
rect 963 2209 1005 2211
rect 894 2194 1005 2209
rect 698 2138 766 2148
rect 698 2105 715 2138
rect 755 2105 766 2138
rect 698 2093 766 2105
rect 698 2091 762 2093
rect 1233 2074 1270 2298
rect 1546 2294 1610 2306
rect 1650 2076 1677 2446
rect 1865 2441 1902 2451
rect 1961 2471 2048 2481
rect 1961 2451 1970 2471
rect 1990 2451 2048 2471
rect 1961 2442 2048 2451
rect 1961 2441 1998 2442
rect 1741 2428 1811 2433
rect 1736 2422 1811 2428
rect 1736 2389 1744 2422
rect 1797 2389 1811 2422
rect 2017 2389 2048 2442
rect 2078 2471 2115 2550
rect 2230 2481 2261 2482
rect 2078 2451 2087 2471
rect 2107 2451 2115 2471
rect 2078 2441 2115 2451
rect 2174 2474 2261 2481
rect 2174 2471 2235 2474
rect 2174 2451 2183 2471
rect 2203 2454 2235 2471
rect 2256 2454 2261 2474
rect 2203 2451 2261 2454
rect 2174 2444 2261 2451
rect 2286 2471 2323 2613
rect 2589 2612 2626 2613
rect 2438 2481 2474 2482
rect 2286 2451 2295 2471
rect 2315 2451 2323 2471
rect 2174 2442 2230 2444
rect 2174 2441 2211 2442
rect 2286 2441 2323 2451
rect 2382 2471 2530 2481
rect 2630 2478 2726 2480
rect 2382 2451 2391 2471
rect 2411 2451 2501 2471
rect 2521 2451 2530 2471
rect 2382 2445 2530 2451
rect 2382 2442 2446 2445
rect 2382 2441 2419 2442
rect 2438 2415 2446 2442
rect 2467 2442 2530 2445
rect 2588 2471 2726 2478
rect 2588 2451 2597 2471
rect 2617 2451 2726 2471
rect 2588 2442 2726 2451
rect 2467 2415 2474 2442
rect 2493 2441 2530 2442
rect 2589 2441 2626 2442
rect 2438 2390 2474 2415
rect 1736 2388 1819 2389
rect 1909 2388 1950 2389
rect 1736 2381 1950 2388
rect 1736 2364 1919 2381
rect 1736 2331 1749 2364
rect 1802 2361 1919 2364
rect 1939 2361 1950 2381
rect 1802 2353 1950 2361
rect 2017 2385 2376 2389
rect 2017 2380 2339 2385
rect 2017 2356 2130 2380
rect 2154 2361 2339 2380
rect 2363 2361 2376 2385
rect 2154 2356 2376 2361
rect 2017 2353 2376 2356
rect 2438 2353 2473 2390
rect 2541 2387 2641 2390
rect 2541 2383 2608 2387
rect 2541 2357 2553 2383
rect 2579 2361 2608 2383
rect 2634 2361 2641 2387
rect 2579 2357 2641 2361
rect 2541 2353 2641 2357
rect 1802 2331 1819 2353
rect 2017 2332 2048 2353
rect 2438 2332 2474 2353
rect 1860 2331 1897 2332
rect 1736 2317 1819 2331
rect 1509 2074 1677 2076
rect 1233 2073 1677 2074
rect 477 2043 1677 2073
rect 1747 2107 1819 2317
rect 1859 2322 1897 2331
rect 1859 2302 1868 2322
rect 1888 2302 1897 2322
rect 1859 2294 1897 2302
rect 1963 2326 2048 2332
rect 2073 2331 2110 2332
rect 1963 2306 1971 2326
rect 1991 2306 2048 2326
rect 1963 2298 2048 2306
rect 2072 2322 2110 2331
rect 2072 2302 2081 2322
rect 2101 2302 2110 2322
rect 1963 2297 1999 2298
rect 2072 2294 2110 2302
rect 2176 2326 2261 2332
rect 2281 2331 2318 2332
rect 2176 2306 2184 2326
rect 2204 2325 2261 2326
rect 2204 2306 2233 2325
rect 2176 2305 2233 2306
rect 2254 2305 2261 2325
rect 2176 2298 2261 2305
rect 2280 2322 2318 2331
rect 2280 2302 2289 2322
rect 2309 2302 2318 2322
rect 2176 2297 2212 2298
rect 2280 2294 2318 2302
rect 2384 2326 2528 2332
rect 2384 2306 2392 2326
rect 2412 2306 2500 2326
rect 2520 2306 2528 2326
rect 2384 2298 2528 2306
rect 2384 2297 2420 2298
rect 2492 2297 2528 2298
rect 2594 2331 2631 2332
rect 2594 2330 2632 2331
rect 2594 2322 2658 2330
rect 2594 2302 2603 2322
rect 2623 2308 2658 2322
rect 2678 2308 2681 2328
rect 2623 2303 2681 2308
rect 2623 2302 2658 2303
rect 1860 2265 1897 2294
rect 1861 2263 1897 2265
rect 2073 2263 2110 2294
rect 1861 2241 2110 2263
rect 1942 2235 2053 2241
rect 1942 2227 1983 2235
rect 1942 2207 1950 2227
rect 1969 2207 1983 2227
rect 1942 2205 1983 2207
rect 2011 2227 2053 2235
rect 2011 2207 2027 2227
rect 2046 2207 2053 2227
rect 2011 2205 2053 2207
rect 1942 2190 2053 2205
rect 1747 2068 1766 2107
rect 1811 2068 1819 2107
rect 1747 2051 1819 2068
rect 2281 2095 2318 2294
rect 2594 2290 2658 2302
rect 2281 2089 2322 2095
rect 2698 2091 2725 2442
rect 2557 2089 2725 2091
rect 2281 2063 2725 2089
rect 477 1996 542 2043
rect 477 1978 500 1996
rect 518 1978 542 1996
rect 1390 2023 1425 2025
rect 1390 2021 1494 2023
rect 2283 2021 2322 2063
rect 2557 2062 2725 2063
rect 1390 2014 2324 2021
rect 1390 2013 1441 2014
rect 1390 1993 1393 2013
rect 1418 1994 1441 2013
rect 1473 1994 2324 2014
rect 1418 1993 2324 1994
rect 1390 1986 2324 1993
rect 1663 1985 2324 1986
rect 477 1957 542 1978
rect 754 1968 794 1971
rect 754 1964 1657 1968
rect 754 1944 1631 1964
rect 1651 1944 1657 1964
rect 754 1941 1657 1944
rect 478 1897 543 1917
rect 478 1879 502 1897
rect 520 1879 543 1897
rect 478 1852 543 1879
rect 754 1852 794 1941
rect 1238 1939 1654 1941
rect 1238 1938 1579 1939
rect 895 1907 1005 1921
rect 895 1904 938 1907
rect 895 1899 899 1904
rect 477 1817 794 1852
rect 817 1877 899 1899
rect 928 1877 938 1904
rect 966 1880 973 1907
rect 1002 1899 1005 1907
rect 1002 1880 1067 1899
rect 966 1877 1067 1880
rect 817 1875 1067 1877
rect 478 1741 543 1817
rect 817 1796 854 1875
rect 895 1862 1005 1875
rect 969 1806 1000 1807
rect 817 1776 826 1796
rect 846 1776 854 1796
rect 817 1766 854 1776
rect 913 1796 1000 1806
rect 913 1776 922 1796
rect 942 1776 1000 1796
rect 913 1767 1000 1776
rect 913 1766 950 1767
rect 478 1723 500 1741
rect 518 1723 543 1741
rect 478 1702 543 1723
rect 691 1721 756 1730
rect 691 1684 701 1721
rect 741 1713 756 1721
rect 969 1714 1000 1767
rect 1030 1796 1067 1875
rect 1182 1806 1213 1807
rect 1030 1776 1039 1796
rect 1059 1776 1067 1796
rect 1030 1766 1067 1776
rect 1126 1799 1213 1806
rect 1126 1796 1187 1799
rect 1126 1776 1135 1796
rect 1155 1779 1187 1796
rect 1208 1779 1213 1799
rect 1155 1776 1213 1779
rect 1126 1769 1213 1776
rect 1238 1796 1275 1938
rect 1541 1937 1578 1938
rect 1390 1806 1426 1807
rect 1238 1776 1247 1796
rect 1267 1776 1275 1796
rect 1126 1767 1182 1769
rect 1126 1766 1163 1767
rect 1238 1766 1275 1776
rect 1334 1796 1482 1806
rect 1582 1803 1678 1805
rect 1334 1776 1343 1796
rect 1363 1776 1453 1796
rect 1473 1776 1482 1796
rect 1334 1770 1482 1776
rect 1334 1767 1398 1770
rect 1334 1766 1371 1767
rect 1390 1740 1398 1767
rect 1419 1767 1482 1770
rect 1540 1796 1678 1803
rect 1540 1776 1549 1796
rect 1569 1776 1678 1796
rect 1540 1767 1678 1776
rect 1419 1740 1426 1767
rect 1445 1766 1482 1767
rect 1541 1766 1578 1767
rect 1390 1715 1426 1740
rect 861 1713 902 1714
rect 741 1706 902 1713
rect 741 1686 871 1706
rect 891 1686 902 1706
rect 741 1684 902 1686
rect 691 1678 902 1684
rect 969 1710 1328 1714
rect 969 1705 1291 1710
rect 969 1681 1082 1705
rect 1106 1686 1291 1705
rect 1315 1686 1328 1710
rect 1106 1681 1328 1686
rect 969 1678 1328 1681
rect 1390 1678 1425 1715
rect 1493 1712 1593 1715
rect 1493 1708 1560 1712
rect 1493 1682 1505 1708
rect 1531 1686 1560 1708
rect 1586 1686 1593 1712
rect 1531 1682 1593 1686
rect 1493 1678 1593 1682
rect 691 1665 758 1678
rect 483 1642 539 1662
rect 483 1624 502 1642
rect 520 1624 539 1642
rect 483 1589 539 1624
rect 445 1511 539 1589
rect 691 1644 705 1665
rect 741 1644 758 1665
rect 969 1657 1000 1678
rect 1390 1657 1426 1678
rect 812 1656 849 1657
rect 691 1637 758 1644
rect 811 1647 849 1656
rect 445 1370 538 1511
rect 691 1485 756 1637
rect 811 1627 820 1647
rect 840 1627 849 1647
rect 811 1619 849 1627
rect 915 1651 1000 1657
rect 1025 1656 1062 1657
rect 915 1631 923 1651
rect 943 1631 1000 1651
rect 915 1623 1000 1631
rect 1024 1647 1062 1656
rect 1024 1627 1033 1647
rect 1053 1627 1062 1647
rect 915 1622 951 1623
rect 1024 1619 1062 1627
rect 1128 1651 1213 1657
rect 1233 1656 1270 1657
rect 1128 1631 1136 1651
rect 1156 1650 1213 1651
rect 1156 1631 1185 1650
rect 1128 1630 1185 1631
rect 1206 1630 1213 1650
rect 1128 1623 1213 1630
rect 1232 1647 1270 1656
rect 1232 1627 1241 1647
rect 1261 1627 1270 1647
rect 1128 1622 1164 1623
rect 1232 1619 1270 1627
rect 1336 1651 1480 1657
rect 1336 1631 1344 1651
rect 1364 1631 1452 1651
rect 1472 1631 1480 1651
rect 1336 1623 1480 1631
rect 1336 1622 1372 1623
rect 1444 1622 1480 1623
rect 1546 1656 1583 1657
rect 1546 1655 1584 1656
rect 1546 1647 1610 1655
rect 1546 1627 1555 1647
rect 1575 1633 1610 1647
rect 1630 1633 1633 1653
rect 1575 1628 1633 1633
rect 1575 1627 1610 1628
rect 812 1590 849 1619
rect 813 1588 849 1590
rect 1025 1588 1062 1619
rect 813 1566 1062 1588
rect 894 1560 1005 1566
rect 894 1552 935 1560
rect 894 1532 902 1552
rect 921 1532 935 1552
rect 894 1530 935 1532
rect 963 1552 1005 1560
rect 963 1532 979 1552
rect 998 1532 1005 1552
rect 963 1530 1005 1532
rect 894 1515 1005 1530
rect 1233 1520 1270 1619
rect 1546 1615 1610 1627
rect 1650 1576 1677 1767
rect 896 1506 1000 1515
rect 684 1475 805 1485
rect 684 1473 753 1475
rect 684 1432 697 1473
rect 734 1434 753 1473
rect 790 1434 805 1475
rect 734 1432 805 1434
rect 684 1414 805 1432
rect 896 1370 1000 1379
rect 1231 1370 1272 1520
rect 445 1368 1272 1370
rect 453 1367 1272 1368
rect 1651 1486 1676 1576
rect 2811 1544 2910 3101
rect 3016 1737 3115 4638
rect 3506 4621 3537 4642
rect 3927 4621 3963 4642
rect 3349 4620 3386 4621
rect 3348 4611 3386 4620
rect 3348 4591 3357 4611
rect 3377 4591 3386 4611
rect 3348 4583 3386 4591
rect 3452 4615 3537 4621
rect 3562 4620 3599 4621
rect 3452 4595 3460 4615
rect 3480 4595 3537 4615
rect 3452 4587 3537 4595
rect 3561 4611 3599 4620
rect 3561 4591 3570 4611
rect 3590 4591 3599 4611
rect 3452 4586 3488 4587
rect 3561 4583 3599 4591
rect 3665 4615 3750 4621
rect 3770 4620 3807 4621
rect 3665 4595 3673 4615
rect 3693 4614 3750 4615
rect 3693 4595 3722 4614
rect 3665 4594 3722 4595
rect 3743 4594 3750 4614
rect 3665 4587 3750 4594
rect 3769 4611 3807 4620
rect 3769 4591 3778 4611
rect 3798 4591 3807 4611
rect 3665 4586 3701 4587
rect 3769 4583 3807 4591
rect 3873 4615 4017 4621
rect 3873 4595 3881 4615
rect 3901 4595 3989 4615
rect 4009 4595 4017 4615
rect 3873 4587 4017 4595
rect 3873 4586 3909 4587
rect 3981 4586 4017 4587
rect 4083 4620 4120 4621
rect 4083 4619 4121 4620
rect 4083 4611 4147 4619
rect 4083 4591 4092 4611
rect 4112 4597 4147 4611
rect 4167 4597 4170 4617
rect 4112 4592 4170 4597
rect 4112 4591 4147 4592
rect 3349 4554 3386 4583
rect 3350 4552 3386 4554
rect 3562 4552 3599 4583
rect 3350 4530 3599 4552
rect 3431 4524 3542 4530
rect 3431 4516 3472 4524
rect 3431 4496 3439 4516
rect 3458 4496 3472 4516
rect 3431 4494 3472 4496
rect 3500 4516 3542 4524
rect 3500 4496 3516 4516
rect 3535 4496 3542 4516
rect 3500 4494 3542 4496
rect 3431 4479 3542 4494
rect 3770 4462 3807 4583
rect 4083 4579 4147 4591
rect 3888 4462 3917 4466
rect 4187 4464 4214 4731
rect 4046 4462 4214 4464
rect 3770 4436 4214 4462
rect 3729 4168 3774 4177
rect 3729 4130 3739 4168
rect 3764 4130 3774 4168
rect 3729 4119 3774 4130
rect 3732 4111 3774 4119
rect 3732 3406 3775 4111
rect 3888 3497 3917 4436
rect 4046 4435 4214 4436
rect 4618 4286 4702 4290
rect 5170 4286 5258 7137
rect 5797 7124 5852 7136
rect 5797 7090 5815 7124
rect 5844 7090 5852 7124
rect 5797 7064 5852 7090
rect 5404 7031 5572 7032
rect 5797 7031 5814 7064
rect 5404 7030 5814 7031
rect 5843 7030 5852 7064
rect 5404 7005 5852 7030
rect 5404 7003 5572 7005
rect 5404 6736 5431 7003
rect 5797 6999 5852 7005
rect 5471 6876 5535 6888
rect 5811 6884 5848 6999
rect 6076 6973 6187 6988
rect 6076 6971 6118 6973
rect 6076 6951 6083 6971
rect 6102 6951 6118 6971
rect 6076 6943 6118 6951
rect 6146 6971 6187 6973
rect 6146 6951 6160 6971
rect 6179 6951 6187 6971
rect 6146 6943 6187 6951
rect 6076 6937 6187 6943
rect 6019 6915 6268 6937
rect 6019 6884 6056 6915
rect 6232 6913 6268 6915
rect 6232 6884 6269 6913
rect 5471 6875 5506 6876
rect 5448 6870 5506 6875
rect 5448 6850 5451 6870
rect 5471 6856 5506 6870
rect 5526 6856 5535 6876
rect 5471 6848 5535 6856
rect 5497 6847 5535 6848
rect 5498 6846 5535 6847
rect 5601 6880 5637 6881
rect 5709 6880 5745 6881
rect 5601 6872 5745 6880
rect 5601 6852 5609 6872
rect 5629 6852 5717 6872
rect 5737 6852 5745 6872
rect 5601 6846 5745 6852
rect 5811 6876 5849 6884
rect 5917 6880 5953 6881
rect 5811 6856 5820 6876
rect 5840 6856 5849 6876
rect 5811 6847 5849 6856
rect 5868 6873 5953 6880
rect 5868 6853 5875 6873
rect 5896 6872 5953 6873
rect 5896 6853 5925 6872
rect 5868 6852 5925 6853
rect 5945 6852 5953 6872
rect 5811 6846 5848 6847
rect 5868 6846 5953 6852
rect 6019 6876 6057 6884
rect 6130 6880 6166 6881
rect 6019 6856 6028 6876
rect 6048 6856 6057 6876
rect 6019 6847 6057 6856
rect 6081 6872 6166 6880
rect 6081 6852 6138 6872
rect 6158 6852 6166 6872
rect 6019 6846 6056 6847
rect 6081 6846 6166 6852
rect 6232 6876 6270 6884
rect 6232 6856 6241 6876
rect 6261 6856 6270 6876
rect 6232 6847 6270 6856
rect 6232 6846 6269 6847
rect 5655 6825 5691 6846
rect 6081 6825 6112 6846
rect 6326 6829 6397 7482
rect 6912 7416 6955 8129
rect 7572 8040 7667 8060
rect 7572 7996 7592 8040
rect 7652 7996 7667 8040
rect 7572 7700 7667 7996
rect 7572 7659 7605 7700
rect 7641 7659 7667 7700
rect 7767 7739 7829 8210
rect 9109 8150 9146 8151
rect 9412 8150 9449 8292
rect 9474 8312 9561 8319
rect 9474 8309 9532 8312
rect 9474 8289 9479 8309
rect 9500 8292 9532 8309
rect 9552 8292 9561 8312
rect 9500 8289 9561 8292
rect 9474 8282 9561 8289
rect 9620 8312 9657 8322
rect 9620 8292 9628 8312
rect 9648 8292 9657 8312
rect 9474 8281 9505 8282
rect 9620 8213 9657 8292
rect 9687 8321 9718 8374
rect 9931 8367 9946 8375
rect 9986 8367 9996 8404
rect 11187 8393 11252 8532
rect 11527 8477 11564 8556
rect 11605 8543 11715 8556
rect 11679 8487 11710 8488
rect 11527 8457 11536 8477
rect 11556 8457 11564 8477
rect 9931 8358 9996 8367
rect 10144 8365 10209 8386
rect 10144 8347 10169 8365
rect 10187 8347 10209 8365
rect 11187 8375 11210 8393
rect 11228 8375 11252 8393
rect 11187 8358 11252 8375
rect 11407 8439 11475 8452
rect 11527 8447 11564 8457
rect 11623 8477 11710 8487
rect 11623 8457 11632 8477
rect 11652 8457 11710 8477
rect 11623 8448 11710 8457
rect 11623 8447 11660 8448
rect 11407 8397 11414 8439
rect 11463 8397 11475 8439
rect 11407 8394 11475 8397
rect 11679 8395 11710 8448
rect 11740 8477 11777 8556
rect 11892 8487 11923 8488
rect 11740 8457 11749 8477
rect 11769 8457 11777 8477
rect 11740 8447 11777 8457
rect 11836 8480 11923 8487
rect 11836 8477 11897 8480
rect 11836 8457 11845 8477
rect 11865 8460 11897 8477
rect 11918 8460 11923 8480
rect 11865 8457 11923 8460
rect 11836 8450 11923 8457
rect 11948 8477 11985 8619
rect 12251 8618 12288 8619
rect 12996 8616 13412 8621
rect 12996 8615 13337 8616
rect 12653 8584 12763 8598
rect 12653 8581 12696 8584
rect 12653 8576 12657 8581
rect 12575 8554 12657 8576
rect 12686 8554 12696 8581
rect 12724 8557 12731 8584
rect 12760 8576 12763 8584
rect 12760 8557 12825 8576
rect 12724 8554 12825 8557
rect 12575 8552 12825 8554
rect 12100 8487 12136 8488
rect 11948 8457 11957 8477
rect 11977 8457 11985 8477
rect 11836 8448 11892 8450
rect 11836 8447 11873 8448
rect 11948 8447 11985 8457
rect 12044 8477 12192 8487
rect 12292 8484 12388 8486
rect 12044 8457 12053 8477
rect 12073 8457 12163 8477
rect 12183 8457 12192 8477
rect 12044 8451 12192 8457
rect 12044 8448 12108 8451
rect 12044 8447 12081 8448
rect 12100 8421 12108 8448
rect 12129 8448 12192 8451
rect 12250 8477 12388 8484
rect 12250 8457 12259 8477
rect 12279 8457 12388 8477
rect 12250 8448 12388 8457
rect 12575 8473 12612 8552
rect 12653 8539 12763 8552
rect 12727 8483 12758 8484
rect 12575 8453 12584 8473
rect 12604 8453 12612 8473
rect 12129 8421 12136 8448
rect 12155 8447 12192 8448
rect 12251 8447 12288 8448
rect 12100 8396 12136 8421
rect 11571 8394 11612 8395
rect 11407 8387 11612 8394
rect 11407 8376 11581 8387
rect 9737 8321 9774 8322
rect 9687 8312 9774 8321
rect 9687 8292 9745 8312
rect 9765 8292 9774 8312
rect 9687 8282 9774 8292
rect 9833 8312 9870 8322
rect 9833 8292 9841 8312
rect 9861 8292 9870 8312
rect 9687 8281 9718 8282
rect 9682 8213 9792 8226
rect 9833 8213 9870 8292
rect 10144 8271 10209 8347
rect 11407 8343 11415 8376
rect 11408 8334 11415 8343
rect 11464 8367 11581 8376
rect 11601 8367 11612 8387
rect 11464 8359 11612 8367
rect 11679 8391 12038 8395
rect 11679 8386 12001 8391
rect 11679 8362 11792 8386
rect 11816 8367 12001 8386
rect 12025 8367 12038 8391
rect 11816 8362 12038 8367
rect 11679 8359 12038 8362
rect 12100 8359 12135 8396
rect 12203 8393 12303 8396
rect 12203 8389 12270 8393
rect 12203 8363 12215 8389
rect 12241 8367 12270 8389
rect 12296 8367 12303 8393
rect 12241 8363 12303 8367
rect 12203 8359 12303 8363
rect 11464 8343 11475 8359
rect 11464 8334 11472 8343
rect 11679 8338 11710 8359
rect 12100 8338 12136 8359
rect 11522 8337 11559 8338
rect 11187 8294 11252 8313
rect 11187 8276 11212 8294
rect 11230 8276 11252 8294
rect 9620 8211 9870 8213
rect 9620 8208 9721 8211
rect 9620 8189 9685 8208
rect 9682 8181 9685 8189
rect 9714 8181 9721 8208
rect 9749 8184 9759 8211
rect 9788 8189 9870 8211
rect 9893 8236 10210 8271
rect 9788 8184 9792 8189
rect 9749 8181 9792 8184
rect 9682 8167 9792 8181
rect 9108 8149 9449 8150
rect 9033 8147 9449 8149
rect 9893 8147 9933 8236
rect 10144 8209 10209 8236
rect 10144 8191 10167 8209
rect 10185 8191 10209 8209
rect 10144 8171 10209 8191
rect 9030 8144 9933 8147
rect 9030 8124 9036 8144
rect 9056 8124 9933 8144
rect 9030 8120 9933 8124
rect 9893 8117 9933 8120
rect 10145 8110 10210 8131
rect 8363 8102 9024 8103
rect 8363 8095 9297 8102
rect 8363 8094 9269 8095
rect 8363 8074 9214 8094
rect 9246 8075 9269 8094
rect 9294 8075 9297 8095
rect 9246 8074 9297 8075
rect 8363 8067 9297 8074
rect 7962 8025 8130 8026
rect 8365 8025 8404 8067
rect 9193 8065 9297 8067
rect 9262 8063 9297 8065
rect 10145 8092 10169 8110
rect 10187 8092 10210 8110
rect 10145 8045 10210 8092
rect 7962 7999 8406 8025
rect 7962 7997 8130 7999
rect 7767 7720 7831 7739
rect 7767 7681 7784 7720
rect 7818 7681 7831 7720
rect 7767 7662 7831 7681
rect 7572 7633 7667 7659
rect 7962 7646 7989 7997
rect 8365 7993 8406 7999
rect 8029 7786 8093 7798
rect 8369 7794 8406 7993
rect 8868 8020 8940 8037
rect 8868 7981 8876 8020
rect 8921 7981 8940 8020
rect 8634 7883 8745 7898
rect 8634 7881 8676 7883
rect 8634 7861 8641 7881
rect 8660 7861 8676 7881
rect 8634 7853 8676 7861
rect 8704 7881 8745 7883
rect 8704 7861 8718 7881
rect 8737 7861 8745 7881
rect 8704 7853 8745 7861
rect 8634 7847 8745 7853
rect 8577 7825 8826 7847
rect 8577 7794 8614 7825
rect 8790 7823 8826 7825
rect 8790 7794 8827 7823
rect 8029 7785 8064 7786
rect 8006 7780 8064 7785
rect 8006 7760 8009 7780
rect 8029 7766 8064 7780
rect 8084 7766 8093 7786
rect 8029 7758 8093 7766
rect 8055 7757 8093 7758
rect 8056 7756 8093 7757
rect 8159 7790 8195 7791
rect 8267 7790 8303 7791
rect 8159 7782 8303 7790
rect 8159 7762 8167 7782
rect 8187 7762 8275 7782
rect 8295 7762 8303 7782
rect 8159 7756 8303 7762
rect 8369 7786 8407 7794
rect 8475 7790 8511 7791
rect 8369 7766 8378 7786
rect 8398 7766 8407 7786
rect 8369 7757 8407 7766
rect 8426 7783 8511 7790
rect 8426 7763 8433 7783
rect 8454 7782 8511 7783
rect 8454 7763 8483 7782
rect 8426 7762 8483 7763
rect 8503 7762 8511 7782
rect 8369 7756 8406 7757
rect 8426 7756 8511 7762
rect 8577 7786 8615 7794
rect 8688 7790 8724 7791
rect 8577 7766 8586 7786
rect 8606 7766 8615 7786
rect 8577 7757 8615 7766
rect 8639 7782 8724 7790
rect 8639 7762 8696 7782
rect 8716 7762 8724 7782
rect 8577 7756 8614 7757
rect 8639 7756 8724 7762
rect 8790 7786 8828 7794
rect 8790 7766 8799 7786
rect 8819 7766 8828 7786
rect 8790 7757 8828 7766
rect 8868 7771 8940 7981
rect 9010 8015 10210 8045
rect 9010 8014 9454 8015
rect 9010 8012 9178 8014
rect 8868 7757 8951 7771
rect 8790 7756 8827 7757
rect 8213 7735 8249 7756
rect 8639 7735 8670 7756
rect 8868 7735 8885 7757
rect 8046 7731 8146 7735
rect 8046 7727 8108 7731
rect 8046 7701 8053 7727
rect 8079 7705 8108 7727
rect 8134 7705 8146 7731
rect 8079 7701 8146 7705
rect 8046 7698 8146 7701
rect 8214 7698 8249 7735
rect 8311 7732 8670 7735
rect 8311 7727 8533 7732
rect 8311 7703 8324 7727
rect 8348 7708 8533 7727
rect 8557 7708 8670 7732
rect 8348 7703 8670 7708
rect 8311 7699 8670 7703
rect 8737 7727 8885 7735
rect 8737 7707 8748 7727
rect 8768 7724 8885 7727
rect 8938 7724 8951 7757
rect 8768 7707 8951 7724
rect 8737 7700 8951 7707
rect 8737 7699 8778 7700
rect 8868 7699 8951 7700
rect 8213 7673 8249 7698
rect 8061 7646 8098 7647
rect 8157 7646 8194 7647
rect 8213 7646 8220 7673
rect 7961 7637 8099 7646
rect 7961 7617 8070 7637
rect 8090 7617 8099 7637
rect 7961 7610 8099 7617
rect 8157 7643 8220 7646
rect 8241 7646 8249 7673
rect 8268 7646 8305 7647
rect 8241 7643 8305 7646
rect 8157 7637 8305 7643
rect 8157 7617 8166 7637
rect 8186 7617 8276 7637
rect 8296 7617 8305 7637
rect 7961 7608 8057 7610
rect 8157 7607 8305 7617
rect 8364 7637 8401 7647
rect 8476 7646 8513 7647
rect 8457 7644 8513 7646
rect 8364 7617 8372 7637
rect 8392 7617 8401 7637
rect 8213 7606 8249 7607
rect 8061 7475 8098 7476
rect 8364 7475 8401 7617
rect 8426 7637 8513 7644
rect 8426 7634 8484 7637
rect 8426 7614 8431 7634
rect 8452 7617 8484 7634
rect 8504 7617 8513 7637
rect 8452 7614 8513 7617
rect 8426 7607 8513 7614
rect 8572 7637 8609 7647
rect 8572 7617 8580 7637
rect 8600 7617 8609 7637
rect 8426 7606 8457 7607
rect 8572 7538 8609 7617
rect 8639 7646 8670 7699
rect 8876 7666 8890 7699
rect 8943 7666 8951 7699
rect 8876 7660 8951 7666
rect 8876 7655 8946 7660
rect 8689 7646 8726 7647
rect 8639 7637 8726 7646
rect 8639 7617 8697 7637
rect 8717 7617 8726 7637
rect 8639 7607 8726 7617
rect 8785 7637 8822 7647
rect 9010 7642 9037 8012
rect 9077 7782 9141 7794
rect 9417 7790 9454 8014
rect 9925 7995 9989 7997
rect 9921 7983 9989 7995
rect 9921 7950 9932 7983
rect 9972 7950 9989 7983
rect 9921 7940 9989 7950
rect 9682 7879 9793 7894
rect 9682 7877 9724 7879
rect 9682 7857 9689 7877
rect 9708 7857 9724 7877
rect 9682 7849 9724 7857
rect 9752 7877 9793 7879
rect 9752 7857 9766 7877
rect 9785 7857 9793 7877
rect 9752 7849 9793 7857
rect 9682 7843 9793 7849
rect 9625 7821 9874 7843
rect 9625 7790 9662 7821
rect 9838 7819 9874 7821
rect 9838 7790 9875 7819
rect 9077 7781 9112 7782
rect 9054 7776 9112 7781
rect 9054 7756 9057 7776
rect 9077 7762 9112 7776
rect 9132 7762 9141 7782
rect 9077 7754 9141 7762
rect 9103 7753 9141 7754
rect 9104 7752 9141 7753
rect 9207 7786 9243 7787
rect 9315 7786 9351 7787
rect 9207 7778 9351 7786
rect 9207 7758 9215 7778
rect 9235 7758 9323 7778
rect 9343 7758 9351 7778
rect 9207 7752 9351 7758
rect 9417 7782 9455 7790
rect 9523 7786 9559 7787
rect 9417 7762 9426 7782
rect 9446 7762 9455 7782
rect 9417 7753 9455 7762
rect 9474 7779 9559 7786
rect 9474 7759 9481 7779
rect 9502 7778 9559 7779
rect 9502 7759 9531 7778
rect 9474 7758 9531 7759
rect 9551 7758 9559 7778
rect 9417 7752 9454 7753
rect 9474 7752 9559 7758
rect 9625 7782 9663 7790
rect 9736 7786 9772 7787
rect 9625 7762 9634 7782
rect 9654 7762 9663 7782
rect 9625 7753 9663 7762
rect 9687 7778 9772 7786
rect 9687 7758 9744 7778
rect 9764 7758 9772 7778
rect 9625 7752 9662 7753
rect 9687 7752 9772 7758
rect 9838 7782 9876 7790
rect 9838 7762 9847 7782
rect 9867 7762 9876 7782
rect 9838 7753 9876 7762
rect 9925 7756 9989 7940
rect 10145 7814 10210 8015
rect 11187 8075 11252 8276
rect 11408 8150 11472 8334
rect 11521 8328 11559 8337
rect 11521 8308 11530 8328
rect 11550 8308 11559 8328
rect 11521 8300 11559 8308
rect 11625 8332 11710 8338
rect 11735 8337 11772 8338
rect 11625 8312 11633 8332
rect 11653 8312 11710 8332
rect 11625 8304 11710 8312
rect 11734 8328 11772 8337
rect 11734 8308 11743 8328
rect 11763 8308 11772 8328
rect 11625 8303 11661 8304
rect 11734 8300 11772 8308
rect 11838 8332 11923 8338
rect 11943 8337 11980 8338
rect 11838 8312 11846 8332
rect 11866 8331 11923 8332
rect 11866 8312 11895 8331
rect 11838 8311 11895 8312
rect 11916 8311 11923 8331
rect 11838 8304 11923 8311
rect 11942 8328 11980 8337
rect 11942 8308 11951 8328
rect 11971 8308 11980 8328
rect 11838 8303 11874 8304
rect 11942 8300 11980 8308
rect 12046 8332 12190 8338
rect 12046 8312 12054 8332
rect 12074 8312 12162 8332
rect 12182 8312 12190 8332
rect 12046 8304 12190 8312
rect 12046 8303 12082 8304
rect 12154 8303 12190 8304
rect 12256 8337 12293 8338
rect 12256 8336 12294 8337
rect 12256 8328 12320 8336
rect 12256 8308 12265 8328
rect 12285 8314 12320 8328
rect 12340 8314 12343 8334
rect 12285 8309 12343 8314
rect 12285 8308 12320 8309
rect 11522 8271 11559 8300
rect 11523 8269 11559 8271
rect 11735 8269 11772 8300
rect 11523 8247 11772 8269
rect 11604 8241 11715 8247
rect 11604 8233 11645 8241
rect 11604 8213 11612 8233
rect 11631 8213 11645 8233
rect 11604 8211 11645 8213
rect 11673 8233 11715 8241
rect 11673 8213 11689 8233
rect 11708 8213 11715 8233
rect 11673 8211 11715 8213
rect 11604 8196 11715 8211
rect 11408 8140 11476 8150
rect 11408 8107 11425 8140
rect 11465 8107 11476 8140
rect 11408 8095 11476 8107
rect 11408 8093 11472 8095
rect 11943 8076 11980 8300
rect 12256 8296 12320 8308
rect 12360 8078 12387 8448
rect 12575 8443 12612 8453
rect 12671 8473 12758 8483
rect 12671 8453 12680 8473
rect 12700 8453 12758 8473
rect 12671 8444 12758 8453
rect 12671 8443 12708 8444
rect 12451 8430 12521 8435
rect 12446 8424 12521 8430
rect 12446 8391 12454 8424
rect 12507 8391 12521 8424
rect 12727 8391 12758 8444
rect 12788 8473 12825 8552
rect 12940 8483 12971 8484
rect 12788 8453 12797 8473
rect 12817 8453 12825 8473
rect 12788 8443 12825 8453
rect 12884 8476 12971 8483
rect 12884 8473 12945 8476
rect 12884 8453 12893 8473
rect 12913 8456 12945 8473
rect 12966 8456 12971 8476
rect 12913 8453 12971 8456
rect 12884 8446 12971 8453
rect 12996 8473 13033 8615
rect 13299 8614 13336 8615
rect 13148 8483 13184 8484
rect 12996 8453 13005 8473
rect 13025 8453 13033 8473
rect 12884 8444 12940 8446
rect 12884 8443 12921 8444
rect 12996 8443 13033 8453
rect 13092 8473 13240 8483
rect 13340 8480 13436 8482
rect 13092 8453 13101 8473
rect 13121 8453 13211 8473
rect 13231 8453 13240 8473
rect 13092 8447 13240 8453
rect 13092 8444 13156 8447
rect 13092 8443 13129 8444
rect 13148 8417 13156 8444
rect 13177 8444 13240 8447
rect 13298 8473 13436 8480
rect 13298 8453 13307 8473
rect 13327 8453 13436 8473
rect 13298 8444 13436 8453
rect 13177 8417 13184 8444
rect 13203 8443 13240 8444
rect 13299 8443 13336 8444
rect 13148 8392 13184 8417
rect 12446 8390 12529 8391
rect 12619 8390 12660 8391
rect 12446 8383 12660 8390
rect 12446 8366 12629 8383
rect 12446 8333 12459 8366
rect 12512 8363 12629 8366
rect 12649 8363 12660 8383
rect 12512 8355 12660 8363
rect 12727 8387 13086 8391
rect 12727 8382 13049 8387
rect 12727 8358 12840 8382
rect 12864 8363 13049 8382
rect 13073 8363 13086 8387
rect 12864 8358 13086 8363
rect 12727 8355 13086 8358
rect 13148 8355 13183 8392
rect 13251 8389 13351 8392
rect 13251 8385 13318 8389
rect 13251 8359 13263 8385
rect 13289 8363 13318 8385
rect 13344 8363 13351 8389
rect 13289 8359 13351 8363
rect 13251 8355 13351 8359
rect 12512 8333 12529 8355
rect 12727 8334 12758 8355
rect 13148 8334 13184 8355
rect 12570 8333 12607 8334
rect 12446 8319 12529 8333
rect 12219 8076 12387 8078
rect 11943 8075 12387 8076
rect 11187 8045 12387 8075
rect 12457 8109 12529 8319
rect 12569 8324 12607 8333
rect 12569 8304 12578 8324
rect 12598 8304 12607 8324
rect 12569 8296 12607 8304
rect 12673 8328 12758 8334
rect 12783 8333 12820 8334
rect 12673 8308 12681 8328
rect 12701 8308 12758 8328
rect 12673 8300 12758 8308
rect 12782 8324 12820 8333
rect 12782 8304 12791 8324
rect 12811 8304 12820 8324
rect 12673 8299 12709 8300
rect 12782 8296 12820 8304
rect 12886 8328 12971 8334
rect 12991 8333 13028 8334
rect 12886 8308 12894 8328
rect 12914 8327 12971 8328
rect 12914 8308 12943 8327
rect 12886 8307 12943 8308
rect 12964 8307 12971 8327
rect 12886 8300 12971 8307
rect 12990 8324 13028 8333
rect 12990 8304 12999 8324
rect 13019 8304 13028 8324
rect 12886 8299 12922 8300
rect 12990 8296 13028 8304
rect 13094 8328 13238 8334
rect 13094 8308 13102 8328
rect 13122 8308 13210 8328
rect 13230 8308 13238 8328
rect 13094 8300 13238 8308
rect 13094 8299 13130 8300
rect 13202 8299 13238 8300
rect 13304 8333 13341 8334
rect 13304 8332 13342 8333
rect 13304 8324 13368 8332
rect 13304 8304 13313 8324
rect 13333 8310 13368 8324
rect 13388 8310 13391 8330
rect 13333 8305 13391 8310
rect 13333 8304 13368 8305
rect 12570 8267 12607 8296
rect 12571 8265 12607 8267
rect 12783 8265 12820 8296
rect 12571 8243 12820 8265
rect 12652 8237 12763 8243
rect 12652 8229 12693 8237
rect 12652 8209 12660 8229
rect 12679 8209 12693 8229
rect 12652 8207 12693 8209
rect 12721 8229 12763 8237
rect 12721 8209 12737 8229
rect 12756 8209 12763 8229
rect 12721 8207 12763 8209
rect 12652 8192 12763 8207
rect 12457 8070 12476 8109
rect 12521 8070 12529 8109
rect 12457 8053 12529 8070
rect 12991 8097 13028 8296
rect 13304 8292 13368 8304
rect 12991 8091 13032 8097
rect 13408 8093 13435 8444
rect 13267 8091 13435 8093
rect 12991 8065 13435 8091
rect 11187 7998 11252 8045
rect 11187 7980 11210 7998
rect 11228 7980 11252 7998
rect 12100 8025 12135 8027
rect 12100 8023 12204 8025
rect 12993 8023 13032 8065
rect 13267 8064 13435 8065
rect 12100 8016 13034 8023
rect 12100 8015 12151 8016
rect 12100 7995 12103 8015
rect 12128 7996 12151 8015
rect 12183 7996 13034 8016
rect 12128 7995 13034 7996
rect 12100 7988 13034 7995
rect 12373 7987 13034 7988
rect 11187 7959 11252 7980
rect 11464 7970 11504 7973
rect 11464 7966 12367 7970
rect 11464 7946 12341 7966
rect 12361 7946 12367 7966
rect 11464 7943 12367 7946
rect 11188 7899 11253 7919
rect 11188 7881 11212 7899
rect 11230 7881 11253 7899
rect 11188 7854 11253 7881
rect 11464 7854 11504 7943
rect 11948 7941 12364 7943
rect 11948 7940 12289 7941
rect 11605 7909 11715 7923
rect 11605 7906 11648 7909
rect 11605 7901 11609 7906
rect 11187 7819 11504 7854
rect 11527 7879 11609 7901
rect 11638 7879 11648 7906
rect 11676 7882 11683 7909
rect 11712 7901 11715 7909
rect 11712 7882 11777 7901
rect 11676 7879 11777 7882
rect 11527 7877 11777 7879
rect 10145 7796 10167 7814
rect 10185 7796 10210 7814
rect 10145 7777 10210 7796
rect 9838 7752 9875 7753
rect 9261 7731 9297 7752
rect 9687 7731 9718 7752
rect 9925 7747 9933 7756
rect 9922 7731 9933 7747
rect 9094 7727 9194 7731
rect 9094 7723 9156 7727
rect 9094 7697 9101 7723
rect 9127 7701 9156 7723
rect 9182 7701 9194 7727
rect 9127 7697 9194 7701
rect 9094 7694 9194 7697
rect 9262 7694 9297 7731
rect 9359 7728 9718 7731
rect 9359 7723 9581 7728
rect 9359 7699 9372 7723
rect 9396 7704 9581 7723
rect 9605 7704 9718 7728
rect 9396 7699 9718 7704
rect 9359 7695 9718 7699
rect 9785 7723 9933 7731
rect 9785 7703 9796 7723
rect 9816 7714 9933 7723
rect 9982 7747 9989 7756
rect 9982 7714 9990 7747
rect 11188 7743 11253 7819
rect 11527 7798 11564 7877
rect 11605 7864 11715 7877
rect 11679 7808 11710 7809
rect 11527 7778 11536 7798
rect 11556 7778 11564 7798
rect 11527 7768 11564 7778
rect 11623 7798 11710 7808
rect 11623 7778 11632 7798
rect 11652 7778 11710 7798
rect 11623 7769 11710 7778
rect 11623 7768 11660 7769
rect 9816 7703 9990 7714
rect 9785 7696 9990 7703
rect 9785 7695 9826 7696
rect 9261 7669 9297 7694
rect 9109 7642 9146 7643
rect 9205 7642 9242 7643
rect 9261 7642 9268 7669
rect 8785 7617 8793 7637
rect 8813 7617 8822 7637
rect 8639 7606 8670 7607
rect 8634 7538 8744 7551
rect 8785 7538 8822 7617
rect 9009 7633 9147 7642
rect 9009 7613 9118 7633
rect 9138 7613 9147 7633
rect 9009 7606 9147 7613
rect 9205 7639 9268 7642
rect 9289 7642 9297 7669
rect 9316 7642 9353 7643
rect 9289 7639 9353 7642
rect 9205 7633 9353 7639
rect 9205 7613 9214 7633
rect 9234 7613 9324 7633
rect 9344 7613 9353 7633
rect 9009 7604 9105 7606
rect 9205 7603 9353 7613
rect 9412 7633 9449 7643
rect 9524 7642 9561 7643
rect 9505 7640 9561 7642
rect 9412 7613 9420 7633
rect 9440 7613 9449 7633
rect 9261 7602 9297 7603
rect 8572 7536 8822 7538
rect 8572 7533 8673 7536
rect 8572 7514 8637 7533
rect 8634 7506 8637 7514
rect 8666 7506 8673 7533
rect 8701 7509 8711 7536
rect 8740 7514 8822 7536
rect 8740 7509 8744 7514
rect 8701 7506 8744 7509
rect 8634 7492 8744 7506
rect 8060 7474 8401 7475
rect 7985 7469 8401 7474
rect 9109 7471 9146 7472
rect 9412 7471 9449 7613
rect 9474 7633 9561 7640
rect 9474 7630 9532 7633
rect 9474 7610 9479 7630
rect 9500 7613 9532 7630
rect 9552 7613 9561 7633
rect 9500 7610 9561 7613
rect 9474 7603 9561 7610
rect 9620 7633 9657 7643
rect 9620 7613 9628 7633
rect 9648 7613 9657 7633
rect 9474 7602 9505 7603
rect 9620 7534 9657 7613
rect 9687 7642 9718 7695
rect 9922 7693 9990 7696
rect 9922 7651 9934 7693
rect 9983 7651 9990 7693
rect 9737 7642 9774 7643
rect 9687 7633 9774 7642
rect 9687 7613 9745 7633
rect 9765 7613 9774 7633
rect 9687 7603 9774 7613
rect 9833 7633 9870 7643
rect 9922 7638 9990 7651
rect 10145 7715 10210 7732
rect 10145 7697 10169 7715
rect 10187 7697 10210 7715
rect 11188 7725 11210 7743
rect 11228 7725 11253 7743
rect 11188 7704 11253 7725
rect 11401 7723 11466 7732
rect 9833 7613 9841 7633
rect 9861 7613 9870 7633
rect 9687 7602 9718 7603
rect 9682 7534 9792 7547
rect 9833 7534 9870 7613
rect 10145 7558 10210 7697
rect 11401 7686 11411 7723
rect 11451 7715 11466 7723
rect 11679 7716 11710 7769
rect 11740 7798 11777 7877
rect 11892 7808 11923 7809
rect 11740 7778 11749 7798
rect 11769 7778 11777 7798
rect 11740 7768 11777 7778
rect 11836 7801 11923 7808
rect 11836 7798 11897 7801
rect 11836 7778 11845 7798
rect 11865 7781 11897 7798
rect 11918 7781 11923 7801
rect 11865 7778 11923 7781
rect 11836 7771 11923 7778
rect 11948 7798 11985 7940
rect 12251 7939 12288 7940
rect 12100 7808 12136 7809
rect 11948 7778 11957 7798
rect 11977 7778 11985 7798
rect 11836 7769 11892 7771
rect 11836 7768 11873 7769
rect 11948 7768 11985 7778
rect 12044 7798 12192 7808
rect 12292 7805 12388 7807
rect 12044 7778 12053 7798
rect 12073 7778 12163 7798
rect 12183 7778 12192 7798
rect 12044 7772 12192 7778
rect 12044 7769 12108 7772
rect 12044 7768 12081 7769
rect 12100 7742 12108 7769
rect 12129 7769 12192 7772
rect 12250 7798 12388 7805
rect 12250 7778 12259 7798
rect 12279 7778 12388 7798
rect 12250 7769 12388 7778
rect 12129 7742 12136 7769
rect 12155 7768 12192 7769
rect 12251 7768 12288 7769
rect 12100 7717 12136 7742
rect 11571 7715 11612 7716
rect 11451 7708 11612 7715
rect 11451 7688 11581 7708
rect 11601 7688 11612 7708
rect 11451 7686 11612 7688
rect 11401 7680 11612 7686
rect 11679 7712 12038 7716
rect 11679 7707 12001 7712
rect 11679 7683 11792 7707
rect 11816 7688 12001 7707
rect 12025 7688 12038 7712
rect 11816 7683 12038 7688
rect 11679 7680 12038 7683
rect 12100 7680 12135 7717
rect 12203 7714 12303 7717
rect 12203 7710 12270 7714
rect 12203 7684 12215 7710
rect 12241 7688 12270 7710
rect 12296 7688 12303 7714
rect 12241 7684 12303 7688
rect 12203 7680 12303 7684
rect 11401 7667 11468 7680
rect 10145 7552 10167 7558
rect 9620 7532 9870 7534
rect 9620 7529 9721 7532
rect 9620 7510 9685 7529
rect 9682 7502 9685 7510
rect 9714 7502 9721 7529
rect 9749 7505 9759 7532
rect 9788 7510 9870 7532
rect 9899 7540 10167 7552
rect 10185 7540 10210 7558
rect 9899 7517 10210 7540
rect 11193 7644 11249 7664
rect 11193 7626 11212 7644
rect 11230 7626 11249 7644
rect 9899 7516 9954 7517
rect 9788 7505 9792 7510
rect 9749 7502 9792 7505
rect 9682 7488 9792 7502
rect 9108 7470 9449 7471
rect 7985 7449 7988 7469
rect 8008 7449 8401 7469
rect 9033 7469 9449 7470
rect 9899 7469 9942 7516
rect 11193 7513 11249 7626
rect 11401 7646 11415 7667
rect 11451 7646 11468 7667
rect 11679 7659 11710 7680
rect 12100 7659 12136 7680
rect 11522 7658 11559 7659
rect 11401 7639 11468 7646
rect 11521 7649 11559 7658
rect 9033 7465 9942 7469
rect 6908 7414 7619 7416
rect 8158 7414 8247 7417
rect 6908 7405 8247 7414
rect 6908 7367 8170 7405
rect 8195 7370 8214 7405
rect 8239 7370 8247 7405
rect 8352 7416 8397 7449
rect 9033 7445 9036 7465
rect 9056 7445 9942 7465
rect 9410 7440 9942 7445
rect 10150 7459 10209 7481
rect 10150 7441 10169 7459
rect 10187 7441 10209 7459
rect 9198 7416 9297 7418
rect 8352 7406 9297 7416
rect 8352 7380 9220 7406
rect 8353 7379 9220 7380
rect 8195 7367 8247 7370
rect 6908 7359 8247 7367
rect 9198 7368 9220 7379
rect 9245 7371 9264 7406
rect 9289 7371 9297 7406
rect 9245 7368 9297 7371
rect 9198 7360 9297 7368
rect 10150 7367 10209 7441
rect 11193 7406 11248 7513
rect 11401 7487 11466 7639
rect 11521 7629 11530 7649
rect 11550 7629 11559 7649
rect 11521 7621 11559 7629
rect 11625 7653 11710 7659
rect 11735 7658 11772 7659
rect 11625 7633 11633 7653
rect 11653 7633 11710 7653
rect 11625 7625 11710 7633
rect 11734 7649 11772 7658
rect 11734 7629 11743 7649
rect 11763 7629 11772 7649
rect 11625 7624 11661 7625
rect 11734 7621 11772 7629
rect 11838 7653 11923 7659
rect 11943 7658 11980 7659
rect 11838 7633 11846 7653
rect 11866 7652 11923 7653
rect 11866 7633 11895 7652
rect 11838 7632 11895 7633
rect 11916 7632 11923 7652
rect 11838 7625 11923 7632
rect 11942 7649 11980 7658
rect 11942 7629 11951 7649
rect 11971 7629 11980 7649
rect 11838 7624 11874 7625
rect 11942 7621 11980 7629
rect 12046 7653 12190 7659
rect 12046 7633 12054 7653
rect 12074 7633 12162 7653
rect 12182 7633 12190 7653
rect 12046 7625 12190 7633
rect 12046 7624 12082 7625
rect 12154 7624 12190 7625
rect 12256 7658 12293 7659
rect 12256 7657 12294 7658
rect 12256 7649 12320 7657
rect 12256 7629 12265 7649
rect 12285 7635 12320 7649
rect 12340 7635 12343 7655
rect 12285 7630 12343 7635
rect 12285 7629 12320 7630
rect 11522 7592 11559 7621
rect 11523 7590 11559 7592
rect 11735 7590 11772 7621
rect 11523 7568 11772 7590
rect 11604 7562 11715 7568
rect 11604 7554 11645 7562
rect 11604 7534 11612 7554
rect 11631 7534 11645 7554
rect 11604 7532 11645 7534
rect 11673 7554 11715 7562
rect 11673 7534 11689 7554
rect 11708 7534 11715 7554
rect 11673 7532 11715 7534
rect 11604 7517 11715 7532
rect 11943 7522 11980 7621
rect 12256 7617 12320 7629
rect 11606 7514 11710 7517
rect 11394 7477 11515 7487
rect 11394 7475 11463 7477
rect 11394 7434 11407 7475
rect 11444 7436 11463 7475
rect 11500 7436 11515 7477
rect 11444 7434 11515 7436
rect 11394 7416 11515 7434
rect 9224 7359 9296 7360
rect 6908 7358 8246 7359
rect 6908 7356 7619 7358
rect 7768 7317 7832 7321
rect 10143 7319 10209 7367
rect 11186 7372 11251 7406
rect 11606 7372 11710 7374
rect 11941 7372 11982 7522
rect 12360 7514 12387 7769
rect 12449 7759 12529 7770
rect 12449 7733 12466 7759
rect 12506 7733 12529 7759
rect 12449 7706 12529 7733
rect 12449 7680 12470 7706
rect 12510 7680 12529 7706
rect 12449 7661 12529 7680
rect 12449 7635 12473 7661
rect 12513 7635 12529 7661
rect 12449 7584 12529 7635
rect 11186 7369 11982 7372
rect 12361 7383 12387 7514
rect 12451 7384 12521 7584
rect 12361 7369 12389 7383
rect 11186 7334 12389 7369
rect 12450 7362 12522 7384
rect 7768 7308 7842 7317
rect 6283 6825 6397 6829
rect 5488 6821 5588 6825
rect 5488 6817 5550 6821
rect 5488 6791 5495 6817
rect 5521 6795 5550 6817
rect 5576 6795 5588 6821
rect 5521 6791 5588 6795
rect 5488 6788 5588 6791
rect 5656 6788 5691 6825
rect 5753 6822 6112 6825
rect 5753 6817 5975 6822
rect 5753 6793 5766 6817
rect 5790 6798 5975 6817
rect 5999 6798 6112 6822
rect 5790 6793 6112 6798
rect 5753 6789 6112 6793
rect 6179 6822 6397 6825
rect 6179 6821 6362 6822
rect 6179 6817 6305 6821
rect 6179 6797 6190 6817
rect 6210 6797 6305 6817
rect 6329 6798 6362 6821
rect 6386 6798 6397 6822
rect 6329 6797 6397 6798
rect 6179 6790 6397 6797
rect 6179 6789 6220 6790
rect 5655 6763 5691 6788
rect 5503 6736 5540 6737
rect 5599 6736 5636 6737
rect 5655 6736 5662 6763
rect 5403 6727 5541 6736
rect 5403 6707 5512 6727
rect 5532 6707 5541 6727
rect 5403 6700 5541 6707
rect 5599 6733 5662 6736
rect 5683 6736 5691 6763
rect 5710 6736 5747 6737
rect 5683 6733 5747 6736
rect 5599 6727 5747 6733
rect 5599 6707 5608 6727
rect 5628 6707 5718 6727
rect 5738 6707 5747 6727
rect 5403 6698 5499 6700
rect 5599 6697 5747 6707
rect 5806 6727 5843 6737
rect 5918 6736 5955 6737
rect 5899 6734 5955 6736
rect 5806 6707 5814 6727
rect 5834 6707 5843 6727
rect 5655 6696 5691 6697
rect 5503 6565 5540 6566
rect 5806 6565 5843 6707
rect 5868 6727 5955 6734
rect 5868 6724 5926 6727
rect 5868 6704 5873 6724
rect 5894 6707 5926 6724
rect 5946 6707 5955 6727
rect 5894 6704 5955 6707
rect 5868 6697 5955 6704
rect 6014 6727 6051 6737
rect 6014 6707 6022 6727
rect 6042 6707 6051 6727
rect 5868 6696 5899 6697
rect 6014 6628 6051 6707
rect 6081 6736 6112 6789
rect 6283 6787 6397 6790
rect 6326 6755 6397 6787
rect 7572 7266 7656 7291
rect 7572 7238 7587 7266
rect 7631 7238 7656 7266
rect 7572 7209 7656 7238
rect 7768 7260 7782 7308
rect 7819 7260 7842 7308
rect 7768 7232 7842 7260
rect 7572 7181 7584 7209
rect 7628 7181 7656 7209
rect 7572 7160 7656 7181
rect 6131 6736 6168 6737
rect 6081 6727 6168 6736
rect 6081 6707 6139 6727
rect 6159 6707 6168 6727
rect 6081 6697 6168 6707
rect 6227 6727 6264 6737
rect 6227 6707 6235 6727
rect 6255 6707 6264 6727
rect 6081 6696 6112 6697
rect 6076 6628 6186 6641
rect 6227 6628 6264 6707
rect 6014 6626 6264 6628
rect 6014 6623 6115 6626
rect 6014 6604 6079 6623
rect 6076 6596 6079 6604
rect 6108 6596 6115 6623
rect 6143 6599 6153 6626
rect 6182 6604 6264 6626
rect 6182 6599 6186 6604
rect 6143 6596 6186 6599
rect 6076 6582 6186 6596
rect 5502 6564 5843 6565
rect 5427 6561 5843 6564
rect 5427 6559 5850 6561
rect 5427 6539 5430 6559
rect 5450 6539 5850 6559
rect 4618 4198 5258 4286
rect 4618 3847 4702 4198
rect 5184 4167 5228 4173
rect 5184 4141 5192 4167
rect 5217 4141 5228 4167
rect 5184 4092 5228 4141
rect 5184 4072 5581 4092
rect 5601 4072 5604 4092
rect 5184 4067 5604 4072
rect 5184 4066 5529 4067
rect 5184 4062 5228 4066
rect 5491 4065 5528 4066
rect 4845 4035 4955 4049
rect 4845 4032 4888 4035
rect 4845 4027 4849 4032
rect 4767 4005 4849 4027
rect 4878 4005 4888 4032
rect 4916 4008 4923 4035
rect 4952 4027 4955 4035
rect 4952 4008 5017 4027
rect 4916 4005 5017 4008
rect 4767 4003 5017 4005
rect 4767 3924 4804 4003
rect 4845 3990 4955 4003
rect 4919 3934 4950 3935
rect 4767 3904 4776 3924
rect 4796 3904 4804 3924
rect 4767 3894 4804 3904
rect 4863 3924 4950 3934
rect 4863 3904 4872 3924
rect 4892 3904 4950 3924
rect 4863 3895 4950 3904
rect 4863 3894 4900 3895
rect 4618 3841 4727 3847
rect 4919 3842 4950 3895
rect 4980 3924 5017 4003
rect 5132 3934 5163 3935
rect 4980 3904 4989 3924
rect 5009 3904 5017 3924
rect 4980 3894 5017 3904
rect 5076 3927 5163 3934
rect 5076 3924 5137 3927
rect 5076 3904 5085 3924
rect 5105 3907 5137 3924
rect 5158 3907 5163 3927
rect 5105 3904 5163 3907
rect 5076 3897 5163 3904
rect 5188 3924 5225 4062
rect 5340 3934 5376 3935
rect 5188 3904 5197 3924
rect 5217 3904 5225 3924
rect 5076 3895 5132 3897
rect 5076 3894 5113 3895
rect 5188 3894 5225 3904
rect 5284 3924 5432 3934
rect 5532 3931 5628 3933
rect 5284 3904 5293 3924
rect 5313 3904 5403 3924
rect 5423 3904 5432 3924
rect 5284 3898 5432 3904
rect 5284 3895 5348 3898
rect 5284 3894 5321 3895
rect 5340 3868 5348 3895
rect 5369 3895 5432 3898
rect 5490 3924 5628 3931
rect 5490 3904 5499 3924
rect 5519 3904 5628 3924
rect 5490 3895 5628 3904
rect 5369 3868 5376 3895
rect 5395 3894 5432 3895
rect 5491 3894 5528 3895
rect 5340 3843 5376 3868
rect 4811 3841 4852 3842
rect 4618 3834 4852 3841
rect 4618 3814 4821 3834
rect 4841 3814 4852 3834
rect 4618 3806 4852 3814
rect 4919 3838 5278 3842
rect 4919 3833 5241 3838
rect 4919 3809 5032 3833
rect 5056 3814 5241 3833
rect 5265 3814 5278 3838
rect 5056 3809 5278 3814
rect 4919 3806 5278 3809
rect 5340 3806 5375 3843
rect 5443 3840 5543 3843
rect 5443 3836 5510 3840
rect 5443 3810 5455 3836
rect 5481 3814 5510 3836
rect 5536 3814 5543 3840
rect 5481 3810 5543 3814
rect 5443 3806 5543 3810
rect 4618 3788 4727 3806
rect 4919 3785 4950 3806
rect 5340 3785 5376 3806
rect 4762 3784 4799 3785
rect 4761 3775 4799 3784
rect 4761 3755 4770 3775
rect 4790 3755 4799 3775
rect 4761 3747 4799 3755
rect 4865 3779 4950 3785
rect 4975 3784 5012 3785
rect 4865 3759 4873 3779
rect 4893 3759 4950 3779
rect 4865 3751 4950 3759
rect 4974 3775 5012 3784
rect 4974 3755 4983 3775
rect 5003 3755 5012 3775
rect 4865 3750 4901 3751
rect 4974 3747 5012 3755
rect 5078 3779 5163 3785
rect 5183 3784 5220 3785
rect 5078 3759 5086 3779
rect 5106 3778 5163 3779
rect 5106 3759 5135 3778
rect 5078 3758 5135 3759
rect 5156 3758 5163 3778
rect 5078 3751 5163 3758
rect 5182 3775 5220 3784
rect 5182 3755 5191 3775
rect 5211 3755 5220 3775
rect 5078 3750 5114 3751
rect 5182 3747 5220 3755
rect 5286 3780 5430 3785
rect 5286 3779 5339 3780
rect 5286 3759 5294 3779
rect 5314 3760 5339 3779
rect 5372 3779 5430 3780
rect 5372 3760 5402 3779
rect 5314 3759 5402 3760
rect 5422 3759 5430 3779
rect 5286 3751 5430 3759
rect 5286 3750 5322 3751
rect 5394 3750 5430 3751
rect 5496 3784 5533 3785
rect 5496 3783 5534 3784
rect 5496 3775 5560 3783
rect 5496 3755 5505 3775
rect 5525 3761 5560 3775
rect 5580 3761 5583 3781
rect 5525 3756 5583 3761
rect 5525 3755 5560 3756
rect 4762 3718 4799 3747
rect 4763 3716 4799 3718
rect 4975 3716 5012 3747
rect 4763 3694 5012 3716
rect 4844 3688 4955 3694
rect 4844 3680 4885 3688
rect 4844 3660 4852 3680
rect 4871 3660 4885 3680
rect 4844 3658 4885 3660
rect 4913 3680 4955 3688
rect 4913 3660 4929 3680
rect 4948 3660 4955 3680
rect 4913 3658 4955 3660
rect 4844 3643 4955 3658
rect 5183 3626 5220 3747
rect 5496 3743 5560 3755
rect 5600 3632 5627 3895
rect 5654 3641 5690 3648
rect 5654 3632 5660 3641
rect 5578 3628 5660 3632
rect 5459 3626 5660 3628
rect 5183 3603 5660 3626
rect 5683 3603 5690 3641
rect 5183 3600 5690 3603
rect 5459 3599 5627 3600
rect 5654 3597 5690 3600
rect 5772 3499 5850 6539
rect 6906 5792 6965 5802
rect 6906 5764 6919 5792
rect 6947 5764 6965 5792
rect 6906 5715 6965 5764
rect 6512 5580 6680 5581
rect 6916 5580 6963 5715
rect 6512 5554 6963 5580
rect 6512 5552 6680 5554
rect 6512 5285 6539 5552
rect 6916 5548 6963 5554
rect 6579 5425 6643 5437
rect 6919 5433 6956 5548
rect 7184 5522 7295 5537
rect 7184 5520 7226 5522
rect 7184 5500 7191 5520
rect 7210 5500 7226 5520
rect 7184 5492 7226 5500
rect 7254 5520 7295 5522
rect 7254 5500 7268 5520
rect 7287 5500 7295 5520
rect 7254 5492 7295 5500
rect 7184 5486 7295 5492
rect 7127 5464 7376 5486
rect 7127 5433 7164 5464
rect 7340 5462 7376 5464
rect 7340 5433 7377 5462
rect 6579 5424 6614 5425
rect 6556 5419 6614 5424
rect 6556 5399 6559 5419
rect 6579 5405 6614 5419
rect 6634 5405 6643 5425
rect 6579 5397 6643 5405
rect 6605 5396 6643 5397
rect 6606 5395 6643 5396
rect 6709 5429 6745 5430
rect 6817 5429 6853 5430
rect 6709 5421 6853 5429
rect 6709 5401 6717 5421
rect 6737 5401 6825 5421
rect 6845 5401 6853 5421
rect 6709 5395 6853 5401
rect 6919 5425 6957 5433
rect 7025 5429 7061 5430
rect 6919 5405 6928 5425
rect 6948 5405 6957 5425
rect 6919 5396 6957 5405
rect 6976 5422 7061 5429
rect 6976 5402 6983 5422
rect 7004 5421 7061 5422
rect 7004 5402 7033 5421
rect 6976 5401 7033 5402
rect 7053 5401 7061 5421
rect 6919 5395 6956 5396
rect 6976 5395 7061 5401
rect 7127 5425 7165 5433
rect 7238 5429 7274 5430
rect 7127 5405 7136 5425
rect 7156 5405 7165 5425
rect 7127 5396 7165 5405
rect 7189 5421 7274 5429
rect 7189 5401 7246 5421
rect 7266 5401 7274 5421
rect 7127 5395 7164 5396
rect 7189 5395 7274 5401
rect 7340 5425 7378 5433
rect 7340 5405 7349 5425
rect 7369 5405 7378 5425
rect 7340 5396 7378 5405
rect 7340 5395 7377 5396
rect 6763 5374 6799 5395
rect 7189 5374 7220 5395
rect 7400 5380 7457 5388
rect 7400 5374 7408 5380
rect 6596 5370 6696 5374
rect 6596 5366 6658 5370
rect 6596 5340 6603 5366
rect 6629 5344 6658 5366
rect 6684 5344 6696 5370
rect 6629 5340 6696 5344
rect 6596 5337 6696 5340
rect 6764 5337 6799 5374
rect 6861 5371 7220 5374
rect 6861 5366 7083 5371
rect 6861 5342 6874 5366
rect 6898 5347 7083 5366
rect 7107 5347 7220 5371
rect 6898 5342 7220 5347
rect 6861 5338 7220 5342
rect 7287 5366 7408 5374
rect 7287 5346 7298 5366
rect 7318 5357 7408 5366
rect 7434 5357 7457 5380
rect 7318 5346 7457 5357
rect 7287 5344 7457 5346
rect 7287 5339 7408 5344
rect 7287 5338 7328 5339
rect 6763 5312 6799 5337
rect 6611 5285 6648 5286
rect 6707 5285 6744 5286
rect 6763 5285 6770 5312
rect 6511 5276 6649 5285
rect 6511 5256 6620 5276
rect 6640 5256 6649 5276
rect 6511 5249 6649 5256
rect 6707 5282 6770 5285
rect 6791 5285 6799 5312
rect 6818 5285 6855 5286
rect 6791 5282 6855 5285
rect 6707 5276 6855 5282
rect 6707 5256 6716 5276
rect 6736 5256 6826 5276
rect 6846 5256 6855 5276
rect 6511 5247 6607 5249
rect 6707 5246 6855 5256
rect 6914 5276 6951 5286
rect 7026 5285 7063 5286
rect 7007 5283 7063 5285
rect 6914 5256 6922 5276
rect 6942 5256 6951 5276
rect 6763 5245 6799 5246
rect 6611 5114 6648 5115
rect 6914 5114 6951 5256
rect 6976 5276 7063 5283
rect 6976 5273 7034 5276
rect 6976 5253 6981 5273
rect 7002 5256 7034 5273
rect 7054 5256 7063 5276
rect 7002 5253 7063 5256
rect 6976 5246 7063 5253
rect 7122 5276 7159 5286
rect 7122 5256 7130 5276
rect 7150 5256 7159 5276
rect 6976 5245 7007 5246
rect 7122 5177 7159 5256
rect 7189 5285 7220 5338
rect 7239 5285 7276 5286
rect 7189 5276 7276 5285
rect 7189 5256 7247 5276
rect 7267 5256 7276 5276
rect 7189 5246 7276 5256
rect 7335 5276 7372 5286
rect 7335 5256 7343 5276
rect 7363 5256 7372 5276
rect 7189 5245 7220 5246
rect 7184 5177 7294 5190
rect 7335 5177 7372 5256
rect 7122 5175 7372 5177
rect 7122 5172 7223 5175
rect 7122 5153 7187 5172
rect 7184 5145 7187 5153
rect 7216 5145 7223 5172
rect 7251 5148 7261 5175
rect 7290 5153 7372 5175
rect 7290 5148 7294 5153
rect 7251 5145 7294 5148
rect 7184 5131 7294 5145
rect 6610 5113 6951 5114
rect 6535 5108 6951 5113
rect 6535 5088 6538 5108
rect 6558 5088 6952 5108
rect 6761 5055 6798 5065
rect 6761 5018 6770 5055
rect 6787 5018 6798 5055
rect 6761 4997 6798 5018
rect 6470 4058 6638 4059
rect 6767 4058 6796 4997
rect 6909 4383 6952 5088
rect 6910 4375 6952 4383
rect 6910 4364 6955 4375
rect 6910 4326 6920 4364
rect 6945 4326 6955 4364
rect 6910 4317 6955 4326
rect 6470 4032 6914 4058
rect 6470 4030 6638 4032
rect 6470 3763 6497 4030
rect 6767 4028 6796 4032
rect 6537 3903 6601 3915
rect 6877 3911 6914 4032
rect 7142 4000 7253 4015
rect 7142 3998 7184 4000
rect 7142 3978 7149 3998
rect 7168 3978 7184 3998
rect 7142 3970 7184 3978
rect 7212 3998 7253 4000
rect 7212 3978 7226 3998
rect 7245 3978 7253 3998
rect 7212 3970 7253 3978
rect 7142 3964 7253 3970
rect 7085 3942 7334 3964
rect 7085 3911 7122 3942
rect 7298 3940 7334 3942
rect 7298 3911 7335 3940
rect 6537 3902 6572 3903
rect 6514 3897 6572 3902
rect 6514 3877 6517 3897
rect 6537 3883 6572 3897
rect 6592 3883 6601 3903
rect 6537 3875 6601 3883
rect 6563 3874 6601 3875
rect 6564 3873 6601 3874
rect 6667 3907 6703 3908
rect 6775 3907 6811 3908
rect 6667 3899 6811 3907
rect 6667 3879 6675 3899
rect 6695 3879 6783 3899
rect 6803 3879 6811 3899
rect 6667 3873 6811 3879
rect 6877 3903 6915 3911
rect 6983 3907 7019 3908
rect 6877 3883 6886 3903
rect 6906 3883 6915 3903
rect 6877 3874 6915 3883
rect 6934 3900 7019 3907
rect 6934 3880 6941 3900
rect 6962 3899 7019 3900
rect 6962 3880 6991 3899
rect 6934 3879 6991 3880
rect 7011 3879 7019 3899
rect 6877 3873 6914 3874
rect 6934 3873 7019 3879
rect 7085 3903 7123 3911
rect 7196 3907 7232 3908
rect 7085 3883 7094 3903
rect 7114 3883 7123 3903
rect 7085 3874 7123 3883
rect 7147 3899 7232 3907
rect 7147 3879 7204 3899
rect 7224 3879 7232 3899
rect 7085 3873 7122 3874
rect 7147 3873 7232 3879
rect 7298 3903 7336 3911
rect 7298 3883 7307 3903
rect 7327 3883 7336 3903
rect 7298 3874 7336 3883
rect 7298 3873 7335 3874
rect 6721 3852 6757 3873
rect 7147 3852 7178 3873
rect 7572 3856 7664 7160
rect 7770 5393 7842 7232
rect 8872 7182 8944 7199
rect 8872 7134 8884 7182
rect 8930 7134 8944 7182
rect 9412 7162 9453 7164
rect 9684 7162 9788 7164
rect 10143 7162 10208 7319
rect 11186 7177 11251 7334
rect 11606 7332 11710 7334
rect 11941 7332 11982 7334
rect 12450 7314 12464 7362
rect 12510 7314 12522 7362
rect 12450 7297 12522 7314
rect 13552 7264 13624 9103
rect 13730 7336 13822 10640
rect 14216 10623 14247 10644
rect 14637 10623 14673 10644
rect 14059 10622 14096 10623
rect 14058 10613 14096 10622
rect 14058 10593 14067 10613
rect 14087 10593 14096 10613
rect 14058 10585 14096 10593
rect 14162 10617 14247 10623
rect 14272 10622 14309 10623
rect 14162 10597 14170 10617
rect 14190 10597 14247 10617
rect 14162 10589 14247 10597
rect 14271 10613 14309 10622
rect 14271 10593 14280 10613
rect 14300 10593 14309 10613
rect 14162 10588 14198 10589
rect 14271 10585 14309 10593
rect 14375 10617 14460 10623
rect 14480 10622 14517 10623
rect 14375 10597 14383 10617
rect 14403 10616 14460 10617
rect 14403 10597 14432 10616
rect 14375 10596 14432 10597
rect 14453 10596 14460 10616
rect 14375 10589 14460 10596
rect 14479 10613 14517 10622
rect 14479 10593 14488 10613
rect 14508 10593 14517 10613
rect 14375 10588 14411 10589
rect 14479 10585 14517 10593
rect 14583 10617 14727 10623
rect 14583 10597 14591 10617
rect 14611 10597 14699 10617
rect 14719 10597 14727 10617
rect 14583 10589 14727 10597
rect 14583 10588 14619 10589
rect 14691 10588 14727 10589
rect 14793 10622 14830 10623
rect 14793 10621 14831 10622
rect 14793 10613 14857 10621
rect 14793 10593 14802 10613
rect 14822 10599 14857 10613
rect 14877 10599 14880 10619
rect 14822 10594 14880 10599
rect 14822 10593 14857 10594
rect 14059 10556 14096 10585
rect 14060 10554 14096 10556
rect 14272 10554 14309 10585
rect 14060 10532 14309 10554
rect 14141 10526 14252 10532
rect 14141 10518 14182 10526
rect 14141 10498 14149 10518
rect 14168 10498 14182 10518
rect 14141 10496 14182 10498
rect 14210 10518 14252 10526
rect 14210 10498 14226 10518
rect 14245 10498 14252 10518
rect 14210 10496 14252 10498
rect 14141 10481 14252 10496
rect 14480 10464 14517 10585
rect 14793 10581 14857 10593
rect 14598 10464 14627 10468
rect 14897 10466 14924 10733
rect 14756 10464 14924 10466
rect 14480 10438 14924 10464
rect 14439 10170 14484 10179
rect 14439 10132 14449 10170
rect 14474 10132 14484 10170
rect 14439 10121 14484 10132
rect 14442 10113 14484 10121
rect 14442 9408 14485 10113
rect 14598 9499 14627 10438
rect 14756 10437 14924 10438
rect 14596 9478 14633 9499
rect 14596 9441 14607 9478
rect 14624 9441 14633 9478
rect 14596 9431 14633 9441
rect 14442 9388 14836 9408
rect 14856 9388 14859 9408
rect 14443 9383 14859 9388
rect 14443 9382 14784 9383
rect 14100 9351 14210 9365
rect 14100 9348 14143 9351
rect 14100 9343 14104 9348
rect 14022 9321 14104 9343
rect 14133 9321 14143 9348
rect 14171 9324 14178 9351
rect 14207 9343 14210 9351
rect 14207 9324 14272 9343
rect 14171 9321 14272 9324
rect 14022 9319 14272 9321
rect 14022 9240 14059 9319
rect 14100 9306 14210 9319
rect 14174 9250 14205 9251
rect 14022 9220 14031 9240
rect 14051 9220 14059 9240
rect 14022 9210 14059 9220
rect 14118 9240 14205 9250
rect 14118 9220 14127 9240
rect 14147 9220 14205 9240
rect 14118 9211 14205 9220
rect 14118 9210 14155 9211
rect 14174 9158 14205 9211
rect 14235 9240 14272 9319
rect 14387 9250 14418 9251
rect 14235 9220 14244 9240
rect 14264 9220 14272 9240
rect 14235 9210 14272 9220
rect 14331 9243 14418 9250
rect 14331 9240 14392 9243
rect 14331 9220 14340 9240
rect 14360 9223 14392 9240
rect 14413 9223 14418 9243
rect 14360 9220 14418 9223
rect 14331 9213 14418 9220
rect 14443 9240 14480 9382
rect 14746 9381 14783 9382
rect 14595 9250 14631 9251
rect 14443 9220 14452 9240
rect 14472 9220 14480 9240
rect 14331 9211 14387 9213
rect 14331 9210 14368 9211
rect 14443 9210 14480 9220
rect 14539 9240 14687 9250
rect 14787 9247 14883 9249
rect 14539 9220 14548 9240
rect 14568 9220 14658 9240
rect 14678 9220 14687 9240
rect 14539 9214 14687 9220
rect 14539 9211 14603 9214
rect 14539 9210 14576 9211
rect 14595 9184 14603 9211
rect 14624 9211 14687 9214
rect 14745 9240 14883 9247
rect 14745 9220 14754 9240
rect 14774 9220 14883 9240
rect 14745 9211 14883 9220
rect 14624 9184 14631 9211
rect 14650 9210 14687 9211
rect 14746 9210 14783 9211
rect 14595 9159 14631 9184
rect 14066 9157 14107 9158
rect 13986 9152 14107 9157
rect 13937 9150 14107 9152
rect 13937 9139 14076 9150
rect 13937 9116 13960 9139
rect 13986 9130 14076 9139
rect 14096 9130 14107 9150
rect 13986 9122 14107 9130
rect 14174 9154 14533 9158
rect 14174 9149 14496 9154
rect 14174 9125 14287 9149
rect 14311 9130 14496 9149
rect 14520 9130 14533 9154
rect 14311 9125 14533 9130
rect 14174 9122 14533 9125
rect 14595 9122 14630 9159
rect 14698 9156 14798 9159
rect 14698 9152 14765 9156
rect 14698 9126 14710 9152
rect 14736 9130 14765 9152
rect 14791 9130 14798 9156
rect 14736 9126 14798 9130
rect 14698 9122 14798 9126
rect 13986 9116 13994 9122
rect 13937 9108 13994 9116
rect 14174 9101 14205 9122
rect 14595 9101 14631 9122
rect 14017 9100 14054 9101
rect 14016 9091 14054 9100
rect 14016 9071 14025 9091
rect 14045 9071 14054 9091
rect 14016 9063 14054 9071
rect 14120 9095 14205 9101
rect 14230 9100 14267 9101
rect 14120 9075 14128 9095
rect 14148 9075 14205 9095
rect 14120 9067 14205 9075
rect 14229 9091 14267 9100
rect 14229 9071 14238 9091
rect 14258 9071 14267 9091
rect 14120 9066 14156 9067
rect 14229 9063 14267 9071
rect 14333 9095 14418 9101
rect 14438 9100 14475 9101
rect 14333 9075 14341 9095
rect 14361 9094 14418 9095
rect 14361 9075 14390 9094
rect 14333 9074 14390 9075
rect 14411 9074 14418 9094
rect 14333 9067 14418 9074
rect 14437 9091 14475 9100
rect 14437 9071 14446 9091
rect 14466 9071 14475 9091
rect 14333 9066 14369 9067
rect 14437 9063 14475 9071
rect 14541 9095 14685 9101
rect 14541 9075 14549 9095
rect 14569 9075 14657 9095
rect 14677 9075 14685 9095
rect 14541 9067 14685 9075
rect 14541 9066 14577 9067
rect 14649 9066 14685 9067
rect 14751 9100 14788 9101
rect 14751 9099 14789 9100
rect 14751 9091 14815 9099
rect 14751 9071 14760 9091
rect 14780 9077 14815 9091
rect 14835 9077 14838 9097
rect 14780 9072 14838 9077
rect 14780 9071 14815 9072
rect 14017 9034 14054 9063
rect 14018 9032 14054 9034
rect 14230 9032 14267 9063
rect 14018 9010 14267 9032
rect 14099 9004 14210 9010
rect 14099 8996 14140 9004
rect 14099 8976 14107 8996
rect 14126 8976 14140 8996
rect 14099 8974 14140 8976
rect 14168 8996 14210 9004
rect 14168 8976 14184 8996
rect 14203 8976 14210 8996
rect 14168 8974 14210 8976
rect 14099 8959 14210 8974
rect 14438 8948 14475 9063
rect 14751 9059 14815 9071
rect 14431 8942 14478 8948
rect 14855 8944 14882 9211
rect 14714 8942 14882 8944
rect 14431 8916 14882 8942
rect 14431 8781 14478 8916
rect 14714 8915 14882 8916
rect 14429 8732 14488 8781
rect 14429 8704 14447 8732
rect 14475 8704 14488 8732
rect 14429 8694 14488 8704
rect 15544 7957 15622 10997
rect 15544 7937 15944 7957
rect 15964 7937 15967 7957
rect 15544 7935 15967 7937
rect 15551 7932 15967 7935
rect 15551 7931 15892 7932
rect 15208 7900 15318 7914
rect 15208 7897 15251 7900
rect 15208 7892 15212 7897
rect 15130 7870 15212 7892
rect 15241 7870 15251 7897
rect 15279 7873 15286 7900
rect 15315 7892 15318 7900
rect 15315 7873 15380 7892
rect 15279 7870 15380 7873
rect 15130 7868 15380 7870
rect 15130 7789 15167 7868
rect 15208 7855 15318 7868
rect 15282 7799 15313 7800
rect 15130 7769 15139 7789
rect 15159 7769 15167 7789
rect 15130 7759 15167 7769
rect 15226 7789 15313 7799
rect 15226 7769 15235 7789
rect 15255 7769 15313 7789
rect 15226 7760 15313 7769
rect 15226 7759 15263 7760
rect 15000 7706 15111 7709
rect 15282 7707 15313 7760
rect 15343 7789 15380 7868
rect 15495 7799 15526 7800
rect 15343 7769 15352 7789
rect 15372 7769 15380 7789
rect 15343 7759 15380 7769
rect 15439 7792 15526 7799
rect 15439 7789 15500 7792
rect 15439 7769 15448 7789
rect 15468 7772 15500 7789
rect 15521 7772 15526 7792
rect 15468 7769 15526 7772
rect 15439 7762 15526 7769
rect 15551 7789 15588 7931
rect 15854 7930 15891 7931
rect 15703 7799 15739 7800
rect 15551 7769 15560 7789
rect 15580 7769 15588 7789
rect 15439 7760 15495 7762
rect 15439 7759 15476 7760
rect 15551 7759 15588 7769
rect 15647 7789 15795 7799
rect 15895 7796 15991 7798
rect 15647 7769 15656 7789
rect 15676 7769 15766 7789
rect 15786 7769 15795 7789
rect 15647 7763 15795 7769
rect 15647 7760 15711 7763
rect 15647 7759 15684 7760
rect 15703 7733 15711 7760
rect 15732 7760 15795 7763
rect 15853 7789 15991 7796
rect 15853 7769 15862 7789
rect 15882 7769 15991 7789
rect 15853 7760 15991 7769
rect 15732 7733 15739 7760
rect 15758 7759 15795 7760
rect 15854 7759 15891 7760
rect 15703 7708 15739 7733
rect 15174 7706 15215 7707
rect 15000 7699 15215 7706
rect 15000 7698 15065 7699
rect 15000 7674 15008 7698
rect 15032 7675 15065 7698
rect 15089 7679 15184 7699
rect 15204 7679 15215 7699
rect 15089 7675 15215 7679
rect 15032 7674 15215 7675
rect 15000 7671 15215 7674
rect 15282 7703 15641 7707
rect 15282 7698 15604 7703
rect 15282 7674 15395 7698
rect 15419 7679 15604 7698
rect 15628 7679 15641 7703
rect 15419 7674 15641 7679
rect 15282 7671 15641 7674
rect 15703 7671 15738 7708
rect 15806 7705 15906 7708
rect 15806 7701 15873 7705
rect 15806 7675 15818 7701
rect 15844 7679 15873 7701
rect 15899 7679 15906 7705
rect 15844 7675 15906 7679
rect 15806 7671 15906 7675
rect 15000 7667 15111 7671
rect 15282 7650 15313 7671
rect 15703 7650 15739 7671
rect 15125 7649 15162 7650
rect 15124 7640 15162 7649
rect 15124 7620 15133 7640
rect 15153 7620 15162 7640
rect 15124 7612 15162 7620
rect 15228 7644 15313 7650
rect 15338 7649 15375 7650
rect 15228 7624 15236 7644
rect 15256 7624 15313 7644
rect 15228 7616 15313 7624
rect 15337 7640 15375 7649
rect 15337 7620 15346 7640
rect 15366 7620 15375 7640
rect 15228 7615 15264 7616
rect 15337 7612 15375 7620
rect 15441 7644 15526 7650
rect 15546 7649 15583 7650
rect 15441 7624 15449 7644
rect 15469 7643 15526 7644
rect 15469 7624 15498 7643
rect 15441 7623 15498 7624
rect 15519 7623 15526 7643
rect 15441 7616 15526 7623
rect 15545 7640 15583 7649
rect 15545 7620 15554 7640
rect 15574 7620 15583 7640
rect 15441 7615 15477 7616
rect 15545 7612 15583 7620
rect 15649 7644 15793 7650
rect 15649 7624 15657 7644
rect 15677 7643 15765 7644
rect 15677 7624 15711 7643
rect 15649 7621 15711 7624
rect 15735 7624 15765 7643
rect 15785 7624 15793 7644
rect 15735 7621 15793 7624
rect 15649 7616 15793 7621
rect 15649 7615 15685 7616
rect 15757 7615 15793 7616
rect 15859 7649 15896 7650
rect 15859 7648 15897 7649
rect 15859 7640 15923 7648
rect 15859 7620 15868 7640
rect 15888 7626 15923 7640
rect 15943 7626 15946 7646
rect 15888 7621 15946 7626
rect 15888 7620 15923 7621
rect 15125 7583 15162 7612
rect 15126 7581 15162 7583
rect 15338 7581 15375 7612
rect 15126 7559 15375 7581
rect 15207 7553 15318 7559
rect 15207 7545 15248 7553
rect 15207 7525 15215 7545
rect 15234 7525 15248 7545
rect 15207 7523 15248 7525
rect 15276 7545 15318 7553
rect 15276 7525 15292 7545
rect 15311 7525 15318 7545
rect 15276 7523 15318 7525
rect 15207 7508 15318 7523
rect 15546 7497 15583 7612
rect 15859 7608 15923 7620
rect 15542 7491 15597 7497
rect 15963 7493 15990 7760
rect 15822 7491 15990 7493
rect 15542 7466 15990 7491
rect 16303 7551 16409 12804
rect 19575 12792 19594 12818
rect 19634 12792 19655 12818
rect 19575 12765 19655 12792
rect 19575 12739 19598 12765
rect 19638 12739 19655 12765
rect 19575 12728 19655 12739
rect 19717 12729 19744 12984
rect 20122 12976 20163 13126
rect 20394 12981 20498 13126
rect 20589 13064 20710 13082
rect 20589 13062 20660 13064
rect 20589 13021 20604 13062
rect 20641 13023 20660 13062
rect 20697 13023 20710 13064
rect 20641 13021 20710 13023
rect 20589 13011 20710 13021
rect 19784 12869 19848 12881
rect 20124 12877 20161 12976
rect 20389 12966 20500 12981
rect 20389 12964 20431 12966
rect 20389 12944 20396 12964
rect 20415 12944 20431 12964
rect 20389 12936 20431 12944
rect 20459 12964 20500 12966
rect 20459 12944 20473 12964
rect 20492 12944 20500 12964
rect 20459 12936 20500 12944
rect 20389 12930 20500 12936
rect 20332 12908 20581 12930
rect 20332 12877 20369 12908
rect 20545 12906 20581 12908
rect 20545 12877 20582 12906
rect 19784 12868 19819 12869
rect 19761 12863 19819 12868
rect 19761 12843 19764 12863
rect 19784 12849 19819 12863
rect 19839 12849 19848 12869
rect 19784 12841 19848 12849
rect 19810 12840 19848 12841
rect 19811 12839 19848 12840
rect 19914 12873 19950 12874
rect 20022 12873 20058 12874
rect 19914 12865 20058 12873
rect 19914 12845 19922 12865
rect 19942 12845 20030 12865
rect 20050 12845 20058 12865
rect 19914 12839 20058 12845
rect 20124 12869 20162 12877
rect 20230 12873 20266 12874
rect 20124 12849 20133 12869
rect 20153 12849 20162 12869
rect 20124 12840 20162 12849
rect 20181 12866 20266 12873
rect 20181 12846 20188 12866
rect 20209 12865 20266 12866
rect 20209 12846 20238 12865
rect 20181 12845 20238 12846
rect 20258 12845 20266 12865
rect 20124 12839 20161 12840
rect 20181 12839 20266 12845
rect 20332 12869 20370 12877
rect 20443 12873 20479 12874
rect 20332 12849 20341 12869
rect 20361 12849 20370 12869
rect 20332 12840 20370 12849
rect 20394 12865 20479 12873
rect 20394 12845 20451 12865
rect 20471 12845 20479 12865
rect 20332 12839 20369 12840
rect 20394 12839 20479 12845
rect 20545 12869 20583 12877
rect 20545 12849 20554 12869
rect 20574 12849 20583 12869
rect 20638 12859 20703 13011
rect 20856 12985 20911 13126
rect 20545 12840 20583 12849
rect 20636 12852 20703 12859
rect 20545 12839 20582 12840
rect 19968 12818 20004 12839
rect 20394 12818 20425 12839
rect 20636 12831 20653 12852
rect 20689 12831 20703 12852
rect 20855 12872 20911 12985
rect 20855 12854 20874 12872
rect 20892 12854 20911 12872
rect 20855 12834 20911 12854
rect 20636 12818 20703 12831
rect 19801 12814 19901 12818
rect 19801 12810 19863 12814
rect 19801 12784 19808 12810
rect 19834 12788 19863 12810
rect 19889 12788 19901 12814
rect 19834 12784 19901 12788
rect 19801 12781 19901 12784
rect 19969 12781 20004 12818
rect 20066 12815 20425 12818
rect 20066 12810 20288 12815
rect 20066 12786 20079 12810
rect 20103 12791 20288 12810
rect 20312 12791 20425 12815
rect 20103 12786 20425 12791
rect 20066 12782 20425 12786
rect 20492 12812 20703 12818
rect 20492 12810 20653 12812
rect 20492 12790 20503 12810
rect 20523 12790 20653 12810
rect 20492 12783 20653 12790
rect 20492 12782 20533 12783
rect 19968 12756 20004 12781
rect 19816 12729 19853 12730
rect 19912 12729 19949 12730
rect 19968 12729 19975 12756
rect 19716 12720 19854 12729
rect 19716 12700 19825 12720
rect 19845 12700 19854 12720
rect 19716 12693 19854 12700
rect 19912 12726 19975 12729
rect 19996 12729 20004 12756
rect 20023 12729 20060 12730
rect 19996 12726 20060 12729
rect 19912 12720 20060 12726
rect 19912 12700 19921 12720
rect 19941 12700 20031 12720
rect 20051 12700 20060 12720
rect 19716 12691 19812 12693
rect 19912 12690 20060 12700
rect 20119 12720 20156 12730
rect 20231 12729 20268 12730
rect 20212 12727 20268 12729
rect 20119 12700 20127 12720
rect 20147 12700 20156 12720
rect 19968 12689 20004 12690
rect 19816 12558 19853 12559
rect 20119 12558 20156 12700
rect 20181 12720 20268 12727
rect 20181 12717 20239 12720
rect 20181 12697 20186 12717
rect 20207 12700 20239 12717
rect 20259 12700 20268 12720
rect 20207 12697 20268 12700
rect 20181 12690 20268 12697
rect 20327 12720 20364 12730
rect 20327 12700 20335 12720
rect 20355 12700 20364 12720
rect 20181 12689 20212 12690
rect 20327 12621 20364 12700
rect 20394 12729 20425 12782
rect 20638 12775 20653 12783
rect 20693 12775 20703 12812
rect 20638 12766 20703 12775
rect 20851 12773 20916 12794
rect 20851 12755 20876 12773
rect 20894 12755 20916 12773
rect 20444 12729 20481 12730
rect 20394 12720 20481 12729
rect 20394 12700 20452 12720
rect 20472 12700 20481 12720
rect 20394 12690 20481 12700
rect 20540 12720 20577 12730
rect 20540 12700 20548 12720
rect 20568 12700 20577 12720
rect 20394 12689 20425 12690
rect 20389 12621 20499 12634
rect 20540 12621 20577 12700
rect 20851 12679 20916 12755
rect 20327 12619 20577 12621
rect 20327 12616 20428 12619
rect 20327 12597 20392 12616
rect 20389 12589 20392 12597
rect 20421 12589 20428 12616
rect 20456 12592 20466 12619
rect 20495 12597 20577 12619
rect 20600 12644 20917 12679
rect 20495 12592 20499 12597
rect 20456 12589 20499 12592
rect 20389 12575 20499 12589
rect 19815 12557 20156 12558
rect 19740 12555 20156 12557
rect 20600 12555 20640 12644
rect 20851 12617 20916 12644
rect 20851 12599 20874 12617
rect 20892 12599 20916 12617
rect 20851 12579 20916 12599
rect 19737 12552 20640 12555
rect 19737 12532 19743 12552
rect 19763 12532 20640 12552
rect 19737 12528 20640 12532
rect 20600 12525 20640 12528
rect 20852 12518 20917 12539
rect 19070 12510 19731 12511
rect 19070 12503 20004 12510
rect 19070 12502 19976 12503
rect 19070 12482 19921 12502
rect 19953 12483 19976 12502
rect 20001 12483 20004 12503
rect 19953 12482 20004 12483
rect 19070 12475 20004 12482
rect 18669 12433 18837 12434
rect 19072 12433 19111 12475
rect 19900 12473 20004 12475
rect 19969 12471 20004 12473
rect 20852 12500 20876 12518
rect 20894 12500 20917 12518
rect 20852 12453 20917 12500
rect 18669 12407 19113 12433
rect 18669 12405 18837 12407
rect 18669 12054 18696 12405
rect 19072 12401 19113 12407
rect 18736 12194 18800 12206
rect 19076 12202 19113 12401
rect 19575 12428 19647 12445
rect 19575 12389 19583 12428
rect 19628 12389 19647 12428
rect 19341 12291 19452 12306
rect 19341 12289 19383 12291
rect 19341 12269 19348 12289
rect 19367 12269 19383 12289
rect 19341 12261 19383 12269
rect 19411 12289 19452 12291
rect 19411 12269 19425 12289
rect 19444 12269 19452 12289
rect 19411 12261 19452 12269
rect 19341 12255 19452 12261
rect 19284 12233 19533 12255
rect 19284 12202 19321 12233
rect 19497 12231 19533 12233
rect 19497 12202 19534 12231
rect 18736 12193 18771 12194
rect 18713 12188 18771 12193
rect 18713 12168 18716 12188
rect 18736 12174 18771 12188
rect 18791 12174 18800 12194
rect 18736 12166 18800 12174
rect 18762 12165 18800 12166
rect 18763 12164 18800 12165
rect 18866 12198 18902 12199
rect 18974 12198 19010 12199
rect 18866 12190 19010 12198
rect 18866 12170 18874 12190
rect 18894 12170 18982 12190
rect 19002 12170 19010 12190
rect 18866 12164 19010 12170
rect 19076 12194 19114 12202
rect 19182 12198 19218 12199
rect 19076 12174 19085 12194
rect 19105 12174 19114 12194
rect 19076 12165 19114 12174
rect 19133 12191 19218 12198
rect 19133 12171 19140 12191
rect 19161 12190 19218 12191
rect 19161 12171 19190 12190
rect 19133 12170 19190 12171
rect 19210 12170 19218 12190
rect 19076 12164 19113 12165
rect 19133 12164 19218 12170
rect 19284 12194 19322 12202
rect 19395 12198 19431 12199
rect 19284 12174 19293 12194
rect 19313 12174 19322 12194
rect 19284 12165 19322 12174
rect 19346 12190 19431 12198
rect 19346 12170 19403 12190
rect 19423 12170 19431 12190
rect 19284 12164 19321 12165
rect 19346 12164 19431 12170
rect 19497 12194 19535 12202
rect 19497 12174 19506 12194
rect 19526 12174 19535 12194
rect 19497 12165 19535 12174
rect 19575 12179 19647 12389
rect 19717 12423 20917 12453
rect 19717 12422 20161 12423
rect 19717 12420 19885 12422
rect 19575 12165 19658 12179
rect 19497 12164 19534 12165
rect 18920 12143 18956 12164
rect 19346 12143 19377 12164
rect 19575 12143 19592 12165
rect 18753 12139 18853 12143
rect 18753 12135 18815 12139
rect 18753 12109 18760 12135
rect 18786 12113 18815 12135
rect 18841 12113 18853 12139
rect 18786 12109 18853 12113
rect 18753 12106 18853 12109
rect 18921 12106 18956 12143
rect 19018 12140 19377 12143
rect 19018 12135 19240 12140
rect 19018 12111 19031 12135
rect 19055 12116 19240 12135
rect 19264 12116 19377 12140
rect 19055 12111 19377 12116
rect 19018 12107 19377 12111
rect 19444 12135 19592 12143
rect 19444 12115 19455 12135
rect 19475 12132 19592 12135
rect 19645 12132 19658 12165
rect 19475 12115 19658 12132
rect 19444 12108 19658 12115
rect 19444 12107 19485 12108
rect 19575 12107 19658 12108
rect 18920 12081 18956 12106
rect 18768 12054 18805 12055
rect 18864 12054 18901 12055
rect 18920 12054 18927 12081
rect 18668 12045 18806 12054
rect 18668 12025 18777 12045
rect 18797 12025 18806 12045
rect 18668 12018 18806 12025
rect 18864 12051 18927 12054
rect 18948 12054 18956 12081
rect 18975 12054 19012 12055
rect 18948 12051 19012 12054
rect 18864 12045 19012 12051
rect 18864 12025 18873 12045
rect 18893 12025 18983 12045
rect 19003 12025 19012 12045
rect 18668 12016 18764 12018
rect 18864 12015 19012 12025
rect 19071 12045 19108 12055
rect 19183 12054 19220 12055
rect 19164 12052 19220 12054
rect 19071 12025 19079 12045
rect 19099 12025 19108 12045
rect 18920 12014 18956 12015
rect 18768 11883 18805 11884
rect 19071 11883 19108 12025
rect 19133 12045 19220 12052
rect 19133 12042 19191 12045
rect 19133 12022 19138 12042
rect 19159 12025 19191 12042
rect 19211 12025 19220 12045
rect 19159 12022 19220 12025
rect 19133 12015 19220 12022
rect 19279 12045 19316 12055
rect 19279 12025 19287 12045
rect 19307 12025 19316 12045
rect 19133 12014 19164 12015
rect 19279 11946 19316 12025
rect 19346 12054 19377 12107
rect 19583 12074 19597 12107
rect 19650 12074 19658 12107
rect 19583 12068 19658 12074
rect 19583 12063 19653 12068
rect 19396 12054 19433 12055
rect 19346 12045 19433 12054
rect 19346 12025 19404 12045
rect 19424 12025 19433 12045
rect 19346 12015 19433 12025
rect 19492 12045 19529 12055
rect 19717 12050 19744 12420
rect 19784 12190 19848 12202
rect 20124 12198 20161 12422
rect 20632 12403 20696 12405
rect 20628 12391 20696 12403
rect 20628 12358 20639 12391
rect 20679 12358 20696 12391
rect 20628 12348 20696 12358
rect 20389 12287 20500 12302
rect 20389 12285 20431 12287
rect 20389 12265 20396 12285
rect 20415 12265 20431 12285
rect 20389 12257 20431 12265
rect 20459 12285 20500 12287
rect 20459 12265 20473 12285
rect 20492 12265 20500 12285
rect 20459 12257 20500 12265
rect 20389 12251 20500 12257
rect 20332 12229 20581 12251
rect 20332 12198 20369 12229
rect 20545 12227 20581 12229
rect 20545 12198 20582 12227
rect 19784 12189 19819 12190
rect 19761 12184 19819 12189
rect 19761 12164 19764 12184
rect 19784 12170 19819 12184
rect 19839 12170 19848 12190
rect 19784 12162 19848 12170
rect 19810 12161 19848 12162
rect 19811 12160 19848 12161
rect 19914 12194 19950 12195
rect 20022 12194 20058 12195
rect 19914 12186 20058 12194
rect 19914 12166 19922 12186
rect 19942 12166 20030 12186
rect 20050 12166 20058 12186
rect 19914 12160 20058 12166
rect 20124 12190 20162 12198
rect 20230 12194 20266 12195
rect 20124 12170 20133 12190
rect 20153 12170 20162 12190
rect 20124 12161 20162 12170
rect 20181 12187 20266 12194
rect 20181 12167 20188 12187
rect 20209 12186 20266 12187
rect 20209 12167 20238 12186
rect 20181 12166 20238 12167
rect 20258 12166 20266 12186
rect 20124 12160 20161 12161
rect 20181 12160 20266 12166
rect 20332 12190 20370 12198
rect 20443 12194 20479 12195
rect 20332 12170 20341 12190
rect 20361 12170 20370 12190
rect 20332 12161 20370 12170
rect 20394 12186 20479 12194
rect 20394 12166 20451 12186
rect 20471 12166 20479 12186
rect 20332 12160 20369 12161
rect 20394 12160 20479 12166
rect 20545 12190 20583 12198
rect 20545 12170 20554 12190
rect 20574 12170 20583 12190
rect 20545 12161 20583 12170
rect 20632 12164 20696 12348
rect 20852 12222 20917 12423
rect 20852 12204 20874 12222
rect 20892 12204 20917 12222
rect 20852 12185 20917 12204
rect 20545 12160 20582 12161
rect 19968 12139 20004 12160
rect 20394 12139 20425 12160
rect 20632 12155 20640 12164
rect 20629 12139 20640 12155
rect 19801 12135 19901 12139
rect 19801 12131 19863 12135
rect 19801 12105 19808 12131
rect 19834 12109 19863 12131
rect 19889 12109 19901 12135
rect 19834 12105 19901 12109
rect 19801 12102 19901 12105
rect 19969 12102 20004 12139
rect 20066 12136 20425 12139
rect 20066 12131 20288 12136
rect 20066 12107 20079 12131
rect 20103 12112 20288 12131
rect 20312 12112 20425 12136
rect 20103 12107 20425 12112
rect 20066 12103 20425 12107
rect 20492 12131 20640 12139
rect 20492 12111 20503 12131
rect 20523 12122 20640 12131
rect 20689 12155 20696 12164
rect 20689 12122 20697 12155
rect 20523 12111 20697 12122
rect 20492 12104 20697 12111
rect 20492 12103 20533 12104
rect 19968 12077 20004 12102
rect 19816 12050 19853 12051
rect 19912 12050 19949 12051
rect 19968 12050 19975 12077
rect 19492 12025 19500 12045
rect 19520 12025 19529 12045
rect 19346 12014 19377 12015
rect 19341 11946 19451 11959
rect 19492 11946 19529 12025
rect 19716 12041 19854 12050
rect 19716 12021 19825 12041
rect 19845 12021 19854 12041
rect 19716 12014 19854 12021
rect 19912 12047 19975 12050
rect 19996 12050 20004 12077
rect 20023 12050 20060 12051
rect 19996 12047 20060 12050
rect 19912 12041 20060 12047
rect 19912 12021 19921 12041
rect 19941 12021 20031 12041
rect 20051 12021 20060 12041
rect 19716 12012 19812 12014
rect 19912 12011 20060 12021
rect 20119 12041 20156 12051
rect 20231 12050 20268 12051
rect 20212 12048 20268 12050
rect 20119 12021 20127 12041
rect 20147 12021 20156 12041
rect 19968 12010 20004 12011
rect 19279 11944 19529 11946
rect 19279 11941 19380 11944
rect 19279 11922 19344 11941
rect 19341 11914 19344 11922
rect 19373 11914 19380 11941
rect 19408 11917 19418 11944
rect 19447 11922 19529 11944
rect 19447 11917 19451 11922
rect 19408 11914 19451 11917
rect 19341 11900 19451 11914
rect 18767 11882 19108 11883
rect 18692 11877 19108 11882
rect 19816 11879 19853 11880
rect 20119 11879 20156 12021
rect 20181 12041 20268 12048
rect 20181 12038 20239 12041
rect 20181 12018 20186 12038
rect 20207 12021 20239 12038
rect 20259 12021 20268 12041
rect 20207 12018 20268 12021
rect 20181 12011 20268 12018
rect 20327 12041 20364 12051
rect 20327 12021 20335 12041
rect 20355 12021 20364 12041
rect 20181 12010 20212 12011
rect 20327 11942 20364 12021
rect 20394 12050 20425 12103
rect 20629 12101 20697 12104
rect 20629 12059 20641 12101
rect 20690 12059 20697 12101
rect 20444 12050 20481 12051
rect 20394 12041 20481 12050
rect 20394 12021 20452 12041
rect 20472 12021 20481 12041
rect 20394 12011 20481 12021
rect 20540 12041 20577 12051
rect 20629 12046 20697 12059
rect 20852 12123 20917 12140
rect 20852 12105 20876 12123
rect 20894 12105 20917 12123
rect 20540 12021 20548 12041
rect 20568 12021 20577 12041
rect 20394 12010 20425 12011
rect 20389 11942 20499 11955
rect 20540 11942 20577 12021
rect 20852 11966 20917 12105
rect 20852 11960 20874 11966
rect 20327 11940 20577 11942
rect 20327 11937 20428 11940
rect 20327 11918 20392 11937
rect 20389 11910 20392 11918
rect 20421 11910 20428 11937
rect 20456 11913 20466 11940
rect 20495 11918 20577 11940
rect 20606 11948 20874 11960
rect 20892 11948 20917 11966
rect 20606 11925 20917 11948
rect 20606 11924 20661 11925
rect 20495 11913 20499 11918
rect 20456 11910 20499 11913
rect 20389 11896 20499 11910
rect 19815 11878 20156 11879
rect 18692 11857 18695 11877
rect 18715 11857 19108 11877
rect 19740 11877 20156 11878
rect 20606 11877 20649 11924
rect 19740 11873 20649 11877
rect 19059 11824 19104 11857
rect 19740 11853 19743 11873
rect 19763 11853 20649 11873
rect 20117 11848 20649 11853
rect 20857 11867 20916 11889
rect 20857 11849 20876 11867
rect 20894 11849 20916 11867
rect 19905 11824 20004 11826
rect 19059 11814 20004 11824
rect 17616 11794 17675 11804
rect 17616 11766 17629 11794
rect 17657 11766 17675 11794
rect 19059 11788 19927 11814
rect 19060 11787 19927 11788
rect 19905 11776 19927 11787
rect 19952 11779 19971 11814
rect 19996 11779 20004 11814
rect 19952 11776 20004 11779
rect 20857 11778 20916 11849
rect 19905 11768 20004 11776
rect 19931 11767 20003 11768
rect 17616 11717 17675 11766
rect 19585 11741 19652 11760
rect 19585 11720 19602 11741
rect 17222 11582 17390 11583
rect 17626 11582 17673 11717
rect 17222 11556 17673 11582
rect 17222 11554 17390 11556
rect 17222 11287 17249 11554
rect 17626 11550 17673 11556
rect 19583 11675 19602 11720
rect 19632 11720 19652 11741
rect 19632 11675 19653 11720
rect 20122 11717 20163 11719
rect 20394 11717 20498 11719
rect 20854 11717 20918 11778
rect 17289 11427 17353 11439
rect 17629 11435 17666 11550
rect 17894 11524 18005 11539
rect 17894 11522 17936 11524
rect 17894 11502 17901 11522
rect 17920 11502 17936 11522
rect 17894 11494 17936 11502
rect 17964 11522 18005 11524
rect 17964 11502 17978 11522
rect 17997 11502 18005 11522
rect 17964 11494 18005 11502
rect 17894 11488 18005 11494
rect 17837 11466 18086 11488
rect 19583 11467 19653 11675
rect 19715 11682 20918 11717
rect 19715 11668 19743 11682
rect 19717 11537 19743 11668
rect 20122 11679 20918 11682
rect 17837 11435 17874 11466
rect 18050 11464 18086 11466
rect 18050 11435 18087 11464
rect 17289 11426 17324 11427
rect 17266 11421 17324 11426
rect 17266 11401 17269 11421
rect 17289 11407 17324 11421
rect 17344 11407 17353 11427
rect 17289 11399 17353 11407
rect 17315 11398 17353 11399
rect 17316 11397 17353 11398
rect 17419 11431 17455 11432
rect 17527 11431 17563 11432
rect 17419 11423 17563 11431
rect 17419 11403 17427 11423
rect 17447 11403 17535 11423
rect 17555 11403 17563 11423
rect 17419 11397 17563 11403
rect 17629 11427 17667 11435
rect 17735 11431 17771 11432
rect 17629 11407 17638 11427
rect 17658 11407 17667 11427
rect 17629 11398 17667 11407
rect 17686 11424 17771 11431
rect 17686 11404 17693 11424
rect 17714 11423 17771 11424
rect 17714 11404 17743 11423
rect 17686 11403 17743 11404
rect 17763 11403 17771 11423
rect 17629 11397 17666 11398
rect 17686 11397 17771 11403
rect 17837 11427 17875 11435
rect 17948 11431 17984 11432
rect 17837 11407 17846 11427
rect 17866 11407 17875 11427
rect 17837 11398 17875 11407
rect 17899 11423 17984 11431
rect 17899 11403 17956 11423
rect 17976 11403 17984 11423
rect 17837 11397 17874 11398
rect 17899 11397 17984 11403
rect 18050 11427 18088 11435
rect 18050 11407 18059 11427
rect 18079 11407 18088 11427
rect 18050 11398 18088 11407
rect 19575 11416 19655 11467
rect 18050 11397 18087 11398
rect 17473 11376 17509 11397
rect 17899 11376 17930 11397
rect 18110 11382 18167 11390
rect 18110 11376 18118 11382
rect 17306 11372 17406 11376
rect 17306 11368 17368 11372
rect 17306 11342 17313 11368
rect 17339 11346 17368 11368
rect 17394 11346 17406 11372
rect 17339 11342 17406 11346
rect 17306 11339 17406 11342
rect 17474 11339 17509 11376
rect 17571 11373 17930 11376
rect 17571 11368 17793 11373
rect 17571 11344 17584 11368
rect 17608 11349 17793 11368
rect 17817 11349 17930 11373
rect 17608 11344 17930 11349
rect 17571 11340 17930 11344
rect 17997 11368 18118 11376
rect 17997 11348 18008 11368
rect 18028 11359 18118 11368
rect 18144 11359 18167 11382
rect 18028 11348 18167 11359
rect 17997 11346 18167 11348
rect 18470 11375 18542 11395
rect 18470 11352 18498 11375
rect 18524 11352 18542 11375
rect 17997 11341 18118 11346
rect 17997 11340 18038 11341
rect 17473 11314 17509 11339
rect 17321 11287 17358 11288
rect 17417 11287 17454 11288
rect 17473 11287 17480 11314
rect 17221 11278 17359 11287
rect 17221 11258 17330 11278
rect 17350 11258 17359 11278
rect 17221 11251 17359 11258
rect 17417 11284 17480 11287
rect 17501 11287 17509 11314
rect 17528 11287 17565 11288
rect 17501 11284 17565 11287
rect 17417 11278 17565 11284
rect 17417 11258 17426 11278
rect 17446 11258 17536 11278
rect 17556 11258 17565 11278
rect 17221 11249 17317 11251
rect 17417 11248 17565 11258
rect 17624 11278 17661 11288
rect 17736 11287 17773 11288
rect 17717 11285 17773 11287
rect 17624 11258 17632 11278
rect 17652 11258 17661 11278
rect 17473 11247 17509 11248
rect 17321 11116 17358 11117
rect 17624 11116 17661 11258
rect 17686 11278 17773 11285
rect 17686 11275 17744 11278
rect 17686 11255 17691 11275
rect 17712 11258 17744 11275
rect 17764 11258 17773 11278
rect 17712 11255 17773 11258
rect 17686 11248 17773 11255
rect 17832 11278 17869 11288
rect 17832 11258 17840 11278
rect 17860 11258 17869 11278
rect 17686 11247 17717 11248
rect 17832 11179 17869 11258
rect 17899 11287 17930 11340
rect 18470 11290 18542 11352
rect 19575 11390 19591 11416
rect 19631 11390 19655 11416
rect 19575 11371 19655 11390
rect 19575 11345 19594 11371
rect 19634 11345 19655 11371
rect 19575 11318 19655 11345
rect 19575 11292 19598 11318
rect 19638 11292 19655 11318
rect 17949 11287 17986 11288
rect 17899 11278 17986 11287
rect 17899 11258 17957 11278
rect 17977 11258 17986 11278
rect 17899 11248 17986 11258
rect 18045 11278 18082 11288
rect 18045 11258 18053 11278
rect 18073 11258 18082 11278
rect 17899 11247 17930 11248
rect 17894 11179 18004 11192
rect 18045 11179 18082 11258
rect 17832 11177 18082 11179
rect 17832 11174 17933 11177
rect 17832 11155 17897 11174
rect 17894 11147 17897 11155
rect 17926 11147 17933 11174
rect 17961 11150 17971 11177
rect 18000 11155 18082 11177
rect 18000 11150 18004 11155
rect 17961 11147 18004 11150
rect 17894 11133 18004 11147
rect 17320 11115 17661 11116
rect 17245 11110 17661 11115
rect 17245 11090 17248 11110
rect 17268 11090 17662 11110
rect 17471 11057 17508 11067
rect 17471 11020 17480 11057
rect 17497 11020 17508 11057
rect 17471 10999 17508 11020
rect 17180 10060 17348 10061
rect 17477 10060 17506 10999
rect 17619 10385 17662 11090
rect 18474 10739 18536 11290
rect 19575 11281 19655 11292
rect 19717 11282 19744 11537
rect 20122 11529 20163 11679
rect 20394 11673 20498 11679
rect 20854 11676 20918 11679
rect 20589 11617 20710 11635
rect 20589 11615 20660 11617
rect 20589 11574 20604 11615
rect 20641 11576 20660 11615
rect 20697 11576 20710 11617
rect 20641 11574 20710 11576
rect 20589 11564 20710 11574
rect 19784 11422 19848 11434
rect 20124 11430 20161 11529
rect 20389 11519 20500 11532
rect 20389 11517 20431 11519
rect 20389 11497 20396 11517
rect 20415 11497 20431 11517
rect 20389 11489 20431 11497
rect 20459 11517 20500 11519
rect 20459 11497 20473 11517
rect 20492 11497 20500 11517
rect 20459 11489 20500 11497
rect 20389 11483 20500 11489
rect 20332 11461 20581 11483
rect 20332 11430 20369 11461
rect 20545 11459 20581 11461
rect 20545 11430 20582 11459
rect 19784 11421 19819 11422
rect 19761 11416 19819 11421
rect 19761 11396 19764 11416
rect 19784 11402 19819 11416
rect 19839 11402 19848 11422
rect 19784 11394 19848 11402
rect 19810 11393 19848 11394
rect 19811 11392 19848 11393
rect 19914 11426 19950 11427
rect 20022 11426 20058 11427
rect 19914 11418 20058 11426
rect 19914 11398 19922 11418
rect 19942 11398 20030 11418
rect 20050 11398 20058 11418
rect 19914 11392 20058 11398
rect 20124 11422 20162 11430
rect 20230 11426 20266 11427
rect 20124 11402 20133 11422
rect 20153 11402 20162 11422
rect 20124 11393 20162 11402
rect 20181 11419 20266 11426
rect 20181 11399 20188 11419
rect 20209 11418 20266 11419
rect 20209 11399 20238 11418
rect 20181 11398 20238 11399
rect 20258 11398 20266 11418
rect 20124 11392 20161 11393
rect 20181 11392 20266 11398
rect 20332 11422 20370 11430
rect 20443 11426 20479 11427
rect 20332 11402 20341 11422
rect 20361 11402 20370 11422
rect 20332 11393 20370 11402
rect 20394 11418 20479 11426
rect 20394 11398 20451 11418
rect 20471 11398 20479 11418
rect 20332 11392 20369 11393
rect 20394 11392 20479 11398
rect 20545 11422 20583 11430
rect 20545 11402 20554 11422
rect 20574 11402 20583 11422
rect 20638 11412 20703 11564
rect 20856 11538 20911 11676
rect 20545 11393 20583 11402
rect 20636 11405 20703 11412
rect 20545 11392 20582 11393
rect 19968 11371 20004 11392
rect 20394 11371 20425 11392
rect 20636 11384 20653 11405
rect 20689 11384 20703 11405
rect 20855 11425 20911 11538
rect 20855 11407 20874 11425
rect 20892 11407 20911 11425
rect 20855 11387 20911 11407
rect 20636 11371 20703 11384
rect 19801 11367 19901 11371
rect 19801 11363 19863 11367
rect 19801 11337 19808 11363
rect 19834 11341 19863 11363
rect 19889 11341 19901 11367
rect 19834 11337 19901 11341
rect 19801 11334 19901 11337
rect 19969 11334 20004 11371
rect 20066 11368 20425 11371
rect 20066 11363 20288 11368
rect 20066 11339 20079 11363
rect 20103 11344 20288 11363
rect 20312 11344 20425 11368
rect 20103 11339 20425 11344
rect 20066 11335 20425 11339
rect 20492 11365 20703 11371
rect 20492 11363 20653 11365
rect 20492 11343 20503 11363
rect 20523 11343 20653 11363
rect 20492 11336 20653 11343
rect 20492 11335 20533 11336
rect 19968 11309 20004 11334
rect 19816 11282 19853 11283
rect 19912 11282 19949 11283
rect 19968 11282 19975 11309
rect 19716 11273 19854 11282
rect 19716 11253 19825 11273
rect 19845 11253 19854 11273
rect 19716 11246 19854 11253
rect 19912 11279 19975 11282
rect 19996 11282 20004 11309
rect 20023 11282 20060 11283
rect 19996 11279 20060 11282
rect 19912 11273 20060 11279
rect 19912 11253 19921 11273
rect 19941 11253 20031 11273
rect 20051 11253 20060 11273
rect 19716 11244 19812 11246
rect 19912 11243 20060 11253
rect 20119 11273 20156 11283
rect 20231 11282 20268 11283
rect 20212 11280 20268 11282
rect 20119 11253 20127 11273
rect 20147 11253 20156 11273
rect 19968 11242 20004 11243
rect 19816 11111 19853 11112
rect 20119 11111 20156 11253
rect 20181 11273 20268 11280
rect 20181 11270 20239 11273
rect 20181 11250 20186 11270
rect 20207 11253 20239 11270
rect 20259 11253 20268 11273
rect 20207 11250 20268 11253
rect 20181 11243 20268 11250
rect 20327 11273 20364 11283
rect 20327 11253 20335 11273
rect 20355 11253 20364 11273
rect 20181 11242 20212 11243
rect 20327 11174 20364 11253
rect 20394 11282 20425 11335
rect 20638 11328 20653 11336
rect 20693 11328 20703 11365
rect 20638 11319 20703 11328
rect 20851 11326 20916 11347
rect 20851 11308 20876 11326
rect 20894 11308 20916 11326
rect 20444 11282 20481 11283
rect 20394 11273 20481 11282
rect 20394 11253 20452 11273
rect 20472 11253 20481 11273
rect 20394 11243 20481 11253
rect 20540 11273 20577 11283
rect 20540 11253 20548 11273
rect 20568 11253 20577 11273
rect 20394 11242 20425 11243
rect 20389 11174 20499 11187
rect 20540 11174 20577 11253
rect 20851 11232 20916 11308
rect 20327 11172 20577 11174
rect 20327 11169 20428 11172
rect 20327 11150 20392 11169
rect 20389 11142 20392 11150
rect 20421 11142 20428 11169
rect 20456 11145 20466 11172
rect 20495 11150 20577 11172
rect 20600 11197 20917 11232
rect 20495 11145 20499 11150
rect 20456 11142 20499 11145
rect 20389 11128 20499 11142
rect 19815 11110 20156 11111
rect 19740 11108 20156 11110
rect 20600 11108 20640 11197
rect 20851 11170 20916 11197
rect 20851 11152 20874 11170
rect 20892 11152 20916 11170
rect 20851 11132 20916 11152
rect 19737 11105 20640 11108
rect 19737 11085 19743 11105
rect 19763 11085 20640 11105
rect 19737 11081 20640 11085
rect 20600 11078 20640 11081
rect 20852 11071 20917 11092
rect 19070 11063 19731 11064
rect 19070 11056 20004 11063
rect 19070 11055 19976 11056
rect 19070 11035 19921 11055
rect 19953 11036 19976 11055
rect 20001 11036 20004 11056
rect 19953 11035 20004 11036
rect 19070 11028 20004 11035
rect 18669 10986 18837 10987
rect 19072 10986 19111 11028
rect 19900 11026 20004 11028
rect 19969 11024 20004 11026
rect 20852 11053 20876 11071
rect 20894 11053 20917 11071
rect 20852 11006 20917 11053
rect 18669 10960 19113 10986
rect 18669 10958 18837 10960
rect 18471 10655 18540 10739
rect 17620 10377 17662 10385
rect 17620 10366 17665 10377
rect 17620 10328 17630 10366
rect 17655 10328 17665 10366
rect 17620 10319 17665 10328
rect 18469 10176 18540 10655
rect 18669 10607 18696 10958
rect 19072 10954 19113 10960
rect 18736 10747 18800 10759
rect 19076 10755 19113 10954
rect 19575 10981 19647 10998
rect 19575 10942 19583 10981
rect 19628 10942 19647 10981
rect 19341 10844 19452 10859
rect 19341 10842 19383 10844
rect 19341 10822 19348 10842
rect 19367 10822 19383 10842
rect 19341 10814 19383 10822
rect 19411 10842 19452 10844
rect 19411 10822 19425 10842
rect 19444 10822 19452 10842
rect 19411 10814 19452 10822
rect 19341 10808 19452 10814
rect 19284 10786 19533 10808
rect 19284 10755 19321 10786
rect 19497 10784 19533 10786
rect 19497 10755 19534 10784
rect 18736 10746 18771 10747
rect 18713 10741 18771 10746
rect 18713 10721 18716 10741
rect 18736 10727 18771 10741
rect 18791 10727 18800 10747
rect 18736 10719 18800 10727
rect 18762 10718 18800 10719
rect 18763 10717 18800 10718
rect 18866 10751 18902 10752
rect 18974 10751 19010 10752
rect 18866 10743 19010 10751
rect 18866 10723 18874 10743
rect 18894 10723 18982 10743
rect 19002 10723 19010 10743
rect 18866 10717 19010 10723
rect 19076 10747 19114 10755
rect 19182 10751 19218 10752
rect 19076 10727 19085 10747
rect 19105 10727 19114 10747
rect 19076 10718 19114 10727
rect 19133 10744 19218 10751
rect 19133 10724 19140 10744
rect 19161 10743 19218 10744
rect 19161 10724 19190 10743
rect 19133 10723 19190 10724
rect 19210 10723 19218 10743
rect 19076 10717 19113 10718
rect 19133 10717 19218 10723
rect 19284 10747 19322 10755
rect 19395 10751 19431 10752
rect 19284 10727 19293 10747
rect 19313 10727 19322 10747
rect 19284 10718 19322 10727
rect 19346 10743 19431 10751
rect 19346 10723 19403 10743
rect 19423 10723 19431 10743
rect 19284 10717 19321 10718
rect 19346 10717 19431 10723
rect 19497 10747 19535 10755
rect 19497 10727 19506 10747
rect 19526 10727 19535 10747
rect 19497 10718 19535 10727
rect 19575 10732 19647 10942
rect 19717 10976 20917 11006
rect 19717 10975 20161 10976
rect 19717 10973 19885 10975
rect 19575 10718 19658 10732
rect 19497 10717 19534 10718
rect 18920 10696 18956 10717
rect 19346 10696 19377 10717
rect 19575 10696 19592 10718
rect 18753 10692 18853 10696
rect 18753 10688 18815 10692
rect 18753 10662 18760 10688
rect 18786 10666 18815 10688
rect 18841 10666 18853 10692
rect 18786 10662 18853 10666
rect 18753 10659 18853 10662
rect 18921 10659 18956 10696
rect 19018 10693 19377 10696
rect 19018 10688 19240 10693
rect 19018 10664 19031 10688
rect 19055 10669 19240 10688
rect 19264 10669 19377 10693
rect 19055 10664 19377 10669
rect 19018 10660 19377 10664
rect 19444 10688 19592 10696
rect 19444 10668 19455 10688
rect 19475 10685 19592 10688
rect 19645 10685 19658 10718
rect 19475 10668 19658 10685
rect 19444 10661 19658 10668
rect 19444 10660 19485 10661
rect 19575 10660 19658 10661
rect 18920 10634 18956 10659
rect 18768 10607 18805 10608
rect 18864 10607 18901 10608
rect 18920 10607 18927 10634
rect 18668 10598 18806 10607
rect 18668 10578 18777 10598
rect 18797 10578 18806 10598
rect 18668 10571 18806 10578
rect 18864 10604 18927 10607
rect 18948 10607 18956 10634
rect 18975 10607 19012 10608
rect 18948 10604 19012 10607
rect 18864 10598 19012 10604
rect 18864 10578 18873 10598
rect 18893 10578 18983 10598
rect 19003 10578 19012 10598
rect 18668 10569 18764 10571
rect 18864 10568 19012 10578
rect 19071 10598 19108 10608
rect 19183 10607 19220 10608
rect 19164 10605 19220 10607
rect 19071 10578 19079 10598
rect 19099 10578 19108 10598
rect 18920 10567 18956 10568
rect 18768 10436 18805 10437
rect 19071 10436 19108 10578
rect 19133 10598 19220 10605
rect 19133 10595 19191 10598
rect 19133 10575 19138 10595
rect 19159 10578 19191 10595
rect 19211 10578 19220 10598
rect 19159 10575 19220 10578
rect 19133 10568 19220 10575
rect 19279 10598 19316 10608
rect 19279 10578 19287 10598
rect 19307 10578 19316 10598
rect 19133 10567 19164 10568
rect 19279 10499 19316 10578
rect 19346 10607 19377 10660
rect 19583 10627 19597 10660
rect 19650 10627 19658 10660
rect 19583 10621 19658 10627
rect 19583 10616 19653 10621
rect 19396 10607 19433 10608
rect 19346 10598 19433 10607
rect 19346 10578 19404 10598
rect 19424 10578 19433 10598
rect 19346 10568 19433 10578
rect 19492 10598 19529 10608
rect 19717 10603 19744 10973
rect 19784 10743 19848 10755
rect 20124 10751 20161 10975
rect 20632 10956 20696 10958
rect 20628 10944 20696 10956
rect 20628 10911 20639 10944
rect 20679 10911 20696 10944
rect 20628 10901 20696 10911
rect 20389 10840 20500 10855
rect 20389 10838 20431 10840
rect 20389 10818 20396 10838
rect 20415 10818 20431 10838
rect 20389 10810 20431 10818
rect 20459 10838 20500 10840
rect 20459 10818 20473 10838
rect 20492 10818 20500 10838
rect 20459 10810 20500 10818
rect 20389 10804 20500 10810
rect 20332 10782 20581 10804
rect 20332 10751 20369 10782
rect 20545 10780 20581 10782
rect 20545 10751 20582 10780
rect 19784 10742 19819 10743
rect 19761 10737 19819 10742
rect 19761 10717 19764 10737
rect 19784 10723 19819 10737
rect 19839 10723 19848 10743
rect 19784 10715 19848 10723
rect 19810 10714 19848 10715
rect 19811 10713 19848 10714
rect 19914 10747 19950 10748
rect 20022 10747 20058 10748
rect 19914 10739 20058 10747
rect 19914 10719 19922 10739
rect 19942 10719 20030 10739
rect 20050 10719 20058 10739
rect 19914 10713 20058 10719
rect 20124 10743 20162 10751
rect 20230 10747 20266 10748
rect 20124 10723 20133 10743
rect 20153 10723 20162 10743
rect 20124 10714 20162 10723
rect 20181 10740 20266 10747
rect 20181 10720 20188 10740
rect 20209 10739 20266 10740
rect 20209 10720 20238 10739
rect 20181 10719 20238 10720
rect 20258 10719 20266 10739
rect 20124 10713 20161 10714
rect 20181 10713 20266 10719
rect 20332 10743 20370 10751
rect 20443 10747 20479 10748
rect 20332 10723 20341 10743
rect 20361 10723 20370 10743
rect 20332 10714 20370 10723
rect 20394 10739 20479 10747
rect 20394 10719 20451 10739
rect 20471 10719 20479 10739
rect 20332 10713 20369 10714
rect 20394 10713 20479 10719
rect 20545 10743 20583 10751
rect 20545 10723 20554 10743
rect 20574 10723 20583 10743
rect 20545 10714 20583 10723
rect 20632 10717 20696 10901
rect 20852 10775 20917 10976
rect 20852 10757 20874 10775
rect 20892 10757 20917 10775
rect 20852 10738 20917 10757
rect 20545 10713 20582 10714
rect 19968 10692 20004 10713
rect 20394 10692 20425 10713
rect 20632 10708 20640 10717
rect 20629 10692 20640 10708
rect 19801 10688 19901 10692
rect 19801 10684 19863 10688
rect 19801 10658 19808 10684
rect 19834 10662 19863 10684
rect 19889 10662 19901 10688
rect 19834 10658 19901 10662
rect 19801 10655 19901 10658
rect 19969 10655 20004 10692
rect 20066 10689 20425 10692
rect 20066 10684 20288 10689
rect 20066 10660 20079 10684
rect 20103 10665 20288 10684
rect 20312 10665 20425 10689
rect 20103 10660 20425 10665
rect 20066 10656 20425 10660
rect 20492 10684 20640 10692
rect 20492 10664 20503 10684
rect 20523 10675 20640 10684
rect 20689 10708 20696 10717
rect 20689 10675 20697 10708
rect 20523 10664 20697 10675
rect 20492 10657 20697 10664
rect 20492 10656 20533 10657
rect 19968 10630 20004 10655
rect 19816 10603 19853 10604
rect 19912 10603 19949 10604
rect 19968 10603 19975 10630
rect 19492 10578 19500 10598
rect 19520 10578 19529 10598
rect 19346 10567 19377 10568
rect 19341 10499 19451 10512
rect 19492 10499 19529 10578
rect 19716 10594 19854 10603
rect 19716 10574 19825 10594
rect 19845 10574 19854 10594
rect 19716 10567 19854 10574
rect 19912 10600 19975 10603
rect 19996 10603 20004 10630
rect 20023 10603 20060 10604
rect 19996 10600 20060 10603
rect 19912 10594 20060 10600
rect 19912 10574 19921 10594
rect 19941 10574 20031 10594
rect 20051 10574 20060 10594
rect 19716 10565 19812 10567
rect 19912 10564 20060 10574
rect 20119 10594 20156 10604
rect 20231 10603 20268 10604
rect 20212 10601 20268 10603
rect 20119 10574 20127 10594
rect 20147 10574 20156 10594
rect 19968 10563 20004 10564
rect 19279 10497 19529 10499
rect 19279 10494 19380 10497
rect 19279 10475 19344 10494
rect 19341 10467 19344 10475
rect 19373 10467 19380 10494
rect 19408 10470 19418 10497
rect 19447 10475 19529 10497
rect 19447 10470 19451 10475
rect 19408 10467 19451 10470
rect 19341 10453 19451 10467
rect 18767 10435 19108 10436
rect 18692 10430 19108 10435
rect 19816 10432 19853 10433
rect 20119 10432 20156 10574
rect 20181 10594 20268 10601
rect 20181 10591 20239 10594
rect 20181 10571 20186 10591
rect 20207 10574 20239 10591
rect 20259 10574 20268 10594
rect 20207 10571 20268 10574
rect 20181 10564 20268 10571
rect 20327 10594 20364 10604
rect 20327 10574 20335 10594
rect 20355 10574 20364 10594
rect 20181 10563 20212 10564
rect 20327 10495 20364 10574
rect 20394 10603 20425 10656
rect 20629 10654 20697 10657
rect 20629 10612 20641 10654
rect 20690 10612 20697 10654
rect 20444 10603 20481 10604
rect 20394 10594 20481 10603
rect 20394 10574 20452 10594
rect 20472 10574 20481 10594
rect 20394 10564 20481 10574
rect 20540 10594 20577 10604
rect 20629 10599 20697 10612
rect 20852 10676 20917 10693
rect 20852 10658 20876 10676
rect 20894 10658 20917 10676
rect 20540 10574 20548 10594
rect 20568 10574 20577 10594
rect 20394 10563 20425 10564
rect 20389 10495 20499 10508
rect 20540 10495 20577 10574
rect 20852 10519 20917 10658
rect 20852 10513 20874 10519
rect 20327 10493 20577 10495
rect 20327 10490 20428 10493
rect 20327 10471 20392 10490
rect 20389 10463 20392 10471
rect 20421 10463 20428 10490
rect 20456 10466 20466 10493
rect 20495 10471 20577 10493
rect 20606 10501 20874 10513
rect 20892 10501 20917 10519
rect 20606 10478 20917 10501
rect 20606 10477 20661 10478
rect 20495 10466 20499 10471
rect 20456 10463 20499 10466
rect 20389 10449 20499 10463
rect 19815 10431 20156 10432
rect 18692 10410 18695 10430
rect 18715 10410 19108 10430
rect 19740 10430 20156 10431
rect 20606 10430 20649 10477
rect 19740 10426 20649 10430
rect 19059 10377 19104 10410
rect 19740 10406 19743 10426
rect 19763 10406 20649 10426
rect 20117 10401 20649 10406
rect 20857 10420 20916 10442
rect 20857 10402 20876 10420
rect 20894 10402 20916 10420
rect 19905 10377 20004 10379
rect 19059 10367 20004 10377
rect 19059 10341 19927 10367
rect 19060 10340 19927 10341
rect 19905 10329 19927 10340
rect 19952 10332 19971 10367
rect 19996 10332 20004 10367
rect 19952 10329 20004 10332
rect 19905 10321 20004 10329
rect 19931 10320 20003 10321
rect 20857 10272 20916 10402
rect 19579 10242 19655 10266
rect 19579 10176 19591 10242
rect 19645 10176 19655 10242
rect 20123 10197 20164 10199
rect 20395 10197 20499 10199
rect 20857 10197 20918 10272
rect 18469 10126 18541 10176
rect 17180 10034 17624 10060
rect 17180 10032 17348 10034
rect 17180 9765 17207 10032
rect 17477 10030 17506 10034
rect 17247 9905 17311 9917
rect 17587 9913 17624 10034
rect 17852 10002 17963 10017
rect 17852 10000 17894 10002
rect 17852 9980 17859 10000
rect 17878 9980 17894 10000
rect 17852 9972 17894 9980
rect 17922 10000 17963 10002
rect 17922 9980 17936 10000
rect 17955 9980 17963 10000
rect 17922 9972 17963 9980
rect 17852 9966 17963 9972
rect 17795 9944 18044 9966
rect 17795 9913 17832 9944
rect 18008 9942 18044 9944
rect 18008 9913 18045 9942
rect 17247 9904 17282 9905
rect 17224 9899 17282 9904
rect 17224 9879 17227 9899
rect 17247 9885 17282 9899
rect 17302 9885 17311 9905
rect 17247 9877 17311 9885
rect 17273 9876 17311 9877
rect 17274 9875 17311 9876
rect 17377 9909 17413 9910
rect 17485 9909 17521 9910
rect 17377 9901 17521 9909
rect 17377 9881 17385 9901
rect 17405 9881 17493 9901
rect 17513 9881 17521 9901
rect 17377 9875 17521 9881
rect 17587 9905 17625 9913
rect 17693 9909 17729 9910
rect 17587 9885 17596 9905
rect 17616 9885 17625 9905
rect 17587 9876 17625 9885
rect 17644 9902 17729 9909
rect 17644 9882 17651 9902
rect 17672 9901 17729 9902
rect 17672 9882 17701 9901
rect 17644 9881 17701 9882
rect 17721 9881 17729 9901
rect 17587 9875 17624 9876
rect 17644 9875 17729 9881
rect 17795 9905 17833 9913
rect 17906 9909 17942 9910
rect 17795 9885 17804 9905
rect 17824 9885 17833 9905
rect 17795 9876 17833 9885
rect 17857 9901 17942 9909
rect 17857 9881 17914 9901
rect 17934 9881 17942 9901
rect 17795 9875 17832 9876
rect 17857 9875 17942 9881
rect 18008 9905 18046 9913
rect 18008 9885 18017 9905
rect 18037 9885 18046 9905
rect 18008 9876 18046 9885
rect 18008 9875 18045 9876
rect 17431 9854 17467 9875
rect 17857 9854 17888 9875
rect 18038 9854 18372 9858
rect 17264 9850 17364 9854
rect 17264 9846 17326 9850
rect 17264 9820 17271 9846
rect 17297 9824 17326 9846
rect 17352 9824 17364 9850
rect 17297 9820 17364 9824
rect 17264 9817 17364 9820
rect 17432 9817 17467 9854
rect 17529 9851 17888 9854
rect 17529 9846 17751 9851
rect 17529 9822 17542 9846
rect 17566 9827 17751 9846
rect 17775 9827 17888 9851
rect 17566 9822 17888 9827
rect 17529 9818 17888 9822
rect 17955 9846 18372 9854
rect 17955 9826 17966 9846
rect 17986 9826 18372 9846
rect 17955 9819 18372 9826
rect 17955 9818 17996 9819
rect 18038 9818 18372 9819
rect 17431 9792 17467 9817
rect 17279 9765 17316 9766
rect 17375 9765 17412 9766
rect 17431 9765 17438 9792
rect 17179 9756 17317 9765
rect 17179 9736 17288 9756
rect 17308 9736 17317 9756
rect 17179 9729 17317 9736
rect 17375 9762 17438 9765
rect 17459 9765 17467 9792
rect 17486 9765 17523 9766
rect 17459 9762 17523 9765
rect 17375 9756 17523 9762
rect 17375 9736 17384 9756
rect 17404 9736 17494 9756
rect 17514 9736 17523 9756
rect 17179 9727 17275 9729
rect 17375 9726 17523 9736
rect 17582 9756 17619 9766
rect 17694 9765 17731 9766
rect 17675 9763 17731 9765
rect 17582 9736 17590 9756
rect 17610 9736 17619 9756
rect 17431 9725 17467 9726
rect 17279 9594 17316 9595
rect 17582 9594 17619 9736
rect 17644 9756 17731 9763
rect 17644 9753 17702 9756
rect 17644 9733 17649 9753
rect 17670 9736 17702 9753
rect 17722 9736 17731 9756
rect 17670 9733 17731 9736
rect 17644 9726 17731 9733
rect 17790 9756 17827 9766
rect 17790 9736 17798 9756
rect 17818 9736 17827 9756
rect 17644 9725 17675 9726
rect 17790 9657 17827 9736
rect 17857 9765 17888 9818
rect 17907 9765 17944 9766
rect 17857 9756 17944 9765
rect 17857 9736 17915 9756
rect 17935 9736 17944 9756
rect 17857 9726 17944 9736
rect 18003 9756 18040 9766
rect 18003 9736 18011 9756
rect 18031 9736 18040 9756
rect 17857 9725 17888 9726
rect 17852 9657 17962 9670
rect 18003 9657 18040 9736
rect 17790 9655 18040 9657
rect 17790 9652 17891 9655
rect 17790 9633 17855 9652
rect 17852 9625 17855 9633
rect 17884 9625 17891 9652
rect 17919 9628 17929 9655
rect 17958 9633 18040 9655
rect 17958 9628 17962 9633
rect 17919 9625 17962 9628
rect 17852 9611 17962 9625
rect 17278 9593 17619 9594
rect 17203 9588 17619 9593
rect 17203 9568 17206 9588
rect 17226 9568 17619 9588
rect 17512 9203 17543 9568
rect 17430 9174 17543 9203
rect 17431 8874 17467 9174
rect 18291 9069 18372 9818
rect 18471 9217 18541 10126
rect 19579 10156 19655 10176
rect 19579 10119 19596 10156
rect 19640 10119 19655 10156
rect 19716 10162 20918 10197
rect 19716 10148 19744 10162
rect 19579 10103 19655 10119
rect 19584 9947 19654 10103
rect 19718 10017 19744 10148
rect 20123 10159 20918 10162
rect 19576 9896 19656 9947
rect 19576 9870 19592 9896
rect 19632 9870 19656 9896
rect 19576 9851 19656 9870
rect 19576 9825 19595 9851
rect 19635 9825 19656 9851
rect 19576 9798 19656 9825
rect 19576 9772 19599 9798
rect 19639 9772 19656 9798
rect 19576 9761 19656 9772
rect 19718 9762 19745 10017
rect 20123 10009 20164 10159
rect 20857 10147 20918 10159
rect 20590 10097 20711 10115
rect 20590 10095 20661 10097
rect 20590 10054 20605 10095
rect 20642 10056 20661 10095
rect 20698 10056 20711 10097
rect 20642 10054 20711 10056
rect 20590 10044 20711 10054
rect 20395 10014 20499 10023
rect 19785 9902 19849 9914
rect 20125 9910 20162 10009
rect 20390 9999 20501 10014
rect 20390 9997 20432 9999
rect 20390 9977 20397 9997
rect 20416 9977 20432 9997
rect 20390 9969 20432 9977
rect 20460 9997 20501 9999
rect 20460 9977 20474 9997
rect 20493 9977 20501 9997
rect 20460 9969 20501 9977
rect 20390 9963 20501 9969
rect 20333 9941 20582 9963
rect 20333 9910 20370 9941
rect 20546 9939 20582 9941
rect 20546 9910 20583 9939
rect 19785 9901 19820 9902
rect 19762 9896 19820 9901
rect 19762 9876 19765 9896
rect 19785 9882 19820 9896
rect 19840 9882 19849 9902
rect 19785 9874 19849 9882
rect 19811 9873 19849 9874
rect 19812 9872 19849 9873
rect 19915 9906 19951 9907
rect 20023 9906 20059 9907
rect 19915 9898 20059 9906
rect 19915 9878 19923 9898
rect 19943 9878 20031 9898
rect 20051 9878 20059 9898
rect 19915 9872 20059 9878
rect 20125 9902 20163 9910
rect 20231 9906 20267 9907
rect 20125 9882 20134 9902
rect 20154 9882 20163 9902
rect 20125 9873 20163 9882
rect 20182 9899 20267 9906
rect 20182 9879 20189 9899
rect 20210 9898 20267 9899
rect 20210 9879 20239 9898
rect 20182 9878 20239 9879
rect 20259 9878 20267 9898
rect 20125 9872 20162 9873
rect 20182 9872 20267 9878
rect 20333 9902 20371 9910
rect 20444 9906 20480 9907
rect 20333 9882 20342 9902
rect 20362 9882 20371 9902
rect 20333 9873 20371 9882
rect 20395 9898 20480 9906
rect 20395 9878 20452 9898
rect 20472 9878 20480 9898
rect 20333 9872 20370 9873
rect 20395 9872 20480 9878
rect 20546 9902 20584 9910
rect 20546 9882 20555 9902
rect 20575 9882 20584 9902
rect 20639 9892 20704 10044
rect 20857 10018 20912 10147
rect 20546 9873 20584 9882
rect 20637 9885 20704 9892
rect 20546 9872 20583 9873
rect 19969 9851 20005 9872
rect 20395 9851 20426 9872
rect 20637 9864 20654 9885
rect 20690 9864 20704 9885
rect 20856 9905 20912 10018
rect 20856 9887 20875 9905
rect 20893 9887 20912 9905
rect 20856 9867 20912 9887
rect 20637 9851 20704 9864
rect 19802 9847 19902 9851
rect 19802 9843 19864 9847
rect 19802 9817 19809 9843
rect 19835 9821 19864 9843
rect 19890 9821 19902 9847
rect 19835 9817 19902 9821
rect 19802 9814 19902 9817
rect 19970 9814 20005 9851
rect 20067 9848 20426 9851
rect 20067 9843 20289 9848
rect 20067 9819 20080 9843
rect 20104 9824 20289 9843
rect 20313 9824 20426 9848
rect 20104 9819 20426 9824
rect 20067 9815 20426 9819
rect 20493 9845 20704 9851
rect 20493 9843 20654 9845
rect 20493 9823 20504 9843
rect 20524 9823 20654 9843
rect 20493 9816 20654 9823
rect 20493 9815 20534 9816
rect 19969 9789 20005 9814
rect 19817 9762 19854 9763
rect 19913 9762 19950 9763
rect 19969 9762 19976 9789
rect 19717 9753 19855 9762
rect 19717 9733 19826 9753
rect 19846 9733 19855 9753
rect 19717 9726 19855 9733
rect 19913 9759 19976 9762
rect 19997 9762 20005 9789
rect 20024 9762 20061 9763
rect 19997 9759 20061 9762
rect 19913 9753 20061 9759
rect 19913 9733 19922 9753
rect 19942 9733 20032 9753
rect 20052 9733 20061 9753
rect 19717 9724 19813 9726
rect 19913 9723 20061 9733
rect 20120 9753 20157 9763
rect 20232 9762 20269 9763
rect 20213 9760 20269 9762
rect 20120 9733 20128 9753
rect 20148 9733 20157 9753
rect 19969 9722 20005 9723
rect 19817 9591 19854 9592
rect 20120 9591 20157 9733
rect 20182 9753 20269 9760
rect 20182 9750 20240 9753
rect 20182 9730 20187 9750
rect 20208 9733 20240 9750
rect 20260 9733 20269 9753
rect 20208 9730 20269 9733
rect 20182 9723 20269 9730
rect 20328 9753 20365 9763
rect 20328 9733 20336 9753
rect 20356 9733 20365 9753
rect 20182 9722 20213 9723
rect 20328 9654 20365 9733
rect 20395 9762 20426 9815
rect 20639 9808 20654 9816
rect 20694 9808 20704 9845
rect 20639 9799 20704 9808
rect 20852 9806 20917 9827
rect 20852 9788 20877 9806
rect 20895 9788 20917 9806
rect 20445 9762 20482 9763
rect 20395 9753 20482 9762
rect 20395 9733 20453 9753
rect 20473 9733 20482 9753
rect 20395 9723 20482 9733
rect 20541 9753 20578 9763
rect 20541 9733 20549 9753
rect 20569 9733 20578 9753
rect 20395 9722 20426 9723
rect 20390 9654 20500 9667
rect 20541 9654 20578 9733
rect 20852 9712 20917 9788
rect 20328 9652 20578 9654
rect 20328 9649 20429 9652
rect 20328 9630 20393 9649
rect 20390 9622 20393 9630
rect 20422 9622 20429 9649
rect 20457 9625 20467 9652
rect 20496 9630 20578 9652
rect 20601 9677 20918 9712
rect 20496 9625 20500 9630
rect 20457 9622 20500 9625
rect 20390 9608 20500 9622
rect 19816 9590 20157 9591
rect 19741 9588 20157 9590
rect 20601 9588 20641 9677
rect 20852 9650 20917 9677
rect 20852 9632 20875 9650
rect 20893 9632 20917 9650
rect 20852 9612 20917 9632
rect 19738 9585 20641 9588
rect 19738 9565 19744 9585
rect 19764 9565 20641 9585
rect 19738 9561 20641 9565
rect 20601 9558 20641 9561
rect 20853 9551 20918 9572
rect 19071 9543 19732 9544
rect 19071 9536 20005 9543
rect 19071 9535 19977 9536
rect 19071 9515 19922 9535
rect 19954 9516 19977 9535
rect 20002 9516 20005 9536
rect 19954 9515 20005 9516
rect 19071 9508 20005 9515
rect 18670 9466 18838 9467
rect 19073 9466 19112 9508
rect 19901 9506 20005 9508
rect 19970 9504 20005 9506
rect 20853 9533 20877 9551
rect 20895 9533 20918 9551
rect 20853 9486 20918 9533
rect 18670 9440 19114 9466
rect 18670 9438 18838 9440
rect 17431 8851 17435 8874
rect 17459 8851 17467 8874
rect 17631 8852 17730 8856
rect 17431 8830 17467 8851
rect 17431 8807 17435 8830
rect 17459 8807 17467 8830
rect 17431 8803 17467 8807
rect 17627 8846 17730 8852
rect 17627 8808 17653 8846
rect 17678 8811 17697 8846
rect 17722 8811 17730 8846
rect 17678 8808 17730 8811
rect 17627 8800 17730 8808
rect 17627 8799 17729 8800
rect 17223 8721 17391 8722
rect 17627 8721 17674 8799
rect 17223 8695 17674 8721
rect 17223 8693 17391 8695
rect 17223 8320 17250 8693
rect 17420 8645 17506 8654
rect 17420 8627 17439 8645
rect 17491 8627 17506 8645
rect 17420 8623 17506 8627
rect 17290 8460 17354 8472
rect 17290 8459 17325 8460
rect 17267 8454 17325 8459
rect 17267 8434 17270 8454
rect 17290 8440 17325 8454
rect 17345 8440 17354 8460
rect 17290 8432 17354 8440
rect 17316 8431 17354 8432
rect 17317 8430 17354 8431
rect 17420 8464 17456 8465
rect 17476 8464 17506 8623
rect 17627 8583 17674 8695
rect 17630 8468 17667 8583
rect 17895 8557 18006 8572
rect 17895 8555 17937 8557
rect 17895 8535 17902 8555
rect 17921 8535 17937 8555
rect 17895 8527 17937 8535
rect 17965 8555 18006 8557
rect 17965 8535 17979 8555
rect 17998 8535 18006 8555
rect 17965 8527 18006 8535
rect 17895 8521 18006 8527
rect 17838 8499 18087 8521
rect 17838 8468 17875 8499
rect 18051 8497 18087 8499
rect 18051 8468 18088 8497
rect 18292 8484 18371 9069
rect 18468 8617 18547 9217
rect 18670 9087 18697 9438
rect 19073 9434 19114 9440
rect 18737 9227 18801 9239
rect 19077 9235 19114 9434
rect 19576 9461 19648 9478
rect 19576 9422 19584 9461
rect 19629 9422 19648 9461
rect 19342 9324 19453 9339
rect 19342 9322 19384 9324
rect 19342 9302 19349 9322
rect 19368 9302 19384 9322
rect 19342 9294 19384 9302
rect 19412 9322 19453 9324
rect 19412 9302 19426 9322
rect 19445 9302 19453 9322
rect 19412 9294 19453 9302
rect 19342 9288 19453 9294
rect 19285 9266 19534 9288
rect 19285 9235 19322 9266
rect 19498 9264 19534 9266
rect 19498 9235 19535 9264
rect 18737 9226 18772 9227
rect 18714 9221 18772 9226
rect 18714 9201 18717 9221
rect 18737 9207 18772 9221
rect 18792 9207 18801 9227
rect 18737 9199 18801 9207
rect 18763 9198 18801 9199
rect 18764 9197 18801 9198
rect 18867 9231 18903 9232
rect 18975 9231 19011 9232
rect 18867 9223 19011 9231
rect 18867 9203 18875 9223
rect 18895 9203 18983 9223
rect 19003 9203 19011 9223
rect 18867 9197 19011 9203
rect 19077 9227 19115 9235
rect 19183 9231 19219 9232
rect 19077 9207 19086 9227
rect 19106 9207 19115 9227
rect 19077 9198 19115 9207
rect 19134 9224 19219 9231
rect 19134 9204 19141 9224
rect 19162 9223 19219 9224
rect 19162 9204 19191 9223
rect 19134 9203 19191 9204
rect 19211 9203 19219 9223
rect 19077 9197 19114 9198
rect 19134 9197 19219 9203
rect 19285 9227 19323 9235
rect 19396 9231 19432 9232
rect 19285 9207 19294 9227
rect 19314 9207 19323 9227
rect 19285 9198 19323 9207
rect 19347 9223 19432 9231
rect 19347 9203 19404 9223
rect 19424 9203 19432 9223
rect 19285 9197 19322 9198
rect 19347 9197 19432 9203
rect 19498 9227 19536 9235
rect 19498 9207 19507 9227
rect 19527 9207 19536 9227
rect 19498 9198 19536 9207
rect 19576 9212 19648 9422
rect 19718 9456 20918 9486
rect 19718 9455 20162 9456
rect 19718 9453 19886 9455
rect 19576 9198 19659 9212
rect 19498 9197 19535 9198
rect 18921 9176 18957 9197
rect 19347 9176 19378 9197
rect 19576 9176 19593 9198
rect 18754 9172 18854 9176
rect 18754 9168 18816 9172
rect 18754 9142 18761 9168
rect 18787 9146 18816 9168
rect 18842 9146 18854 9172
rect 18787 9142 18854 9146
rect 18754 9139 18854 9142
rect 18922 9139 18957 9176
rect 19019 9173 19378 9176
rect 19019 9168 19241 9173
rect 19019 9144 19032 9168
rect 19056 9149 19241 9168
rect 19265 9149 19378 9173
rect 19056 9144 19378 9149
rect 19019 9140 19378 9144
rect 19445 9168 19593 9176
rect 19445 9148 19456 9168
rect 19476 9165 19593 9168
rect 19646 9165 19659 9198
rect 19476 9148 19659 9165
rect 19445 9141 19659 9148
rect 19445 9140 19486 9141
rect 19576 9140 19659 9141
rect 18921 9114 18957 9139
rect 18769 9087 18806 9088
rect 18865 9087 18902 9088
rect 18921 9087 18928 9114
rect 18669 9078 18807 9087
rect 18669 9058 18778 9078
rect 18798 9058 18807 9078
rect 18669 9051 18807 9058
rect 18865 9084 18928 9087
rect 18949 9087 18957 9114
rect 18976 9087 19013 9088
rect 18949 9084 19013 9087
rect 18865 9078 19013 9084
rect 18865 9058 18874 9078
rect 18894 9058 18984 9078
rect 19004 9058 19013 9078
rect 18669 9049 18765 9051
rect 18865 9048 19013 9058
rect 19072 9078 19109 9088
rect 19184 9087 19221 9088
rect 19165 9085 19221 9087
rect 19072 9058 19080 9078
rect 19100 9058 19109 9078
rect 18921 9047 18957 9048
rect 18769 8916 18806 8917
rect 19072 8916 19109 9058
rect 19134 9078 19221 9085
rect 19134 9075 19192 9078
rect 19134 9055 19139 9075
rect 19160 9058 19192 9075
rect 19212 9058 19221 9078
rect 19160 9055 19221 9058
rect 19134 9048 19221 9055
rect 19280 9078 19317 9088
rect 19280 9058 19288 9078
rect 19308 9058 19317 9078
rect 19134 9047 19165 9048
rect 19280 8979 19317 9058
rect 19347 9087 19378 9140
rect 19584 9107 19598 9140
rect 19651 9107 19659 9140
rect 19584 9101 19659 9107
rect 19584 9096 19654 9101
rect 19397 9087 19434 9088
rect 19347 9078 19434 9087
rect 19347 9058 19405 9078
rect 19425 9058 19434 9078
rect 19347 9048 19434 9058
rect 19493 9078 19530 9088
rect 19718 9083 19745 9453
rect 19785 9223 19849 9235
rect 20125 9231 20162 9455
rect 20633 9436 20697 9438
rect 20629 9424 20697 9436
rect 20629 9391 20640 9424
rect 20680 9391 20697 9424
rect 20629 9381 20697 9391
rect 20390 9320 20501 9335
rect 20390 9318 20432 9320
rect 20390 9298 20397 9318
rect 20416 9298 20432 9318
rect 20390 9290 20432 9298
rect 20460 9318 20501 9320
rect 20460 9298 20474 9318
rect 20493 9298 20501 9318
rect 20460 9290 20501 9298
rect 20390 9284 20501 9290
rect 20333 9262 20582 9284
rect 20333 9231 20370 9262
rect 20546 9260 20582 9262
rect 20546 9231 20583 9260
rect 19785 9222 19820 9223
rect 19762 9217 19820 9222
rect 19762 9197 19765 9217
rect 19785 9203 19820 9217
rect 19840 9203 19849 9223
rect 19785 9195 19849 9203
rect 19811 9194 19849 9195
rect 19812 9193 19849 9194
rect 19915 9227 19951 9228
rect 20023 9227 20059 9228
rect 19915 9219 20059 9227
rect 19915 9199 19923 9219
rect 19943 9199 20031 9219
rect 20051 9199 20059 9219
rect 19915 9193 20059 9199
rect 20125 9223 20163 9231
rect 20231 9227 20267 9228
rect 20125 9203 20134 9223
rect 20154 9203 20163 9223
rect 20125 9194 20163 9203
rect 20182 9220 20267 9227
rect 20182 9200 20189 9220
rect 20210 9219 20267 9220
rect 20210 9200 20239 9219
rect 20182 9199 20239 9200
rect 20259 9199 20267 9219
rect 20125 9193 20162 9194
rect 20182 9193 20267 9199
rect 20333 9223 20371 9231
rect 20444 9227 20480 9228
rect 20333 9203 20342 9223
rect 20362 9203 20371 9223
rect 20333 9194 20371 9203
rect 20395 9219 20480 9227
rect 20395 9199 20452 9219
rect 20472 9199 20480 9219
rect 20333 9193 20370 9194
rect 20395 9193 20480 9199
rect 20546 9223 20584 9231
rect 20546 9203 20555 9223
rect 20575 9203 20584 9223
rect 20546 9194 20584 9203
rect 20633 9197 20697 9381
rect 20853 9255 20918 9456
rect 20853 9237 20875 9255
rect 20893 9237 20918 9255
rect 20853 9218 20918 9237
rect 20546 9193 20583 9194
rect 19969 9172 20005 9193
rect 20395 9172 20426 9193
rect 20633 9188 20641 9197
rect 20630 9172 20641 9188
rect 19802 9168 19902 9172
rect 19802 9164 19864 9168
rect 19802 9138 19809 9164
rect 19835 9142 19864 9164
rect 19890 9142 19902 9168
rect 19835 9138 19902 9142
rect 19802 9135 19902 9138
rect 19970 9135 20005 9172
rect 20067 9169 20426 9172
rect 20067 9164 20289 9169
rect 20067 9140 20080 9164
rect 20104 9145 20289 9164
rect 20313 9145 20426 9169
rect 20104 9140 20426 9145
rect 20067 9136 20426 9140
rect 20493 9164 20641 9172
rect 20493 9144 20504 9164
rect 20524 9155 20641 9164
rect 20690 9188 20697 9197
rect 20690 9155 20698 9188
rect 20524 9144 20698 9155
rect 20493 9137 20698 9144
rect 20493 9136 20534 9137
rect 19969 9110 20005 9135
rect 19817 9083 19854 9084
rect 19913 9083 19950 9084
rect 19969 9083 19976 9110
rect 19493 9058 19501 9078
rect 19521 9058 19530 9078
rect 19347 9047 19378 9048
rect 19342 8979 19452 8992
rect 19493 8979 19530 9058
rect 19717 9074 19855 9083
rect 19717 9054 19826 9074
rect 19846 9054 19855 9074
rect 19717 9047 19855 9054
rect 19913 9080 19976 9083
rect 19997 9083 20005 9110
rect 20024 9083 20061 9084
rect 19997 9080 20061 9083
rect 19913 9074 20061 9080
rect 19913 9054 19922 9074
rect 19942 9054 20032 9074
rect 20052 9054 20061 9074
rect 19717 9045 19813 9047
rect 19913 9044 20061 9054
rect 20120 9074 20157 9084
rect 20232 9083 20269 9084
rect 20213 9081 20269 9083
rect 20120 9054 20128 9074
rect 20148 9054 20157 9074
rect 19969 9043 20005 9044
rect 19280 8977 19530 8979
rect 19280 8974 19381 8977
rect 19280 8955 19345 8974
rect 19342 8947 19345 8955
rect 19374 8947 19381 8974
rect 19409 8950 19419 8977
rect 19448 8955 19530 8977
rect 19448 8950 19452 8955
rect 19409 8947 19452 8950
rect 19342 8933 19452 8947
rect 18768 8915 19109 8916
rect 18693 8910 19109 8915
rect 19817 8912 19854 8913
rect 20120 8912 20157 9054
rect 20182 9074 20269 9081
rect 20182 9071 20240 9074
rect 20182 9051 20187 9071
rect 20208 9054 20240 9071
rect 20260 9054 20269 9074
rect 20208 9051 20269 9054
rect 20182 9044 20269 9051
rect 20328 9074 20365 9084
rect 20328 9054 20336 9074
rect 20356 9054 20365 9074
rect 20182 9043 20213 9044
rect 20328 8975 20365 9054
rect 20395 9083 20426 9136
rect 20630 9134 20698 9137
rect 20630 9092 20642 9134
rect 20691 9092 20698 9134
rect 20445 9083 20482 9084
rect 20395 9074 20482 9083
rect 20395 9054 20453 9074
rect 20473 9054 20482 9074
rect 20395 9044 20482 9054
rect 20541 9074 20578 9084
rect 20630 9079 20698 9092
rect 20853 9156 20918 9173
rect 20853 9138 20877 9156
rect 20895 9138 20918 9156
rect 20541 9054 20549 9074
rect 20569 9054 20578 9074
rect 20395 9043 20426 9044
rect 20390 8975 20500 8988
rect 20541 8975 20578 9054
rect 20853 8999 20918 9138
rect 20853 8993 20875 8999
rect 20328 8973 20578 8975
rect 20328 8970 20429 8973
rect 20328 8951 20393 8970
rect 20390 8943 20393 8951
rect 20422 8943 20429 8970
rect 20457 8946 20467 8973
rect 20496 8951 20578 8973
rect 20607 8981 20875 8993
rect 20893 8981 20918 8999
rect 20607 8958 20918 8981
rect 20607 8957 20662 8958
rect 20496 8946 20500 8951
rect 20457 8943 20500 8946
rect 20390 8929 20500 8943
rect 19816 8911 20157 8912
rect 18693 8890 18696 8910
rect 18716 8890 19109 8910
rect 19741 8910 20157 8911
rect 20607 8910 20650 8957
rect 19741 8906 20650 8910
rect 19060 8857 19105 8890
rect 19741 8886 19744 8906
rect 19764 8886 20650 8906
rect 20118 8881 20650 8886
rect 20858 8900 20917 8922
rect 20858 8882 20877 8900
rect 20895 8882 20917 8900
rect 19906 8857 20005 8859
rect 19060 8847 20005 8857
rect 19060 8821 19928 8847
rect 19061 8820 19928 8821
rect 19906 8809 19928 8820
rect 19953 8812 19972 8847
rect 19997 8812 20005 8847
rect 19953 8809 20005 8812
rect 20858 8811 20917 8882
rect 19906 8801 20005 8809
rect 19932 8800 20004 8801
rect 19586 8774 19653 8793
rect 19586 8753 19603 8774
rect 18467 8575 18547 8617
rect 19584 8708 19603 8753
rect 19633 8753 19653 8774
rect 19633 8708 19654 8753
rect 20123 8750 20164 8752
rect 20395 8750 20499 8752
rect 20855 8750 20919 8811
rect 17528 8464 17564 8465
rect 17420 8456 17564 8464
rect 17420 8436 17428 8456
rect 17448 8436 17536 8456
rect 17556 8436 17564 8456
rect 17420 8430 17564 8436
rect 17630 8460 17668 8468
rect 17736 8464 17772 8465
rect 17630 8440 17639 8460
rect 17659 8440 17668 8460
rect 17630 8431 17668 8440
rect 17687 8457 17772 8464
rect 17687 8437 17694 8457
rect 17715 8456 17772 8457
rect 17715 8437 17744 8456
rect 17687 8436 17744 8437
rect 17764 8436 17772 8456
rect 17630 8430 17667 8431
rect 17687 8430 17772 8436
rect 17838 8460 17876 8468
rect 17949 8464 17985 8465
rect 17838 8440 17847 8460
rect 17867 8440 17876 8460
rect 17838 8431 17876 8440
rect 17900 8456 17985 8464
rect 17900 8436 17957 8456
rect 17977 8436 17985 8456
rect 17838 8430 17875 8431
rect 17900 8430 17985 8436
rect 18051 8460 18089 8468
rect 18051 8440 18060 8460
rect 18080 8440 18089 8460
rect 18051 8431 18089 8440
rect 18289 8448 18375 8484
rect 18051 8430 18088 8431
rect 17474 8409 17510 8430
rect 17900 8409 17931 8430
rect 18127 8409 18173 8413
rect 17307 8405 17407 8409
rect 17307 8401 17369 8405
rect 17307 8375 17314 8401
rect 17340 8379 17369 8401
rect 17395 8379 17407 8405
rect 17340 8375 17407 8379
rect 17307 8372 17407 8375
rect 17475 8372 17510 8409
rect 17572 8406 17931 8409
rect 17572 8401 17794 8406
rect 17572 8377 17585 8401
rect 17609 8382 17794 8401
rect 17818 8382 17931 8406
rect 17609 8377 17931 8382
rect 17572 8373 17931 8377
rect 17998 8401 18173 8409
rect 17998 8381 18009 8401
rect 18029 8381 18173 8401
rect 18289 8407 18306 8448
rect 18360 8407 18375 8448
rect 18289 8388 18375 8407
rect 17998 8374 18173 8381
rect 17998 8373 18039 8374
rect 17474 8347 17510 8372
rect 17322 8320 17359 8321
rect 17418 8320 17455 8321
rect 17474 8320 17481 8347
rect 17222 8311 17360 8320
rect 17222 8291 17331 8311
rect 17351 8291 17360 8311
rect 17222 8284 17360 8291
rect 17418 8317 17481 8320
rect 17502 8320 17510 8347
rect 17529 8320 17566 8321
rect 17502 8317 17566 8320
rect 17418 8311 17566 8317
rect 17418 8291 17427 8311
rect 17447 8291 17537 8311
rect 17557 8291 17566 8311
rect 17222 8282 17318 8284
rect 17418 8281 17566 8291
rect 17625 8311 17662 8321
rect 17737 8320 17774 8321
rect 17718 8318 17774 8320
rect 17625 8291 17633 8311
rect 17653 8291 17662 8311
rect 17474 8280 17510 8281
rect 17322 8149 17359 8150
rect 17625 8149 17662 8291
rect 17687 8311 17774 8318
rect 17687 8308 17745 8311
rect 17687 8288 17692 8308
rect 17713 8291 17745 8308
rect 17765 8291 17774 8311
rect 17713 8288 17774 8291
rect 17687 8281 17774 8288
rect 17833 8311 17870 8321
rect 17833 8291 17841 8311
rect 17861 8291 17870 8311
rect 17687 8280 17718 8281
rect 17833 8212 17870 8291
rect 17900 8320 17931 8373
rect 17950 8320 17987 8321
rect 17900 8311 17987 8320
rect 17900 8291 17958 8311
rect 17978 8291 17987 8311
rect 17900 8281 17987 8291
rect 18046 8311 18083 8321
rect 18046 8291 18054 8311
rect 18074 8291 18083 8311
rect 17900 8280 17931 8281
rect 17895 8212 18005 8225
rect 18046 8212 18083 8291
rect 18127 8291 18173 8374
rect 18467 8291 18542 8575
rect 19584 8500 19654 8708
rect 19716 8715 20919 8750
rect 19716 8701 19744 8715
rect 19718 8570 19744 8701
rect 20123 8712 20919 8715
rect 19576 8449 19656 8500
rect 19576 8423 19592 8449
rect 19632 8423 19656 8449
rect 19576 8404 19656 8423
rect 19576 8378 19595 8404
rect 19635 8378 19656 8404
rect 19576 8351 19656 8378
rect 19576 8325 19599 8351
rect 19639 8325 19656 8351
rect 19576 8314 19656 8325
rect 19718 8315 19745 8570
rect 20123 8562 20164 8712
rect 20395 8706 20499 8712
rect 20855 8709 20919 8712
rect 20590 8650 20711 8668
rect 20590 8648 20661 8650
rect 20590 8607 20605 8648
rect 20642 8609 20661 8648
rect 20698 8609 20711 8650
rect 20642 8607 20711 8609
rect 20590 8597 20711 8607
rect 19785 8455 19849 8467
rect 20125 8463 20162 8562
rect 20390 8552 20501 8565
rect 20390 8550 20432 8552
rect 20390 8530 20397 8550
rect 20416 8530 20432 8550
rect 20390 8522 20432 8530
rect 20460 8550 20501 8552
rect 20460 8530 20474 8550
rect 20493 8530 20501 8550
rect 20460 8522 20501 8530
rect 20390 8516 20501 8522
rect 20333 8494 20582 8516
rect 20333 8463 20370 8494
rect 20546 8492 20582 8494
rect 20546 8463 20583 8492
rect 19785 8454 19820 8455
rect 19762 8449 19820 8454
rect 19762 8429 19765 8449
rect 19785 8435 19820 8449
rect 19840 8435 19849 8455
rect 19785 8427 19849 8435
rect 19811 8426 19849 8427
rect 19812 8425 19849 8426
rect 19915 8459 19951 8460
rect 20023 8459 20059 8460
rect 19915 8451 20059 8459
rect 19915 8431 19923 8451
rect 19943 8431 20031 8451
rect 20051 8431 20059 8451
rect 19915 8425 20059 8431
rect 20125 8455 20163 8463
rect 20231 8459 20267 8460
rect 20125 8435 20134 8455
rect 20154 8435 20163 8455
rect 20125 8426 20163 8435
rect 20182 8452 20267 8459
rect 20182 8432 20189 8452
rect 20210 8451 20267 8452
rect 20210 8432 20239 8451
rect 20182 8431 20239 8432
rect 20259 8431 20267 8451
rect 20125 8425 20162 8426
rect 20182 8425 20267 8431
rect 20333 8455 20371 8463
rect 20444 8459 20480 8460
rect 20333 8435 20342 8455
rect 20362 8435 20371 8455
rect 20333 8426 20371 8435
rect 20395 8451 20480 8459
rect 20395 8431 20452 8451
rect 20472 8431 20480 8451
rect 20333 8425 20370 8426
rect 20395 8425 20480 8431
rect 20546 8455 20584 8463
rect 20546 8435 20555 8455
rect 20575 8435 20584 8455
rect 20639 8445 20704 8597
rect 20857 8571 20912 8709
rect 20546 8426 20584 8435
rect 20637 8438 20704 8445
rect 20546 8425 20583 8426
rect 19969 8404 20005 8425
rect 20395 8404 20426 8425
rect 20637 8417 20654 8438
rect 20690 8417 20704 8438
rect 20856 8458 20912 8571
rect 20856 8440 20875 8458
rect 20893 8440 20912 8458
rect 20856 8420 20912 8440
rect 20637 8404 20704 8417
rect 19802 8400 19902 8404
rect 19802 8396 19864 8400
rect 19802 8370 19809 8396
rect 19835 8374 19864 8396
rect 19890 8374 19902 8400
rect 19835 8370 19902 8374
rect 19802 8367 19902 8370
rect 19970 8367 20005 8404
rect 20067 8401 20426 8404
rect 20067 8396 20289 8401
rect 20067 8372 20080 8396
rect 20104 8377 20289 8396
rect 20313 8377 20426 8401
rect 20104 8372 20426 8377
rect 20067 8368 20426 8372
rect 20493 8398 20704 8404
rect 20493 8396 20654 8398
rect 20493 8376 20504 8396
rect 20524 8376 20654 8396
rect 20493 8369 20654 8376
rect 20493 8368 20534 8369
rect 19969 8342 20005 8367
rect 19817 8315 19854 8316
rect 19913 8315 19950 8316
rect 19969 8315 19976 8342
rect 18127 8256 18542 8291
rect 19717 8306 19855 8315
rect 19717 8286 19826 8306
rect 19846 8286 19855 8306
rect 19717 8279 19855 8286
rect 19913 8312 19976 8315
rect 19997 8315 20005 8342
rect 20024 8315 20061 8316
rect 19997 8312 20061 8315
rect 19913 8306 20061 8312
rect 19913 8286 19922 8306
rect 19942 8286 20032 8306
rect 20052 8286 20061 8306
rect 19717 8277 19813 8279
rect 19913 8276 20061 8286
rect 20120 8306 20157 8316
rect 20232 8315 20269 8316
rect 20213 8313 20269 8315
rect 20120 8286 20128 8306
rect 20148 8286 20157 8306
rect 19969 8275 20005 8276
rect 18127 8255 18173 8256
rect 17833 8210 18083 8212
rect 17833 8207 17934 8210
rect 17833 8188 17898 8207
rect 17895 8180 17898 8188
rect 17927 8180 17934 8207
rect 17962 8183 17972 8210
rect 18001 8188 18083 8210
rect 18467 8204 18542 8256
rect 18001 8183 18005 8188
rect 17962 8180 18005 8183
rect 17895 8166 18005 8180
rect 17321 8148 17662 8149
rect 17246 8143 17662 8148
rect 17246 8123 17249 8143
rect 17269 8123 17663 8143
rect 16303 7476 17109 7551
rect 15542 7432 15551 7466
rect 15580 7465 15990 7466
rect 15580 7432 15597 7465
rect 15822 7464 15990 7465
rect 15542 7406 15597 7432
rect 15542 7372 15550 7406
rect 15579 7372 15597 7406
rect 15542 7360 15597 7372
rect 13738 7315 13822 7336
rect 13738 7287 13766 7315
rect 13810 7287 13822 7315
rect 13552 7236 13626 7264
rect 13552 7188 13575 7236
rect 13612 7188 13626 7236
rect 13738 7258 13822 7287
rect 13738 7230 13763 7258
rect 13807 7230 13822 7258
rect 13738 7205 13822 7230
rect 15878 7219 15966 7223
rect 13552 7179 13626 7188
rect 8872 7112 8944 7134
rect 9005 7127 10208 7162
rect 9005 7113 9033 7127
rect 8873 6912 8943 7112
rect 9007 6982 9033 7113
rect 9412 7124 10208 7127
rect 8865 6861 8945 6912
rect 8865 6835 8881 6861
rect 8921 6835 8945 6861
rect 8865 6816 8945 6835
rect 8865 6790 8884 6816
rect 8924 6790 8945 6816
rect 8865 6763 8945 6790
rect 8865 6737 8888 6763
rect 8928 6737 8945 6763
rect 8865 6726 8945 6737
rect 9007 6727 9034 6982
rect 9412 6974 9453 7124
rect 9684 7122 9788 7124
rect 10143 7090 10208 7124
rect 11185 7129 11251 7177
rect 13562 7175 13626 7179
rect 15878 7202 16142 7219
rect 15878 7148 16058 7202
rect 16121 7148 16142 7202
rect 13775 7138 14486 7140
rect 13148 7137 14486 7138
rect 12098 7136 12170 7137
rect 9879 7062 10000 7080
rect 9879 7060 9950 7062
rect 9879 7019 9894 7060
rect 9931 7021 9950 7060
rect 9987 7021 10000 7062
rect 9931 7019 10000 7021
rect 9879 7009 10000 7019
rect 9684 6979 9788 6982
rect 9074 6867 9138 6879
rect 9414 6875 9451 6974
rect 9679 6964 9790 6979
rect 9679 6962 9721 6964
rect 9679 6942 9686 6962
rect 9705 6942 9721 6962
rect 9679 6934 9721 6942
rect 9749 6962 9790 6964
rect 9749 6942 9763 6962
rect 9782 6942 9790 6962
rect 9749 6934 9790 6942
rect 9679 6928 9790 6934
rect 9622 6906 9871 6928
rect 9622 6875 9659 6906
rect 9835 6904 9871 6906
rect 9835 6875 9872 6904
rect 9074 6866 9109 6867
rect 9051 6861 9109 6866
rect 9051 6841 9054 6861
rect 9074 6847 9109 6861
rect 9129 6847 9138 6867
rect 9074 6839 9138 6847
rect 9100 6838 9138 6839
rect 9101 6837 9138 6838
rect 9204 6871 9240 6872
rect 9312 6871 9348 6872
rect 9204 6863 9348 6871
rect 9204 6843 9212 6863
rect 9232 6843 9320 6863
rect 9340 6843 9348 6863
rect 9204 6837 9348 6843
rect 9414 6867 9452 6875
rect 9520 6871 9556 6872
rect 9414 6847 9423 6867
rect 9443 6847 9452 6867
rect 9414 6838 9452 6847
rect 9471 6864 9556 6871
rect 9471 6844 9478 6864
rect 9499 6863 9556 6864
rect 9499 6844 9528 6863
rect 9471 6843 9528 6844
rect 9548 6843 9556 6863
rect 9414 6837 9451 6838
rect 9471 6837 9556 6843
rect 9622 6867 9660 6875
rect 9733 6871 9769 6872
rect 9622 6847 9631 6867
rect 9651 6847 9660 6867
rect 9622 6838 9660 6847
rect 9684 6863 9769 6871
rect 9684 6843 9741 6863
rect 9761 6843 9769 6863
rect 9622 6837 9659 6838
rect 9684 6837 9769 6843
rect 9835 6867 9873 6875
rect 9835 6847 9844 6867
rect 9864 6847 9873 6867
rect 9928 6857 9993 7009
rect 10146 6983 10201 7090
rect 11185 7055 11244 7129
rect 12097 7128 12196 7136
rect 12097 7125 12149 7128
rect 12097 7090 12105 7125
rect 12130 7090 12149 7125
rect 12174 7117 12196 7128
rect 13147 7129 14486 7137
rect 13147 7126 13199 7129
rect 12174 7116 13041 7117
rect 12174 7090 13042 7116
rect 12097 7080 13042 7090
rect 12097 7078 12196 7080
rect 11185 7037 11207 7055
rect 11225 7037 11244 7055
rect 11185 7015 11244 7037
rect 11452 7051 11984 7056
rect 11452 7031 12338 7051
rect 12358 7031 12361 7051
rect 12997 7047 13042 7080
rect 13147 7091 13155 7126
rect 13180 7091 13199 7126
rect 13224 7091 14486 7129
rect 13147 7082 14486 7091
rect 13147 7079 13236 7082
rect 13775 7080 14486 7082
rect 15878 7131 16142 7148
rect 11452 7027 12361 7031
rect 9835 6838 9873 6847
rect 9926 6850 9993 6857
rect 9835 6837 9872 6838
rect 9258 6816 9294 6837
rect 9684 6816 9715 6837
rect 9926 6829 9943 6850
rect 9979 6829 9993 6850
rect 10145 6870 10201 6983
rect 11452 6980 11495 7027
rect 11945 7026 12361 7027
rect 12993 7027 13386 7047
rect 13406 7027 13409 7047
rect 11945 7025 12286 7026
rect 11602 6994 11712 7008
rect 11602 6991 11645 6994
rect 11602 6986 11606 6991
rect 11440 6979 11495 6980
rect 10145 6852 10164 6870
rect 10182 6852 10201 6870
rect 10145 6832 10201 6852
rect 11184 6956 11495 6979
rect 11184 6938 11209 6956
rect 11227 6944 11495 6956
rect 11524 6964 11606 6986
rect 11635 6964 11645 6991
rect 11673 6967 11680 6994
rect 11709 6986 11712 6994
rect 11709 6967 11774 6986
rect 11673 6964 11774 6967
rect 11524 6962 11774 6964
rect 11227 6938 11249 6944
rect 9926 6816 9993 6829
rect 9091 6812 9191 6816
rect 9091 6808 9153 6812
rect 9091 6782 9098 6808
rect 9124 6786 9153 6808
rect 9179 6786 9191 6812
rect 9124 6782 9191 6786
rect 9091 6779 9191 6782
rect 9259 6779 9294 6816
rect 9356 6813 9715 6816
rect 9356 6808 9578 6813
rect 9356 6784 9369 6808
rect 9393 6789 9578 6808
rect 9602 6789 9715 6813
rect 9393 6784 9715 6789
rect 9356 6780 9715 6784
rect 9782 6810 9993 6816
rect 9782 6808 9943 6810
rect 9782 6788 9793 6808
rect 9813 6788 9943 6808
rect 9782 6781 9943 6788
rect 9782 6780 9823 6781
rect 9258 6754 9294 6779
rect 9106 6727 9143 6728
rect 9202 6727 9239 6728
rect 9258 6727 9265 6754
rect 9006 6718 9144 6727
rect 9006 6698 9115 6718
rect 9135 6698 9144 6718
rect 9006 6691 9144 6698
rect 9202 6724 9265 6727
rect 9286 6727 9294 6754
rect 9313 6727 9350 6728
rect 9286 6724 9350 6727
rect 9202 6718 9350 6724
rect 9202 6698 9211 6718
rect 9231 6698 9321 6718
rect 9341 6698 9350 6718
rect 9006 6689 9102 6691
rect 9202 6688 9350 6698
rect 9409 6718 9446 6728
rect 9521 6727 9558 6728
rect 9502 6725 9558 6727
rect 9409 6698 9417 6718
rect 9437 6698 9446 6718
rect 9258 6687 9294 6688
rect 9106 6556 9143 6557
rect 9409 6556 9446 6698
rect 9471 6718 9558 6725
rect 9471 6715 9529 6718
rect 9471 6695 9476 6715
rect 9497 6698 9529 6715
rect 9549 6698 9558 6718
rect 9497 6695 9558 6698
rect 9471 6688 9558 6695
rect 9617 6718 9654 6728
rect 9617 6698 9625 6718
rect 9645 6698 9654 6718
rect 9471 6687 9502 6688
rect 9617 6619 9654 6698
rect 9684 6727 9715 6780
rect 9928 6773 9943 6781
rect 9983 6773 9993 6810
rect 11184 6799 11249 6938
rect 11524 6883 11561 6962
rect 11602 6949 11712 6962
rect 11676 6893 11707 6894
rect 11524 6863 11533 6883
rect 11553 6863 11561 6883
rect 9928 6764 9993 6773
rect 10141 6771 10206 6792
rect 10141 6753 10166 6771
rect 10184 6753 10206 6771
rect 11184 6781 11207 6799
rect 11225 6781 11249 6799
rect 11184 6764 11249 6781
rect 11404 6845 11472 6858
rect 11524 6853 11561 6863
rect 11620 6883 11707 6893
rect 11620 6863 11629 6883
rect 11649 6863 11707 6883
rect 11620 6854 11707 6863
rect 11620 6853 11657 6854
rect 11404 6803 11411 6845
rect 11460 6803 11472 6845
rect 11404 6800 11472 6803
rect 11676 6801 11707 6854
rect 11737 6883 11774 6962
rect 11889 6893 11920 6894
rect 11737 6863 11746 6883
rect 11766 6863 11774 6883
rect 11737 6853 11774 6863
rect 11833 6886 11920 6893
rect 11833 6883 11894 6886
rect 11833 6863 11842 6883
rect 11862 6866 11894 6883
rect 11915 6866 11920 6886
rect 11862 6863 11920 6866
rect 11833 6856 11920 6863
rect 11945 6883 11982 7025
rect 12248 7024 12285 7025
rect 12993 7022 13409 7027
rect 12993 7021 13334 7022
rect 12650 6990 12760 7004
rect 12650 6987 12693 6990
rect 12650 6982 12654 6987
rect 12572 6960 12654 6982
rect 12683 6960 12693 6987
rect 12721 6963 12728 6990
rect 12757 6982 12760 6990
rect 12757 6963 12822 6982
rect 12721 6960 12822 6963
rect 12572 6958 12822 6960
rect 12097 6893 12133 6894
rect 11945 6863 11954 6883
rect 11974 6863 11982 6883
rect 11833 6854 11889 6856
rect 11833 6853 11870 6854
rect 11945 6853 11982 6863
rect 12041 6883 12189 6893
rect 12289 6890 12385 6892
rect 12041 6863 12050 6883
rect 12070 6863 12160 6883
rect 12180 6863 12189 6883
rect 12041 6857 12189 6863
rect 12041 6854 12105 6857
rect 12041 6853 12078 6854
rect 12097 6827 12105 6854
rect 12126 6854 12189 6857
rect 12247 6883 12385 6890
rect 12247 6863 12256 6883
rect 12276 6863 12385 6883
rect 12247 6854 12385 6863
rect 12572 6879 12609 6958
rect 12650 6945 12760 6958
rect 12724 6889 12755 6890
rect 12572 6859 12581 6879
rect 12601 6859 12609 6879
rect 12126 6827 12133 6854
rect 12152 6853 12189 6854
rect 12248 6853 12285 6854
rect 12097 6802 12133 6827
rect 11568 6800 11609 6801
rect 11404 6793 11609 6800
rect 11404 6782 11578 6793
rect 9734 6727 9771 6728
rect 9684 6718 9771 6727
rect 9684 6698 9742 6718
rect 9762 6698 9771 6718
rect 9684 6688 9771 6698
rect 9830 6718 9867 6728
rect 9830 6698 9838 6718
rect 9858 6698 9867 6718
rect 9684 6687 9715 6688
rect 9679 6619 9789 6632
rect 9830 6619 9867 6698
rect 10141 6677 10206 6753
rect 11404 6749 11412 6782
rect 11405 6740 11412 6749
rect 11461 6773 11578 6782
rect 11598 6773 11609 6793
rect 11461 6765 11609 6773
rect 11676 6797 12035 6801
rect 11676 6792 11998 6797
rect 11676 6768 11789 6792
rect 11813 6773 11998 6792
rect 12022 6773 12035 6797
rect 11813 6768 12035 6773
rect 11676 6765 12035 6768
rect 12097 6765 12132 6802
rect 12200 6799 12300 6802
rect 12200 6795 12267 6799
rect 12200 6769 12212 6795
rect 12238 6773 12267 6795
rect 12293 6773 12300 6799
rect 12238 6769 12300 6773
rect 12200 6765 12300 6769
rect 11461 6749 11472 6765
rect 11461 6740 11469 6749
rect 11676 6744 11707 6765
rect 12097 6744 12133 6765
rect 11519 6743 11556 6744
rect 11184 6700 11249 6719
rect 11184 6682 11209 6700
rect 11227 6682 11249 6700
rect 9617 6617 9867 6619
rect 9617 6614 9718 6617
rect 9617 6595 9682 6614
rect 9679 6587 9682 6595
rect 9711 6587 9718 6614
rect 9746 6590 9756 6617
rect 9785 6595 9867 6617
rect 9890 6642 10207 6677
rect 9785 6590 9789 6595
rect 9746 6587 9789 6590
rect 9679 6573 9789 6587
rect 9105 6555 9446 6556
rect 9030 6553 9446 6555
rect 9890 6553 9930 6642
rect 10141 6615 10206 6642
rect 10141 6597 10164 6615
rect 10182 6597 10206 6615
rect 10141 6577 10206 6597
rect 9027 6550 9930 6553
rect 9027 6530 9033 6550
rect 9053 6530 9930 6550
rect 9027 6526 9930 6530
rect 9890 6523 9930 6526
rect 10142 6516 10207 6537
rect 8360 6508 9021 6509
rect 8360 6501 9294 6508
rect 8360 6500 9266 6501
rect 8360 6480 9211 6500
rect 9243 6481 9266 6500
rect 9291 6481 9294 6501
rect 9243 6480 9294 6481
rect 8360 6473 9294 6480
rect 7959 6431 8127 6432
rect 8362 6431 8401 6473
rect 9190 6471 9294 6473
rect 9259 6469 9294 6471
rect 10142 6498 10166 6516
rect 10184 6498 10207 6516
rect 10142 6451 10207 6498
rect 7959 6405 8403 6431
rect 7959 6403 8127 6405
rect 7959 6052 7986 6403
rect 8362 6399 8403 6405
rect 8026 6192 8090 6204
rect 8366 6200 8403 6399
rect 8865 6426 8937 6443
rect 8865 6387 8873 6426
rect 8918 6387 8937 6426
rect 8631 6289 8742 6304
rect 8631 6287 8673 6289
rect 8631 6267 8638 6287
rect 8657 6267 8673 6287
rect 8631 6259 8673 6267
rect 8701 6287 8742 6289
rect 8701 6267 8715 6287
rect 8734 6267 8742 6287
rect 8701 6259 8742 6267
rect 8631 6253 8742 6259
rect 8574 6231 8823 6253
rect 8574 6200 8611 6231
rect 8787 6229 8823 6231
rect 8787 6200 8824 6229
rect 8026 6191 8061 6192
rect 8003 6186 8061 6191
rect 8003 6166 8006 6186
rect 8026 6172 8061 6186
rect 8081 6172 8090 6192
rect 8026 6164 8090 6172
rect 8052 6163 8090 6164
rect 8053 6162 8090 6163
rect 8156 6196 8192 6197
rect 8264 6196 8300 6197
rect 8156 6188 8300 6196
rect 8156 6168 8164 6188
rect 8184 6168 8272 6188
rect 8292 6168 8300 6188
rect 8156 6162 8300 6168
rect 8366 6192 8404 6200
rect 8472 6196 8508 6197
rect 8366 6172 8375 6192
rect 8395 6172 8404 6192
rect 8366 6163 8404 6172
rect 8423 6189 8508 6196
rect 8423 6169 8430 6189
rect 8451 6188 8508 6189
rect 8451 6169 8480 6188
rect 8423 6168 8480 6169
rect 8500 6168 8508 6188
rect 8366 6162 8403 6163
rect 8423 6162 8508 6168
rect 8574 6192 8612 6200
rect 8685 6196 8721 6197
rect 8574 6172 8583 6192
rect 8603 6172 8612 6192
rect 8574 6163 8612 6172
rect 8636 6188 8721 6196
rect 8636 6168 8693 6188
rect 8713 6168 8721 6188
rect 8574 6162 8611 6163
rect 8636 6162 8721 6168
rect 8787 6192 8825 6200
rect 8787 6172 8796 6192
rect 8816 6172 8825 6192
rect 8787 6163 8825 6172
rect 8865 6177 8937 6387
rect 9007 6421 10207 6451
rect 9007 6420 9451 6421
rect 9007 6418 9175 6420
rect 8865 6163 8948 6177
rect 8787 6162 8824 6163
rect 8210 6141 8246 6162
rect 8636 6141 8667 6162
rect 8865 6141 8882 6163
rect 8043 6137 8143 6141
rect 8043 6133 8105 6137
rect 8043 6107 8050 6133
rect 8076 6111 8105 6133
rect 8131 6111 8143 6137
rect 8076 6107 8143 6111
rect 8043 6104 8143 6107
rect 8211 6104 8246 6141
rect 8308 6138 8667 6141
rect 8308 6133 8530 6138
rect 8308 6109 8321 6133
rect 8345 6114 8530 6133
rect 8554 6114 8667 6138
rect 8345 6109 8667 6114
rect 8308 6105 8667 6109
rect 8734 6133 8882 6141
rect 8734 6113 8745 6133
rect 8765 6130 8882 6133
rect 8935 6130 8948 6163
rect 8765 6113 8948 6130
rect 8734 6106 8948 6113
rect 8734 6105 8775 6106
rect 8865 6105 8948 6106
rect 8210 6079 8246 6104
rect 8058 6052 8095 6053
rect 8154 6052 8191 6053
rect 8210 6052 8217 6079
rect 7958 6043 8096 6052
rect 7958 6023 8067 6043
rect 8087 6023 8096 6043
rect 7958 6016 8096 6023
rect 8154 6049 8217 6052
rect 8238 6052 8246 6079
rect 8265 6052 8302 6053
rect 8238 6049 8302 6052
rect 8154 6043 8302 6049
rect 8154 6023 8163 6043
rect 8183 6023 8273 6043
rect 8293 6023 8302 6043
rect 7958 6014 8054 6016
rect 8154 6013 8302 6023
rect 8361 6043 8398 6053
rect 8473 6052 8510 6053
rect 8454 6050 8510 6052
rect 8361 6023 8369 6043
rect 8389 6023 8398 6043
rect 8210 6012 8246 6013
rect 8058 5881 8095 5882
rect 8361 5881 8398 6023
rect 8423 6043 8510 6050
rect 8423 6040 8481 6043
rect 8423 6020 8428 6040
rect 8449 6023 8481 6040
rect 8501 6023 8510 6043
rect 8449 6020 8510 6023
rect 8423 6013 8510 6020
rect 8569 6043 8606 6053
rect 8569 6023 8577 6043
rect 8597 6023 8606 6043
rect 8423 6012 8454 6013
rect 8569 5944 8606 6023
rect 8636 6052 8667 6105
rect 8873 6072 8887 6105
rect 8940 6072 8948 6105
rect 8873 6066 8948 6072
rect 8873 6061 8943 6066
rect 8686 6052 8723 6053
rect 8636 6043 8723 6052
rect 8636 6023 8694 6043
rect 8714 6023 8723 6043
rect 8636 6013 8723 6023
rect 8782 6043 8819 6053
rect 9007 6048 9034 6418
rect 9074 6188 9138 6200
rect 9414 6196 9451 6420
rect 9922 6401 9986 6403
rect 9918 6389 9986 6401
rect 9918 6356 9929 6389
rect 9969 6356 9986 6389
rect 9918 6346 9986 6356
rect 9679 6285 9790 6300
rect 9679 6283 9721 6285
rect 9679 6263 9686 6283
rect 9705 6263 9721 6283
rect 9679 6255 9721 6263
rect 9749 6283 9790 6285
rect 9749 6263 9763 6283
rect 9782 6263 9790 6283
rect 9749 6255 9790 6263
rect 9679 6249 9790 6255
rect 9622 6227 9871 6249
rect 9622 6196 9659 6227
rect 9835 6225 9871 6227
rect 9835 6196 9872 6225
rect 9074 6187 9109 6188
rect 9051 6182 9109 6187
rect 9051 6162 9054 6182
rect 9074 6168 9109 6182
rect 9129 6168 9138 6188
rect 9074 6160 9138 6168
rect 9100 6159 9138 6160
rect 9101 6158 9138 6159
rect 9204 6192 9240 6193
rect 9312 6192 9348 6193
rect 9204 6184 9348 6192
rect 9204 6164 9212 6184
rect 9232 6164 9320 6184
rect 9340 6164 9348 6184
rect 9204 6158 9348 6164
rect 9414 6188 9452 6196
rect 9520 6192 9556 6193
rect 9414 6168 9423 6188
rect 9443 6168 9452 6188
rect 9414 6159 9452 6168
rect 9471 6185 9556 6192
rect 9471 6165 9478 6185
rect 9499 6184 9556 6185
rect 9499 6165 9528 6184
rect 9471 6164 9528 6165
rect 9548 6164 9556 6184
rect 9414 6158 9451 6159
rect 9471 6158 9556 6164
rect 9622 6188 9660 6196
rect 9733 6192 9769 6193
rect 9622 6168 9631 6188
rect 9651 6168 9660 6188
rect 9622 6159 9660 6168
rect 9684 6184 9769 6192
rect 9684 6164 9741 6184
rect 9761 6164 9769 6184
rect 9622 6158 9659 6159
rect 9684 6158 9769 6164
rect 9835 6188 9873 6196
rect 9835 6168 9844 6188
rect 9864 6168 9873 6188
rect 9835 6159 9873 6168
rect 9922 6162 9986 6346
rect 10142 6220 10207 6421
rect 11184 6481 11249 6682
rect 11405 6556 11469 6740
rect 11518 6734 11556 6743
rect 11518 6714 11527 6734
rect 11547 6714 11556 6734
rect 11518 6706 11556 6714
rect 11622 6738 11707 6744
rect 11732 6743 11769 6744
rect 11622 6718 11630 6738
rect 11650 6718 11707 6738
rect 11622 6710 11707 6718
rect 11731 6734 11769 6743
rect 11731 6714 11740 6734
rect 11760 6714 11769 6734
rect 11622 6709 11658 6710
rect 11731 6706 11769 6714
rect 11835 6738 11920 6744
rect 11940 6743 11977 6744
rect 11835 6718 11843 6738
rect 11863 6737 11920 6738
rect 11863 6718 11892 6737
rect 11835 6717 11892 6718
rect 11913 6717 11920 6737
rect 11835 6710 11920 6717
rect 11939 6734 11977 6743
rect 11939 6714 11948 6734
rect 11968 6714 11977 6734
rect 11835 6709 11871 6710
rect 11939 6706 11977 6714
rect 12043 6738 12187 6744
rect 12043 6718 12051 6738
rect 12071 6718 12159 6738
rect 12179 6718 12187 6738
rect 12043 6710 12187 6718
rect 12043 6709 12079 6710
rect 12151 6709 12187 6710
rect 12253 6743 12290 6744
rect 12253 6742 12291 6743
rect 12253 6734 12317 6742
rect 12253 6714 12262 6734
rect 12282 6720 12317 6734
rect 12337 6720 12340 6740
rect 12282 6715 12340 6720
rect 12282 6714 12317 6715
rect 11519 6677 11556 6706
rect 11520 6675 11556 6677
rect 11732 6675 11769 6706
rect 11520 6653 11769 6675
rect 11601 6647 11712 6653
rect 11601 6639 11642 6647
rect 11601 6619 11609 6639
rect 11628 6619 11642 6639
rect 11601 6617 11642 6619
rect 11670 6639 11712 6647
rect 11670 6619 11686 6639
rect 11705 6619 11712 6639
rect 11670 6617 11712 6619
rect 11601 6602 11712 6617
rect 11405 6546 11473 6556
rect 11405 6513 11422 6546
rect 11462 6513 11473 6546
rect 11405 6501 11473 6513
rect 11405 6499 11469 6501
rect 11940 6482 11977 6706
rect 12253 6702 12317 6714
rect 12357 6484 12384 6854
rect 12572 6849 12609 6859
rect 12668 6879 12755 6889
rect 12668 6859 12677 6879
rect 12697 6859 12755 6879
rect 12668 6850 12755 6859
rect 12668 6849 12705 6850
rect 12448 6836 12518 6841
rect 12443 6830 12518 6836
rect 12443 6797 12451 6830
rect 12504 6797 12518 6830
rect 12724 6797 12755 6850
rect 12785 6879 12822 6958
rect 12937 6889 12968 6890
rect 12785 6859 12794 6879
rect 12814 6859 12822 6879
rect 12785 6849 12822 6859
rect 12881 6882 12968 6889
rect 12881 6879 12942 6882
rect 12881 6859 12890 6879
rect 12910 6862 12942 6879
rect 12963 6862 12968 6882
rect 12910 6859 12968 6862
rect 12881 6852 12968 6859
rect 12993 6879 13030 7021
rect 13296 7020 13333 7021
rect 13145 6889 13181 6890
rect 12993 6859 13002 6879
rect 13022 6859 13030 6879
rect 12881 6850 12937 6852
rect 12881 6849 12918 6850
rect 12993 6849 13030 6859
rect 13089 6879 13237 6889
rect 13337 6886 13433 6888
rect 13089 6859 13098 6879
rect 13118 6859 13208 6879
rect 13228 6859 13237 6879
rect 13089 6853 13237 6859
rect 13089 6850 13153 6853
rect 13089 6849 13126 6850
rect 13145 6823 13153 6850
rect 13174 6850 13237 6853
rect 13295 6879 13433 6886
rect 13295 6859 13304 6879
rect 13324 6859 13433 6879
rect 13295 6850 13433 6859
rect 13174 6823 13181 6850
rect 13200 6849 13237 6850
rect 13296 6849 13333 6850
rect 13145 6798 13181 6823
rect 12443 6796 12526 6797
rect 12616 6796 12657 6797
rect 12443 6789 12657 6796
rect 12443 6772 12626 6789
rect 12443 6739 12456 6772
rect 12509 6769 12626 6772
rect 12646 6769 12657 6789
rect 12509 6761 12657 6769
rect 12724 6793 13083 6797
rect 12724 6788 13046 6793
rect 12724 6764 12837 6788
rect 12861 6769 13046 6788
rect 13070 6769 13083 6793
rect 12861 6764 13083 6769
rect 12724 6761 13083 6764
rect 13145 6761 13180 6798
rect 13248 6795 13348 6798
rect 13248 6791 13315 6795
rect 13248 6765 13260 6791
rect 13286 6769 13315 6791
rect 13341 6769 13348 6795
rect 13286 6765 13348 6769
rect 13248 6761 13348 6765
rect 12509 6739 12526 6761
rect 12724 6740 12755 6761
rect 13145 6740 13181 6761
rect 12567 6739 12604 6740
rect 12443 6725 12526 6739
rect 12216 6482 12384 6484
rect 11940 6481 12384 6482
rect 11184 6451 12384 6481
rect 12454 6515 12526 6725
rect 12566 6730 12604 6739
rect 12566 6710 12575 6730
rect 12595 6710 12604 6730
rect 12566 6702 12604 6710
rect 12670 6734 12755 6740
rect 12780 6739 12817 6740
rect 12670 6714 12678 6734
rect 12698 6714 12755 6734
rect 12670 6706 12755 6714
rect 12779 6730 12817 6739
rect 12779 6710 12788 6730
rect 12808 6710 12817 6730
rect 12670 6705 12706 6706
rect 12779 6702 12817 6710
rect 12883 6734 12968 6740
rect 12988 6739 13025 6740
rect 12883 6714 12891 6734
rect 12911 6733 12968 6734
rect 12911 6714 12940 6733
rect 12883 6713 12940 6714
rect 12961 6713 12968 6733
rect 12883 6706 12968 6713
rect 12987 6730 13025 6739
rect 12987 6710 12996 6730
rect 13016 6710 13025 6730
rect 12883 6705 12919 6706
rect 12987 6702 13025 6710
rect 13091 6734 13235 6740
rect 13091 6714 13099 6734
rect 13119 6714 13207 6734
rect 13227 6714 13235 6734
rect 13091 6706 13235 6714
rect 13091 6705 13127 6706
rect 13199 6705 13235 6706
rect 13301 6739 13338 6740
rect 13301 6738 13339 6739
rect 13301 6730 13365 6738
rect 13301 6710 13310 6730
rect 13330 6716 13365 6730
rect 13385 6716 13388 6736
rect 13330 6711 13388 6716
rect 13330 6710 13365 6711
rect 12567 6673 12604 6702
rect 12568 6671 12604 6673
rect 12780 6671 12817 6702
rect 12568 6649 12817 6671
rect 12649 6643 12760 6649
rect 12649 6635 12690 6643
rect 12649 6615 12657 6635
rect 12676 6615 12690 6635
rect 12649 6613 12690 6615
rect 12718 6635 12760 6643
rect 12718 6615 12734 6635
rect 12753 6615 12760 6635
rect 12718 6613 12760 6615
rect 12649 6598 12760 6613
rect 12454 6476 12473 6515
rect 12518 6476 12526 6515
rect 12454 6459 12526 6476
rect 12988 6503 13025 6702
rect 13301 6698 13365 6710
rect 12988 6497 13029 6503
rect 13405 6499 13432 6850
rect 13727 6837 13822 6863
rect 13563 6815 13627 6834
rect 13563 6776 13576 6815
rect 13610 6776 13627 6815
rect 13563 6757 13627 6776
rect 13264 6497 13432 6499
rect 12988 6471 13432 6497
rect 11184 6404 11249 6451
rect 11184 6386 11207 6404
rect 11225 6386 11249 6404
rect 12097 6431 12132 6433
rect 12097 6429 12201 6431
rect 12990 6429 13029 6471
rect 13264 6470 13432 6471
rect 12097 6422 13031 6429
rect 12097 6421 12148 6422
rect 12097 6401 12100 6421
rect 12125 6402 12148 6421
rect 12180 6402 13031 6422
rect 12125 6401 13031 6402
rect 12097 6394 13031 6401
rect 12370 6393 13031 6394
rect 11184 6365 11249 6386
rect 11461 6376 11501 6379
rect 11461 6372 12364 6376
rect 11461 6352 12338 6372
rect 12358 6352 12364 6372
rect 11461 6349 12364 6352
rect 11185 6305 11250 6325
rect 11185 6287 11209 6305
rect 11227 6287 11250 6305
rect 11185 6260 11250 6287
rect 11461 6260 11501 6349
rect 11945 6347 12361 6349
rect 11945 6346 12286 6347
rect 11602 6315 11712 6329
rect 11602 6312 11645 6315
rect 11602 6307 11606 6312
rect 11184 6225 11501 6260
rect 11524 6285 11606 6307
rect 11635 6285 11645 6312
rect 11673 6288 11680 6315
rect 11709 6307 11712 6315
rect 11709 6288 11774 6307
rect 11673 6285 11774 6288
rect 11524 6283 11774 6285
rect 10142 6202 10164 6220
rect 10182 6202 10207 6220
rect 10142 6183 10207 6202
rect 9835 6158 9872 6159
rect 9258 6137 9294 6158
rect 9684 6137 9715 6158
rect 9922 6153 9930 6162
rect 9919 6137 9930 6153
rect 9091 6133 9191 6137
rect 9091 6129 9153 6133
rect 9091 6103 9098 6129
rect 9124 6107 9153 6129
rect 9179 6107 9191 6133
rect 9124 6103 9191 6107
rect 9091 6100 9191 6103
rect 9259 6100 9294 6137
rect 9356 6134 9715 6137
rect 9356 6129 9578 6134
rect 9356 6105 9369 6129
rect 9393 6110 9578 6129
rect 9602 6110 9715 6134
rect 9393 6105 9715 6110
rect 9356 6101 9715 6105
rect 9782 6129 9930 6137
rect 9782 6109 9793 6129
rect 9813 6120 9930 6129
rect 9979 6153 9986 6162
rect 9979 6120 9987 6153
rect 11185 6149 11250 6225
rect 11524 6204 11561 6283
rect 11602 6270 11712 6283
rect 11676 6214 11707 6215
rect 11524 6184 11533 6204
rect 11553 6184 11561 6204
rect 11524 6174 11561 6184
rect 11620 6204 11707 6214
rect 11620 6184 11629 6204
rect 11649 6184 11707 6204
rect 11620 6175 11707 6184
rect 11620 6174 11657 6175
rect 9813 6109 9987 6120
rect 9782 6102 9987 6109
rect 9782 6101 9823 6102
rect 9258 6075 9294 6100
rect 9106 6048 9143 6049
rect 9202 6048 9239 6049
rect 9258 6048 9265 6075
rect 8782 6023 8790 6043
rect 8810 6023 8819 6043
rect 8636 6012 8667 6013
rect 8631 5944 8741 5957
rect 8782 5944 8819 6023
rect 9006 6039 9144 6048
rect 9006 6019 9115 6039
rect 9135 6019 9144 6039
rect 9006 6012 9144 6019
rect 9202 6045 9265 6048
rect 9286 6048 9294 6075
rect 9313 6048 9350 6049
rect 9286 6045 9350 6048
rect 9202 6039 9350 6045
rect 9202 6019 9211 6039
rect 9231 6019 9321 6039
rect 9341 6019 9350 6039
rect 9006 6010 9102 6012
rect 9202 6009 9350 6019
rect 9409 6039 9446 6049
rect 9521 6048 9558 6049
rect 9502 6046 9558 6048
rect 9409 6019 9417 6039
rect 9437 6019 9446 6039
rect 9258 6008 9294 6009
rect 8569 5942 8819 5944
rect 8569 5939 8670 5942
rect 8569 5920 8634 5939
rect 8631 5912 8634 5920
rect 8663 5912 8670 5939
rect 8698 5915 8708 5942
rect 8737 5920 8819 5942
rect 8737 5915 8741 5920
rect 8698 5912 8741 5915
rect 8631 5898 8741 5912
rect 8057 5880 8398 5881
rect 7982 5875 8398 5880
rect 9106 5877 9143 5878
rect 9409 5877 9446 6019
rect 9471 6039 9558 6046
rect 9471 6036 9529 6039
rect 9471 6016 9476 6036
rect 9497 6019 9529 6036
rect 9549 6019 9558 6039
rect 9497 6016 9558 6019
rect 9471 6009 9558 6016
rect 9617 6039 9654 6049
rect 9617 6019 9625 6039
rect 9645 6019 9654 6039
rect 9471 6008 9502 6009
rect 9617 5940 9654 6019
rect 9684 6048 9715 6101
rect 9919 6099 9987 6102
rect 9919 6057 9931 6099
rect 9980 6057 9987 6099
rect 9734 6048 9771 6049
rect 9684 6039 9771 6048
rect 9684 6019 9742 6039
rect 9762 6019 9771 6039
rect 9684 6009 9771 6019
rect 9830 6039 9867 6049
rect 9919 6044 9987 6057
rect 10142 6121 10207 6138
rect 10142 6103 10166 6121
rect 10184 6103 10207 6121
rect 11185 6131 11207 6149
rect 11225 6131 11250 6149
rect 11185 6110 11250 6131
rect 11398 6129 11463 6138
rect 9830 6019 9838 6039
rect 9858 6019 9867 6039
rect 9684 6008 9715 6009
rect 9679 5940 9789 5953
rect 9830 5940 9867 6019
rect 10142 5964 10207 6103
rect 11398 6092 11408 6129
rect 11448 6121 11463 6129
rect 11676 6122 11707 6175
rect 11737 6204 11774 6283
rect 11889 6214 11920 6215
rect 11737 6184 11746 6204
rect 11766 6184 11774 6204
rect 11737 6174 11774 6184
rect 11833 6207 11920 6214
rect 11833 6204 11894 6207
rect 11833 6184 11842 6204
rect 11862 6187 11894 6204
rect 11915 6187 11920 6207
rect 11862 6184 11920 6187
rect 11833 6177 11920 6184
rect 11945 6204 11982 6346
rect 12248 6345 12285 6346
rect 13565 6286 13627 6757
rect 13727 6796 13753 6837
rect 13789 6796 13822 6837
rect 13727 6500 13822 6796
rect 13727 6456 13742 6500
rect 13802 6456 13822 6500
rect 13727 6436 13822 6456
rect 14439 6367 14482 7080
rect 14439 6347 14833 6367
rect 14853 6347 14856 6367
rect 14440 6342 14856 6347
rect 14440 6341 14781 6342
rect 14097 6310 14207 6324
rect 14097 6307 14140 6310
rect 14097 6302 14101 6307
rect 13560 6234 13635 6286
rect 14019 6280 14101 6302
rect 14130 6280 14140 6307
rect 14168 6283 14175 6310
rect 14204 6302 14207 6310
rect 14204 6283 14269 6302
rect 14168 6280 14269 6283
rect 14019 6278 14269 6280
rect 13929 6234 13975 6235
rect 12097 6214 12133 6215
rect 11945 6184 11954 6204
rect 11974 6184 11982 6204
rect 11833 6175 11889 6177
rect 11833 6174 11870 6175
rect 11945 6174 11982 6184
rect 12041 6204 12189 6214
rect 12289 6211 12385 6213
rect 12041 6184 12050 6204
rect 12070 6184 12160 6204
rect 12180 6184 12189 6204
rect 12041 6178 12189 6184
rect 12041 6175 12105 6178
rect 12041 6174 12078 6175
rect 12097 6148 12105 6175
rect 12126 6175 12189 6178
rect 12247 6204 12385 6211
rect 12247 6184 12256 6204
rect 12276 6184 12385 6204
rect 12247 6175 12385 6184
rect 13560 6199 13975 6234
rect 12126 6148 12133 6175
rect 12152 6174 12189 6175
rect 12248 6174 12285 6175
rect 12097 6123 12133 6148
rect 11568 6121 11609 6122
rect 11448 6114 11609 6121
rect 11448 6094 11578 6114
rect 11598 6094 11609 6114
rect 11448 6092 11609 6094
rect 11398 6086 11609 6092
rect 11676 6118 12035 6122
rect 11676 6113 11998 6118
rect 11676 6089 11789 6113
rect 11813 6094 11998 6113
rect 12022 6094 12035 6118
rect 11813 6089 12035 6094
rect 11676 6086 12035 6089
rect 12097 6086 12132 6123
rect 12200 6120 12300 6123
rect 12200 6116 12267 6120
rect 12200 6090 12212 6116
rect 12238 6094 12267 6116
rect 12293 6094 12300 6120
rect 12238 6090 12300 6094
rect 12200 6086 12300 6090
rect 11398 6073 11465 6086
rect 10142 5958 10164 5964
rect 9617 5938 9867 5940
rect 9617 5935 9718 5938
rect 9617 5916 9682 5935
rect 9679 5908 9682 5916
rect 9711 5908 9718 5935
rect 9746 5911 9756 5938
rect 9785 5916 9867 5938
rect 9896 5946 10164 5958
rect 10182 5946 10207 5964
rect 9896 5923 10207 5946
rect 11190 6050 11246 6070
rect 11190 6032 11209 6050
rect 11227 6032 11246 6050
rect 9896 5922 9951 5923
rect 9785 5911 9789 5916
rect 9746 5908 9789 5911
rect 9679 5894 9789 5908
rect 9105 5876 9446 5877
rect 7982 5855 7985 5875
rect 8005 5855 8398 5875
rect 9030 5875 9446 5876
rect 9896 5875 9939 5922
rect 11190 5919 11246 6032
rect 11398 6052 11412 6073
rect 11448 6052 11465 6073
rect 11676 6065 11707 6086
rect 12097 6065 12133 6086
rect 11519 6064 11556 6065
rect 11398 6045 11465 6052
rect 11518 6055 11556 6064
rect 9030 5871 9939 5875
rect 8349 5822 8394 5855
rect 9030 5851 9033 5871
rect 9053 5851 9939 5871
rect 9407 5846 9939 5851
rect 10147 5865 10206 5887
rect 10147 5847 10166 5865
rect 10184 5847 10206 5865
rect 9195 5822 9294 5824
rect 8349 5812 9294 5822
rect 8349 5786 9217 5812
rect 8350 5785 9217 5786
rect 9195 5774 9217 5785
rect 9242 5777 9261 5812
rect 9286 5777 9294 5812
rect 9242 5774 9294 5777
rect 10147 5776 10206 5847
rect 11190 5781 11245 5919
rect 11398 5893 11463 6045
rect 11518 6035 11527 6055
rect 11547 6035 11556 6055
rect 11518 6027 11556 6035
rect 11622 6059 11707 6065
rect 11732 6064 11769 6065
rect 11622 6039 11630 6059
rect 11650 6039 11707 6059
rect 11622 6031 11707 6039
rect 11731 6055 11769 6064
rect 11731 6035 11740 6055
rect 11760 6035 11769 6055
rect 11622 6030 11658 6031
rect 11731 6027 11769 6035
rect 11835 6059 11920 6065
rect 11940 6064 11977 6065
rect 11835 6039 11843 6059
rect 11863 6058 11920 6059
rect 11863 6039 11892 6058
rect 11835 6038 11892 6039
rect 11913 6038 11920 6058
rect 11835 6031 11920 6038
rect 11939 6055 11977 6064
rect 11939 6035 11948 6055
rect 11968 6035 11977 6055
rect 11835 6030 11871 6031
rect 11939 6027 11977 6035
rect 12043 6059 12187 6065
rect 12043 6039 12051 6059
rect 12071 6039 12159 6059
rect 12179 6039 12187 6059
rect 12043 6031 12187 6039
rect 12043 6030 12079 6031
rect 12151 6030 12187 6031
rect 12253 6064 12290 6065
rect 12253 6063 12291 6064
rect 12253 6055 12317 6063
rect 12253 6035 12262 6055
rect 12282 6041 12317 6055
rect 12337 6041 12340 6061
rect 12282 6036 12340 6041
rect 12282 6035 12317 6036
rect 11519 5998 11556 6027
rect 11520 5996 11556 5998
rect 11732 5996 11769 6027
rect 11520 5974 11769 5996
rect 11601 5968 11712 5974
rect 11601 5960 11642 5968
rect 11601 5940 11609 5960
rect 11628 5940 11642 5960
rect 11601 5938 11642 5940
rect 11670 5960 11712 5968
rect 11670 5940 11686 5960
rect 11705 5940 11712 5960
rect 11670 5938 11712 5940
rect 11601 5925 11712 5938
rect 11940 5928 11977 6027
rect 12253 6023 12317 6035
rect 11391 5883 11512 5893
rect 11391 5881 11460 5883
rect 11391 5840 11404 5881
rect 11441 5842 11460 5881
rect 11497 5842 11512 5883
rect 11441 5840 11512 5842
rect 11391 5822 11512 5840
rect 11183 5778 11247 5781
rect 11603 5778 11707 5784
rect 11938 5778 11979 5928
rect 12357 5920 12384 6175
rect 12446 6165 12526 6176
rect 12446 6139 12463 6165
rect 12503 6139 12526 6165
rect 12446 6112 12526 6139
rect 12446 6086 12467 6112
rect 12507 6086 12526 6112
rect 12446 6067 12526 6086
rect 12446 6041 12470 6067
rect 12510 6041 12526 6067
rect 12446 5990 12526 6041
rect 9195 5766 9294 5774
rect 9221 5765 9293 5766
rect 8875 5739 8942 5758
rect 8875 5718 8892 5739
rect 8873 5673 8892 5718
rect 8922 5718 8942 5739
rect 8922 5673 8943 5718
rect 9412 5715 9453 5717
rect 9684 5715 9788 5717
rect 10144 5715 10208 5776
rect 8873 5465 8943 5673
rect 9005 5680 10208 5715
rect 9005 5666 9033 5680
rect 9007 5535 9033 5666
rect 9412 5677 10208 5680
rect 11183 5775 11979 5778
rect 12358 5789 12384 5920
rect 12358 5775 12386 5789
rect 11183 5740 12386 5775
rect 12448 5782 12518 5990
rect 13560 5915 13635 6199
rect 13929 6116 13975 6199
rect 14019 6199 14056 6278
rect 14097 6265 14207 6278
rect 14171 6209 14202 6210
rect 14019 6179 14028 6199
rect 14048 6179 14056 6199
rect 14019 6169 14056 6179
rect 14115 6199 14202 6209
rect 14115 6179 14124 6199
rect 14144 6179 14202 6199
rect 14115 6170 14202 6179
rect 14115 6169 14152 6170
rect 14171 6117 14202 6170
rect 14232 6199 14269 6278
rect 14384 6209 14415 6210
rect 14232 6179 14241 6199
rect 14261 6179 14269 6199
rect 14232 6169 14269 6179
rect 14328 6202 14415 6209
rect 14328 6199 14389 6202
rect 14328 6179 14337 6199
rect 14357 6182 14389 6199
rect 14410 6182 14415 6202
rect 14357 6179 14415 6182
rect 14328 6172 14415 6179
rect 14440 6199 14477 6341
rect 14743 6340 14780 6341
rect 14592 6209 14628 6210
rect 14440 6179 14449 6199
rect 14469 6179 14477 6199
rect 14328 6170 14384 6172
rect 14328 6169 14365 6170
rect 14440 6169 14477 6179
rect 14536 6199 14684 6209
rect 14784 6206 14880 6208
rect 14536 6179 14545 6199
rect 14565 6179 14655 6199
rect 14675 6179 14684 6199
rect 14536 6173 14684 6179
rect 14536 6170 14600 6173
rect 14536 6169 14573 6170
rect 14592 6143 14600 6170
rect 14621 6170 14684 6173
rect 14742 6199 14880 6206
rect 14742 6179 14751 6199
rect 14771 6179 14880 6199
rect 14742 6170 14880 6179
rect 14621 6143 14628 6170
rect 14647 6169 14684 6170
rect 14743 6169 14780 6170
rect 14592 6118 14628 6143
rect 14063 6116 14104 6117
rect 13929 6109 14104 6116
rect 13727 6083 13813 6102
rect 13727 6042 13742 6083
rect 13796 6042 13813 6083
rect 13929 6089 14073 6109
rect 14093 6089 14104 6109
rect 13929 6081 14104 6089
rect 14171 6113 14530 6117
rect 14171 6108 14493 6113
rect 14171 6084 14284 6108
rect 14308 6089 14493 6108
rect 14517 6089 14530 6113
rect 14308 6084 14530 6089
rect 14171 6081 14530 6084
rect 14592 6081 14627 6118
rect 14695 6115 14795 6118
rect 14695 6111 14762 6115
rect 14695 6085 14707 6111
rect 14733 6089 14762 6111
rect 14788 6089 14795 6115
rect 14733 6085 14795 6089
rect 14695 6081 14795 6085
rect 13929 6077 13975 6081
rect 14171 6060 14202 6081
rect 14592 6060 14628 6081
rect 14014 6059 14051 6060
rect 13727 6006 13813 6042
rect 14013 6050 14051 6059
rect 14013 6030 14022 6050
rect 14042 6030 14051 6050
rect 14013 6022 14051 6030
rect 14117 6054 14202 6060
rect 14227 6059 14264 6060
rect 14117 6034 14125 6054
rect 14145 6034 14202 6054
rect 14117 6026 14202 6034
rect 14226 6050 14264 6059
rect 14226 6030 14235 6050
rect 14255 6030 14264 6050
rect 14117 6025 14153 6026
rect 14226 6022 14264 6030
rect 14330 6054 14415 6060
rect 14435 6059 14472 6060
rect 14330 6034 14338 6054
rect 14358 6053 14415 6054
rect 14358 6034 14387 6053
rect 14330 6033 14387 6034
rect 14408 6033 14415 6053
rect 14330 6026 14415 6033
rect 14434 6050 14472 6059
rect 14434 6030 14443 6050
rect 14463 6030 14472 6050
rect 14330 6025 14366 6026
rect 14434 6022 14472 6030
rect 14538 6054 14682 6060
rect 14538 6034 14546 6054
rect 14566 6034 14654 6054
rect 14674 6034 14682 6054
rect 14538 6026 14682 6034
rect 14538 6025 14574 6026
rect 11183 5679 11247 5740
rect 11603 5738 11707 5740
rect 11938 5738 11979 5740
rect 12448 5737 12469 5782
rect 12449 5716 12469 5737
rect 12499 5737 12518 5782
rect 13555 5873 13635 5915
rect 12499 5716 12516 5737
rect 12449 5697 12516 5716
rect 12098 5689 12170 5690
rect 12097 5681 12196 5689
rect 7760 5373 7842 5393
rect 7760 5350 7788 5373
rect 7814 5350 7842 5373
rect 7760 5288 7842 5350
rect 7764 5253 7842 5288
rect 8865 5414 8945 5465
rect 8865 5388 8881 5414
rect 8921 5388 8945 5414
rect 8865 5369 8945 5388
rect 8865 5343 8884 5369
rect 8924 5343 8945 5369
rect 8865 5316 8945 5343
rect 8865 5290 8888 5316
rect 8928 5290 8945 5316
rect 8865 5279 8945 5290
rect 9007 5280 9034 5535
rect 9412 5527 9453 5677
rect 9684 5671 9788 5677
rect 10144 5674 10208 5677
rect 9879 5615 10000 5633
rect 9879 5613 9950 5615
rect 9879 5572 9894 5613
rect 9931 5574 9950 5613
rect 9987 5574 10000 5615
rect 9931 5572 10000 5574
rect 9879 5562 10000 5572
rect 9074 5420 9138 5432
rect 9414 5428 9451 5527
rect 9679 5517 9790 5530
rect 9679 5515 9721 5517
rect 9679 5495 9686 5515
rect 9705 5495 9721 5515
rect 9679 5487 9721 5495
rect 9749 5515 9790 5517
rect 9749 5495 9763 5515
rect 9782 5495 9790 5515
rect 9749 5487 9790 5495
rect 9679 5481 9790 5487
rect 9622 5459 9871 5481
rect 9622 5428 9659 5459
rect 9835 5457 9871 5459
rect 9835 5428 9872 5457
rect 9074 5419 9109 5420
rect 9051 5414 9109 5419
rect 9051 5394 9054 5414
rect 9074 5400 9109 5414
rect 9129 5400 9138 5420
rect 9074 5392 9138 5400
rect 9100 5391 9138 5392
rect 9101 5390 9138 5391
rect 9204 5424 9240 5425
rect 9312 5424 9348 5425
rect 9204 5416 9348 5424
rect 9204 5396 9212 5416
rect 9232 5396 9320 5416
rect 9340 5396 9348 5416
rect 9204 5390 9348 5396
rect 9414 5420 9452 5428
rect 9520 5424 9556 5425
rect 9414 5400 9423 5420
rect 9443 5400 9452 5420
rect 9414 5391 9452 5400
rect 9471 5417 9556 5424
rect 9471 5397 9478 5417
rect 9499 5416 9556 5417
rect 9499 5397 9528 5416
rect 9471 5396 9528 5397
rect 9548 5396 9556 5416
rect 9414 5390 9451 5391
rect 9471 5390 9556 5396
rect 9622 5420 9660 5428
rect 9733 5424 9769 5425
rect 9622 5400 9631 5420
rect 9651 5400 9660 5420
rect 9622 5391 9660 5400
rect 9684 5416 9769 5424
rect 9684 5396 9741 5416
rect 9761 5396 9769 5416
rect 9622 5390 9659 5391
rect 9684 5390 9769 5396
rect 9835 5420 9873 5428
rect 9835 5400 9844 5420
rect 9864 5400 9873 5420
rect 9928 5410 9993 5562
rect 10146 5536 10201 5674
rect 11185 5608 11244 5679
rect 12097 5678 12149 5681
rect 12097 5643 12105 5678
rect 12130 5643 12149 5678
rect 12174 5670 12196 5681
rect 12174 5669 13041 5670
rect 12174 5643 13042 5669
rect 12097 5633 13042 5643
rect 12097 5631 12196 5633
rect 11185 5590 11207 5608
rect 11225 5590 11244 5608
rect 11185 5568 11244 5590
rect 11452 5604 11984 5609
rect 11452 5584 12338 5604
rect 12358 5584 12361 5604
rect 12997 5600 13042 5633
rect 11452 5580 12361 5584
rect 9835 5391 9873 5400
rect 9926 5403 9993 5410
rect 9835 5390 9872 5391
rect 9258 5369 9294 5390
rect 9684 5369 9715 5390
rect 9926 5382 9943 5403
rect 9979 5382 9993 5403
rect 10145 5423 10201 5536
rect 11452 5533 11495 5580
rect 11945 5579 12361 5580
rect 12993 5580 13386 5600
rect 13406 5580 13409 5600
rect 11945 5578 12286 5579
rect 11602 5547 11712 5561
rect 11602 5544 11645 5547
rect 11602 5539 11606 5544
rect 11440 5532 11495 5533
rect 10145 5405 10164 5423
rect 10182 5405 10201 5423
rect 10145 5385 10201 5405
rect 11184 5509 11495 5532
rect 11184 5491 11209 5509
rect 11227 5497 11495 5509
rect 11524 5517 11606 5539
rect 11635 5517 11645 5544
rect 11673 5520 11680 5547
rect 11709 5539 11712 5547
rect 11709 5520 11774 5539
rect 11673 5517 11774 5520
rect 11524 5515 11774 5517
rect 11227 5491 11249 5497
rect 9926 5369 9993 5382
rect 9091 5365 9191 5369
rect 9091 5361 9153 5365
rect 9091 5335 9098 5361
rect 9124 5339 9153 5361
rect 9179 5339 9191 5365
rect 9124 5335 9191 5339
rect 9091 5332 9191 5335
rect 9259 5332 9294 5369
rect 9356 5366 9715 5369
rect 9356 5361 9578 5366
rect 9356 5337 9369 5361
rect 9393 5342 9578 5361
rect 9602 5342 9715 5366
rect 9393 5337 9715 5342
rect 9356 5333 9715 5337
rect 9782 5363 9993 5369
rect 9782 5361 9943 5363
rect 9782 5341 9793 5361
rect 9813 5341 9943 5361
rect 9782 5334 9943 5341
rect 9782 5333 9823 5334
rect 9258 5307 9294 5332
rect 9106 5280 9143 5281
rect 9202 5280 9239 5281
rect 9258 5280 9265 5307
rect 9006 5271 9144 5280
rect 7764 4737 7826 5253
rect 9006 5251 9115 5271
rect 9135 5251 9144 5271
rect 9006 5244 9144 5251
rect 9202 5277 9265 5280
rect 9286 5280 9294 5307
rect 9313 5280 9350 5281
rect 9286 5277 9350 5280
rect 9202 5271 9350 5277
rect 9202 5251 9211 5271
rect 9231 5251 9321 5271
rect 9341 5251 9350 5271
rect 9006 5242 9102 5244
rect 9202 5241 9350 5251
rect 9409 5271 9446 5281
rect 9521 5280 9558 5281
rect 9502 5278 9558 5280
rect 9409 5251 9417 5271
rect 9437 5251 9446 5271
rect 9258 5240 9294 5241
rect 9106 5109 9143 5110
rect 9409 5109 9446 5251
rect 9471 5271 9558 5278
rect 9471 5268 9529 5271
rect 9471 5248 9476 5268
rect 9497 5251 9529 5268
rect 9549 5251 9558 5271
rect 9497 5248 9558 5251
rect 9471 5241 9558 5248
rect 9617 5271 9654 5281
rect 9617 5251 9625 5271
rect 9645 5251 9654 5271
rect 9471 5240 9502 5241
rect 9617 5172 9654 5251
rect 9684 5280 9715 5333
rect 9928 5326 9943 5334
rect 9983 5326 9993 5363
rect 11184 5352 11249 5491
rect 11524 5436 11561 5515
rect 11602 5502 11712 5515
rect 11676 5446 11707 5447
rect 11524 5416 11533 5436
rect 11553 5416 11561 5436
rect 9928 5317 9993 5326
rect 10141 5324 10206 5345
rect 10141 5306 10166 5324
rect 10184 5306 10206 5324
rect 11184 5334 11207 5352
rect 11225 5334 11249 5352
rect 11184 5317 11249 5334
rect 11404 5398 11472 5411
rect 11524 5406 11561 5416
rect 11620 5436 11707 5446
rect 11620 5416 11629 5436
rect 11649 5416 11707 5436
rect 11620 5407 11707 5416
rect 11620 5406 11657 5407
rect 11404 5356 11411 5398
rect 11460 5356 11472 5398
rect 11404 5353 11472 5356
rect 11676 5354 11707 5407
rect 11737 5436 11774 5515
rect 11889 5446 11920 5447
rect 11737 5416 11746 5436
rect 11766 5416 11774 5436
rect 11737 5406 11774 5416
rect 11833 5439 11920 5446
rect 11833 5436 11894 5439
rect 11833 5416 11842 5436
rect 11862 5419 11894 5436
rect 11915 5419 11920 5439
rect 11862 5416 11920 5419
rect 11833 5409 11920 5416
rect 11945 5436 11982 5578
rect 12248 5577 12285 5578
rect 12993 5575 13409 5580
rect 12993 5574 13334 5575
rect 12650 5543 12760 5557
rect 12650 5540 12693 5543
rect 12650 5535 12654 5540
rect 12572 5513 12654 5535
rect 12683 5513 12693 5540
rect 12721 5516 12728 5543
rect 12757 5535 12760 5543
rect 12757 5516 12822 5535
rect 12721 5513 12822 5516
rect 12572 5511 12822 5513
rect 12097 5446 12133 5447
rect 11945 5416 11954 5436
rect 11974 5416 11982 5436
rect 11833 5407 11889 5409
rect 11833 5406 11870 5407
rect 11945 5406 11982 5416
rect 12041 5436 12189 5446
rect 12289 5443 12385 5445
rect 12041 5416 12050 5436
rect 12070 5416 12160 5436
rect 12180 5416 12189 5436
rect 12041 5410 12189 5416
rect 12041 5407 12105 5410
rect 12041 5406 12078 5407
rect 12097 5380 12105 5407
rect 12126 5407 12189 5410
rect 12247 5436 12385 5443
rect 12247 5416 12256 5436
rect 12276 5416 12385 5436
rect 12247 5407 12385 5416
rect 12572 5432 12609 5511
rect 12650 5498 12760 5511
rect 12724 5442 12755 5443
rect 12572 5412 12581 5432
rect 12601 5412 12609 5432
rect 12126 5380 12133 5407
rect 12152 5406 12189 5407
rect 12248 5406 12285 5407
rect 12097 5355 12133 5380
rect 11568 5353 11609 5354
rect 11404 5346 11609 5353
rect 11404 5335 11578 5346
rect 9734 5280 9771 5281
rect 9684 5271 9771 5280
rect 9684 5251 9742 5271
rect 9762 5251 9771 5271
rect 9684 5241 9771 5251
rect 9830 5271 9867 5281
rect 9830 5251 9838 5271
rect 9858 5251 9867 5271
rect 9684 5240 9715 5241
rect 9679 5172 9789 5185
rect 9830 5172 9867 5251
rect 10141 5230 10206 5306
rect 11404 5302 11412 5335
rect 11405 5293 11412 5302
rect 11461 5326 11578 5335
rect 11598 5326 11609 5346
rect 11461 5318 11609 5326
rect 11676 5350 12035 5354
rect 11676 5345 11998 5350
rect 11676 5321 11789 5345
rect 11813 5326 11998 5345
rect 12022 5326 12035 5350
rect 11813 5321 12035 5326
rect 11676 5318 12035 5321
rect 12097 5318 12132 5355
rect 12200 5352 12300 5355
rect 12200 5348 12267 5352
rect 12200 5322 12212 5348
rect 12238 5326 12267 5348
rect 12293 5326 12300 5352
rect 12238 5322 12300 5326
rect 12200 5318 12300 5322
rect 11461 5302 11472 5318
rect 11461 5293 11469 5302
rect 11676 5297 11707 5318
rect 12097 5297 12133 5318
rect 11519 5296 11556 5297
rect 11184 5253 11249 5272
rect 11184 5235 11209 5253
rect 11227 5235 11249 5253
rect 9617 5170 9867 5172
rect 9617 5167 9718 5170
rect 9617 5148 9682 5167
rect 9679 5140 9682 5148
rect 9711 5140 9718 5167
rect 9746 5143 9756 5170
rect 9785 5148 9867 5170
rect 9890 5195 10207 5230
rect 9785 5143 9789 5148
rect 9746 5140 9789 5143
rect 9679 5126 9789 5140
rect 9105 5108 9446 5109
rect 9030 5106 9446 5108
rect 9890 5106 9930 5195
rect 10141 5168 10206 5195
rect 10141 5150 10164 5168
rect 10182 5150 10206 5168
rect 10141 5130 10206 5150
rect 9027 5103 9930 5106
rect 9027 5083 9033 5103
rect 9053 5083 9930 5103
rect 9027 5079 9930 5083
rect 9890 5076 9930 5079
rect 10142 5069 10207 5090
rect 8360 5061 9021 5062
rect 8360 5054 9294 5061
rect 8360 5053 9266 5054
rect 8360 5033 9211 5053
rect 9243 5034 9266 5053
rect 9291 5034 9294 5054
rect 9243 5033 9294 5034
rect 8360 5026 9294 5033
rect 7959 4984 8127 4985
rect 8362 4984 8401 5026
rect 9190 5024 9294 5026
rect 9259 5022 9294 5024
rect 10142 5051 10166 5069
rect 10184 5051 10207 5069
rect 10142 5004 10207 5051
rect 7959 4958 8403 4984
rect 7959 4956 8127 4958
rect 7761 4653 7830 4737
rect 7759 4174 7830 4653
rect 7959 4605 7986 4956
rect 8362 4952 8403 4958
rect 8026 4745 8090 4757
rect 8366 4753 8403 4952
rect 8865 4979 8937 4996
rect 8865 4940 8873 4979
rect 8918 4940 8937 4979
rect 8631 4842 8742 4857
rect 8631 4840 8673 4842
rect 8631 4820 8638 4840
rect 8657 4820 8673 4840
rect 8631 4812 8673 4820
rect 8701 4840 8742 4842
rect 8701 4820 8715 4840
rect 8734 4820 8742 4840
rect 8701 4812 8742 4820
rect 8631 4806 8742 4812
rect 8574 4784 8823 4806
rect 8574 4753 8611 4784
rect 8787 4782 8823 4784
rect 8787 4753 8824 4782
rect 8026 4744 8061 4745
rect 8003 4739 8061 4744
rect 8003 4719 8006 4739
rect 8026 4725 8061 4739
rect 8081 4725 8090 4745
rect 8026 4717 8090 4725
rect 8052 4716 8090 4717
rect 8053 4715 8090 4716
rect 8156 4749 8192 4750
rect 8264 4749 8300 4750
rect 8156 4741 8300 4749
rect 8156 4721 8164 4741
rect 8184 4721 8272 4741
rect 8292 4721 8300 4741
rect 8156 4715 8300 4721
rect 8366 4745 8404 4753
rect 8472 4749 8508 4750
rect 8366 4725 8375 4745
rect 8395 4725 8404 4745
rect 8366 4716 8404 4725
rect 8423 4742 8508 4749
rect 8423 4722 8430 4742
rect 8451 4741 8508 4742
rect 8451 4722 8480 4741
rect 8423 4721 8480 4722
rect 8500 4721 8508 4741
rect 8366 4715 8403 4716
rect 8423 4715 8508 4721
rect 8574 4745 8612 4753
rect 8685 4749 8721 4750
rect 8574 4725 8583 4745
rect 8603 4725 8612 4745
rect 8574 4716 8612 4725
rect 8636 4741 8721 4749
rect 8636 4721 8693 4741
rect 8713 4721 8721 4741
rect 8574 4715 8611 4716
rect 8636 4715 8721 4721
rect 8787 4745 8825 4753
rect 8787 4725 8796 4745
rect 8816 4725 8825 4745
rect 8787 4716 8825 4725
rect 8865 4730 8937 4940
rect 9007 4974 10207 5004
rect 9007 4973 9451 4974
rect 9007 4971 9175 4973
rect 8865 4716 8948 4730
rect 8787 4715 8824 4716
rect 8210 4694 8246 4715
rect 8636 4694 8667 4715
rect 8865 4694 8882 4716
rect 8043 4690 8143 4694
rect 8043 4686 8105 4690
rect 8043 4660 8050 4686
rect 8076 4664 8105 4686
rect 8131 4664 8143 4690
rect 8076 4660 8143 4664
rect 8043 4657 8143 4660
rect 8211 4657 8246 4694
rect 8308 4691 8667 4694
rect 8308 4686 8530 4691
rect 8308 4662 8321 4686
rect 8345 4667 8530 4686
rect 8554 4667 8667 4691
rect 8345 4662 8667 4667
rect 8308 4658 8667 4662
rect 8734 4686 8882 4694
rect 8734 4666 8745 4686
rect 8765 4683 8882 4686
rect 8935 4683 8948 4716
rect 8765 4666 8948 4683
rect 8734 4659 8948 4666
rect 8734 4658 8775 4659
rect 8865 4658 8948 4659
rect 8210 4632 8246 4657
rect 8058 4605 8095 4606
rect 8154 4605 8191 4606
rect 8210 4605 8217 4632
rect 7958 4596 8096 4605
rect 7958 4576 8067 4596
rect 8087 4576 8096 4596
rect 7958 4569 8096 4576
rect 8154 4602 8217 4605
rect 8238 4605 8246 4632
rect 8265 4605 8302 4606
rect 8238 4602 8302 4605
rect 8154 4596 8302 4602
rect 8154 4576 8163 4596
rect 8183 4576 8273 4596
rect 8293 4576 8302 4596
rect 7958 4567 8054 4569
rect 8154 4566 8302 4576
rect 8361 4596 8398 4606
rect 8473 4605 8510 4606
rect 8454 4603 8510 4605
rect 8361 4576 8369 4596
rect 8389 4576 8398 4596
rect 8210 4565 8246 4566
rect 8058 4434 8095 4435
rect 8361 4434 8398 4576
rect 8423 4596 8510 4603
rect 8423 4593 8481 4596
rect 8423 4573 8428 4593
rect 8449 4576 8481 4593
rect 8501 4576 8510 4596
rect 8449 4573 8510 4576
rect 8423 4566 8510 4573
rect 8569 4596 8606 4606
rect 8569 4576 8577 4596
rect 8597 4576 8606 4596
rect 8423 4565 8454 4566
rect 8569 4497 8606 4576
rect 8636 4605 8667 4658
rect 8873 4625 8887 4658
rect 8940 4625 8948 4658
rect 8873 4619 8948 4625
rect 8873 4614 8943 4619
rect 8686 4605 8723 4606
rect 8636 4596 8723 4605
rect 8636 4576 8694 4596
rect 8714 4576 8723 4596
rect 8636 4566 8723 4576
rect 8782 4596 8819 4606
rect 9007 4601 9034 4971
rect 9074 4741 9138 4753
rect 9414 4749 9451 4973
rect 9922 4954 9986 4956
rect 9918 4942 9986 4954
rect 9918 4909 9929 4942
rect 9969 4909 9986 4942
rect 9918 4899 9986 4909
rect 9679 4838 9790 4853
rect 9679 4836 9721 4838
rect 9679 4816 9686 4836
rect 9705 4816 9721 4836
rect 9679 4808 9721 4816
rect 9749 4836 9790 4838
rect 9749 4816 9763 4836
rect 9782 4816 9790 4836
rect 9749 4808 9790 4816
rect 9679 4802 9790 4808
rect 9622 4780 9871 4802
rect 9622 4749 9659 4780
rect 9835 4778 9871 4780
rect 9835 4749 9872 4778
rect 9074 4740 9109 4741
rect 9051 4735 9109 4740
rect 9051 4715 9054 4735
rect 9074 4721 9109 4735
rect 9129 4721 9138 4741
rect 9074 4713 9138 4721
rect 9100 4712 9138 4713
rect 9101 4711 9138 4712
rect 9204 4745 9240 4746
rect 9312 4745 9348 4746
rect 9204 4737 9348 4745
rect 9204 4717 9212 4737
rect 9232 4717 9320 4737
rect 9340 4717 9348 4737
rect 9204 4711 9348 4717
rect 9414 4741 9452 4749
rect 9520 4745 9556 4746
rect 9414 4721 9423 4741
rect 9443 4721 9452 4741
rect 9414 4712 9452 4721
rect 9471 4738 9556 4745
rect 9471 4718 9478 4738
rect 9499 4737 9556 4738
rect 9499 4718 9528 4737
rect 9471 4717 9528 4718
rect 9548 4717 9556 4737
rect 9414 4711 9451 4712
rect 9471 4711 9556 4717
rect 9622 4741 9660 4749
rect 9733 4745 9769 4746
rect 9622 4721 9631 4741
rect 9651 4721 9660 4741
rect 9622 4712 9660 4721
rect 9684 4737 9769 4745
rect 9684 4717 9741 4737
rect 9761 4717 9769 4737
rect 9622 4711 9659 4712
rect 9684 4711 9769 4717
rect 9835 4741 9873 4749
rect 9835 4721 9844 4741
rect 9864 4721 9873 4741
rect 9835 4712 9873 4721
rect 9922 4715 9986 4899
rect 10142 4773 10207 4974
rect 11184 5034 11249 5235
rect 11405 5109 11469 5293
rect 11518 5287 11556 5296
rect 11518 5267 11527 5287
rect 11547 5267 11556 5287
rect 11518 5259 11556 5267
rect 11622 5291 11707 5297
rect 11732 5296 11769 5297
rect 11622 5271 11630 5291
rect 11650 5271 11707 5291
rect 11622 5263 11707 5271
rect 11731 5287 11769 5296
rect 11731 5267 11740 5287
rect 11760 5267 11769 5287
rect 11622 5262 11658 5263
rect 11731 5259 11769 5267
rect 11835 5291 11920 5297
rect 11940 5296 11977 5297
rect 11835 5271 11843 5291
rect 11863 5290 11920 5291
rect 11863 5271 11892 5290
rect 11835 5270 11892 5271
rect 11913 5270 11920 5290
rect 11835 5263 11920 5270
rect 11939 5287 11977 5296
rect 11939 5267 11948 5287
rect 11968 5267 11977 5287
rect 11835 5262 11871 5263
rect 11939 5259 11977 5267
rect 12043 5291 12187 5297
rect 12043 5271 12051 5291
rect 12071 5271 12159 5291
rect 12179 5271 12187 5291
rect 12043 5263 12187 5271
rect 12043 5262 12079 5263
rect 12151 5262 12187 5263
rect 12253 5296 12290 5297
rect 12253 5295 12291 5296
rect 12253 5287 12317 5295
rect 12253 5267 12262 5287
rect 12282 5273 12317 5287
rect 12337 5273 12340 5293
rect 12282 5268 12340 5273
rect 12282 5267 12317 5268
rect 11519 5230 11556 5259
rect 11520 5228 11556 5230
rect 11732 5228 11769 5259
rect 11520 5206 11769 5228
rect 11601 5200 11712 5206
rect 11601 5192 11642 5200
rect 11601 5172 11609 5192
rect 11628 5172 11642 5192
rect 11601 5170 11642 5172
rect 11670 5192 11712 5200
rect 11670 5172 11686 5192
rect 11705 5172 11712 5192
rect 11670 5170 11712 5172
rect 11601 5155 11712 5170
rect 11405 5099 11473 5109
rect 11405 5066 11422 5099
rect 11462 5066 11473 5099
rect 11405 5054 11473 5066
rect 11405 5052 11469 5054
rect 11940 5035 11977 5259
rect 12253 5255 12317 5267
rect 12357 5037 12384 5407
rect 12572 5402 12609 5412
rect 12668 5432 12755 5442
rect 12668 5412 12677 5432
rect 12697 5412 12755 5432
rect 12668 5403 12755 5412
rect 12668 5402 12705 5403
rect 12448 5389 12518 5394
rect 12443 5383 12518 5389
rect 12443 5350 12451 5383
rect 12504 5350 12518 5383
rect 12724 5350 12755 5403
rect 12785 5432 12822 5511
rect 12937 5442 12968 5443
rect 12785 5412 12794 5432
rect 12814 5412 12822 5432
rect 12785 5402 12822 5412
rect 12881 5435 12968 5442
rect 12881 5432 12942 5435
rect 12881 5412 12890 5432
rect 12910 5415 12942 5432
rect 12963 5415 12968 5435
rect 12910 5412 12968 5415
rect 12881 5405 12968 5412
rect 12993 5432 13030 5574
rect 13296 5573 13333 5574
rect 13145 5442 13181 5443
rect 12993 5412 13002 5432
rect 13022 5412 13030 5432
rect 12881 5403 12937 5405
rect 12881 5402 12918 5403
rect 12993 5402 13030 5412
rect 13089 5432 13237 5442
rect 13337 5439 13433 5441
rect 13089 5412 13098 5432
rect 13118 5412 13208 5432
rect 13228 5412 13237 5432
rect 13089 5406 13237 5412
rect 13089 5403 13153 5406
rect 13089 5402 13126 5403
rect 13145 5376 13153 5403
rect 13174 5403 13237 5406
rect 13295 5432 13433 5439
rect 13295 5412 13304 5432
rect 13324 5412 13433 5432
rect 13295 5403 13433 5412
rect 13174 5376 13181 5403
rect 13200 5402 13237 5403
rect 13296 5402 13333 5403
rect 13145 5351 13181 5376
rect 12443 5349 12526 5350
rect 12616 5349 12657 5350
rect 12443 5342 12657 5349
rect 12443 5325 12626 5342
rect 12443 5292 12456 5325
rect 12509 5322 12626 5325
rect 12646 5322 12657 5342
rect 12509 5314 12657 5322
rect 12724 5346 13083 5350
rect 12724 5341 13046 5346
rect 12724 5317 12837 5341
rect 12861 5322 13046 5341
rect 13070 5322 13083 5346
rect 12861 5317 13083 5322
rect 12724 5314 13083 5317
rect 13145 5314 13180 5351
rect 13248 5348 13348 5351
rect 13248 5344 13315 5348
rect 13248 5318 13260 5344
rect 13286 5322 13315 5344
rect 13341 5322 13348 5348
rect 13286 5318 13348 5322
rect 13248 5314 13348 5318
rect 12509 5292 12526 5314
rect 12724 5293 12755 5314
rect 13145 5293 13181 5314
rect 12567 5292 12604 5293
rect 12443 5278 12526 5292
rect 12216 5035 12384 5037
rect 11940 5034 12384 5035
rect 11184 5004 12384 5034
rect 12454 5068 12526 5278
rect 12566 5283 12604 5292
rect 12566 5263 12575 5283
rect 12595 5263 12604 5283
rect 12566 5255 12604 5263
rect 12670 5287 12755 5293
rect 12780 5292 12817 5293
rect 12670 5267 12678 5287
rect 12698 5267 12755 5287
rect 12670 5259 12755 5267
rect 12779 5283 12817 5292
rect 12779 5263 12788 5283
rect 12808 5263 12817 5283
rect 12670 5258 12706 5259
rect 12779 5255 12817 5263
rect 12883 5287 12968 5293
rect 12988 5292 13025 5293
rect 12883 5267 12891 5287
rect 12911 5286 12968 5287
rect 12911 5267 12940 5286
rect 12883 5266 12940 5267
rect 12961 5266 12968 5286
rect 12883 5259 12968 5266
rect 12987 5283 13025 5292
rect 12987 5263 12996 5283
rect 13016 5263 13025 5283
rect 12883 5258 12919 5259
rect 12987 5255 13025 5263
rect 13091 5287 13235 5293
rect 13091 5267 13099 5287
rect 13119 5267 13207 5287
rect 13227 5267 13235 5287
rect 13091 5259 13235 5267
rect 13091 5258 13127 5259
rect 13199 5258 13235 5259
rect 13301 5292 13338 5293
rect 13301 5291 13339 5292
rect 13301 5283 13365 5291
rect 13301 5263 13310 5283
rect 13330 5269 13365 5283
rect 13385 5269 13388 5289
rect 13330 5264 13388 5269
rect 13330 5263 13365 5264
rect 12567 5226 12604 5255
rect 12568 5224 12604 5226
rect 12780 5224 12817 5255
rect 12568 5202 12817 5224
rect 12649 5196 12760 5202
rect 12649 5188 12690 5196
rect 12649 5168 12657 5188
rect 12676 5168 12690 5188
rect 12649 5166 12690 5168
rect 12718 5188 12760 5196
rect 12718 5168 12734 5188
rect 12753 5168 12760 5188
rect 12718 5166 12760 5168
rect 12649 5151 12760 5166
rect 12454 5029 12473 5068
rect 12518 5029 12526 5068
rect 12454 5012 12526 5029
rect 12988 5056 13025 5255
rect 13301 5251 13365 5263
rect 12988 5050 13029 5056
rect 13405 5052 13432 5403
rect 13555 5273 13634 5873
rect 13731 5421 13810 6006
rect 14014 5993 14051 6022
rect 14015 5991 14051 5993
rect 14227 5991 14264 6022
rect 14015 5969 14264 5991
rect 14096 5963 14207 5969
rect 14096 5955 14137 5963
rect 14096 5935 14104 5955
rect 14123 5935 14137 5955
rect 14096 5933 14137 5935
rect 14165 5955 14207 5963
rect 14165 5935 14181 5955
rect 14200 5935 14207 5955
rect 14165 5933 14207 5935
rect 14096 5918 14207 5933
rect 14435 5907 14472 6022
rect 14428 5795 14475 5907
rect 14596 5867 14626 6026
rect 14646 6025 14682 6026
rect 14748 6059 14785 6060
rect 14748 6058 14786 6059
rect 14748 6050 14812 6058
rect 14748 6030 14757 6050
rect 14777 6036 14812 6050
rect 14832 6036 14835 6056
rect 14777 6031 14835 6036
rect 14777 6030 14812 6031
rect 14748 6018 14812 6030
rect 14596 5863 14682 5867
rect 14596 5845 14611 5863
rect 14663 5845 14682 5863
rect 14596 5836 14682 5845
rect 14852 5797 14879 6170
rect 14711 5795 14879 5797
rect 14428 5769 14879 5795
rect 14428 5691 14475 5769
rect 14711 5768 14879 5769
rect 14373 5690 14475 5691
rect 14372 5682 14475 5690
rect 14372 5679 14424 5682
rect 14372 5644 14380 5679
rect 14405 5644 14424 5679
rect 14449 5644 14475 5682
rect 14372 5638 14475 5644
rect 14635 5683 14671 5687
rect 14635 5660 14643 5683
rect 14667 5660 14671 5683
rect 14635 5639 14671 5660
rect 14372 5634 14471 5638
rect 14635 5616 14643 5639
rect 14667 5616 14671 5639
rect 13264 5050 13432 5052
rect 12988 5024 13432 5050
rect 11184 4957 11249 5004
rect 11184 4939 11207 4957
rect 11225 4939 11249 4957
rect 12097 4984 12132 4986
rect 12097 4982 12201 4984
rect 12990 4982 13029 5024
rect 13264 5023 13432 5024
rect 12097 4975 13031 4982
rect 12097 4974 12148 4975
rect 12097 4954 12100 4974
rect 12125 4955 12148 4974
rect 12180 4955 13031 4975
rect 12125 4954 13031 4955
rect 12097 4947 13031 4954
rect 12370 4946 13031 4947
rect 11184 4918 11249 4939
rect 11461 4929 11501 4932
rect 11461 4925 12364 4929
rect 11461 4905 12338 4925
rect 12358 4905 12364 4925
rect 11461 4902 12364 4905
rect 11185 4858 11250 4878
rect 11185 4840 11209 4858
rect 11227 4840 11250 4858
rect 11185 4813 11250 4840
rect 11461 4813 11501 4902
rect 11945 4900 12361 4902
rect 11945 4899 12286 4900
rect 11602 4868 11712 4882
rect 11602 4865 11645 4868
rect 11602 4860 11606 4865
rect 11184 4778 11501 4813
rect 11524 4838 11606 4860
rect 11635 4838 11645 4865
rect 11673 4841 11680 4868
rect 11709 4860 11712 4868
rect 11709 4841 11774 4860
rect 11673 4838 11774 4841
rect 11524 4836 11774 4838
rect 10142 4755 10164 4773
rect 10182 4755 10207 4773
rect 10142 4736 10207 4755
rect 9835 4711 9872 4712
rect 9258 4690 9294 4711
rect 9684 4690 9715 4711
rect 9922 4706 9930 4715
rect 9919 4690 9930 4706
rect 9091 4686 9191 4690
rect 9091 4682 9153 4686
rect 9091 4656 9098 4682
rect 9124 4660 9153 4682
rect 9179 4660 9191 4686
rect 9124 4656 9191 4660
rect 9091 4653 9191 4656
rect 9259 4653 9294 4690
rect 9356 4687 9715 4690
rect 9356 4682 9578 4687
rect 9356 4658 9369 4682
rect 9393 4663 9578 4682
rect 9602 4663 9715 4687
rect 9393 4658 9715 4663
rect 9356 4654 9715 4658
rect 9782 4682 9930 4690
rect 9782 4662 9793 4682
rect 9813 4673 9930 4682
rect 9979 4706 9986 4715
rect 9979 4673 9987 4706
rect 11185 4702 11250 4778
rect 11524 4757 11561 4836
rect 11602 4823 11712 4836
rect 11676 4767 11707 4768
rect 11524 4737 11533 4757
rect 11553 4737 11561 4757
rect 11524 4727 11561 4737
rect 11620 4757 11707 4767
rect 11620 4737 11629 4757
rect 11649 4737 11707 4757
rect 11620 4728 11707 4737
rect 11620 4727 11657 4728
rect 9813 4662 9987 4673
rect 9782 4655 9987 4662
rect 9782 4654 9823 4655
rect 9258 4628 9294 4653
rect 9106 4601 9143 4602
rect 9202 4601 9239 4602
rect 9258 4601 9265 4628
rect 8782 4576 8790 4596
rect 8810 4576 8819 4596
rect 8636 4565 8667 4566
rect 8631 4497 8741 4510
rect 8782 4497 8819 4576
rect 9006 4592 9144 4601
rect 9006 4572 9115 4592
rect 9135 4572 9144 4592
rect 9006 4565 9144 4572
rect 9202 4598 9265 4601
rect 9286 4601 9294 4628
rect 9313 4601 9350 4602
rect 9286 4598 9350 4601
rect 9202 4592 9350 4598
rect 9202 4572 9211 4592
rect 9231 4572 9321 4592
rect 9341 4572 9350 4592
rect 9006 4563 9102 4565
rect 9202 4562 9350 4572
rect 9409 4592 9446 4602
rect 9521 4601 9558 4602
rect 9502 4599 9558 4601
rect 9409 4572 9417 4592
rect 9437 4572 9446 4592
rect 9258 4561 9294 4562
rect 8569 4495 8819 4497
rect 8569 4492 8670 4495
rect 8569 4473 8634 4492
rect 8631 4465 8634 4473
rect 8663 4465 8670 4492
rect 8698 4468 8708 4495
rect 8737 4473 8819 4495
rect 8737 4468 8741 4473
rect 8698 4465 8741 4468
rect 8631 4451 8741 4465
rect 8057 4433 8398 4434
rect 7982 4428 8398 4433
rect 9106 4430 9143 4431
rect 9409 4430 9446 4572
rect 9471 4592 9558 4599
rect 9471 4589 9529 4592
rect 9471 4569 9476 4589
rect 9497 4572 9529 4589
rect 9549 4572 9558 4592
rect 9497 4569 9558 4572
rect 9471 4562 9558 4569
rect 9617 4592 9654 4602
rect 9617 4572 9625 4592
rect 9645 4572 9654 4592
rect 9471 4561 9502 4562
rect 9617 4493 9654 4572
rect 9684 4601 9715 4654
rect 9919 4652 9987 4655
rect 9919 4610 9931 4652
rect 9980 4610 9987 4652
rect 9734 4601 9771 4602
rect 9684 4592 9771 4601
rect 9684 4572 9742 4592
rect 9762 4572 9771 4592
rect 9684 4562 9771 4572
rect 9830 4592 9867 4602
rect 9919 4597 9987 4610
rect 10142 4674 10207 4691
rect 10142 4656 10166 4674
rect 10184 4656 10207 4674
rect 11185 4684 11207 4702
rect 11225 4684 11250 4702
rect 11185 4663 11250 4684
rect 11398 4682 11463 4691
rect 9830 4572 9838 4592
rect 9858 4572 9867 4592
rect 9684 4561 9715 4562
rect 9679 4493 9789 4506
rect 9830 4493 9867 4572
rect 10142 4517 10207 4656
rect 11398 4645 11408 4682
rect 11448 4674 11463 4682
rect 11676 4675 11707 4728
rect 11737 4757 11774 4836
rect 11889 4767 11920 4768
rect 11737 4737 11746 4757
rect 11766 4737 11774 4757
rect 11737 4727 11774 4737
rect 11833 4760 11920 4767
rect 11833 4757 11894 4760
rect 11833 4737 11842 4757
rect 11862 4740 11894 4757
rect 11915 4740 11920 4760
rect 11862 4737 11920 4740
rect 11833 4730 11920 4737
rect 11945 4757 11982 4899
rect 12248 4898 12285 4899
rect 12097 4767 12133 4768
rect 11945 4737 11954 4757
rect 11974 4737 11982 4757
rect 11833 4728 11889 4730
rect 11833 4727 11870 4728
rect 11945 4727 11982 4737
rect 12041 4757 12189 4767
rect 12289 4764 12385 4766
rect 12041 4737 12050 4757
rect 12070 4737 12160 4757
rect 12180 4737 12189 4757
rect 12041 4731 12189 4737
rect 12041 4728 12105 4731
rect 12041 4727 12078 4728
rect 12097 4701 12105 4728
rect 12126 4728 12189 4731
rect 12247 4757 12385 4764
rect 12247 4737 12256 4757
rect 12276 4737 12385 4757
rect 12247 4728 12385 4737
rect 12126 4701 12133 4728
rect 12152 4727 12189 4728
rect 12248 4727 12285 4728
rect 12097 4676 12133 4701
rect 11568 4674 11609 4675
rect 11448 4667 11609 4674
rect 11448 4647 11578 4667
rect 11598 4647 11609 4667
rect 11448 4645 11609 4647
rect 11398 4639 11609 4645
rect 11676 4671 12035 4675
rect 11676 4666 11998 4671
rect 11676 4642 11789 4666
rect 11813 4647 11998 4666
rect 12022 4647 12035 4671
rect 11813 4642 12035 4647
rect 11676 4639 12035 4642
rect 12097 4639 12132 4676
rect 12200 4673 12300 4676
rect 12200 4669 12267 4673
rect 12200 4643 12212 4669
rect 12238 4647 12267 4669
rect 12293 4647 12300 4673
rect 12238 4643 12300 4647
rect 12200 4639 12300 4643
rect 11398 4626 11465 4639
rect 10142 4511 10164 4517
rect 9617 4491 9867 4493
rect 9617 4488 9718 4491
rect 9617 4469 9682 4488
rect 9679 4461 9682 4469
rect 9711 4461 9718 4488
rect 9746 4464 9756 4491
rect 9785 4469 9867 4491
rect 9896 4499 10164 4511
rect 10182 4499 10207 4517
rect 9896 4476 10207 4499
rect 11190 4603 11246 4623
rect 11190 4585 11209 4603
rect 11227 4585 11246 4603
rect 9896 4475 9951 4476
rect 9785 4464 9789 4469
rect 9746 4461 9789 4464
rect 9679 4447 9789 4461
rect 9105 4429 9446 4430
rect 7982 4408 7985 4428
rect 8005 4408 8398 4428
rect 9030 4428 9446 4429
rect 9896 4428 9939 4475
rect 11190 4472 11246 4585
rect 11398 4605 11412 4626
rect 11448 4605 11465 4626
rect 11676 4618 11707 4639
rect 12097 4618 12133 4639
rect 11519 4617 11556 4618
rect 11398 4598 11465 4605
rect 11518 4608 11556 4617
rect 9030 4424 9939 4428
rect 8349 4375 8394 4408
rect 9030 4404 9033 4424
rect 9053 4404 9939 4424
rect 9407 4399 9939 4404
rect 10147 4418 10206 4440
rect 10147 4400 10166 4418
rect 10184 4400 10206 4418
rect 9195 4375 9294 4377
rect 8349 4365 9294 4375
rect 8349 4339 9217 4365
rect 8350 4338 9217 4339
rect 9195 4327 9217 4338
rect 9242 4330 9261 4365
rect 9286 4330 9294 4365
rect 9242 4327 9294 4330
rect 9195 4319 9294 4327
rect 9221 4318 9293 4319
rect 10147 4270 10206 4400
rect 11190 4343 11245 4472
rect 11398 4446 11463 4598
rect 11518 4588 11527 4608
rect 11547 4588 11556 4608
rect 11518 4580 11556 4588
rect 11622 4612 11707 4618
rect 11732 4617 11769 4618
rect 11622 4592 11630 4612
rect 11650 4592 11707 4612
rect 11622 4584 11707 4592
rect 11731 4608 11769 4617
rect 11731 4588 11740 4608
rect 11760 4588 11769 4608
rect 11622 4583 11658 4584
rect 11731 4580 11769 4588
rect 11835 4612 11920 4618
rect 11940 4617 11977 4618
rect 11835 4592 11843 4612
rect 11863 4611 11920 4612
rect 11863 4592 11892 4611
rect 11835 4591 11892 4592
rect 11913 4591 11920 4611
rect 11835 4584 11920 4591
rect 11939 4608 11977 4617
rect 11939 4588 11948 4608
rect 11968 4588 11977 4608
rect 11835 4583 11871 4584
rect 11939 4580 11977 4588
rect 12043 4612 12187 4618
rect 12043 4592 12051 4612
rect 12071 4592 12159 4612
rect 12179 4592 12187 4612
rect 12043 4584 12187 4592
rect 12043 4583 12079 4584
rect 12151 4583 12187 4584
rect 12253 4617 12290 4618
rect 12253 4616 12291 4617
rect 12253 4608 12317 4616
rect 12253 4588 12262 4608
rect 12282 4594 12317 4608
rect 12337 4594 12340 4614
rect 12282 4589 12340 4594
rect 12282 4588 12317 4589
rect 11519 4551 11556 4580
rect 11520 4549 11556 4551
rect 11732 4549 11769 4580
rect 11520 4527 11769 4549
rect 11601 4521 11712 4527
rect 11601 4513 11642 4521
rect 11601 4493 11609 4513
rect 11628 4493 11642 4513
rect 11601 4491 11642 4493
rect 11670 4513 11712 4521
rect 11670 4493 11686 4513
rect 11705 4493 11712 4513
rect 11670 4491 11712 4493
rect 11601 4476 11712 4491
rect 11940 4481 11977 4580
rect 12253 4576 12317 4588
rect 11603 4467 11707 4476
rect 11391 4436 11512 4446
rect 11391 4434 11460 4436
rect 11391 4393 11404 4434
rect 11441 4395 11460 4434
rect 11497 4395 11512 4436
rect 11441 4393 11512 4395
rect 11391 4375 11512 4393
rect 11184 4331 11245 4343
rect 11938 4331 11979 4481
rect 12357 4473 12384 4728
rect 12446 4718 12526 4729
rect 12446 4692 12463 4718
rect 12503 4692 12526 4718
rect 12446 4665 12526 4692
rect 12446 4639 12467 4665
rect 12507 4639 12526 4665
rect 12446 4620 12526 4639
rect 12446 4594 12470 4620
rect 12510 4594 12526 4620
rect 12446 4543 12526 4594
rect 11184 4328 11979 4331
rect 12358 4342 12384 4473
rect 12448 4387 12518 4543
rect 12447 4371 12523 4387
rect 12358 4328 12386 4342
rect 11184 4293 12386 4328
rect 12447 4334 12462 4371
rect 12506 4334 12523 4371
rect 12447 4314 12523 4334
rect 13561 4364 13631 5273
rect 13730 4752 13811 5421
rect 14635 5316 14671 5616
rect 14559 5287 14672 5316
rect 14559 4922 14590 5287
rect 14483 4902 14876 4922
rect 14896 4902 14899 4922
rect 14483 4897 14899 4902
rect 14483 4896 14824 4897
rect 14140 4865 14250 4879
rect 14140 4862 14183 4865
rect 14140 4857 14144 4862
rect 14062 4835 14144 4857
rect 14173 4835 14183 4862
rect 14211 4838 14218 4865
rect 14247 4857 14250 4865
rect 14247 4838 14312 4857
rect 14211 4835 14312 4838
rect 14062 4833 14312 4835
rect 14062 4754 14099 4833
rect 14140 4820 14250 4833
rect 14214 4764 14245 4765
rect 13724 4672 13823 4752
rect 14062 4734 14071 4754
rect 14091 4734 14099 4754
rect 14062 4724 14099 4734
rect 14158 4754 14245 4764
rect 14158 4734 14167 4754
rect 14187 4734 14245 4754
rect 14158 4725 14245 4734
rect 14158 4724 14195 4725
rect 14214 4672 14245 4725
rect 14275 4754 14312 4833
rect 14427 4764 14458 4765
rect 14275 4734 14284 4754
rect 14304 4734 14312 4754
rect 14275 4724 14312 4734
rect 14371 4757 14458 4764
rect 14371 4754 14432 4757
rect 14371 4734 14380 4754
rect 14400 4737 14432 4754
rect 14453 4737 14458 4757
rect 14400 4734 14458 4737
rect 14371 4727 14458 4734
rect 14483 4754 14520 4896
rect 14786 4895 14823 4896
rect 14635 4764 14671 4765
rect 14483 4734 14492 4754
rect 14512 4734 14520 4754
rect 14371 4725 14427 4727
rect 14371 4724 14408 4725
rect 14483 4724 14520 4734
rect 14579 4754 14727 4764
rect 14827 4761 14923 4763
rect 14579 4734 14588 4754
rect 14608 4734 14698 4754
rect 14718 4734 14727 4754
rect 14579 4728 14727 4734
rect 14579 4725 14643 4728
rect 14579 4724 14616 4725
rect 14635 4698 14643 4725
rect 14664 4725 14727 4728
rect 14785 4754 14923 4761
rect 14785 4734 14794 4754
rect 14814 4734 14923 4754
rect 14785 4725 14923 4734
rect 14664 4698 14671 4725
rect 14690 4724 14727 4725
rect 14786 4724 14823 4725
rect 14635 4673 14671 4698
rect 13724 4671 14064 4672
rect 14106 4671 14147 4672
rect 13724 4664 14147 4671
rect 13724 4644 14116 4664
rect 14136 4644 14147 4664
rect 13724 4636 14147 4644
rect 14214 4668 14573 4672
rect 14214 4663 14536 4668
rect 14214 4639 14327 4663
rect 14351 4644 14536 4663
rect 14560 4644 14573 4668
rect 14351 4639 14573 4644
rect 14214 4636 14573 4639
rect 14635 4636 14670 4673
rect 14738 4670 14838 4673
rect 14738 4666 14805 4670
rect 14738 4640 14750 4666
rect 14776 4644 14805 4666
rect 14831 4644 14838 4670
rect 14776 4640 14838 4644
rect 14738 4636 14838 4640
rect 13724 4632 14064 4636
rect 13561 4314 13633 4364
rect 8869 4240 8945 4264
rect 8869 4174 8881 4240
rect 8935 4174 8945 4240
rect 9413 4195 9454 4197
rect 9685 4195 9789 4197
rect 10147 4195 10208 4270
rect 11184 4218 11245 4293
rect 11603 4291 11707 4293
rect 11938 4291 11979 4293
rect 12447 4248 12457 4314
rect 12511 4248 12523 4314
rect 12447 4224 12523 4248
rect 7759 4124 7831 4174
rect 7328 3852 7664 3856
rect 6554 3848 6654 3852
rect 6554 3844 6616 3848
rect 6554 3818 6561 3844
rect 6587 3822 6616 3844
rect 6642 3822 6654 3848
rect 6587 3818 6654 3822
rect 6554 3815 6654 3818
rect 6722 3815 6757 3852
rect 6819 3849 7178 3852
rect 6819 3844 7041 3849
rect 6819 3820 6832 3844
rect 6856 3825 7041 3844
rect 7065 3825 7178 3849
rect 6856 3820 7178 3825
rect 6819 3816 7178 3820
rect 7245 3844 7664 3852
rect 7245 3824 7256 3844
rect 7276 3824 7664 3844
rect 7245 3817 7664 3824
rect 7245 3816 7286 3817
rect 7328 3816 7664 3817
rect 6721 3790 6757 3815
rect 6569 3763 6606 3764
rect 6665 3763 6702 3764
rect 6721 3763 6728 3790
rect 6469 3754 6607 3763
rect 6469 3734 6578 3754
rect 6598 3734 6607 3754
rect 6469 3727 6607 3734
rect 6665 3760 6728 3763
rect 6749 3763 6757 3790
rect 6776 3763 6813 3764
rect 6749 3760 6813 3763
rect 6665 3754 6813 3760
rect 6665 3734 6674 3754
rect 6694 3734 6784 3754
rect 6804 3734 6813 3754
rect 6469 3725 6565 3727
rect 6665 3724 6813 3734
rect 6872 3754 6909 3764
rect 6984 3763 7021 3764
rect 6965 3761 7021 3763
rect 6872 3734 6880 3754
rect 6900 3734 6909 3754
rect 6721 3723 6757 3724
rect 6569 3592 6606 3593
rect 6872 3592 6909 3734
rect 6934 3754 7021 3761
rect 6934 3751 6992 3754
rect 6934 3731 6939 3751
rect 6960 3734 6992 3751
rect 7012 3734 7021 3754
rect 6960 3731 7021 3734
rect 6934 3724 7021 3731
rect 7080 3754 7117 3764
rect 7080 3734 7088 3754
rect 7108 3734 7117 3754
rect 6934 3723 6965 3724
rect 7080 3655 7117 3734
rect 7147 3763 7178 3816
rect 7572 3780 7664 3816
rect 7197 3763 7234 3764
rect 7147 3754 7234 3763
rect 7147 3734 7205 3754
rect 7225 3734 7234 3754
rect 7147 3724 7234 3734
rect 7293 3754 7330 3764
rect 7293 3734 7301 3754
rect 7321 3734 7330 3754
rect 7147 3723 7178 3724
rect 7142 3655 7252 3668
rect 7293 3655 7330 3734
rect 7080 3653 7330 3655
rect 7080 3650 7181 3653
rect 7080 3631 7145 3650
rect 7142 3623 7145 3631
rect 7174 3623 7181 3650
rect 7209 3626 7219 3653
rect 7248 3631 7330 3653
rect 7248 3626 7252 3631
rect 7209 3623 7252 3626
rect 7142 3609 7252 3623
rect 6568 3591 6909 3592
rect 6493 3586 6909 3591
rect 6493 3566 6496 3586
rect 6516 3566 6909 3586
rect 6653 3522 6758 3525
rect 6652 3499 6758 3522
rect 5772 3497 6273 3499
rect 6414 3497 6763 3499
rect 3886 3476 3923 3497
rect 3886 3439 3897 3476
rect 3914 3439 3923 3476
rect 5772 3491 6763 3497
rect 5772 3486 6724 3491
rect 5772 3465 6683 3486
rect 6703 3470 6724 3486
rect 6744 3470 6763 3491
rect 6703 3465 6763 3470
rect 5772 3440 6763 3465
rect 6248 3439 6430 3440
rect 3886 3429 3923 3439
rect 3732 3386 4126 3406
rect 4146 3386 4149 3406
rect 3733 3381 4149 3386
rect 3733 3380 4074 3381
rect 3390 3349 3500 3363
rect 3390 3346 3433 3349
rect 3390 3341 3394 3346
rect 3312 3319 3394 3341
rect 3423 3319 3433 3346
rect 3461 3322 3468 3349
rect 3497 3341 3500 3349
rect 3497 3322 3562 3341
rect 3461 3319 3562 3322
rect 3312 3317 3562 3319
rect 3312 3238 3349 3317
rect 3390 3304 3500 3317
rect 3464 3248 3495 3249
rect 3312 3218 3321 3238
rect 3341 3218 3349 3238
rect 3312 3208 3349 3218
rect 3408 3238 3495 3248
rect 3408 3218 3417 3238
rect 3437 3218 3495 3238
rect 3408 3209 3495 3218
rect 3408 3208 3445 3209
rect 3464 3156 3495 3209
rect 3525 3238 3562 3317
rect 3677 3248 3708 3249
rect 3525 3218 3534 3238
rect 3554 3218 3562 3238
rect 3525 3208 3562 3218
rect 3621 3241 3708 3248
rect 3621 3238 3682 3241
rect 3621 3218 3630 3238
rect 3650 3221 3682 3238
rect 3703 3221 3708 3241
rect 3650 3218 3708 3221
rect 3621 3211 3708 3218
rect 3733 3238 3770 3380
rect 4036 3379 4073 3380
rect 3885 3248 3921 3249
rect 3733 3218 3742 3238
rect 3762 3218 3770 3238
rect 3621 3209 3677 3211
rect 3621 3208 3658 3209
rect 3733 3208 3770 3218
rect 3829 3238 3977 3248
rect 4077 3245 4173 3247
rect 3829 3218 3838 3238
rect 3858 3218 3948 3238
rect 3968 3218 3977 3238
rect 3829 3212 3977 3218
rect 3829 3209 3893 3212
rect 3829 3208 3866 3209
rect 3885 3182 3893 3209
rect 3914 3209 3977 3212
rect 4035 3238 4173 3245
rect 4035 3218 4044 3238
rect 4064 3218 4173 3238
rect 4035 3209 4173 3218
rect 6802 3210 6833 3566
rect 3914 3182 3921 3209
rect 3940 3208 3977 3209
rect 4036 3208 4073 3209
rect 3885 3157 3921 3182
rect 3356 3155 3397 3156
rect 3276 3150 3397 3155
rect 3227 3148 3397 3150
rect 3227 3137 3366 3148
rect 3227 3114 3250 3137
rect 3276 3128 3366 3137
rect 3386 3128 3397 3148
rect 3276 3120 3397 3128
rect 3464 3152 3823 3156
rect 3464 3147 3786 3152
rect 3464 3123 3577 3147
rect 3601 3128 3786 3147
rect 3810 3128 3823 3152
rect 3601 3123 3823 3128
rect 3464 3120 3823 3123
rect 3885 3120 3920 3157
rect 3988 3154 4088 3157
rect 3988 3150 4055 3154
rect 3988 3124 4000 3150
rect 4026 3128 4055 3150
rect 4081 3128 4088 3154
rect 4026 3124 4088 3128
rect 3988 3120 4088 3124
rect 3276 3114 3284 3120
rect 3227 3106 3284 3114
rect 3464 3099 3495 3120
rect 3885 3099 3921 3120
rect 3307 3098 3344 3099
rect 3306 3089 3344 3098
rect 3306 3069 3315 3089
rect 3335 3069 3344 3089
rect 3306 3061 3344 3069
rect 3410 3093 3495 3099
rect 3520 3098 3557 3099
rect 3410 3073 3418 3093
rect 3438 3073 3495 3093
rect 3410 3065 3495 3073
rect 3519 3089 3557 3098
rect 3519 3069 3528 3089
rect 3548 3069 3557 3089
rect 3410 3064 3446 3065
rect 3519 3061 3557 3069
rect 3623 3093 3708 3099
rect 3728 3098 3765 3099
rect 3623 3073 3631 3093
rect 3651 3092 3708 3093
rect 3651 3073 3680 3092
rect 3623 3072 3680 3073
rect 3701 3072 3708 3092
rect 3623 3065 3708 3072
rect 3727 3089 3765 3098
rect 3727 3069 3736 3089
rect 3756 3069 3765 3089
rect 3623 3064 3659 3065
rect 3727 3061 3765 3069
rect 3831 3093 3975 3099
rect 3831 3073 3839 3093
rect 3859 3073 3947 3093
rect 3967 3073 3975 3093
rect 3831 3065 3975 3073
rect 3831 3064 3867 3065
rect 3939 3064 3975 3065
rect 4041 3098 4078 3099
rect 4041 3097 4079 3098
rect 4041 3089 4105 3097
rect 4041 3069 4050 3089
rect 4070 3075 4105 3089
rect 4125 3075 4128 3095
rect 4070 3070 4128 3075
rect 4070 3069 4105 3070
rect 3307 3032 3344 3061
rect 3308 3030 3344 3032
rect 3520 3030 3557 3061
rect 3308 3008 3557 3030
rect 3389 3002 3500 3008
rect 3389 2994 3430 3002
rect 3389 2974 3397 2994
rect 3416 2974 3430 2994
rect 3389 2972 3430 2974
rect 3458 2994 3500 3002
rect 3458 2974 3474 2994
rect 3493 2974 3500 2994
rect 3458 2972 3500 2974
rect 3389 2957 3500 2972
rect 3728 2946 3765 3061
rect 4041 3057 4105 3069
rect 3721 2940 3768 2946
rect 4145 2942 4172 3209
rect 6720 3181 6833 3210
rect 4004 2940 4172 2942
rect 3721 2914 4172 2940
rect 3721 2779 3768 2914
rect 4004 2913 4172 2914
rect 6721 2872 6757 3181
rect 7581 3067 7662 3780
rect 7761 3215 7831 4124
rect 8869 4154 8945 4174
rect 8869 4117 8886 4154
rect 8930 4117 8945 4154
rect 9006 4160 10208 4195
rect 9006 4146 9034 4160
rect 8869 4101 8945 4117
rect 8874 3945 8944 4101
rect 9008 4015 9034 4146
rect 9413 4157 10208 4160
rect 8866 3894 8946 3945
rect 8866 3868 8882 3894
rect 8922 3868 8946 3894
rect 8866 3849 8946 3868
rect 8866 3823 8885 3849
rect 8925 3823 8946 3849
rect 8866 3796 8946 3823
rect 8866 3770 8889 3796
rect 8929 3770 8946 3796
rect 8866 3759 8946 3770
rect 9008 3760 9035 4015
rect 9413 4007 9454 4157
rect 10147 4145 10208 4157
rect 9880 4095 10001 4113
rect 9880 4093 9951 4095
rect 9880 4052 9895 4093
rect 9932 4054 9951 4093
rect 9988 4054 10001 4095
rect 9932 4052 10001 4054
rect 9880 4042 10001 4052
rect 9685 4012 9789 4021
rect 9075 3900 9139 3912
rect 9415 3908 9452 4007
rect 9680 3997 9791 4012
rect 9680 3995 9722 3997
rect 9680 3975 9687 3995
rect 9706 3975 9722 3995
rect 9680 3967 9722 3975
rect 9750 3995 9791 3997
rect 9750 3975 9764 3995
rect 9783 3975 9791 3995
rect 9750 3967 9791 3975
rect 9680 3961 9791 3967
rect 9623 3939 9872 3961
rect 9623 3908 9660 3939
rect 9836 3937 9872 3939
rect 9836 3908 9873 3937
rect 9075 3899 9110 3900
rect 9052 3894 9110 3899
rect 9052 3874 9055 3894
rect 9075 3880 9110 3894
rect 9130 3880 9139 3900
rect 9075 3872 9139 3880
rect 9101 3871 9139 3872
rect 9102 3870 9139 3871
rect 9205 3904 9241 3905
rect 9313 3904 9349 3905
rect 9205 3896 9349 3904
rect 9205 3876 9213 3896
rect 9233 3876 9321 3896
rect 9341 3876 9349 3896
rect 9205 3870 9349 3876
rect 9415 3900 9453 3908
rect 9521 3904 9557 3905
rect 9415 3880 9424 3900
rect 9444 3880 9453 3900
rect 9415 3871 9453 3880
rect 9472 3897 9557 3904
rect 9472 3877 9479 3897
rect 9500 3896 9557 3897
rect 9500 3877 9529 3896
rect 9472 3876 9529 3877
rect 9549 3876 9557 3896
rect 9415 3870 9452 3871
rect 9472 3870 9557 3876
rect 9623 3900 9661 3908
rect 9734 3904 9770 3905
rect 9623 3880 9632 3900
rect 9652 3880 9661 3900
rect 9623 3871 9661 3880
rect 9685 3896 9770 3904
rect 9685 3876 9742 3896
rect 9762 3876 9770 3896
rect 9623 3870 9660 3871
rect 9685 3870 9770 3876
rect 9836 3900 9874 3908
rect 9836 3880 9845 3900
rect 9865 3880 9874 3900
rect 9929 3890 9994 4042
rect 10147 4016 10202 4145
rect 11186 4088 11245 4218
rect 12099 4169 12171 4170
rect 12098 4161 12197 4169
rect 12098 4158 12150 4161
rect 12098 4123 12106 4158
rect 12131 4123 12150 4158
rect 12175 4150 12197 4161
rect 12175 4149 13042 4150
rect 12175 4123 13043 4149
rect 12098 4113 13043 4123
rect 12098 4111 12197 4113
rect 11186 4070 11208 4088
rect 11226 4070 11245 4088
rect 11186 4048 11245 4070
rect 11453 4084 11985 4089
rect 11453 4064 12339 4084
rect 12359 4064 12362 4084
rect 12998 4080 13043 4113
rect 11453 4060 12362 4064
rect 9836 3871 9874 3880
rect 9927 3883 9994 3890
rect 9836 3870 9873 3871
rect 9259 3849 9295 3870
rect 9685 3849 9716 3870
rect 9927 3862 9944 3883
rect 9980 3862 9994 3883
rect 10146 3903 10202 4016
rect 11453 4013 11496 4060
rect 11946 4059 12362 4060
rect 12994 4060 13387 4080
rect 13407 4060 13410 4080
rect 11946 4058 12287 4059
rect 11603 4027 11713 4041
rect 11603 4024 11646 4027
rect 11603 4019 11607 4024
rect 11441 4012 11496 4013
rect 10146 3885 10165 3903
rect 10183 3885 10202 3903
rect 10146 3865 10202 3885
rect 11185 3989 11496 4012
rect 11185 3971 11210 3989
rect 11228 3977 11496 3989
rect 11525 3997 11607 4019
rect 11636 3997 11646 4024
rect 11674 4000 11681 4027
rect 11710 4019 11713 4027
rect 11710 4000 11775 4019
rect 11674 3997 11775 4000
rect 11525 3995 11775 3997
rect 11228 3971 11250 3977
rect 9927 3849 9994 3862
rect 9092 3845 9192 3849
rect 9092 3841 9154 3845
rect 9092 3815 9099 3841
rect 9125 3819 9154 3841
rect 9180 3819 9192 3845
rect 9125 3815 9192 3819
rect 9092 3812 9192 3815
rect 9260 3812 9295 3849
rect 9357 3846 9716 3849
rect 9357 3841 9579 3846
rect 9357 3817 9370 3841
rect 9394 3822 9579 3841
rect 9603 3822 9716 3846
rect 9394 3817 9716 3822
rect 9357 3813 9716 3817
rect 9783 3843 9994 3849
rect 9783 3841 9944 3843
rect 9783 3821 9794 3841
rect 9814 3821 9944 3841
rect 9783 3814 9944 3821
rect 9783 3813 9824 3814
rect 9259 3787 9295 3812
rect 9107 3760 9144 3761
rect 9203 3760 9240 3761
rect 9259 3760 9266 3787
rect 9007 3751 9145 3760
rect 9007 3731 9116 3751
rect 9136 3731 9145 3751
rect 9007 3724 9145 3731
rect 9203 3757 9266 3760
rect 9287 3760 9295 3787
rect 9314 3760 9351 3761
rect 9287 3757 9351 3760
rect 9203 3751 9351 3757
rect 9203 3731 9212 3751
rect 9232 3731 9322 3751
rect 9342 3731 9351 3751
rect 9007 3722 9103 3724
rect 9203 3721 9351 3731
rect 9410 3751 9447 3761
rect 9522 3760 9559 3761
rect 9503 3758 9559 3760
rect 9410 3731 9418 3751
rect 9438 3731 9447 3751
rect 9259 3720 9295 3721
rect 9107 3589 9144 3590
rect 9410 3589 9447 3731
rect 9472 3751 9559 3758
rect 9472 3748 9530 3751
rect 9472 3728 9477 3748
rect 9498 3731 9530 3748
rect 9550 3731 9559 3751
rect 9498 3728 9559 3731
rect 9472 3721 9559 3728
rect 9618 3751 9655 3761
rect 9618 3731 9626 3751
rect 9646 3731 9655 3751
rect 9472 3720 9503 3721
rect 9618 3652 9655 3731
rect 9685 3760 9716 3813
rect 9929 3806 9944 3814
rect 9984 3806 9994 3843
rect 11185 3832 11250 3971
rect 11525 3916 11562 3995
rect 11603 3982 11713 3995
rect 11677 3926 11708 3927
rect 11525 3896 11534 3916
rect 11554 3896 11562 3916
rect 9929 3797 9994 3806
rect 10142 3804 10207 3825
rect 10142 3786 10167 3804
rect 10185 3786 10207 3804
rect 11185 3814 11208 3832
rect 11226 3814 11250 3832
rect 11185 3797 11250 3814
rect 11405 3878 11473 3891
rect 11525 3886 11562 3896
rect 11621 3916 11708 3926
rect 11621 3896 11630 3916
rect 11650 3896 11708 3916
rect 11621 3887 11708 3896
rect 11621 3886 11658 3887
rect 11405 3836 11412 3878
rect 11461 3836 11473 3878
rect 11405 3833 11473 3836
rect 11677 3834 11708 3887
rect 11738 3916 11775 3995
rect 11890 3926 11921 3927
rect 11738 3896 11747 3916
rect 11767 3896 11775 3916
rect 11738 3886 11775 3896
rect 11834 3919 11921 3926
rect 11834 3916 11895 3919
rect 11834 3896 11843 3916
rect 11863 3899 11895 3916
rect 11916 3899 11921 3919
rect 11863 3896 11921 3899
rect 11834 3889 11921 3896
rect 11946 3916 11983 4058
rect 12249 4057 12286 4058
rect 12994 4055 13410 4060
rect 12994 4054 13335 4055
rect 12651 4023 12761 4037
rect 12651 4020 12694 4023
rect 12651 4015 12655 4020
rect 12573 3993 12655 4015
rect 12684 3993 12694 4020
rect 12722 3996 12729 4023
rect 12758 4015 12761 4023
rect 12758 3996 12823 4015
rect 12722 3993 12823 3996
rect 12573 3991 12823 3993
rect 12098 3926 12134 3927
rect 11946 3896 11955 3916
rect 11975 3896 11983 3916
rect 11834 3887 11890 3889
rect 11834 3886 11871 3887
rect 11946 3886 11983 3896
rect 12042 3916 12190 3926
rect 12290 3923 12386 3925
rect 12042 3896 12051 3916
rect 12071 3896 12161 3916
rect 12181 3896 12190 3916
rect 12042 3890 12190 3896
rect 12042 3887 12106 3890
rect 12042 3886 12079 3887
rect 12098 3860 12106 3887
rect 12127 3887 12190 3890
rect 12248 3916 12386 3923
rect 12248 3896 12257 3916
rect 12277 3896 12386 3916
rect 12248 3887 12386 3896
rect 12573 3912 12610 3991
rect 12651 3978 12761 3991
rect 12725 3922 12756 3923
rect 12573 3892 12582 3912
rect 12602 3892 12610 3912
rect 12127 3860 12134 3887
rect 12153 3886 12190 3887
rect 12249 3886 12286 3887
rect 12098 3835 12134 3860
rect 11569 3833 11610 3834
rect 11405 3826 11610 3833
rect 11405 3815 11579 3826
rect 9735 3760 9772 3761
rect 9685 3751 9772 3760
rect 9685 3731 9743 3751
rect 9763 3731 9772 3751
rect 9685 3721 9772 3731
rect 9831 3751 9868 3761
rect 9831 3731 9839 3751
rect 9859 3731 9868 3751
rect 9685 3720 9716 3721
rect 9680 3652 9790 3665
rect 9831 3652 9868 3731
rect 10142 3710 10207 3786
rect 11405 3782 11413 3815
rect 11406 3773 11413 3782
rect 11462 3806 11579 3815
rect 11599 3806 11610 3826
rect 11462 3798 11610 3806
rect 11677 3830 12036 3834
rect 11677 3825 11999 3830
rect 11677 3801 11790 3825
rect 11814 3806 11999 3825
rect 12023 3806 12036 3830
rect 11814 3801 12036 3806
rect 11677 3798 12036 3801
rect 12098 3798 12133 3835
rect 12201 3832 12301 3835
rect 12201 3828 12268 3832
rect 12201 3802 12213 3828
rect 12239 3806 12268 3828
rect 12294 3806 12301 3832
rect 12239 3802 12301 3806
rect 12201 3798 12301 3802
rect 11462 3782 11473 3798
rect 11462 3773 11470 3782
rect 11677 3777 11708 3798
rect 12098 3777 12134 3798
rect 11520 3776 11557 3777
rect 11185 3733 11250 3752
rect 11185 3715 11210 3733
rect 11228 3715 11250 3733
rect 9618 3650 9868 3652
rect 9618 3647 9719 3650
rect 9618 3628 9683 3647
rect 9680 3620 9683 3628
rect 9712 3620 9719 3647
rect 9747 3623 9757 3650
rect 9786 3628 9868 3650
rect 9891 3675 10208 3710
rect 9786 3623 9790 3628
rect 9747 3620 9790 3623
rect 9680 3606 9790 3620
rect 9106 3588 9447 3589
rect 9031 3586 9447 3588
rect 9891 3586 9931 3675
rect 10142 3648 10207 3675
rect 10142 3630 10165 3648
rect 10183 3630 10207 3648
rect 10142 3610 10207 3630
rect 9028 3583 9931 3586
rect 9028 3563 9034 3583
rect 9054 3563 9931 3583
rect 9028 3559 9931 3563
rect 9891 3556 9931 3559
rect 10143 3549 10208 3570
rect 8361 3541 9022 3542
rect 8361 3534 9295 3541
rect 8361 3533 9267 3534
rect 8361 3513 9212 3533
rect 9244 3514 9267 3533
rect 9292 3514 9295 3534
rect 9244 3513 9295 3514
rect 8361 3506 9295 3513
rect 7960 3464 8128 3465
rect 8363 3464 8402 3506
rect 9191 3504 9295 3506
rect 9260 3502 9295 3504
rect 10143 3531 10167 3549
rect 10185 3531 10208 3549
rect 10143 3484 10208 3531
rect 7960 3438 8404 3464
rect 7960 3436 8128 3438
rect 6721 2849 6725 2872
rect 6749 2849 6757 2872
rect 6921 2850 7020 2854
rect 6721 2828 6757 2849
rect 6721 2805 6725 2828
rect 6749 2805 6757 2828
rect 6721 2801 6757 2805
rect 6917 2844 7020 2850
rect 6917 2806 6943 2844
rect 6968 2809 6987 2844
rect 7012 2809 7020 2844
rect 6968 2806 7020 2809
rect 6917 2798 7020 2806
rect 6917 2797 7019 2798
rect 3719 2730 3778 2779
rect 3719 2702 3737 2730
rect 3765 2702 3778 2730
rect 3719 2692 3778 2702
rect 6513 2719 6681 2720
rect 6917 2719 6964 2797
rect 6513 2693 6964 2719
rect 6513 2691 6681 2693
rect 6513 2318 6540 2691
rect 6710 2643 6796 2652
rect 6710 2625 6729 2643
rect 6781 2625 6796 2643
rect 6710 2621 6796 2625
rect 6580 2458 6644 2470
rect 6580 2457 6615 2458
rect 6557 2452 6615 2457
rect 6557 2432 6560 2452
rect 6580 2438 6615 2452
rect 6635 2438 6644 2458
rect 6580 2430 6644 2438
rect 6606 2429 6644 2430
rect 6607 2428 6644 2429
rect 6710 2462 6746 2463
rect 6766 2462 6796 2621
rect 6917 2581 6964 2693
rect 6920 2466 6957 2581
rect 7185 2555 7296 2570
rect 7185 2553 7227 2555
rect 7185 2533 7192 2553
rect 7211 2533 7227 2553
rect 7185 2525 7227 2533
rect 7255 2553 7296 2555
rect 7255 2533 7269 2553
rect 7288 2533 7296 2553
rect 7255 2525 7296 2533
rect 7185 2519 7296 2525
rect 7128 2497 7377 2519
rect 7128 2466 7165 2497
rect 7341 2495 7377 2497
rect 7341 2466 7378 2495
rect 7582 2482 7661 3067
rect 7758 2615 7837 3215
rect 7960 3085 7987 3436
rect 8363 3432 8404 3438
rect 8027 3225 8091 3237
rect 8367 3233 8404 3432
rect 8866 3459 8938 3476
rect 8866 3420 8874 3459
rect 8919 3420 8938 3459
rect 8632 3322 8743 3337
rect 8632 3320 8674 3322
rect 8632 3300 8639 3320
rect 8658 3300 8674 3320
rect 8632 3292 8674 3300
rect 8702 3320 8743 3322
rect 8702 3300 8716 3320
rect 8735 3300 8743 3320
rect 8702 3292 8743 3300
rect 8632 3286 8743 3292
rect 8575 3264 8824 3286
rect 8575 3233 8612 3264
rect 8788 3262 8824 3264
rect 8788 3233 8825 3262
rect 8027 3224 8062 3225
rect 8004 3219 8062 3224
rect 8004 3199 8007 3219
rect 8027 3205 8062 3219
rect 8082 3205 8091 3225
rect 8027 3197 8091 3205
rect 8053 3196 8091 3197
rect 8054 3195 8091 3196
rect 8157 3229 8193 3230
rect 8265 3229 8301 3230
rect 8157 3221 8301 3229
rect 8157 3201 8165 3221
rect 8185 3201 8273 3221
rect 8293 3201 8301 3221
rect 8157 3195 8301 3201
rect 8367 3225 8405 3233
rect 8473 3229 8509 3230
rect 8367 3205 8376 3225
rect 8396 3205 8405 3225
rect 8367 3196 8405 3205
rect 8424 3222 8509 3229
rect 8424 3202 8431 3222
rect 8452 3221 8509 3222
rect 8452 3202 8481 3221
rect 8424 3201 8481 3202
rect 8501 3201 8509 3221
rect 8367 3195 8404 3196
rect 8424 3195 8509 3201
rect 8575 3225 8613 3233
rect 8686 3229 8722 3230
rect 8575 3205 8584 3225
rect 8604 3205 8613 3225
rect 8575 3196 8613 3205
rect 8637 3221 8722 3229
rect 8637 3201 8694 3221
rect 8714 3201 8722 3221
rect 8575 3195 8612 3196
rect 8637 3195 8722 3201
rect 8788 3225 8826 3233
rect 8788 3205 8797 3225
rect 8817 3205 8826 3225
rect 8788 3196 8826 3205
rect 8866 3210 8938 3420
rect 9008 3454 10208 3484
rect 9008 3453 9452 3454
rect 9008 3451 9176 3453
rect 8866 3196 8949 3210
rect 8788 3195 8825 3196
rect 8211 3174 8247 3195
rect 8637 3174 8668 3195
rect 8866 3174 8883 3196
rect 8044 3170 8144 3174
rect 8044 3166 8106 3170
rect 8044 3140 8051 3166
rect 8077 3144 8106 3166
rect 8132 3144 8144 3170
rect 8077 3140 8144 3144
rect 8044 3137 8144 3140
rect 8212 3137 8247 3174
rect 8309 3171 8668 3174
rect 8309 3166 8531 3171
rect 8309 3142 8322 3166
rect 8346 3147 8531 3166
rect 8555 3147 8668 3171
rect 8346 3142 8668 3147
rect 8309 3138 8668 3142
rect 8735 3166 8883 3174
rect 8735 3146 8746 3166
rect 8766 3163 8883 3166
rect 8936 3163 8949 3196
rect 8766 3146 8949 3163
rect 8735 3139 8949 3146
rect 8735 3138 8776 3139
rect 8866 3138 8949 3139
rect 8211 3112 8247 3137
rect 8059 3085 8096 3086
rect 8155 3085 8192 3086
rect 8211 3085 8218 3112
rect 7959 3076 8097 3085
rect 7959 3056 8068 3076
rect 8088 3056 8097 3076
rect 7959 3049 8097 3056
rect 8155 3082 8218 3085
rect 8239 3085 8247 3112
rect 8266 3085 8303 3086
rect 8239 3082 8303 3085
rect 8155 3076 8303 3082
rect 8155 3056 8164 3076
rect 8184 3056 8274 3076
rect 8294 3056 8303 3076
rect 7959 3047 8055 3049
rect 8155 3046 8303 3056
rect 8362 3076 8399 3086
rect 8474 3085 8511 3086
rect 8455 3083 8511 3085
rect 8362 3056 8370 3076
rect 8390 3056 8399 3076
rect 8211 3045 8247 3046
rect 8059 2914 8096 2915
rect 8362 2914 8399 3056
rect 8424 3076 8511 3083
rect 8424 3073 8482 3076
rect 8424 3053 8429 3073
rect 8450 3056 8482 3073
rect 8502 3056 8511 3076
rect 8450 3053 8511 3056
rect 8424 3046 8511 3053
rect 8570 3076 8607 3086
rect 8570 3056 8578 3076
rect 8598 3056 8607 3076
rect 8424 3045 8455 3046
rect 8570 2977 8607 3056
rect 8637 3085 8668 3138
rect 8874 3105 8888 3138
rect 8941 3105 8949 3138
rect 8874 3099 8949 3105
rect 8874 3094 8944 3099
rect 8687 3085 8724 3086
rect 8637 3076 8724 3085
rect 8637 3056 8695 3076
rect 8715 3056 8724 3076
rect 8637 3046 8724 3056
rect 8783 3076 8820 3086
rect 9008 3081 9035 3451
rect 9075 3221 9139 3233
rect 9415 3229 9452 3453
rect 9923 3434 9987 3436
rect 9919 3422 9987 3434
rect 9919 3389 9930 3422
rect 9970 3389 9987 3422
rect 9919 3379 9987 3389
rect 9680 3318 9791 3333
rect 9680 3316 9722 3318
rect 9680 3296 9687 3316
rect 9706 3296 9722 3316
rect 9680 3288 9722 3296
rect 9750 3316 9791 3318
rect 9750 3296 9764 3316
rect 9783 3296 9791 3316
rect 9750 3288 9791 3296
rect 9680 3282 9791 3288
rect 9623 3260 9872 3282
rect 9623 3229 9660 3260
rect 9836 3258 9872 3260
rect 9836 3229 9873 3258
rect 9075 3220 9110 3221
rect 9052 3215 9110 3220
rect 9052 3195 9055 3215
rect 9075 3201 9110 3215
rect 9130 3201 9139 3221
rect 9075 3193 9139 3201
rect 9101 3192 9139 3193
rect 9102 3191 9139 3192
rect 9205 3225 9241 3226
rect 9313 3225 9349 3226
rect 9205 3217 9349 3225
rect 9205 3197 9213 3217
rect 9233 3197 9321 3217
rect 9341 3197 9349 3217
rect 9205 3191 9349 3197
rect 9415 3221 9453 3229
rect 9521 3225 9557 3226
rect 9415 3201 9424 3221
rect 9444 3201 9453 3221
rect 9415 3192 9453 3201
rect 9472 3218 9557 3225
rect 9472 3198 9479 3218
rect 9500 3217 9557 3218
rect 9500 3198 9529 3217
rect 9472 3197 9529 3198
rect 9549 3197 9557 3217
rect 9415 3191 9452 3192
rect 9472 3191 9557 3197
rect 9623 3221 9661 3229
rect 9734 3225 9770 3226
rect 9623 3201 9632 3221
rect 9652 3201 9661 3221
rect 9623 3192 9661 3201
rect 9685 3217 9770 3225
rect 9685 3197 9742 3217
rect 9762 3197 9770 3217
rect 9623 3191 9660 3192
rect 9685 3191 9770 3197
rect 9836 3221 9874 3229
rect 9836 3201 9845 3221
rect 9865 3201 9874 3221
rect 9836 3192 9874 3201
rect 9923 3195 9987 3379
rect 10143 3253 10208 3454
rect 11185 3514 11250 3715
rect 11406 3589 11470 3773
rect 11519 3767 11557 3776
rect 11519 3747 11528 3767
rect 11548 3747 11557 3767
rect 11519 3739 11557 3747
rect 11623 3771 11708 3777
rect 11733 3776 11770 3777
rect 11623 3751 11631 3771
rect 11651 3751 11708 3771
rect 11623 3743 11708 3751
rect 11732 3767 11770 3776
rect 11732 3747 11741 3767
rect 11761 3747 11770 3767
rect 11623 3742 11659 3743
rect 11732 3739 11770 3747
rect 11836 3771 11921 3777
rect 11941 3776 11978 3777
rect 11836 3751 11844 3771
rect 11864 3770 11921 3771
rect 11864 3751 11893 3770
rect 11836 3750 11893 3751
rect 11914 3750 11921 3770
rect 11836 3743 11921 3750
rect 11940 3767 11978 3776
rect 11940 3747 11949 3767
rect 11969 3747 11978 3767
rect 11836 3742 11872 3743
rect 11940 3739 11978 3747
rect 12044 3771 12188 3777
rect 12044 3751 12052 3771
rect 12072 3751 12160 3771
rect 12180 3751 12188 3771
rect 12044 3743 12188 3751
rect 12044 3742 12080 3743
rect 12152 3742 12188 3743
rect 12254 3776 12291 3777
rect 12254 3775 12292 3776
rect 12254 3767 12318 3775
rect 12254 3747 12263 3767
rect 12283 3753 12318 3767
rect 12338 3753 12341 3773
rect 12283 3748 12341 3753
rect 12283 3747 12318 3748
rect 11520 3710 11557 3739
rect 11521 3708 11557 3710
rect 11733 3708 11770 3739
rect 11521 3686 11770 3708
rect 11602 3680 11713 3686
rect 11602 3672 11643 3680
rect 11602 3652 11610 3672
rect 11629 3652 11643 3672
rect 11602 3650 11643 3652
rect 11671 3672 11713 3680
rect 11671 3652 11687 3672
rect 11706 3652 11713 3672
rect 11671 3650 11713 3652
rect 11602 3635 11713 3650
rect 11406 3579 11474 3589
rect 11406 3546 11423 3579
rect 11463 3546 11474 3579
rect 11406 3534 11474 3546
rect 11406 3532 11470 3534
rect 11941 3515 11978 3739
rect 12254 3735 12318 3747
rect 12358 3517 12385 3887
rect 12573 3882 12610 3892
rect 12669 3912 12756 3922
rect 12669 3892 12678 3912
rect 12698 3892 12756 3912
rect 12669 3883 12756 3892
rect 12669 3882 12706 3883
rect 12449 3869 12519 3874
rect 12444 3863 12519 3869
rect 12444 3830 12452 3863
rect 12505 3830 12519 3863
rect 12725 3830 12756 3883
rect 12786 3912 12823 3991
rect 12938 3922 12969 3923
rect 12786 3892 12795 3912
rect 12815 3892 12823 3912
rect 12786 3882 12823 3892
rect 12882 3915 12969 3922
rect 12882 3912 12943 3915
rect 12882 3892 12891 3912
rect 12911 3895 12943 3912
rect 12964 3895 12969 3915
rect 12911 3892 12969 3895
rect 12882 3885 12969 3892
rect 12994 3912 13031 4054
rect 13297 4053 13334 4054
rect 13146 3922 13182 3923
rect 12994 3892 13003 3912
rect 13023 3892 13031 3912
rect 12882 3883 12938 3885
rect 12882 3882 12919 3883
rect 12994 3882 13031 3892
rect 13090 3912 13238 3922
rect 13338 3919 13434 3921
rect 13090 3892 13099 3912
rect 13119 3892 13209 3912
rect 13229 3892 13238 3912
rect 13090 3886 13238 3892
rect 13090 3883 13154 3886
rect 13090 3882 13127 3883
rect 13146 3856 13154 3883
rect 13175 3883 13238 3886
rect 13296 3912 13434 3919
rect 13296 3892 13305 3912
rect 13325 3892 13434 3912
rect 13296 3883 13434 3892
rect 13175 3856 13182 3883
rect 13201 3882 13238 3883
rect 13297 3882 13334 3883
rect 13146 3831 13182 3856
rect 12444 3829 12527 3830
rect 12617 3829 12658 3830
rect 12444 3822 12658 3829
rect 12444 3805 12627 3822
rect 12444 3772 12457 3805
rect 12510 3802 12627 3805
rect 12647 3802 12658 3822
rect 12510 3794 12658 3802
rect 12725 3826 13084 3830
rect 12725 3821 13047 3826
rect 12725 3797 12838 3821
rect 12862 3802 13047 3821
rect 13071 3802 13084 3826
rect 12862 3797 13084 3802
rect 12725 3794 13084 3797
rect 13146 3794 13181 3831
rect 13249 3828 13349 3831
rect 13249 3824 13316 3828
rect 13249 3798 13261 3824
rect 13287 3802 13316 3824
rect 13342 3802 13349 3828
rect 13287 3798 13349 3802
rect 13249 3794 13349 3798
rect 12510 3772 12527 3794
rect 12725 3773 12756 3794
rect 13146 3773 13182 3794
rect 12568 3772 12605 3773
rect 12444 3758 12527 3772
rect 12217 3515 12385 3517
rect 11941 3514 12385 3515
rect 11185 3484 12385 3514
rect 12455 3548 12527 3758
rect 12567 3763 12605 3772
rect 12567 3743 12576 3763
rect 12596 3743 12605 3763
rect 12567 3735 12605 3743
rect 12671 3767 12756 3773
rect 12781 3772 12818 3773
rect 12671 3747 12679 3767
rect 12699 3747 12756 3767
rect 12671 3739 12756 3747
rect 12780 3763 12818 3772
rect 12780 3743 12789 3763
rect 12809 3743 12818 3763
rect 12671 3738 12707 3739
rect 12780 3735 12818 3743
rect 12884 3767 12969 3773
rect 12989 3772 13026 3773
rect 12884 3747 12892 3767
rect 12912 3766 12969 3767
rect 12912 3747 12941 3766
rect 12884 3746 12941 3747
rect 12962 3746 12969 3766
rect 12884 3739 12969 3746
rect 12988 3763 13026 3772
rect 12988 3743 12997 3763
rect 13017 3743 13026 3763
rect 12884 3738 12920 3739
rect 12988 3735 13026 3743
rect 13092 3767 13236 3773
rect 13092 3747 13100 3767
rect 13120 3747 13208 3767
rect 13228 3747 13236 3767
rect 13092 3739 13236 3747
rect 13092 3738 13128 3739
rect 13200 3738 13236 3739
rect 13302 3772 13339 3773
rect 13302 3771 13340 3772
rect 13302 3763 13366 3771
rect 13302 3743 13311 3763
rect 13331 3749 13366 3763
rect 13386 3749 13389 3769
rect 13331 3744 13389 3749
rect 13331 3743 13366 3744
rect 12568 3706 12605 3735
rect 12569 3704 12605 3706
rect 12781 3704 12818 3735
rect 12569 3682 12818 3704
rect 12650 3676 12761 3682
rect 12650 3668 12691 3676
rect 12650 3648 12658 3668
rect 12677 3648 12691 3668
rect 12650 3646 12691 3648
rect 12719 3668 12761 3676
rect 12719 3648 12735 3668
rect 12754 3648 12761 3668
rect 12719 3646 12761 3648
rect 12650 3631 12761 3646
rect 12455 3509 12474 3548
rect 12519 3509 12527 3548
rect 12455 3492 12527 3509
rect 12989 3536 13026 3735
rect 13302 3731 13366 3743
rect 12989 3530 13030 3536
rect 13406 3532 13433 3883
rect 13562 3835 13633 4314
rect 13562 3751 13631 3835
rect 13265 3530 13433 3532
rect 12989 3504 13433 3530
rect 11185 3437 11250 3484
rect 11185 3419 11208 3437
rect 11226 3419 11250 3437
rect 12098 3464 12133 3466
rect 12098 3462 12202 3464
rect 12991 3462 13030 3504
rect 13265 3503 13433 3504
rect 12098 3455 13032 3462
rect 12098 3454 12149 3455
rect 12098 3434 12101 3454
rect 12126 3435 12149 3454
rect 12181 3435 13032 3455
rect 12126 3434 13032 3435
rect 12098 3427 13032 3434
rect 12371 3426 13032 3427
rect 11185 3398 11250 3419
rect 11462 3409 11502 3412
rect 11462 3405 12365 3409
rect 11462 3385 12339 3405
rect 12359 3385 12365 3405
rect 11462 3382 12365 3385
rect 11186 3338 11251 3358
rect 11186 3320 11210 3338
rect 11228 3320 11251 3338
rect 11186 3293 11251 3320
rect 11462 3293 11502 3382
rect 11946 3380 12362 3382
rect 11946 3379 12287 3380
rect 11603 3348 11713 3362
rect 11603 3345 11646 3348
rect 11603 3340 11607 3345
rect 11185 3258 11502 3293
rect 11525 3318 11607 3340
rect 11636 3318 11646 3345
rect 11674 3321 11681 3348
rect 11710 3340 11713 3348
rect 11710 3321 11775 3340
rect 11674 3318 11775 3321
rect 11525 3316 11775 3318
rect 10143 3235 10165 3253
rect 10183 3235 10208 3253
rect 10143 3216 10208 3235
rect 9836 3191 9873 3192
rect 9259 3170 9295 3191
rect 9685 3170 9716 3191
rect 9923 3186 9931 3195
rect 9920 3170 9931 3186
rect 9092 3166 9192 3170
rect 9092 3162 9154 3166
rect 9092 3136 9099 3162
rect 9125 3140 9154 3162
rect 9180 3140 9192 3166
rect 9125 3136 9192 3140
rect 9092 3133 9192 3136
rect 9260 3133 9295 3170
rect 9357 3167 9716 3170
rect 9357 3162 9579 3167
rect 9357 3138 9370 3162
rect 9394 3143 9579 3162
rect 9603 3143 9716 3167
rect 9394 3138 9716 3143
rect 9357 3134 9716 3138
rect 9783 3162 9931 3170
rect 9783 3142 9794 3162
rect 9814 3153 9931 3162
rect 9980 3186 9987 3195
rect 9980 3153 9988 3186
rect 11186 3182 11251 3258
rect 11525 3237 11562 3316
rect 11603 3303 11713 3316
rect 11677 3247 11708 3248
rect 11525 3217 11534 3237
rect 11554 3217 11562 3237
rect 11525 3207 11562 3217
rect 11621 3237 11708 3247
rect 11621 3217 11630 3237
rect 11650 3217 11708 3237
rect 11621 3208 11708 3217
rect 11621 3207 11658 3208
rect 9814 3142 9988 3153
rect 9783 3135 9988 3142
rect 9783 3134 9824 3135
rect 9259 3108 9295 3133
rect 9107 3081 9144 3082
rect 9203 3081 9240 3082
rect 9259 3081 9266 3108
rect 8783 3056 8791 3076
rect 8811 3056 8820 3076
rect 8637 3045 8668 3046
rect 8632 2977 8742 2990
rect 8783 2977 8820 3056
rect 9007 3072 9145 3081
rect 9007 3052 9116 3072
rect 9136 3052 9145 3072
rect 9007 3045 9145 3052
rect 9203 3078 9266 3081
rect 9287 3081 9295 3108
rect 9314 3081 9351 3082
rect 9287 3078 9351 3081
rect 9203 3072 9351 3078
rect 9203 3052 9212 3072
rect 9232 3052 9322 3072
rect 9342 3052 9351 3072
rect 9007 3043 9103 3045
rect 9203 3042 9351 3052
rect 9410 3072 9447 3082
rect 9522 3081 9559 3082
rect 9503 3079 9559 3081
rect 9410 3052 9418 3072
rect 9438 3052 9447 3072
rect 9259 3041 9295 3042
rect 8570 2975 8820 2977
rect 8570 2972 8671 2975
rect 8570 2953 8635 2972
rect 8632 2945 8635 2953
rect 8664 2945 8671 2972
rect 8699 2948 8709 2975
rect 8738 2953 8820 2975
rect 8738 2948 8742 2953
rect 8699 2945 8742 2948
rect 8632 2931 8742 2945
rect 8058 2913 8399 2914
rect 7983 2908 8399 2913
rect 9107 2910 9144 2911
rect 9410 2910 9447 3052
rect 9472 3072 9559 3079
rect 9472 3069 9530 3072
rect 9472 3049 9477 3069
rect 9498 3052 9530 3069
rect 9550 3052 9559 3072
rect 9498 3049 9559 3052
rect 9472 3042 9559 3049
rect 9618 3072 9655 3082
rect 9618 3052 9626 3072
rect 9646 3052 9655 3072
rect 9472 3041 9503 3042
rect 9618 2973 9655 3052
rect 9685 3081 9716 3134
rect 9920 3132 9988 3135
rect 9920 3090 9932 3132
rect 9981 3090 9988 3132
rect 9735 3081 9772 3082
rect 9685 3072 9772 3081
rect 9685 3052 9743 3072
rect 9763 3052 9772 3072
rect 9685 3042 9772 3052
rect 9831 3072 9868 3082
rect 9920 3077 9988 3090
rect 10143 3154 10208 3171
rect 10143 3136 10167 3154
rect 10185 3136 10208 3154
rect 11186 3164 11208 3182
rect 11226 3164 11251 3182
rect 11186 3143 11251 3164
rect 11399 3162 11464 3171
rect 9831 3052 9839 3072
rect 9859 3052 9868 3072
rect 9685 3041 9716 3042
rect 9680 2973 9790 2986
rect 9831 2973 9868 3052
rect 10143 2997 10208 3136
rect 11399 3125 11409 3162
rect 11449 3154 11464 3162
rect 11677 3155 11708 3208
rect 11738 3237 11775 3316
rect 11890 3247 11921 3248
rect 11738 3217 11747 3237
rect 11767 3217 11775 3237
rect 11738 3207 11775 3217
rect 11834 3240 11921 3247
rect 11834 3237 11895 3240
rect 11834 3217 11843 3237
rect 11863 3220 11895 3237
rect 11916 3220 11921 3240
rect 11863 3217 11921 3220
rect 11834 3210 11921 3217
rect 11946 3237 11983 3379
rect 12249 3378 12286 3379
rect 12098 3247 12134 3248
rect 11946 3217 11955 3237
rect 11975 3217 11983 3237
rect 11834 3208 11890 3210
rect 11834 3207 11871 3208
rect 11946 3207 11983 3217
rect 12042 3237 12190 3247
rect 12290 3244 12386 3246
rect 12042 3217 12051 3237
rect 12071 3217 12161 3237
rect 12181 3217 12190 3237
rect 12042 3211 12190 3217
rect 12042 3208 12106 3211
rect 12042 3207 12079 3208
rect 12098 3181 12106 3208
rect 12127 3208 12190 3211
rect 12248 3237 12386 3244
rect 13566 3239 13628 3751
rect 12248 3217 12257 3237
rect 12277 3217 12386 3237
rect 12248 3208 12386 3217
rect 12127 3181 12134 3208
rect 12153 3207 12190 3208
rect 12249 3207 12286 3208
rect 12098 3156 12134 3181
rect 11569 3154 11610 3155
rect 11449 3147 11610 3154
rect 11449 3127 11579 3147
rect 11599 3127 11610 3147
rect 11449 3125 11610 3127
rect 11399 3119 11610 3125
rect 11677 3151 12036 3155
rect 11677 3146 11999 3151
rect 11677 3122 11790 3146
rect 11814 3127 11999 3146
rect 12023 3127 12036 3151
rect 11814 3122 12036 3127
rect 11677 3119 12036 3122
rect 12098 3119 12133 3156
rect 12201 3153 12301 3156
rect 12201 3149 12268 3153
rect 12201 3123 12213 3149
rect 12239 3127 12268 3149
rect 12294 3127 12301 3153
rect 12239 3123 12301 3127
rect 12201 3119 12301 3123
rect 11399 3106 11466 3119
rect 10143 2991 10165 2997
rect 9618 2971 9868 2973
rect 9618 2968 9719 2971
rect 9618 2949 9683 2968
rect 9680 2941 9683 2949
rect 9712 2941 9719 2968
rect 9747 2944 9757 2971
rect 9786 2949 9868 2971
rect 9897 2979 10165 2991
rect 10183 2979 10208 2997
rect 9897 2956 10208 2979
rect 11191 3083 11247 3103
rect 11191 3065 11210 3083
rect 11228 3065 11247 3083
rect 9897 2955 9952 2956
rect 9786 2944 9790 2949
rect 9747 2941 9790 2944
rect 9680 2927 9790 2941
rect 9106 2909 9447 2910
rect 7983 2888 7986 2908
rect 8006 2888 8399 2908
rect 9031 2908 9447 2909
rect 9897 2908 9940 2955
rect 11191 2952 11247 3065
rect 11399 3085 11413 3106
rect 11449 3085 11466 3106
rect 11677 3098 11708 3119
rect 12098 3098 12134 3119
rect 11520 3097 11557 3098
rect 11399 3078 11466 3085
rect 11519 3088 11557 3097
rect 9031 2904 9940 2908
rect 8350 2855 8395 2888
rect 9031 2884 9034 2904
rect 9054 2884 9940 2904
rect 9408 2879 9940 2884
rect 10148 2898 10207 2920
rect 10148 2880 10167 2898
rect 10185 2880 10207 2898
rect 9196 2855 9295 2857
rect 8350 2845 9295 2855
rect 8350 2819 9218 2845
rect 8351 2818 9218 2819
rect 9196 2807 9218 2818
rect 9243 2810 9262 2845
rect 9287 2810 9295 2845
rect 9243 2807 9295 2810
rect 10148 2809 10207 2880
rect 11191 2814 11246 2952
rect 11399 2926 11464 3078
rect 11519 3068 11528 3088
rect 11548 3068 11557 3088
rect 11519 3060 11557 3068
rect 11623 3092 11708 3098
rect 11733 3097 11770 3098
rect 11623 3072 11631 3092
rect 11651 3072 11708 3092
rect 11623 3064 11708 3072
rect 11732 3088 11770 3097
rect 11732 3068 11741 3088
rect 11761 3068 11770 3088
rect 11623 3063 11659 3064
rect 11732 3060 11770 3068
rect 11836 3092 11921 3098
rect 11941 3097 11978 3098
rect 11836 3072 11844 3092
rect 11864 3091 11921 3092
rect 11864 3072 11893 3091
rect 11836 3071 11893 3072
rect 11914 3071 11921 3091
rect 11836 3064 11921 3071
rect 11940 3088 11978 3097
rect 11940 3068 11949 3088
rect 11969 3068 11978 3088
rect 11836 3063 11872 3064
rect 11940 3060 11978 3068
rect 12044 3092 12188 3098
rect 12044 3072 12052 3092
rect 12072 3072 12160 3092
rect 12180 3072 12188 3092
rect 12044 3064 12188 3072
rect 12044 3063 12080 3064
rect 12152 3063 12188 3064
rect 12254 3097 12291 3098
rect 12254 3096 12292 3097
rect 12254 3088 12318 3096
rect 12254 3068 12263 3088
rect 12283 3074 12318 3088
rect 12338 3074 12341 3094
rect 12283 3069 12341 3074
rect 12283 3068 12318 3069
rect 11520 3031 11557 3060
rect 11521 3029 11557 3031
rect 11733 3029 11770 3060
rect 11521 3007 11770 3029
rect 11602 3001 11713 3007
rect 11602 2993 11643 3001
rect 11602 2973 11610 2993
rect 11629 2973 11643 2993
rect 11602 2971 11643 2973
rect 11671 2993 11713 3001
rect 11671 2973 11687 2993
rect 11706 2973 11713 2993
rect 11671 2971 11713 2973
rect 11602 2958 11713 2971
rect 11941 2961 11978 3060
rect 12254 3056 12318 3068
rect 11392 2916 11513 2926
rect 11392 2914 11461 2916
rect 11392 2873 11405 2914
rect 11442 2875 11461 2914
rect 11498 2875 11513 2916
rect 11442 2873 11513 2875
rect 11392 2855 11513 2873
rect 11184 2811 11248 2814
rect 11604 2811 11708 2817
rect 11939 2811 11980 2961
rect 12358 2953 12385 3208
rect 12447 3198 12527 3209
rect 12447 3172 12464 3198
rect 12504 3172 12527 3198
rect 12447 3145 12527 3172
rect 13570 3200 13628 3239
rect 13570 3165 13632 3200
rect 12447 3119 12468 3145
rect 12508 3119 12527 3145
rect 12447 3100 12527 3119
rect 12447 3074 12471 3100
rect 12511 3074 12527 3100
rect 12447 3023 12527 3074
rect 13519 3138 13632 3165
rect 13519 3136 13578 3138
rect 13519 3105 13533 3136
rect 13558 3115 13578 3136
rect 13604 3115 13632 3138
rect 13558 3105 13632 3115
rect 13519 3095 13632 3105
rect 9196 2799 9295 2807
rect 9222 2798 9294 2799
rect 8876 2772 8943 2791
rect 8876 2751 8893 2772
rect 7757 2573 7837 2615
rect 8874 2706 8893 2751
rect 8923 2751 8943 2772
rect 8923 2706 8944 2751
rect 9413 2748 9454 2750
rect 9685 2748 9789 2750
rect 10145 2748 10209 2809
rect 6818 2462 6854 2463
rect 6710 2454 6854 2462
rect 6710 2434 6718 2454
rect 6738 2434 6826 2454
rect 6846 2434 6854 2454
rect 6710 2428 6854 2434
rect 6920 2458 6958 2466
rect 7026 2462 7062 2463
rect 6920 2438 6929 2458
rect 6949 2438 6958 2458
rect 6920 2429 6958 2438
rect 6977 2455 7062 2462
rect 6977 2435 6984 2455
rect 7005 2454 7062 2455
rect 7005 2435 7034 2454
rect 6977 2434 7034 2435
rect 7054 2434 7062 2454
rect 6920 2428 6957 2429
rect 6977 2428 7062 2434
rect 7128 2458 7166 2466
rect 7239 2462 7275 2463
rect 7128 2438 7137 2458
rect 7157 2438 7166 2458
rect 7128 2429 7166 2438
rect 7190 2454 7275 2462
rect 7190 2434 7247 2454
rect 7267 2434 7275 2454
rect 7128 2428 7165 2429
rect 7190 2428 7275 2434
rect 7341 2458 7379 2466
rect 7341 2438 7350 2458
rect 7370 2438 7379 2458
rect 7341 2429 7379 2438
rect 7579 2446 7665 2482
rect 7341 2428 7378 2429
rect 6764 2407 6800 2428
rect 7190 2407 7221 2428
rect 7417 2407 7463 2411
rect 6597 2403 6697 2407
rect 6597 2399 6659 2403
rect 6597 2373 6604 2399
rect 6630 2377 6659 2399
rect 6685 2377 6697 2403
rect 6630 2373 6697 2377
rect 6597 2370 6697 2373
rect 6765 2370 6800 2407
rect 6862 2404 7221 2407
rect 6862 2399 7084 2404
rect 6862 2375 6875 2399
rect 6899 2380 7084 2399
rect 7108 2380 7221 2404
rect 6899 2375 7221 2380
rect 6862 2371 7221 2375
rect 7288 2399 7463 2407
rect 7288 2379 7299 2399
rect 7319 2379 7463 2399
rect 7579 2405 7596 2446
rect 7650 2405 7665 2446
rect 7579 2386 7665 2405
rect 7288 2372 7463 2379
rect 7288 2371 7329 2372
rect 6764 2345 6800 2370
rect 6612 2318 6649 2319
rect 6708 2318 6745 2319
rect 6764 2318 6771 2345
rect 6512 2309 6650 2318
rect 6512 2289 6621 2309
rect 6641 2289 6650 2309
rect 6512 2282 6650 2289
rect 6708 2315 6771 2318
rect 6792 2318 6800 2345
rect 6819 2318 6856 2319
rect 6792 2315 6856 2318
rect 6708 2309 6856 2315
rect 6708 2289 6717 2309
rect 6737 2289 6827 2309
rect 6847 2289 6856 2309
rect 6512 2280 6608 2282
rect 6708 2279 6856 2289
rect 6915 2309 6952 2319
rect 7027 2318 7064 2319
rect 7008 2316 7064 2318
rect 6915 2289 6923 2309
rect 6943 2289 6952 2309
rect 6764 2278 6800 2279
rect 6612 2147 6649 2148
rect 6915 2147 6952 2289
rect 6977 2309 7064 2316
rect 6977 2306 7035 2309
rect 6977 2286 6982 2306
rect 7003 2289 7035 2306
rect 7055 2289 7064 2309
rect 7003 2286 7064 2289
rect 6977 2279 7064 2286
rect 7123 2309 7160 2319
rect 7123 2289 7131 2309
rect 7151 2289 7160 2309
rect 6977 2278 7008 2279
rect 7123 2210 7160 2289
rect 7190 2318 7221 2371
rect 7240 2318 7277 2319
rect 7190 2309 7277 2318
rect 7190 2289 7248 2309
rect 7268 2289 7277 2309
rect 7190 2279 7277 2289
rect 7336 2309 7373 2319
rect 7336 2289 7344 2309
rect 7364 2289 7373 2309
rect 7190 2278 7221 2279
rect 7185 2210 7295 2223
rect 7336 2210 7373 2289
rect 7417 2289 7463 2372
rect 7757 2289 7832 2573
rect 8874 2498 8944 2706
rect 9006 2713 10209 2748
rect 9006 2699 9034 2713
rect 9008 2568 9034 2699
rect 9413 2710 10209 2713
rect 11184 2808 11980 2811
rect 12359 2822 12385 2953
rect 12359 2808 12387 2822
rect 11184 2773 12387 2808
rect 12449 2815 12519 3023
rect 11184 2712 11248 2773
rect 11604 2771 11708 2773
rect 11939 2771 11980 2773
rect 12449 2770 12470 2815
rect 12450 2749 12470 2770
rect 12500 2770 12519 2815
rect 12500 2749 12517 2770
rect 12450 2730 12517 2749
rect 12099 2722 12171 2723
rect 12098 2714 12197 2722
rect 8866 2447 8946 2498
rect 8866 2421 8882 2447
rect 8922 2421 8946 2447
rect 8866 2402 8946 2421
rect 8866 2376 8885 2402
rect 8925 2376 8946 2402
rect 8866 2349 8946 2376
rect 8866 2323 8889 2349
rect 8929 2323 8946 2349
rect 8866 2312 8946 2323
rect 9008 2313 9035 2568
rect 9413 2560 9454 2710
rect 9685 2704 9789 2710
rect 10145 2707 10209 2710
rect 9880 2648 10001 2666
rect 9880 2646 9951 2648
rect 9880 2605 9895 2646
rect 9932 2607 9951 2646
rect 9988 2607 10001 2648
rect 9932 2605 10001 2607
rect 9880 2595 10001 2605
rect 9075 2453 9139 2465
rect 9415 2461 9452 2560
rect 9680 2550 9791 2563
rect 9680 2548 9722 2550
rect 9680 2528 9687 2548
rect 9706 2528 9722 2548
rect 9680 2520 9722 2528
rect 9750 2548 9791 2550
rect 9750 2528 9764 2548
rect 9783 2528 9791 2548
rect 9750 2520 9791 2528
rect 9680 2514 9791 2520
rect 9623 2492 9872 2514
rect 9623 2461 9660 2492
rect 9836 2490 9872 2492
rect 9836 2461 9873 2490
rect 9075 2452 9110 2453
rect 9052 2447 9110 2452
rect 9052 2427 9055 2447
rect 9075 2433 9110 2447
rect 9130 2433 9139 2453
rect 9075 2425 9139 2433
rect 9101 2424 9139 2425
rect 9102 2423 9139 2424
rect 9205 2457 9241 2458
rect 9313 2457 9349 2458
rect 9205 2449 9349 2457
rect 9205 2429 9213 2449
rect 9233 2429 9321 2449
rect 9341 2429 9349 2449
rect 9205 2423 9349 2429
rect 9415 2453 9453 2461
rect 9521 2457 9557 2458
rect 9415 2433 9424 2453
rect 9444 2433 9453 2453
rect 9415 2424 9453 2433
rect 9472 2450 9557 2457
rect 9472 2430 9479 2450
rect 9500 2449 9557 2450
rect 9500 2430 9529 2449
rect 9472 2429 9529 2430
rect 9549 2429 9557 2449
rect 9415 2423 9452 2424
rect 9472 2423 9557 2429
rect 9623 2453 9661 2461
rect 9734 2457 9770 2458
rect 9623 2433 9632 2453
rect 9652 2433 9661 2453
rect 9623 2424 9661 2433
rect 9685 2449 9770 2457
rect 9685 2429 9742 2449
rect 9762 2429 9770 2449
rect 9623 2423 9660 2424
rect 9685 2423 9770 2429
rect 9836 2453 9874 2461
rect 9836 2433 9845 2453
rect 9865 2433 9874 2453
rect 9929 2443 9994 2595
rect 10147 2569 10202 2707
rect 11186 2641 11245 2712
rect 12098 2711 12150 2714
rect 12098 2676 12106 2711
rect 12131 2676 12150 2711
rect 12175 2703 12197 2714
rect 12175 2702 13042 2703
rect 12175 2676 13043 2702
rect 12098 2666 13043 2676
rect 12098 2664 12197 2666
rect 11186 2623 11208 2641
rect 11226 2623 11245 2641
rect 11186 2601 11245 2623
rect 11453 2637 11985 2642
rect 11453 2617 12339 2637
rect 12359 2617 12362 2637
rect 12998 2633 13043 2666
rect 11453 2613 12362 2617
rect 9836 2424 9874 2433
rect 9927 2436 9994 2443
rect 9836 2423 9873 2424
rect 9259 2402 9295 2423
rect 9685 2402 9716 2423
rect 9927 2415 9944 2436
rect 9980 2415 9994 2436
rect 10146 2456 10202 2569
rect 11453 2566 11496 2613
rect 11946 2612 12362 2613
rect 12994 2613 13387 2633
rect 13407 2613 13410 2633
rect 11946 2611 12287 2612
rect 11603 2580 11713 2594
rect 11603 2577 11646 2580
rect 11603 2572 11607 2577
rect 11441 2565 11496 2566
rect 10146 2438 10165 2456
rect 10183 2438 10202 2456
rect 10146 2418 10202 2438
rect 11185 2542 11496 2565
rect 11185 2524 11210 2542
rect 11228 2530 11496 2542
rect 11525 2550 11607 2572
rect 11636 2550 11646 2577
rect 11674 2553 11681 2580
rect 11710 2572 11713 2580
rect 11710 2553 11775 2572
rect 11674 2550 11775 2553
rect 11525 2548 11775 2550
rect 11228 2524 11250 2530
rect 9927 2402 9994 2415
rect 9092 2398 9192 2402
rect 9092 2394 9154 2398
rect 9092 2368 9099 2394
rect 9125 2372 9154 2394
rect 9180 2372 9192 2398
rect 9125 2368 9192 2372
rect 9092 2365 9192 2368
rect 9260 2365 9295 2402
rect 9357 2399 9716 2402
rect 9357 2394 9579 2399
rect 9357 2370 9370 2394
rect 9394 2375 9579 2394
rect 9603 2375 9716 2399
rect 9394 2370 9716 2375
rect 9357 2366 9716 2370
rect 9783 2396 9994 2402
rect 9783 2394 9944 2396
rect 9783 2374 9794 2394
rect 9814 2374 9944 2394
rect 9783 2367 9944 2374
rect 9783 2366 9824 2367
rect 9259 2340 9295 2365
rect 9107 2313 9144 2314
rect 9203 2313 9240 2314
rect 9259 2313 9266 2340
rect 7417 2254 7832 2289
rect 9007 2304 9145 2313
rect 9007 2284 9116 2304
rect 9136 2284 9145 2304
rect 9007 2277 9145 2284
rect 9203 2310 9266 2313
rect 9287 2313 9295 2340
rect 9314 2313 9351 2314
rect 9287 2310 9351 2313
rect 9203 2304 9351 2310
rect 9203 2284 9212 2304
rect 9232 2284 9322 2304
rect 9342 2284 9351 2304
rect 9007 2275 9103 2277
rect 9203 2274 9351 2284
rect 9410 2304 9447 2314
rect 9522 2313 9559 2314
rect 9503 2311 9559 2313
rect 9410 2284 9418 2304
rect 9438 2284 9447 2304
rect 9259 2273 9295 2274
rect 7417 2253 7463 2254
rect 7123 2208 7373 2210
rect 7123 2205 7224 2208
rect 7123 2186 7188 2205
rect 7185 2178 7188 2186
rect 7217 2178 7224 2205
rect 7252 2181 7262 2208
rect 7291 2186 7373 2208
rect 7757 2202 7832 2254
rect 7291 2181 7295 2186
rect 7252 2178 7295 2181
rect 7185 2164 7295 2178
rect 6611 2146 6952 2147
rect 6536 2141 6952 2146
rect 6536 2121 6539 2141
rect 6559 2121 6953 2141
rect 3016 1712 6084 1737
rect 3016 1647 5879 1712
rect 6010 1647 6084 1712
rect 3016 1630 6084 1647
rect 6910 1617 6953 2121
rect 7570 2032 7665 2052
rect 7570 1988 7590 2032
rect 7650 1988 7665 2032
rect 7570 1692 7665 1988
rect 7570 1651 7603 1692
rect 7639 1651 7665 1692
rect 7765 1731 7827 2202
rect 9107 2142 9144 2143
rect 9410 2142 9447 2284
rect 9472 2304 9559 2311
rect 9472 2301 9530 2304
rect 9472 2281 9477 2301
rect 9498 2284 9530 2301
rect 9550 2284 9559 2304
rect 9498 2281 9559 2284
rect 9472 2274 9559 2281
rect 9618 2304 9655 2314
rect 9618 2284 9626 2304
rect 9646 2284 9655 2304
rect 9472 2273 9503 2274
rect 9618 2205 9655 2284
rect 9685 2313 9716 2366
rect 9929 2359 9944 2367
rect 9984 2359 9994 2396
rect 11185 2385 11250 2524
rect 11525 2469 11562 2548
rect 11603 2535 11713 2548
rect 11677 2479 11708 2480
rect 11525 2449 11534 2469
rect 11554 2449 11562 2469
rect 9929 2350 9994 2359
rect 10142 2357 10207 2378
rect 10142 2339 10167 2357
rect 10185 2339 10207 2357
rect 11185 2367 11208 2385
rect 11226 2367 11250 2385
rect 11185 2350 11250 2367
rect 11405 2431 11473 2444
rect 11525 2439 11562 2449
rect 11621 2469 11708 2479
rect 11621 2449 11630 2469
rect 11650 2449 11708 2469
rect 11621 2440 11708 2449
rect 11621 2439 11658 2440
rect 11405 2389 11412 2431
rect 11461 2389 11473 2431
rect 11405 2386 11473 2389
rect 11677 2387 11708 2440
rect 11738 2469 11775 2548
rect 11890 2479 11921 2480
rect 11738 2449 11747 2469
rect 11767 2449 11775 2469
rect 11738 2439 11775 2449
rect 11834 2472 11921 2479
rect 11834 2469 11895 2472
rect 11834 2449 11843 2469
rect 11863 2452 11895 2469
rect 11916 2452 11921 2472
rect 11863 2449 11921 2452
rect 11834 2442 11921 2449
rect 11946 2469 11983 2611
rect 12249 2610 12286 2611
rect 12994 2608 13410 2613
rect 12994 2607 13335 2608
rect 12651 2576 12761 2590
rect 12651 2573 12694 2576
rect 12651 2568 12655 2573
rect 12573 2546 12655 2568
rect 12684 2546 12694 2573
rect 12722 2549 12729 2576
rect 12758 2568 12761 2576
rect 12758 2549 12823 2568
rect 12722 2546 12823 2549
rect 12573 2544 12823 2546
rect 12098 2479 12134 2480
rect 11946 2449 11955 2469
rect 11975 2449 11983 2469
rect 11834 2440 11890 2442
rect 11834 2439 11871 2440
rect 11946 2439 11983 2449
rect 12042 2469 12190 2479
rect 12290 2476 12386 2478
rect 12042 2449 12051 2469
rect 12071 2449 12161 2469
rect 12181 2449 12190 2469
rect 12042 2443 12190 2449
rect 12042 2440 12106 2443
rect 12042 2439 12079 2440
rect 12098 2413 12106 2440
rect 12127 2440 12190 2443
rect 12248 2469 12386 2476
rect 12248 2449 12257 2469
rect 12277 2449 12386 2469
rect 12248 2440 12386 2449
rect 12573 2465 12610 2544
rect 12651 2531 12761 2544
rect 12725 2475 12756 2476
rect 12573 2445 12582 2465
rect 12602 2445 12610 2465
rect 12127 2413 12134 2440
rect 12153 2439 12190 2440
rect 12249 2439 12286 2440
rect 12098 2388 12134 2413
rect 11569 2386 11610 2387
rect 11405 2379 11610 2386
rect 11405 2368 11579 2379
rect 9735 2313 9772 2314
rect 9685 2304 9772 2313
rect 9685 2284 9743 2304
rect 9763 2284 9772 2304
rect 9685 2274 9772 2284
rect 9831 2304 9868 2314
rect 9831 2284 9839 2304
rect 9859 2284 9868 2304
rect 9685 2273 9716 2274
rect 9680 2205 9790 2218
rect 9831 2205 9868 2284
rect 10142 2263 10207 2339
rect 11405 2335 11413 2368
rect 11406 2326 11413 2335
rect 11462 2359 11579 2368
rect 11599 2359 11610 2379
rect 11462 2351 11610 2359
rect 11677 2383 12036 2387
rect 11677 2378 11999 2383
rect 11677 2354 11790 2378
rect 11814 2359 11999 2378
rect 12023 2359 12036 2383
rect 11814 2354 12036 2359
rect 11677 2351 12036 2354
rect 12098 2351 12133 2388
rect 12201 2385 12301 2388
rect 12201 2381 12268 2385
rect 12201 2355 12213 2381
rect 12239 2359 12268 2381
rect 12294 2359 12301 2385
rect 12239 2355 12301 2359
rect 12201 2351 12301 2355
rect 11462 2335 11473 2351
rect 11462 2326 11470 2335
rect 11677 2330 11708 2351
rect 12098 2330 12134 2351
rect 11520 2329 11557 2330
rect 11185 2286 11250 2305
rect 11185 2268 11210 2286
rect 11228 2268 11250 2286
rect 9618 2203 9868 2205
rect 9618 2200 9719 2203
rect 9618 2181 9683 2200
rect 9680 2173 9683 2181
rect 9712 2173 9719 2200
rect 9747 2176 9757 2203
rect 9786 2181 9868 2203
rect 9891 2228 10208 2263
rect 9786 2176 9790 2181
rect 9747 2173 9790 2176
rect 9680 2159 9790 2173
rect 9106 2141 9447 2142
rect 9031 2139 9447 2141
rect 9891 2139 9931 2228
rect 10142 2201 10207 2228
rect 10142 2183 10165 2201
rect 10183 2183 10207 2201
rect 10142 2163 10207 2183
rect 9028 2136 9931 2139
rect 9028 2116 9034 2136
rect 9054 2116 9931 2136
rect 9028 2112 9931 2116
rect 9891 2109 9931 2112
rect 10143 2102 10208 2123
rect 8361 2094 9022 2095
rect 8361 2087 9295 2094
rect 8361 2086 9267 2087
rect 8361 2066 9212 2086
rect 9244 2067 9267 2086
rect 9292 2067 9295 2087
rect 9244 2066 9295 2067
rect 8361 2059 9295 2066
rect 7960 2017 8128 2018
rect 8363 2017 8402 2059
rect 9191 2057 9295 2059
rect 9260 2055 9295 2057
rect 10143 2084 10167 2102
rect 10185 2084 10208 2102
rect 10143 2037 10208 2084
rect 7960 1991 8404 2017
rect 7960 1989 8128 1991
rect 7765 1712 7829 1731
rect 7765 1673 7782 1712
rect 7816 1673 7829 1712
rect 7765 1654 7829 1673
rect 7570 1625 7665 1651
rect 7960 1638 7987 1989
rect 8363 1985 8404 1991
rect 8027 1778 8091 1790
rect 8367 1786 8404 1985
rect 8866 2012 8938 2029
rect 8866 1973 8874 2012
rect 8919 1973 8938 2012
rect 8632 1875 8743 1890
rect 8632 1873 8674 1875
rect 8632 1853 8639 1873
rect 8658 1853 8674 1873
rect 8632 1845 8674 1853
rect 8702 1873 8743 1875
rect 8702 1853 8716 1873
rect 8735 1853 8743 1873
rect 8702 1845 8743 1853
rect 8632 1839 8743 1845
rect 8575 1817 8824 1839
rect 8575 1786 8612 1817
rect 8788 1815 8824 1817
rect 8788 1786 8825 1815
rect 8027 1777 8062 1778
rect 8004 1772 8062 1777
rect 8004 1752 8007 1772
rect 8027 1758 8062 1772
rect 8082 1758 8091 1778
rect 8027 1750 8091 1758
rect 8053 1749 8091 1750
rect 8054 1748 8091 1749
rect 8157 1782 8193 1783
rect 8265 1782 8301 1783
rect 8157 1774 8301 1782
rect 8157 1754 8165 1774
rect 8185 1754 8273 1774
rect 8293 1754 8301 1774
rect 8157 1748 8301 1754
rect 8367 1778 8405 1786
rect 8473 1782 8509 1783
rect 8367 1758 8376 1778
rect 8396 1758 8405 1778
rect 8367 1749 8405 1758
rect 8424 1775 8509 1782
rect 8424 1755 8431 1775
rect 8452 1774 8509 1775
rect 8452 1755 8481 1774
rect 8424 1754 8481 1755
rect 8501 1754 8509 1774
rect 8367 1748 8404 1749
rect 8424 1748 8509 1754
rect 8575 1778 8613 1786
rect 8686 1782 8722 1783
rect 8575 1758 8584 1778
rect 8604 1758 8613 1778
rect 8575 1749 8613 1758
rect 8637 1774 8722 1782
rect 8637 1754 8694 1774
rect 8714 1754 8722 1774
rect 8575 1748 8612 1749
rect 8637 1748 8722 1754
rect 8788 1778 8826 1786
rect 8788 1758 8797 1778
rect 8817 1758 8826 1778
rect 8788 1749 8826 1758
rect 8866 1763 8938 1973
rect 9008 2007 10208 2037
rect 9008 2006 9452 2007
rect 9008 2004 9176 2006
rect 8866 1749 8949 1763
rect 8788 1748 8825 1749
rect 8211 1727 8247 1748
rect 8637 1727 8668 1748
rect 8866 1727 8883 1749
rect 8044 1723 8144 1727
rect 8044 1719 8106 1723
rect 8044 1693 8051 1719
rect 8077 1697 8106 1719
rect 8132 1697 8144 1723
rect 8077 1693 8144 1697
rect 8044 1690 8144 1693
rect 8212 1690 8247 1727
rect 8309 1724 8668 1727
rect 8309 1719 8531 1724
rect 8309 1695 8322 1719
rect 8346 1700 8531 1719
rect 8555 1700 8668 1724
rect 8346 1695 8668 1700
rect 8309 1691 8668 1695
rect 8735 1719 8883 1727
rect 8735 1699 8746 1719
rect 8766 1716 8883 1719
rect 8936 1716 8949 1749
rect 8766 1699 8949 1716
rect 8735 1692 8949 1699
rect 8735 1691 8776 1692
rect 8866 1691 8949 1692
rect 8211 1665 8247 1690
rect 8059 1638 8096 1639
rect 8155 1638 8192 1639
rect 8211 1638 8218 1665
rect 7959 1629 8097 1638
rect 2771 1531 2928 1544
rect 2771 1527 2932 1531
rect 1651 1381 1677 1486
rect 2771 1420 2812 1527
rect 2912 1420 2932 1527
rect 2771 1391 2932 1420
rect 6908 1408 6957 1617
rect 7959 1609 8068 1629
rect 8088 1609 8097 1629
rect 7959 1602 8097 1609
rect 8155 1635 8218 1638
rect 8239 1638 8247 1665
rect 8266 1638 8303 1639
rect 8239 1635 8303 1638
rect 8155 1629 8303 1635
rect 8155 1609 8164 1629
rect 8184 1609 8274 1629
rect 8294 1609 8303 1629
rect 7959 1600 8055 1602
rect 8155 1599 8303 1609
rect 8362 1629 8399 1639
rect 8474 1638 8511 1639
rect 8455 1636 8511 1638
rect 8362 1609 8370 1629
rect 8390 1609 8399 1629
rect 8211 1598 8247 1599
rect 8059 1467 8096 1468
rect 8362 1467 8399 1609
rect 8424 1629 8511 1636
rect 8424 1626 8482 1629
rect 8424 1606 8429 1626
rect 8450 1609 8482 1626
rect 8502 1609 8511 1629
rect 8450 1606 8511 1609
rect 8424 1599 8511 1606
rect 8570 1629 8607 1639
rect 8570 1609 8578 1629
rect 8598 1609 8607 1629
rect 8424 1598 8455 1599
rect 8570 1530 8607 1609
rect 8637 1638 8668 1691
rect 8874 1658 8888 1691
rect 8941 1658 8949 1691
rect 8874 1652 8949 1658
rect 8874 1647 8944 1652
rect 8687 1638 8724 1639
rect 8637 1629 8724 1638
rect 8637 1609 8695 1629
rect 8715 1609 8724 1629
rect 8637 1599 8724 1609
rect 8783 1629 8820 1639
rect 9008 1634 9035 2004
rect 9075 1774 9139 1786
rect 9415 1782 9452 2006
rect 9923 1987 9987 1989
rect 9919 1975 9987 1987
rect 9919 1942 9930 1975
rect 9970 1942 9987 1975
rect 9919 1932 9987 1942
rect 9680 1871 9791 1886
rect 9680 1869 9722 1871
rect 9680 1849 9687 1869
rect 9706 1849 9722 1869
rect 9680 1841 9722 1849
rect 9750 1869 9791 1871
rect 9750 1849 9764 1869
rect 9783 1849 9791 1869
rect 9750 1841 9791 1849
rect 9680 1835 9791 1841
rect 9623 1813 9872 1835
rect 9623 1782 9660 1813
rect 9836 1811 9872 1813
rect 9836 1782 9873 1811
rect 9075 1773 9110 1774
rect 9052 1768 9110 1773
rect 9052 1748 9055 1768
rect 9075 1754 9110 1768
rect 9130 1754 9139 1774
rect 9075 1746 9139 1754
rect 9101 1745 9139 1746
rect 9102 1744 9139 1745
rect 9205 1778 9241 1779
rect 9313 1778 9349 1779
rect 9205 1770 9349 1778
rect 9205 1750 9213 1770
rect 9233 1750 9321 1770
rect 9341 1750 9349 1770
rect 9205 1744 9349 1750
rect 9415 1774 9453 1782
rect 9521 1778 9557 1779
rect 9415 1754 9424 1774
rect 9444 1754 9453 1774
rect 9415 1745 9453 1754
rect 9472 1771 9557 1778
rect 9472 1751 9479 1771
rect 9500 1770 9557 1771
rect 9500 1751 9529 1770
rect 9472 1750 9529 1751
rect 9549 1750 9557 1770
rect 9415 1744 9452 1745
rect 9472 1744 9557 1750
rect 9623 1774 9661 1782
rect 9734 1778 9770 1779
rect 9623 1754 9632 1774
rect 9652 1754 9661 1774
rect 9623 1745 9661 1754
rect 9685 1770 9770 1778
rect 9685 1750 9742 1770
rect 9762 1750 9770 1770
rect 9623 1744 9660 1745
rect 9685 1744 9770 1750
rect 9836 1774 9874 1782
rect 9836 1754 9845 1774
rect 9865 1754 9874 1774
rect 9836 1745 9874 1754
rect 9923 1748 9987 1932
rect 10143 1806 10208 2007
rect 11185 2067 11250 2268
rect 11406 2142 11470 2326
rect 11519 2320 11557 2329
rect 11519 2300 11528 2320
rect 11548 2300 11557 2320
rect 11519 2292 11557 2300
rect 11623 2324 11708 2330
rect 11733 2329 11770 2330
rect 11623 2304 11631 2324
rect 11651 2304 11708 2324
rect 11623 2296 11708 2304
rect 11732 2320 11770 2329
rect 11732 2300 11741 2320
rect 11761 2300 11770 2320
rect 11623 2295 11659 2296
rect 11732 2292 11770 2300
rect 11836 2324 11921 2330
rect 11941 2329 11978 2330
rect 11836 2304 11844 2324
rect 11864 2323 11921 2324
rect 11864 2304 11893 2323
rect 11836 2303 11893 2304
rect 11914 2303 11921 2323
rect 11836 2296 11921 2303
rect 11940 2320 11978 2329
rect 11940 2300 11949 2320
rect 11969 2300 11978 2320
rect 11836 2295 11872 2296
rect 11940 2292 11978 2300
rect 12044 2324 12188 2330
rect 12044 2304 12052 2324
rect 12072 2304 12160 2324
rect 12180 2304 12188 2324
rect 12044 2296 12188 2304
rect 12044 2295 12080 2296
rect 12152 2295 12188 2296
rect 12254 2329 12291 2330
rect 12254 2328 12292 2329
rect 12254 2320 12318 2328
rect 12254 2300 12263 2320
rect 12283 2306 12318 2320
rect 12338 2306 12341 2326
rect 12283 2301 12341 2306
rect 12283 2300 12318 2301
rect 11520 2263 11557 2292
rect 11521 2261 11557 2263
rect 11733 2261 11770 2292
rect 11521 2239 11770 2261
rect 11602 2233 11713 2239
rect 11602 2225 11643 2233
rect 11602 2205 11610 2225
rect 11629 2205 11643 2225
rect 11602 2203 11643 2205
rect 11671 2225 11713 2233
rect 11671 2205 11687 2225
rect 11706 2205 11713 2225
rect 11671 2203 11713 2205
rect 11602 2188 11713 2203
rect 11406 2132 11474 2142
rect 11406 2099 11423 2132
rect 11463 2099 11474 2132
rect 11406 2087 11474 2099
rect 11406 2085 11470 2087
rect 11941 2068 11978 2292
rect 12254 2288 12318 2300
rect 12358 2070 12385 2440
rect 12573 2435 12610 2445
rect 12669 2465 12756 2475
rect 12669 2445 12678 2465
rect 12698 2445 12756 2465
rect 12669 2436 12756 2445
rect 12669 2435 12706 2436
rect 12449 2422 12519 2427
rect 12444 2416 12519 2422
rect 12444 2383 12452 2416
rect 12505 2383 12519 2416
rect 12725 2383 12756 2436
rect 12786 2465 12823 2544
rect 12938 2475 12969 2476
rect 12786 2445 12795 2465
rect 12815 2445 12823 2465
rect 12786 2435 12823 2445
rect 12882 2468 12969 2475
rect 12882 2465 12943 2468
rect 12882 2445 12891 2465
rect 12911 2448 12943 2465
rect 12964 2448 12969 2468
rect 12911 2445 12969 2448
rect 12882 2438 12969 2445
rect 12994 2465 13031 2607
rect 13297 2606 13334 2607
rect 13146 2475 13182 2476
rect 12994 2445 13003 2465
rect 13023 2445 13031 2465
rect 12882 2436 12938 2438
rect 12882 2435 12919 2436
rect 12994 2435 13031 2445
rect 13090 2465 13238 2475
rect 13338 2472 13434 2474
rect 13090 2445 13099 2465
rect 13119 2445 13209 2465
rect 13229 2445 13238 2465
rect 13090 2439 13238 2445
rect 13090 2436 13154 2439
rect 13090 2435 13127 2436
rect 13146 2409 13154 2436
rect 13175 2436 13238 2439
rect 13296 2465 13434 2472
rect 13296 2445 13305 2465
rect 13325 2445 13434 2465
rect 13296 2436 13434 2445
rect 13175 2409 13182 2436
rect 13201 2435 13238 2436
rect 13297 2435 13334 2436
rect 13146 2384 13182 2409
rect 12444 2382 12527 2383
rect 12617 2382 12658 2383
rect 12444 2375 12658 2382
rect 12444 2358 12627 2375
rect 12444 2325 12457 2358
rect 12510 2355 12627 2358
rect 12647 2355 12658 2375
rect 12510 2347 12658 2355
rect 12725 2379 13084 2383
rect 12725 2374 13047 2379
rect 12725 2350 12838 2374
rect 12862 2355 13047 2374
rect 13071 2355 13084 2379
rect 12862 2350 13084 2355
rect 12725 2347 13084 2350
rect 13146 2347 13181 2384
rect 13249 2381 13349 2384
rect 13249 2377 13316 2381
rect 13249 2351 13261 2377
rect 13287 2355 13316 2377
rect 13342 2355 13349 2381
rect 13287 2351 13349 2355
rect 13249 2347 13349 2351
rect 12510 2325 12527 2347
rect 12725 2326 12756 2347
rect 13146 2326 13182 2347
rect 12568 2325 12605 2326
rect 12444 2311 12527 2325
rect 12217 2068 12385 2070
rect 11941 2067 12385 2068
rect 11185 2037 12385 2067
rect 12455 2101 12527 2311
rect 12567 2316 12605 2325
rect 12567 2296 12576 2316
rect 12596 2296 12605 2316
rect 12567 2288 12605 2296
rect 12671 2320 12756 2326
rect 12781 2325 12818 2326
rect 12671 2300 12679 2320
rect 12699 2300 12756 2320
rect 12671 2292 12756 2300
rect 12780 2316 12818 2325
rect 12780 2296 12789 2316
rect 12809 2296 12818 2316
rect 12671 2291 12707 2292
rect 12780 2288 12818 2296
rect 12884 2320 12969 2326
rect 12989 2325 13026 2326
rect 12884 2300 12892 2320
rect 12912 2319 12969 2320
rect 12912 2300 12941 2319
rect 12884 2299 12941 2300
rect 12962 2299 12969 2319
rect 12884 2292 12969 2299
rect 12988 2316 13026 2325
rect 12988 2296 12997 2316
rect 13017 2296 13026 2316
rect 12884 2291 12920 2292
rect 12988 2288 13026 2296
rect 13092 2320 13236 2326
rect 13092 2300 13100 2320
rect 13120 2300 13208 2320
rect 13228 2300 13236 2320
rect 13092 2292 13236 2300
rect 13092 2291 13128 2292
rect 13200 2291 13236 2292
rect 13302 2325 13339 2326
rect 13302 2324 13340 2325
rect 13302 2316 13366 2324
rect 13302 2296 13311 2316
rect 13331 2302 13366 2316
rect 13386 2302 13389 2322
rect 13331 2297 13389 2302
rect 13331 2296 13366 2297
rect 12568 2259 12605 2288
rect 12569 2257 12605 2259
rect 12781 2257 12818 2288
rect 12569 2235 12818 2257
rect 12650 2229 12761 2235
rect 12650 2221 12691 2229
rect 12650 2201 12658 2221
rect 12677 2201 12691 2221
rect 12650 2199 12691 2201
rect 12719 2221 12761 2229
rect 12719 2201 12735 2221
rect 12754 2201 12761 2221
rect 12719 2199 12761 2201
rect 12650 2184 12761 2199
rect 12455 2062 12474 2101
rect 12519 2062 12527 2101
rect 12455 2045 12527 2062
rect 12989 2089 13026 2288
rect 13302 2284 13366 2296
rect 12989 2083 13030 2089
rect 13406 2085 13433 2436
rect 13265 2083 13433 2085
rect 12989 2057 13433 2083
rect 11185 1990 11250 2037
rect 11185 1972 11208 1990
rect 11226 1972 11250 1990
rect 12098 2017 12133 2019
rect 12098 2015 12202 2017
rect 12991 2015 13030 2057
rect 13265 2056 13433 2057
rect 12098 2008 13032 2015
rect 12098 2007 12149 2008
rect 12098 1987 12101 2007
rect 12126 1988 12149 2007
rect 12181 1988 13032 2008
rect 12126 1987 13032 1988
rect 12098 1980 13032 1987
rect 12371 1979 13032 1980
rect 11185 1951 11250 1972
rect 11462 1962 11502 1965
rect 11462 1958 12365 1962
rect 11462 1938 12339 1958
rect 12359 1938 12365 1958
rect 11462 1935 12365 1938
rect 11186 1891 11251 1911
rect 11186 1873 11210 1891
rect 11228 1873 11251 1891
rect 11186 1846 11251 1873
rect 11462 1846 11502 1935
rect 11946 1933 12362 1935
rect 11946 1932 12287 1933
rect 11603 1901 11713 1915
rect 11603 1898 11646 1901
rect 11603 1893 11607 1898
rect 11185 1811 11502 1846
rect 11525 1871 11607 1893
rect 11636 1871 11646 1898
rect 11674 1874 11681 1901
rect 11710 1893 11713 1901
rect 11710 1874 11775 1893
rect 11674 1871 11775 1874
rect 11525 1869 11775 1871
rect 10143 1788 10165 1806
rect 10183 1788 10208 1806
rect 10143 1769 10208 1788
rect 9836 1744 9873 1745
rect 9259 1723 9295 1744
rect 9685 1723 9716 1744
rect 9923 1739 9931 1748
rect 9920 1723 9931 1739
rect 9092 1719 9192 1723
rect 9092 1715 9154 1719
rect 9092 1689 9099 1715
rect 9125 1693 9154 1715
rect 9180 1693 9192 1719
rect 9125 1689 9192 1693
rect 9092 1686 9192 1689
rect 9260 1686 9295 1723
rect 9357 1720 9716 1723
rect 9357 1715 9579 1720
rect 9357 1691 9370 1715
rect 9394 1696 9579 1715
rect 9603 1696 9716 1720
rect 9394 1691 9716 1696
rect 9357 1687 9716 1691
rect 9783 1715 9931 1723
rect 9783 1695 9794 1715
rect 9814 1706 9931 1715
rect 9980 1739 9987 1748
rect 9980 1706 9988 1739
rect 11186 1735 11251 1811
rect 11525 1790 11562 1869
rect 11603 1856 11713 1869
rect 11677 1800 11708 1801
rect 11525 1770 11534 1790
rect 11554 1770 11562 1790
rect 11525 1760 11562 1770
rect 11621 1790 11708 1800
rect 11621 1770 11630 1790
rect 11650 1770 11708 1790
rect 11621 1761 11708 1770
rect 11621 1760 11658 1761
rect 9814 1695 9988 1706
rect 9783 1688 9988 1695
rect 9783 1687 9824 1688
rect 9259 1661 9295 1686
rect 9107 1634 9144 1635
rect 9203 1634 9240 1635
rect 9259 1634 9266 1661
rect 8783 1609 8791 1629
rect 8811 1609 8820 1629
rect 8637 1598 8668 1599
rect 8632 1530 8742 1543
rect 8783 1530 8820 1609
rect 9007 1625 9145 1634
rect 9007 1605 9116 1625
rect 9136 1605 9145 1625
rect 9007 1598 9145 1605
rect 9203 1631 9266 1634
rect 9287 1634 9295 1661
rect 9314 1634 9351 1635
rect 9287 1631 9351 1634
rect 9203 1625 9351 1631
rect 9203 1605 9212 1625
rect 9232 1605 9322 1625
rect 9342 1605 9351 1625
rect 9007 1596 9103 1598
rect 9203 1595 9351 1605
rect 9410 1625 9447 1635
rect 9522 1634 9559 1635
rect 9503 1632 9559 1634
rect 9410 1605 9418 1625
rect 9438 1605 9447 1625
rect 9259 1594 9295 1595
rect 8570 1528 8820 1530
rect 8570 1525 8671 1528
rect 8570 1506 8635 1525
rect 8632 1498 8635 1506
rect 8664 1498 8671 1525
rect 8699 1501 8709 1528
rect 8738 1506 8820 1528
rect 8738 1501 8742 1506
rect 8699 1498 8742 1501
rect 8632 1484 8742 1498
rect 8058 1466 8399 1467
rect 7983 1461 8399 1466
rect 9107 1463 9144 1464
rect 9410 1463 9447 1605
rect 9472 1625 9559 1632
rect 9472 1622 9530 1625
rect 9472 1602 9477 1622
rect 9498 1605 9530 1622
rect 9550 1605 9559 1625
rect 9498 1602 9559 1605
rect 9472 1595 9559 1602
rect 9618 1625 9655 1635
rect 9618 1605 9626 1625
rect 9646 1605 9655 1625
rect 9472 1594 9503 1595
rect 9618 1526 9655 1605
rect 9685 1634 9716 1687
rect 9920 1685 9988 1688
rect 9920 1643 9932 1685
rect 9981 1643 9988 1685
rect 9735 1634 9772 1635
rect 9685 1625 9772 1634
rect 9685 1605 9743 1625
rect 9763 1605 9772 1625
rect 9685 1595 9772 1605
rect 9831 1625 9868 1635
rect 9920 1630 9988 1643
rect 10143 1707 10208 1724
rect 10143 1689 10167 1707
rect 10185 1689 10208 1707
rect 11186 1717 11208 1735
rect 11226 1717 11251 1735
rect 11186 1696 11251 1717
rect 11399 1715 11464 1724
rect 9831 1605 9839 1625
rect 9859 1605 9868 1625
rect 9685 1594 9716 1595
rect 9680 1526 9790 1539
rect 9831 1526 9868 1605
rect 10143 1550 10208 1689
rect 11399 1678 11409 1715
rect 11449 1707 11464 1715
rect 11677 1708 11708 1761
rect 11738 1790 11775 1869
rect 11890 1800 11921 1801
rect 11738 1770 11747 1790
rect 11767 1770 11775 1790
rect 11738 1760 11775 1770
rect 11834 1793 11921 1800
rect 11834 1790 11895 1793
rect 11834 1770 11843 1790
rect 11863 1773 11895 1790
rect 11916 1773 11921 1793
rect 11863 1770 11921 1773
rect 11834 1763 11921 1770
rect 11946 1790 11983 1932
rect 12249 1931 12286 1932
rect 12098 1800 12134 1801
rect 11946 1770 11955 1790
rect 11975 1770 11983 1790
rect 11834 1761 11890 1763
rect 11834 1760 11871 1761
rect 11946 1760 11983 1770
rect 12042 1790 12190 1800
rect 12290 1797 12386 1799
rect 12042 1770 12051 1790
rect 12071 1770 12161 1790
rect 12181 1770 12190 1790
rect 12042 1764 12190 1770
rect 12042 1761 12106 1764
rect 12042 1760 12079 1761
rect 12098 1734 12106 1761
rect 12127 1761 12190 1764
rect 12248 1790 12386 1797
rect 12248 1770 12257 1790
rect 12277 1770 12386 1790
rect 12248 1761 12386 1770
rect 12127 1734 12134 1761
rect 12153 1760 12190 1761
rect 12249 1760 12286 1761
rect 12098 1709 12134 1734
rect 11569 1707 11610 1708
rect 11449 1700 11610 1707
rect 11449 1680 11579 1700
rect 11599 1680 11610 1700
rect 11449 1678 11610 1680
rect 11399 1672 11610 1678
rect 11677 1704 12036 1708
rect 11677 1699 11999 1704
rect 11677 1675 11790 1699
rect 11814 1680 11999 1699
rect 12023 1680 12036 1704
rect 11814 1675 12036 1680
rect 11677 1672 12036 1675
rect 12098 1672 12133 1709
rect 12201 1706 12301 1709
rect 12201 1702 12268 1706
rect 12201 1676 12213 1702
rect 12239 1680 12268 1702
rect 12294 1680 12301 1706
rect 12239 1676 12301 1680
rect 12201 1672 12301 1676
rect 11399 1659 11466 1672
rect 11191 1636 11247 1656
rect 11191 1618 11210 1636
rect 11228 1618 11247 1636
rect 11191 1583 11247 1618
rect 10143 1544 10165 1550
rect 9618 1524 9868 1526
rect 9618 1521 9719 1524
rect 9618 1502 9683 1521
rect 9680 1494 9683 1502
rect 9712 1494 9719 1521
rect 9747 1497 9757 1524
rect 9786 1502 9868 1524
rect 9897 1532 10165 1544
rect 10183 1532 10208 1550
rect 9897 1509 10208 1532
rect 9897 1508 9952 1509
rect 9786 1497 9790 1502
rect 9747 1494 9790 1497
rect 9680 1480 9790 1494
rect 9106 1462 9447 1463
rect 7983 1441 7986 1461
rect 8006 1441 8399 1461
rect 9031 1461 9447 1462
rect 9897 1461 9940 1508
rect 11153 1505 11247 1583
rect 11399 1638 11413 1659
rect 11449 1638 11466 1659
rect 11677 1651 11708 1672
rect 12098 1651 12134 1672
rect 11520 1650 11557 1651
rect 11399 1631 11466 1638
rect 11519 1641 11557 1650
rect 9031 1457 9940 1461
rect 1651 1367 1679 1381
rect 2775 1378 2932 1391
rect 6906 1406 7723 1408
rect 8156 1406 8245 1409
rect 6906 1397 8245 1406
rect 453 1332 1679 1367
rect 6906 1359 8168 1397
rect 8193 1362 8212 1397
rect 8237 1362 8245 1397
rect 8350 1408 8395 1441
rect 9031 1437 9034 1457
rect 9054 1437 9940 1457
rect 9408 1432 9940 1437
rect 10148 1451 10207 1473
rect 10148 1433 10167 1451
rect 10185 1433 10207 1451
rect 9196 1408 9295 1410
rect 8350 1398 9295 1408
rect 8350 1372 9218 1398
rect 8351 1371 9218 1372
rect 8193 1359 8245 1362
rect 6906 1351 8245 1359
rect 9196 1360 9218 1371
rect 9243 1363 9262 1398
rect 9287 1363 9295 1398
rect 9243 1360 9295 1363
rect 9196 1352 9295 1360
rect 9222 1351 9294 1352
rect 6906 1350 8244 1351
rect 6906 1348 7723 1350
rect 7497 1344 7723 1348
rect 453 1256 538 1332
rect 896 1330 1000 1332
rect 1231 1330 1272 1332
rect 10148 1256 10207 1433
rect 11153 1364 11246 1505
rect 11399 1479 11464 1631
rect 11519 1621 11528 1641
rect 11548 1621 11557 1641
rect 11519 1613 11557 1621
rect 11623 1645 11708 1651
rect 11733 1650 11770 1651
rect 11623 1625 11631 1645
rect 11651 1625 11708 1645
rect 11623 1617 11708 1625
rect 11732 1641 11770 1650
rect 11732 1621 11741 1641
rect 11761 1621 11770 1641
rect 11623 1616 11659 1617
rect 11732 1613 11770 1621
rect 11836 1645 11921 1651
rect 11941 1650 11978 1651
rect 11836 1625 11844 1645
rect 11864 1644 11921 1645
rect 11864 1625 11893 1644
rect 11836 1624 11893 1625
rect 11914 1624 11921 1644
rect 11836 1617 11921 1624
rect 11940 1641 11978 1650
rect 11940 1621 11949 1641
rect 11969 1621 11978 1641
rect 11836 1616 11872 1617
rect 11940 1613 11978 1621
rect 12044 1645 12188 1651
rect 12044 1625 12052 1645
rect 12072 1625 12160 1645
rect 12180 1625 12188 1645
rect 12044 1617 12188 1625
rect 12044 1616 12080 1617
rect 12152 1616 12188 1617
rect 12254 1650 12291 1651
rect 12254 1649 12292 1650
rect 12254 1641 12318 1649
rect 12254 1621 12263 1641
rect 12283 1627 12318 1641
rect 12338 1627 12341 1647
rect 12283 1622 12341 1627
rect 12283 1621 12318 1622
rect 11520 1584 11557 1613
rect 11521 1582 11557 1584
rect 11733 1582 11770 1613
rect 11521 1560 11770 1582
rect 11602 1554 11713 1560
rect 11602 1546 11643 1554
rect 11602 1526 11610 1546
rect 11629 1526 11643 1546
rect 11602 1524 11643 1526
rect 11671 1546 11713 1554
rect 11671 1526 11687 1546
rect 11706 1526 11713 1546
rect 11671 1524 11713 1526
rect 11602 1509 11713 1524
rect 11941 1514 11978 1613
rect 12254 1609 12318 1621
rect 12358 1570 12385 1761
rect 11604 1500 11708 1509
rect 11392 1469 11513 1479
rect 11392 1467 11461 1469
rect 11392 1426 11405 1467
rect 11442 1428 11461 1467
rect 11498 1428 11513 1469
rect 11442 1426 11513 1428
rect 11392 1408 11513 1426
rect 11604 1364 11708 1373
rect 11939 1364 11980 1514
rect 11153 1362 11980 1364
rect 11161 1361 11980 1362
rect 12359 1480 12384 1570
rect 13519 1538 13618 3095
rect 13724 1731 13823 4632
rect 14214 4615 14245 4636
rect 14635 4615 14671 4636
rect 14057 4614 14094 4615
rect 14056 4605 14094 4614
rect 14056 4585 14065 4605
rect 14085 4585 14094 4605
rect 14056 4577 14094 4585
rect 14160 4609 14245 4615
rect 14270 4614 14307 4615
rect 14160 4589 14168 4609
rect 14188 4589 14245 4609
rect 14160 4581 14245 4589
rect 14269 4605 14307 4614
rect 14269 4585 14278 4605
rect 14298 4585 14307 4605
rect 14160 4580 14196 4581
rect 14269 4577 14307 4585
rect 14373 4609 14458 4615
rect 14478 4614 14515 4615
rect 14373 4589 14381 4609
rect 14401 4608 14458 4609
rect 14401 4589 14430 4608
rect 14373 4588 14430 4589
rect 14451 4588 14458 4608
rect 14373 4581 14458 4588
rect 14477 4605 14515 4614
rect 14477 4585 14486 4605
rect 14506 4585 14515 4605
rect 14373 4580 14409 4581
rect 14477 4577 14515 4585
rect 14581 4609 14725 4615
rect 14581 4589 14589 4609
rect 14609 4589 14697 4609
rect 14717 4589 14725 4609
rect 14581 4581 14725 4589
rect 14581 4580 14617 4581
rect 14689 4580 14725 4581
rect 14791 4614 14828 4615
rect 14791 4613 14829 4614
rect 14791 4605 14855 4613
rect 14791 4585 14800 4605
rect 14820 4591 14855 4605
rect 14875 4591 14878 4611
rect 14820 4586 14878 4591
rect 14820 4585 14855 4586
rect 14057 4548 14094 4577
rect 14058 4546 14094 4548
rect 14270 4546 14307 4577
rect 14058 4524 14307 4546
rect 14139 4518 14250 4524
rect 14139 4510 14180 4518
rect 14139 4490 14147 4510
rect 14166 4490 14180 4510
rect 14139 4488 14180 4490
rect 14208 4510 14250 4518
rect 14208 4490 14224 4510
rect 14243 4490 14250 4510
rect 14208 4488 14250 4490
rect 14139 4473 14250 4488
rect 14478 4456 14515 4577
rect 14791 4573 14855 4585
rect 14596 4456 14625 4460
rect 14895 4458 14922 4725
rect 14754 4456 14922 4458
rect 14478 4430 14922 4456
rect 14437 4162 14482 4171
rect 14437 4124 14447 4162
rect 14472 4124 14482 4162
rect 14437 4113 14482 4124
rect 14440 4105 14482 4113
rect 14440 3400 14483 4105
rect 14596 3491 14625 4430
rect 14754 4429 14922 4430
rect 15326 4280 15410 4284
rect 15878 4280 15966 7131
rect 16505 7118 16560 7130
rect 16505 7084 16523 7118
rect 16552 7084 16560 7118
rect 16505 7058 16560 7084
rect 16112 7025 16280 7026
rect 16505 7025 16522 7058
rect 16112 7024 16522 7025
rect 16551 7024 16560 7058
rect 16112 6999 16560 7024
rect 16112 6997 16280 6999
rect 16112 6730 16139 6997
rect 16505 6993 16560 6999
rect 16179 6870 16243 6882
rect 16519 6878 16556 6993
rect 16784 6967 16895 6982
rect 16784 6965 16826 6967
rect 16784 6945 16791 6965
rect 16810 6945 16826 6965
rect 16784 6937 16826 6945
rect 16854 6965 16895 6967
rect 16854 6945 16868 6965
rect 16887 6945 16895 6965
rect 16854 6937 16895 6945
rect 16784 6931 16895 6937
rect 16727 6909 16976 6931
rect 16727 6878 16764 6909
rect 16940 6907 16976 6909
rect 16940 6878 16977 6907
rect 16179 6869 16214 6870
rect 16156 6864 16214 6869
rect 16156 6844 16159 6864
rect 16179 6850 16214 6864
rect 16234 6850 16243 6870
rect 16179 6842 16243 6850
rect 16205 6841 16243 6842
rect 16206 6840 16243 6841
rect 16309 6874 16345 6875
rect 16417 6874 16453 6875
rect 16309 6866 16453 6874
rect 16309 6846 16317 6866
rect 16337 6846 16425 6866
rect 16445 6846 16453 6866
rect 16309 6840 16453 6846
rect 16519 6870 16557 6878
rect 16625 6874 16661 6875
rect 16519 6850 16528 6870
rect 16548 6850 16557 6870
rect 16519 6841 16557 6850
rect 16576 6867 16661 6874
rect 16576 6847 16583 6867
rect 16604 6866 16661 6867
rect 16604 6847 16633 6866
rect 16576 6846 16633 6847
rect 16653 6846 16661 6866
rect 16519 6840 16556 6841
rect 16576 6840 16661 6846
rect 16727 6870 16765 6878
rect 16838 6874 16874 6875
rect 16727 6850 16736 6870
rect 16756 6850 16765 6870
rect 16727 6841 16765 6850
rect 16789 6866 16874 6874
rect 16789 6846 16846 6866
rect 16866 6846 16874 6866
rect 16727 6840 16764 6841
rect 16789 6840 16874 6846
rect 16940 6870 16978 6878
rect 16940 6850 16949 6870
rect 16969 6850 16978 6870
rect 16940 6841 16978 6850
rect 16940 6840 16977 6841
rect 16363 6819 16399 6840
rect 16789 6819 16820 6840
rect 17034 6823 17105 7476
rect 17620 7410 17663 8123
rect 18280 8034 18375 8054
rect 18280 7990 18300 8034
rect 18360 7990 18375 8034
rect 18280 7694 18375 7990
rect 18280 7653 18313 7694
rect 18349 7653 18375 7694
rect 18475 7733 18537 8204
rect 19817 8144 19854 8145
rect 20120 8144 20157 8286
rect 20182 8306 20269 8313
rect 20182 8303 20240 8306
rect 20182 8283 20187 8303
rect 20208 8286 20240 8303
rect 20260 8286 20269 8306
rect 20208 8283 20269 8286
rect 20182 8276 20269 8283
rect 20328 8306 20365 8316
rect 20328 8286 20336 8306
rect 20356 8286 20365 8306
rect 20182 8275 20213 8276
rect 20328 8207 20365 8286
rect 20395 8315 20426 8368
rect 20639 8361 20654 8369
rect 20694 8361 20704 8398
rect 20639 8352 20704 8361
rect 20852 8359 20917 8380
rect 20852 8341 20877 8359
rect 20895 8341 20917 8359
rect 20445 8315 20482 8316
rect 20395 8306 20482 8315
rect 20395 8286 20453 8306
rect 20473 8286 20482 8306
rect 20395 8276 20482 8286
rect 20541 8306 20578 8316
rect 20541 8286 20549 8306
rect 20569 8286 20578 8306
rect 20395 8275 20426 8276
rect 20390 8207 20500 8220
rect 20541 8207 20578 8286
rect 20852 8265 20917 8341
rect 20328 8205 20578 8207
rect 20328 8202 20429 8205
rect 20328 8183 20393 8202
rect 20390 8175 20393 8183
rect 20422 8175 20429 8202
rect 20457 8178 20467 8205
rect 20496 8183 20578 8205
rect 20601 8230 20918 8265
rect 20496 8178 20500 8183
rect 20457 8175 20500 8178
rect 20390 8161 20500 8175
rect 19816 8143 20157 8144
rect 19741 8141 20157 8143
rect 20601 8141 20641 8230
rect 20852 8203 20917 8230
rect 20852 8185 20875 8203
rect 20893 8185 20917 8203
rect 20852 8165 20917 8185
rect 19738 8138 20641 8141
rect 19738 8118 19744 8138
rect 19764 8118 20641 8138
rect 19738 8114 20641 8118
rect 20601 8111 20641 8114
rect 20853 8104 20918 8125
rect 19071 8096 19732 8097
rect 19071 8089 20005 8096
rect 19071 8088 19977 8089
rect 19071 8068 19922 8088
rect 19954 8069 19977 8088
rect 20002 8069 20005 8089
rect 19954 8068 20005 8069
rect 19071 8061 20005 8068
rect 18670 8019 18838 8020
rect 19073 8019 19112 8061
rect 19901 8059 20005 8061
rect 19970 8057 20005 8059
rect 20853 8086 20877 8104
rect 20895 8086 20918 8104
rect 20853 8039 20918 8086
rect 18670 7993 19114 8019
rect 18670 7991 18838 7993
rect 18475 7714 18539 7733
rect 18475 7675 18492 7714
rect 18526 7675 18539 7714
rect 18475 7656 18539 7675
rect 18280 7627 18375 7653
rect 18670 7640 18697 7991
rect 19073 7987 19114 7993
rect 18737 7780 18801 7792
rect 19077 7788 19114 7987
rect 19576 8014 19648 8031
rect 19576 7975 19584 8014
rect 19629 7975 19648 8014
rect 19342 7877 19453 7892
rect 19342 7875 19384 7877
rect 19342 7855 19349 7875
rect 19368 7855 19384 7875
rect 19342 7847 19384 7855
rect 19412 7875 19453 7877
rect 19412 7855 19426 7875
rect 19445 7855 19453 7875
rect 19412 7847 19453 7855
rect 19342 7841 19453 7847
rect 19285 7819 19534 7841
rect 19285 7788 19322 7819
rect 19498 7817 19534 7819
rect 19498 7788 19535 7817
rect 18737 7779 18772 7780
rect 18714 7774 18772 7779
rect 18714 7754 18717 7774
rect 18737 7760 18772 7774
rect 18792 7760 18801 7780
rect 18737 7752 18801 7760
rect 18763 7751 18801 7752
rect 18764 7750 18801 7751
rect 18867 7784 18903 7785
rect 18975 7784 19011 7785
rect 18867 7776 19011 7784
rect 18867 7756 18875 7776
rect 18895 7756 18983 7776
rect 19003 7756 19011 7776
rect 18867 7750 19011 7756
rect 19077 7780 19115 7788
rect 19183 7784 19219 7785
rect 19077 7760 19086 7780
rect 19106 7760 19115 7780
rect 19077 7751 19115 7760
rect 19134 7777 19219 7784
rect 19134 7757 19141 7777
rect 19162 7776 19219 7777
rect 19162 7757 19191 7776
rect 19134 7756 19191 7757
rect 19211 7756 19219 7776
rect 19077 7750 19114 7751
rect 19134 7750 19219 7756
rect 19285 7780 19323 7788
rect 19396 7784 19432 7785
rect 19285 7760 19294 7780
rect 19314 7760 19323 7780
rect 19285 7751 19323 7760
rect 19347 7776 19432 7784
rect 19347 7756 19404 7776
rect 19424 7756 19432 7776
rect 19285 7750 19322 7751
rect 19347 7750 19432 7756
rect 19498 7780 19536 7788
rect 19498 7760 19507 7780
rect 19527 7760 19536 7780
rect 19498 7751 19536 7760
rect 19576 7765 19648 7975
rect 19718 8009 20918 8039
rect 19718 8008 20162 8009
rect 19718 8006 19886 8008
rect 19576 7751 19659 7765
rect 19498 7750 19535 7751
rect 18921 7729 18957 7750
rect 19347 7729 19378 7750
rect 19576 7729 19593 7751
rect 18754 7725 18854 7729
rect 18754 7721 18816 7725
rect 18754 7695 18761 7721
rect 18787 7699 18816 7721
rect 18842 7699 18854 7725
rect 18787 7695 18854 7699
rect 18754 7692 18854 7695
rect 18922 7692 18957 7729
rect 19019 7726 19378 7729
rect 19019 7721 19241 7726
rect 19019 7697 19032 7721
rect 19056 7702 19241 7721
rect 19265 7702 19378 7726
rect 19056 7697 19378 7702
rect 19019 7693 19378 7697
rect 19445 7721 19593 7729
rect 19445 7701 19456 7721
rect 19476 7718 19593 7721
rect 19646 7718 19659 7751
rect 19476 7701 19659 7718
rect 19445 7694 19659 7701
rect 19445 7693 19486 7694
rect 19576 7693 19659 7694
rect 18921 7667 18957 7692
rect 18769 7640 18806 7641
rect 18865 7640 18902 7641
rect 18921 7640 18928 7667
rect 18669 7631 18807 7640
rect 18669 7611 18778 7631
rect 18798 7611 18807 7631
rect 18669 7604 18807 7611
rect 18865 7637 18928 7640
rect 18949 7640 18957 7667
rect 18976 7640 19013 7641
rect 18949 7637 19013 7640
rect 18865 7631 19013 7637
rect 18865 7611 18874 7631
rect 18894 7611 18984 7631
rect 19004 7611 19013 7631
rect 18669 7602 18765 7604
rect 18865 7601 19013 7611
rect 19072 7631 19109 7641
rect 19184 7640 19221 7641
rect 19165 7638 19221 7640
rect 19072 7611 19080 7631
rect 19100 7611 19109 7631
rect 18921 7600 18957 7601
rect 18769 7469 18806 7470
rect 19072 7469 19109 7611
rect 19134 7631 19221 7638
rect 19134 7628 19192 7631
rect 19134 7608 19139 7628
rect 19160 7611 19192 7628
rect 19212 7611 19221 7631
rect 19160 7608 19221 7611
rect 19134 7601 19221 7608
rect 19280 7631 19317 7641
rect 19280 7611 19288 7631
rect 19308 7611 19317 7631
rect 19134 7600 19165 7601
rect 19280 7532 19317 7611
rect 19347 7640 19378 7693
rect 19584 7660 19598 7693
rect 19651 7660 19659 7693
rect 19584 7654 19659 7660
rect 19584 7649 19654 7654
rect 19397 7640 19434 7641
rect 19347 7631 19434 7640
rect 19347 7611 19405 7631
rect 19425 7611 19434 7631
rect 19347 7601 19434 7611
rect 19493 7631 19530 7641
rect 19718 7636 19745 8006
rect 19785 7776 19849 7788
rect 20125 7784 20162 8008
rect 20633 7989 20697 7991
rect 20629 7977 20697 7989
rect 20629 7944 20640 7977
rect 20680 7944 20697 7977
rect 20629 7934 20697 7944
rect 20390 7873 20501 7888
rect 20390 7871 20432 7873
rect 20390 7851 20397 7871
rect 20416 7851 20432 7871
rect 20390 7843 20432 7851
rect 20460 7871 20501 7873
rect 20460 7851 20474 7871
rect 20493 7851 20501 7871
rect 20460 7843 20501 7851
rect 20390 7837 20501 7843
rect 20333 7815 20582 7837
rect 20333 7784 20370 7815
rect 20546 7813 20582 7815
rect 20546 7784 20583 7813
rect 19785 7775 19820 7776
rect 19762 7770 19820 7775
rect 19762 7750 19765 7770
rect 19785 7756 19820 7770
rect 19840 7756 19849 7776
rect 19785 7748 19849 7756
rect 19811 7747 19849 7748
rect 19812 7746 19849 7747
rect 19915 7780 19951 7781
rect 20023 7780 20059 7781
rect 19915 7772 20059 7780
rect 19915 7752 19923 7772
rect 19943 7752 20031 7772
rect 20051 7752 20059 7772
rect 19915 7746 20059 7752
rect 20125 7776 20163 7784
rect 20231 7780 20267 7781
rect 20125 7756 20134 7776
rect 20154 7756 20163 7776
rect 20125 7747 20163 7756
rect 20182 7773 20267 7780
rect 20182 7753 20189 7773
rect 20210 7772 20267 7773
rect 20210 7753 20239 7772
rect 20182 7752 20239 7753
rect 20259 7752 20267 7772
rect 20125 7746 20162 7747
rect 20182 7746 20267 7752
rect 20333 7776 20371 7784
rect 20444 7780 20480 7781
rect 20333 7756 20342 7776
rect 20362 7756 20371 7776
rect 20333 7747 20371 7756
rect 20395 7772 20480 7780
rect 20395 7752 20452 7772
rect 20472 7752 20480 7772
rect 20333 7746 20370 7747
rect 20395 7746 20480 7752
rect 20546 7776 20584 7784
rect 20546 7756 20555 7776
rect 20575 7756 20584 7776
rect 20546 7747 20584 7756
rect 20633 7750 20697 7934
rect 20853 7808 20918 8009
rect 20853 7790 20875 7808
rect 20893 7790 20918 7808
rect 20853 7771 20918 7790
rect 20546 7746 20583 7747
rect 19969 7725 20005 7746
rect 20395 7725 20426 7746
rect 20633 7741 20641 7750
rect 20630 7725 20641 7741
rect 19802 7721 19902 7725
rect 19802 7717 19864 7721
rect 19802 7691 19809 7717
rect 19835 7695 19864 7717
rect 19890 7695 19902 7721
rect 19835 7691 19902 7695
rect 19802 7688 19902 7691
rect 19970 7688 20005 7725
rect 20067 7722 20426 7725
rect 20067 7717 20289 7722
rect 20067 7693 20080 7717
rect 20104 7698 20289 7717
rect 20313 7698 20426 7722
rect 20104 7693 20426 7698
rect 20067 7689 20426 7693
rect 20493 7717 20641 7725
rect 20493 7697 20504 7717
rect 20524 7708 20641 7717
rect 20690 7741 20697 7750
rect 20690 7708 20698 7741
rect 20524 7697 20698 7708
rect 20493 7690 20698 7697
rect 20493 7689 20534 7690
rect 19969 7663 20005 7688
rect 19817 7636 19854 7637
rect 19913 7636 19950 7637
rect 19969 7636 19976 7663
rect 19493 7611 19501 7631
rect 19521 7611 19530 7631
rect 19347 7600 19378 7601
rect 19342 7532 19452 7545
rect 19493 7532 19530 7611
rect 19717 7627 19855 7636
rect 19717 7607 19826 7627
rect 19846 7607 19855 7627
rect 19717 7600 19855 7607
rect 19913 7633 19976 7636
rect 19997 7636 20005 7663
rect 20024 7636 20061 7637
rect 19997 7633 20061 7636
rect 19913 7627 20061 7633
rect 19913 7607 19922 7627
rect 19942 7607 20032 7627
rect 20052 7607 20061 7627
rect 19717 7598 19813 7600
rect 19913 7597 20061 7607
rect 20120 7627 20157 7637
rect 20232 7636 20269 7637
rect 20213 7634 20269 7636
rect 20120 7607 20128 7627
rect 20148 7607 20157 7627
rect 19969 7596 20005 7597
rect 19280 7530 19530 7532
rect 19280 7527 19381 7530
rect 19280 7508 19345 7527
rect 19342 7500 19345 7508
rect 19374 7500 19381 7527
rect 19409 7503 19419 7530
rect 19448 7508 19530 7530
rect 19448 7503 19452 7508
rect 19409 7500 19452 7503
rect 19342 7486 19452 7500
rect 18768 7468 19109 7469
rect 18693 7463 19109 7468
rect 19817 7465 19854 7466
rect 20120 7465 20157 7607
rect 20182 7627 20269 7634
rect 20182 7624 20240 7627
rect 20182 7604 20187 7624
rect 20208 7607 20240 7624
rect 20260 7607 20269 7627
rect 20208 7604 20269 7607
rect 20182 7597 20269 7604
rect 20328 7627 20365 7637
rect 20328 7607 20336 7627
rect 20356 7607 20365 7627
rect 20182 7596 20213 7597
rect 20328 7528 20365 7607
rect 20395 7636 20426 7689
rect 20630 7687 20698 7690
rect 20630 7645 20642 7687
rect 20691 7645 20698 7687
rect 20445 7636 20482 7637
rect 20395 7627 20482 7636
rect 20395 7607 20453 7627
rect 20473 7607 20482 7627
rect 20395 7597 20482 7607
rect 20541 7627 20578 7637
rect 20630 7632 20698 7645
rect 20853 7709 20918 7726
rect 20853 7691 20877 7709
rect 20895 7691 20918 7709
rect 20541 7607 20549 7627
rect 20569 7607 20578 7627
rect 20395 7596 20426 7597
rect 20390 7528 20500 7541
rect 20541 7528 20578 7607
rect 20853 7552 20918 7691
rect 20853 7546 20875 7552
rect 20328 7526 20578 7528
rect 20328 7523 20429 7526
rect 20328 7504 20393 7523
rect 20390 7496 20393 7504
rect 20422 7496 20429 7523
rect 20457 7499 20467 7526
rect 20496 7504 20578 7526
rect 20607 7534 20875 7546
rect 20893 7534 20918 7552
rect 20607 7511 20918 7534
rect 20607 7510 20662 7511
rect 20496 7499 20500 7504
rect 20457 7496 20500 7499
rect 20390 7482 20500 7496
rect 19816 7464 20157 7465
rect 18693 7443 18696 7463
rect 18716 7443 19109 7463
rect 19741 7463 20157 7464
rect 20607 7463 20650 7510
rect 19741 7459 20650 7463
rect 17616 7408 18327 7410
rect 18866 7408 18955 7411
rect 17616 7399 18955 7408
rect 17616 7361 18878 7399
rect 18903 7364 18922 7399
rect 18947 7364 18955 7399
rect 19060 7410 19105 7443
rect 19741 7439 19744 7459
rect 19764 7439 20650 7459
rect 20118 7434 20650 7439
rect 20858 7453 20917 7475
rect 20858 7435 20877 7453
rect 20895 7435 20917 7453
rect 19906 7410 20005 7412
rect 19060 7400 20005 7410
rect 19060 7374 19928 7400
rect 19061 7373 19928 7374
rect 18903 7361 18955 7364
rect 17616 7353 18955 7361
rect 19906 7362 19928 7373
rect 19953 7365 19972 7400
rect 19997 7365 20005 7400
rect 19953 7362 20005 7365
rect 19906 7354 20005 7362
rect 20858 7361 20917 7435
rect 19932 7353 20004 7354
rect 17616 7352 18954 7353
rect 17616 7350 18327 7352
rect 18476 7311 18540 7315
rect 20851 7313 20917 7361
rect 18476 7302 18550 7311
rect 16991 6819 17105 6823
rect 16196 6815 16296 6819
rect 16196 6811 16258 6815
rect 16196 6785 16203 6811
rect 16229 6789 16258 6811
rect 16284 6789 16296 6815
rect 16229 6785 16296 6789
rect 16196 6782 16296 6785
rect 16364 6782 16399 6819
rect 16461 6816 16820 6819
rect 16461 6811 16683 6816
rect 16461 6787 16474 6811
rect 16498 6792 16683 6811
rect 16707 6792 16820 6816
rect 16498 6787 16820 6792
rect 16461 6783 16820 6787
rect 16887 6816 17105 6819
rect 16887 6815 17070 6816
rect 16887 6811 17013 6815
rect 16887 6791 16898 6811
rect 16918 6791 17013 6811
rect 17037 6792 17070 6815
rect 17094 6792 17105 6816
rect 17037 6791 17105 6792
rect 16887 6784 17105 6791
rect 16887 6783 16928 6784
rect 16363 6757 16399 6782
rect 16211 6730 16248 6731
rect 16307 6730 16344 6731
rect 16363 6730 16370 6757
rect 16111 6721 16249 6730
rect 16111 6701 16220 6721
rect 16240 6701 16249 6721
rect 16111 6694 16249 6701
rect 16307 6727 16370 6730
rect 16391 6730 16399 6757
rect 16418 6730 16455 6731
rect 16391 6727 16455 6730
rect 16307 6721 16455 6727
rect 16307 6701 16316 6721
rect 16336 6701 16426 6721
rect 16446 6701 16455 6721
rect 16111 6692 16207 6694
rect 16307 6691 16455 6701
rect 16514 6721 16551 6731
rect 16626 6730 16663 6731
rect 16607 6728 16663 6730
rect 16514 6701 16522 6721
rect 16542 6701 16551 6721
rect 16363 6690 16399 6691
rect 16211 6559 16248 6560
rect 16514 6559 16551 6701
rect 16576 6721 16663 6728
rect 16576 6718 16634 6721
rect 16576 6698 16581 6718
rect 16602 6701 16634 6718
rect 16654 6701 16663 6721
rect 16602 6698 16663 6701
rect 16576 6691 16663 6698
rect 16722 6721 16759 6731
rect 16722 6701 16730 6721
rect 16750 6701 16759 6721
rect 16576 6690 16607 6691
rect 16722 6622 16759 6701
rect 16789 6730 16820 6783
rect 16991 6781 17105 6784
rect 17034 6749 17105 6781
rect 18280 7260 18364 7285
rect 18280 7232 18295 7260
rect 18339 7232 18364 7260
rect 18280 7203 18364 7232
rect 18476 7254 18490 7302
rect 18527 7254 18550 7302
rect 18476 7226 18550 7254
rect 18280 7175 18292 7203
rect 18336 7175 18364 7203
rect 18280 7154 18364 7175
rect 16839 6730 16876 6731
rect 16789 6721 16876 6730
rect 16789 6701 16847 6721
rect 16867 6701 16876 6721
rect 16789 6691 16876 6701
rect 16935 6721 16972 6731
rect 16935 6701 16943 6721
rect 16963 6701 16972 6721
rect 16789 6690 16820 6691
rect 16784 6622 16894 6635
rect 16935 6622 16972 6701
rect 16722 6620 16972 6622
rect 16722 6617 16823 6620
rect 16722 6598 16787 6617
rect 16784 6590 16787 6598
rect 16816 6590 16823 6617
rect 16851 6593 16861 6620
rect 16890 6598 16972 6620
rect 16890 6593 16894 6598
rect 16851 6590 16894 6593
rect 16784 6576 16894 6590
rect 16210 6558 16551 6559
rect 16135 6555 16551 6558
rect 16135 6553 16558 6555
rect 16135 6533 16138 6553
rect 16158 6533 16558 6553
rect 15326 4192 15966 4280
rect 15326 3841 15410 4192
rect 15892 4161 15936 4167
rect 15892 4135 15900 4161
rect 15925 4135 15936 4161
rect 15892 4086 15936 4135
rect 15892 4066 16289 4086
rect 16309 4066 16312 4086
rect 15892 4061 16312 4066
rect 15892 4060 16237 4061
rect 15892 4056 15936 4060
rect 16199 4059 16236 4060
rect 15553 4029 15663 4043
rect 15553 4026 15596 4029
rect 15553 4021 15557 4026
rect 15475 3999 15557 4021
rect 15586 3999 15596 4026
rect 15624 4002 15631 4029
rect 15660 4021 15663 4029
rect 15660 4002 15725 4021
rect 15624 3999 15725 4002
rect 15475 3997 15725 3999
rect 15475 3918 15512 3997
rect 15553 3984 15663 3997
rect 15627 3928 15658 3929
rect 15475 3898 15484 3918
rect 15504 3898 15512 3918
rect 15475 3888 15512 3898
rect 15571 3918 15658 3928
rect 15571 3898 15580 3918
rect 15600 3898 15658 3918
rect 15571 3889 15658 3898
rect 15571 3888 15608 3889
rect 15326 3835 15435 3841
rect 15627 3836 15658 3889
rect 15688 3918 15725 3997
rect 15840 3928 15871 3929
rect 15688 3898 15697 3918
rect 15717 3898 15725 3918
rect 15688 3888 15725 3898
rect 15784 3921 15871 3928
rect 15784 3918 15845 3921
rect 15784 3898 15793 3918
rect 15813 3901 15845 3918
rect 15866 3901 15871 3921
rect 15813 3898 15871 3901
rect 15784 3891 15871 3898
rect 15896 3918 15933 4056
rect 16048 3928 16084 3929
rect 15896 3898 15905 3918
rect 15925 3898 15933 3918
rect 15784 3889 15840 3891
rect 15784 3888 15821 3889
rect 15896 3888 15933 3898
rect 15992 3918 16140 3928
rect 16240 3925 16336 3927
rect 15992 3898 16001 3918
rect 16021 3898 16111 3918
rect 16131 3898 16140 3918
rect 15992 3892 16140 3898
rect 15992 3889 16056 3892
rect 15992 3888 16029 3889
rect 16048 3862 16056 3889
rect 16077 3889 16140 3892
rect 16198 3918 16336 3925
rect 16198 3898 16207 3918
rect 16227 3898 16336 3918
rect 16198 3889 16336 3898
rect 16077 3862 16084 3889
rect 16103 3888 16140 3889
rect 16199 3888 16236 3889
rect 16048 3837 16084 3862
rect 15519 3835 15560 3836
rect 15326 3828 15560 3835
rect 15326 3808 15529 3828
rect 15549 3808 15560 3828
rect 15326 3800 15560 3808
rect 15627 3832 15986 3836
rect 15627 3827 15949 3832
rect 15627 3803 15740 3827
rect 15764 3808 15949 3827
rect 15973 3808 15986 3832
rect 15764 3803 15986 3808
rect 15627 3800 15986 3803
rect 16048 3800 16083 3837
rect 16151 3834 16251 3837
rect 16151 3830 16218 3834
rect 16151 3804 16163 3830
rect 16189 3808 16218 3830
rect 16244 3808 16251 3834
rect 16189 3804 16251 3808
rect 16151 3800 16251 3804
rect 15326 3782 15435 3800
rect 15627 3779 15658 3800
rect 16048 3779 16084 3800
rect 15470 3778 15507 3779
rect 15469 3769 15507 3778
rect 15469 3749 15478 3769
rect 15498 3749 15507 3769
rect 15469 3741 15507 3749
rect 15573 3773 15658 3779
rect 15683 3778 15720 3779
rect 15573 3753 15581 3773
rect 15601 3753 15658 3773
rect 15573 3745 15658 3753
rect 15682 3769 15720 3778
rect 15682 3749 15691 3769
rect 15711 3749 15720 3769
rect 15573 3744 15609 3745
rect 15682 3741 15720 3749
rect 15786 3773 15871 3779
rect 15891 3778 15928 3779
rect 15786 3753 15794 3773
rect 15814 3772 15871 3773
rect 15814 3753 15843 3772
rect 15786 3752 15843 3753
rect 15864 3752 15871 3772
rect 15786 3745 15871 3752
rect 15890 3769 15928 3778
rect 15890 3749 15899 3769
rect 15919 3749 15928 3769
rect 15786 3744 15822 3745
rect 15890 3741 15928 3749
rect 15994 3774 16138 3779
rect 15994 3773 16047 3774
rect 15994 3753 16002 3773
rect 16022 3754 16047 3773
rect 16080 3773 16138 3774
rect 16080 3754 16110 3773
rect 16022 3753 16110 3754
rect 16130 3753 16138 3773
rect 15994 3745 16138 3753
rect 15994 3744 16030 3745
rect 16102 3744 16138 3745
rect 16204 3778 16241 3779
rect 16204 3777 16242 3778
rect 16204 3769 16268 3777
rect 16204 3749 16213 3769
rect 16233 3755 16268 3769
rect 16288 3755 16291 3775
rect 16233 3750 16291 3755
rect 16233 3749 16268 3750
rect 15470 3712 15507 3741
rect 15471 3710 15507 3712
rect 15683 3710 15720 3741
rect 15471 3688 15720 3710
rect 15552 3682 15663 3688
rect 15552 3674 15593 3682
rect 15552 3654 15560 3674
rect 15579 3654 15593 3674
rect 15552 3652 15593 3654
rect 15621 3674 15663 3682
rect 15621 3654 15637 3674
rect 15656 3654 15663 3674
rect 15621 3652 15663 3654
rect 15552 3637 15663 3652
rect 15891 3620 15928 3741
rect 16204 3737 16268 3749
rect 16308 3626 16335 3889
rect 16362 3635 16398 3642
rect 16362 3626 16368 3635
rect 16286 3622 16368 3626
rect 16167 3620 16368 3622
rect 15891 3597 16368 3620
rect 16391 3597 16398 3635
rect 15891 3594 16398 3597
rect 16167 3593 16335 3594
rect 16362 3591 16398 3594
rect 16480 3493 16558 6533
rect 17614 5786 17673 5796
rect 17614 5758 17627 5786
rect 17655 5758 17673 5786
rect 17614 5709 17673 5758
rect 17220 5574 17388 5575
rect 17624 5574 17671 5709
rect 17220 5548 17671 5574
rect 17220 5546 17388 5548
rect 17220 5279 17247 5546
rect 17624 5542 17671 5548
rect 17287 5419 17351 5431
rect 17627 5427 17664 5542
rect 17892 5516 18003 5531
rect 17892 5514 17934 5516
rect 17892 5494 17899 5514
rect 17918 5494 17934 5514
rect 17892 5486 17934 5494
rect 17962 5514 18003 5516
rect 17962 5494 17976 5514
rect 17995 5494 18003 5514
rect 17962 5486 18003 5494
rect 17892 5480 18003 5486
rect 17835 5458 18084 5480
rect 17835 5427 17872 5458
rect 18048 5456 18084 5458
rect 18048 5427 18085 5456
rect 17287 5418 17322 5419
rect 17264 5413 17322 5418
rect 17264 5393 17267 5413
rect 17287 5399 17322 5413
rect 17342 5399 17351 5419
rect 17287 5391 17351 5399
rect 17313 5390 17351 5391
rect 17314 5389 17351 5390
rect 17417 5423 17453 5424
rect 17525 5423 17561 5424
rect 17417 5415 17561 5423
rect 17417 5395 17425 5415
rect 17445 5395 17533 5415
rect 17553 5395 17561 5415
rect 17417 5389 17561 5395
rect 17627 5419 17665 5427
rect 17733 5423 17769 5424
rect 17627 5399 17636 5419
rect 17656 5399 17665 5419
rect 17627 5390 17665 5399
rect 17684 5416 17769 5423
rect 17684 5396 17691 5416
rect 17712 5415 17769 5416
rect 17712 5396 17741 5415
rect 17684 5395 17741 5396
rect 17761 5395 17769 5415
rect 17627 5389 17664 5390
rect 17684 5389 17769 5395
rect 17835 5419 17873 5427
rect 17946 5423 17982 5424
rect 17835 5399 17844 5419
rect 17864 5399 17873 5419
rect 17835 5390 17873 5399
rect 17897 5415 17982 5423
rect 17897 5395 17954 5415
rect 17974 5395 17982 5415
rect 17835 5389 17872 5390
rect 17897 5389 17982 5395
rect 18048 5419 18086 5427
rect 18048 5399 18057 5419
rect 18077 5399 18086 5419
rect 18048 5390 18086 5399
rect 18048 5389 18085 5390
rect 17471 5368 17507 5389
rect 17897 5368 17928 5389
rect 18108 5374 18165 5382
rect 18108 5368 18116 5374
rect 17304 5364 17404 5368
rect 17304 5360 17366 5364
rect 17304 5334 17311 5360
rect 17337 5338 17366 5360
rect 17392 5338 17404 5364
rect 17337 5334 17404 5338
rect 17304 5331 17404 5334
rect 17472 5331 17507 5368
rect 17569 5365 17928 5368
rect 17569 5360 17791 5365
rect 17569 5336 17582 5360
rect 17606 5341 17791 5360
rect 17815 5341 17928 5365
rect 17606 5336 17928 5341
rect 17569 5332 17928 5336
rect 17995 5360 18116 5368
rect 17995 5340 18006 5360
rect 18026 5351 18116 5360
rect 18142 5351 18165 5374
rect 18026 5340 18165 5351
rect 17995 5338 18165 5340
rect 17995 5333 18116 5338
rect 17995 5332 18036 5333
rect 17471 5306 17507 5331
rect 17319 5279 17356 5280
rect 17415 5279 17452 5280
rect 17471 5279 17478 5306
rect 17219 5270 17357 5279
rect 17219 5250 17328 5270
rect 17348 5250 17357 5270
rect 17219 5243 17357 5250
rect 17415 5276 17478 5279
rect 17499 5279 17507 5306
rect 17526 5279 17563 5280
rect 17499 5276 17563 5279
rect 17415 5270 17563 5276
rect 17415 5250 17424 5270
rect 17444 5250 17534 5270
rect 17554 5250 17563 5270
rect 17219 5241 17315 5243
rect 17415 5240 17563 5250
rect 17622 5270 17659 5280
rect 17734 5279 17771 5280
rect 17715 5277 17771 5279
rect 17622 5250 17630 5270
rect 17650 5250 17659 5270
rect 17471 5239 17507 5240
rect 17319 5108 17356 5109
rect 17622 5108 17659 5250
rect 17684 5270 17771 5277
rect 17684 5267 17742 5270
rect 17684 5247 17689 5267
rect 17710 5250 17742 5267
rect 17762 5250 17771 5270
rect 17710 5247 17771 5250
rect 17684 5240 17771 5247
rect 17830 5270 17867 5280
rect 17830 5250 17838 5270
rect 17858 5250 17867 5270
rect 17684 5239 17715 5240
rect 17830 5171 17867 5250
rect 17897 5279 17928 5332
rect 17947 5279 17984 5280
rect 17897 5270 17984 5279
rect 17897 5250 17955 5270
rect 17975 5250 17984 5270
rect 17897 5240 17984 5250
rect 18043 5270 18080 5280
rect 18043 5250 18051 5270
rect 18071 5250 18080 5270
rect 17897 5239 17928 5240
rect 17892 5171 18002 5184
rect 18043 5171 18080 5250
rect 17830 5169 18080 5171
rect 17830 5166 17931 5169
rect 17830 5147 17895 5166
rect 17892 5139 17895 5147
rect 17924 5139 17931 5166
rect 17959 5142 17969 5169
rect 17998 5147 18080 5169
rect 17998 5142 18002 5147
rect 17959 5139 18002 5142
rect 17892 5125 18002 5139
rect 17318 5107 17659 5108
rect 17243 5102 17659 5107
rect 17243 5082 17246 5102
rect 17266 5082 17660 5102
rect 17469 5049 17506 5059
rect 17469 5012 17478 5049
rect 17495 5012 17506 5049
rect 17469 4991 17506 5012
rect 17178 4052 17346 4053
rect 17475 4052 17504 4991
rect 17617 4377 17660 5082
rect 17618 4369 17660 4377
rect 17618 4358 17663 4369
rect 17618 4320 17628 4358
rect 17653 4320 17663 4358
rect 17618 4311 17663 4320
rect 17178 4026 17622 4052
rect 17178 4024 17346 4026
rect 17178 3757 17205 4024
rect 17475 4022 17504 4026
rect 17245 3897 17309 3909
rect 17585 3905 17622 4026
rect 17850 3994 17961 4009
rect 17850 3992 17892 3994
rect 17850 3972 17857 3992
rect 17876 3972 17892 3992
rect 17850 3964 17892 3972
rect 17920 3992 17961 3994
rect 17920 3972 17934 3992
rect 17953 3972 17961 3992
rect 17920 3964 17961 3972
rect 17850 3958 17961 3964
rect 17793 3936 18042 3958
rect 17793 3905 17830 3936
rect 18006 3934 18042 3936
rect 18006 3905 18043 3934
rect 17245 3896 17280 3897
rect 17222 3891 17280 3896
rect 17222 3871 17225 3891
rect 17245 3877 17280 3891
rect 17300 3877 17309 3897
rect 17245 3869 17309 3877
rect 17271 3868 17309 3869
rect 17272 3867 17309 3868
rect 17375 3901 17411 3902
rect 17483 3901 17519 3902
rect 17375 3893 17519 3901
rect 17375 3873 17383 3893
rect 17403 3873 17491 3893
rect 17511 3873 17519 3893
rect 17375 3867 17519 3873
rect 17585 3897 17623 3905
rect 17691 3901 17727 3902
rect 17585 3877 17594 3897
rect 17614 3877 17623 3897
rect 17585 3868 17623 3877
rect 17642 3894 17727 3901
rect 17642 3874 17649 3894
rect 17670 3893 17727 3894
rect 17670 3874 17699 3893
rect 17642 3873 17699 3874
rect 17719 3873 17727 3893
rect 17585 3867 17622 3868
rect 17642 3867 17727 3873
rect 17793 3897 17831 3905
rect 17904 3901 17940 3902
rect 17793 3877 17802 3897
rect 17822 3877 17831 3897
rect 17793 3868 17831 3877
rect 17855 3893 17940 3901
rect 17855 3873 17912 3893
rect 17932 3873 17940 3893
rect 17793 3867 17830 3868
rect 17855 3867 17940 3873
rect 18006 3897 18044 3905
rect 18006 3877 18015 3897
rect 18035 3877 18044 3897
rect 18006 3868 18044 3877
rect 18006 3867 18043 3868
rect 17429 3846 17465 3867
rect 17855 3846 17886 3867
rect 18280 3850 18372 7154
rect 18478 5387 18550 7226
rect 19580 7176 19652 7193
rect 19580 7128 19592 7176
rect 19638 7128 19652 7176
rect 20120 7156 20161 7158
rect 20392 7156 20496 7158
rect 20851 7156 20916 7313
rect 19580 7106 19652 7128
rect 19713 7121 20916 7156
rect 19713 7107 19741 7121
rect 19581 6906 19651 7106
rect 19715 6976 19741 7107
rect 20120 7118 20916 7121
rect 19573 6855 19653 6906
rect 19573 6829 19589 6855
rect 19629 6829 19653 6855
rect 19573 6810 19653 6829
rect 19573 6784 19592 6810
rect 19632 6784 19653 6810
rect 19573 6757 19653 6784
rect 19573 6731 19596 6757
rect 19636 6731 19653 6757
rect 19573 6720 19653 6731
rect 19715 6721 19742 6976
rect 20120 6968 20161 7118
rect 20392 7116 20496 7118
rect 20851 7084 20916 7118
rect 20587 7056 20708 7074
rect 20587 7054 20658 7056
rect 20587 7013 20602 7054
rect 20639 7015 20658 7054
rect 20695 7015 20708 7056
rect 20639 7013 20708 7015
rect 20587 7003 20708 7013
rect 20392 6973 20496 6976
rect 19782 6861 19846 6873
rect 20122 6869 20159 6968
rect 20387 6958 20498 6973
rect 20387 6956 20429 6958
rect 20387 6936 20394 6956
rect 20413 6936 20429 6956
rect 20387 6928 20429 6936
rect 20457 6956 20498 6958
rect 20457 6936 20471 6956
rect 20490 6936 20498 6956
rect 20457 6928 20498 6936
rect 20387 6922 20498 6928
rect 20330 6900 20579 6922
rect 20330 6869 20367 6900
rect 20543 6898 20579 6900
rect 20543 6869 20580 6898
rect 19782 6860 19817 6861
rect 19759 6855 19817 6860
rect 19759 6835 19762 6855
rect 19782 6841 19817 6855
rect 19837 6841 19846 6861
rect 19782 6833 19846 6841
rect 19808 6832 19846 6833
rect 19809 6831 19846 6832
rect 19912 6865 19948 6866
rect 20020 6865 20056 6866
rect 19912 6857 20056 6865
rect 19912 6837 19920 6857
rect 19940 6837 20028 6857
rect 20048 6837 20056 6857
rect 19912 6831 20056 6837
rect 20122 6861 20160 6869
rect 20228 6865 20264 6866
rect 20122 6841 20131 6861
rect 20151 6841 20160 6861
rect 20122 6832 20160 6841
rect 20179 6858 20264 6865
rect 20179 6838 20186 6858
rect 20207 6857 20264 6858
rect 20207 6838 20236 6857
rect 20179 6837 20236 6838
rect 20256 6837 20264 6857
rect 20122 6831 20159 6832
rect 20179 6831 20264 6837
rect 20330 6861 20368 6869
rect 20441 6865 20477 6866
rect 20330 6841 20339 6861
rect 20359 6841 20368 6861
rect 20330 6832 20368 6841
rect 20392 6857 20477 6865
rect 20392 6837 20449 6857
rect 20469 6837 20477 6857
rect 20330 6831 20367 6832
rect 20392 6831 20477 6837
rect 20543 6861 20581 6869
rect 20543 6841 20552 6861
rect 20572 6841 20581 6861
rect 20636 6851 20701 7003
rect 20854 6977 20909 7084
rect 20543 6832 20581 6841
rect 20634 6844 20701 6851
rect 20543 6831 20580 6832
rect 19966 6810 20002 6831
rect 20392 6810 20423 6831
rect 20634 6823 20651 6844
rect 20687 6823 20701 6844
rect 20853 6864 20909 6977
rect 20853 6846 20872 6864
rect 20890 6846 20909 6864
rect 20853 6826 20909 6846
rect 20634 6810 20701 6823
rect 19799 6806 19899 6810
rect 19799 6802 19861 6806
rect 19799 6776 19806 6802
rect 19832 6780 19861 6802
rect 19887 6780 19899 6806
rect 19832 6776 19899 6780
rect 19799 6773 19899 6776
rect 19967 6773 20002 6810
rect 20064 6807 20423 6810
rect 20064 6802 20286 6807
rect 20064 6778 20077 6802
rect 20101 6783 20286 6802
rect 20310 6783 20423 6807
rect 20101 6778 20423 6783
rect 20064 6774 20423 6778
rect 20490 6804 20701 6810
rect 20490 6802 20651 6804
rect 20490 6782 20501 6802
rect 20521 6782 20651 6802
rect 20490 6775 20651 6782
rect 20490 6774 20531 6775
rect 19966 6748 20002 6773
rect 19814 6721 19851 6722
rect 19910 6721 19947 6722
rect 19966 6721 19973 6748
rect 19714 6712 19852 6721
rect 19714 6692 19823 6712
rect 19843 6692 19852 6712
rect 19714 6685 19852 6692
rect 19910 6718 19973 6721
rect 19994 6721 20002 6748
rect 20021 6721 20058 6722
rect 19994 6718 20058 6721
rect 19910 6712 20058 6718
rect 19910 6692 19919 6712
rect 19939 6692 20029 6712
rect 20049 6692 20058 6712
rect 19714 6683 19810 6685
rect 19910 6682 20058 6692
rect 20117 6712 20154 6722
rect 20229 6721 20266 6722
rect 20210 6719 20266 6721
rect 20117 6692 20125 6712
rect 20145 6692 20154 6712
rect 19966 6681 20002 6682
rect 19814 6550 19851 6551
rect 20117 6550 20154 6692
rect 20179 6712 20266 6719
rect 20179 6709 20237 6712
rect 20179 6689 20184 6709
rect 20205 6692 20237 6709
rect 20257 6692 20266 6712
rect 20205 6689 20266 6692
rect 20179 6682 20266 6689
rect 20325 6712 20362 6722
rect 20325 6692 20333 6712
rect 20353 6692 20362 6712
rect 20179 6681 20210 6682
rect 20325 6613 20362 6692
rect 20392 6721 20423 6774
rect 20636 6767 20651 6775
rect 20691 6767 20701 6804
rect 20636 6758 20701 6767
rect 20849 6765 20914 6786
rect 20849 6747 20874 6765
rect 20892 6747 20914 6765
rect 20442 6721 20479 6722
rect 20392 6712 20479 6721
rect 20392 6692 20450 6712
rect 20470 6692 20479 6712
rect 20392 6682 20479 6692
rect 20538 6712 20575 6722
rect 20538 6692 20546 6712
rect 20566 6692 20575 6712
rect 20392 6681 20423 6682
rect 20387 6613 20497 6626
rect 20538 6613 20575 6692
rect 20849 6671 20914 6747
rect 20325 6611 20575 6613
rect 20325 6608 20426 6611
rect 20325 6589 20390 6608
rect 20387 6581 20390 6589
rect 20419 6581 20426 6608
rect 20454 6584 20464 6611
rect 20493 6589 20575 6611
rect 20598 6636 20915 6671
rect 20493 6584 20497 6589
rect 20454 6581 20497 6584
rect 20387 6567 20497 6581
rect 19813 6549 20154 6550
rect 19738 6547 20154 6549
rect 20598 6547 20638 6636
rect 20849 6609 20914 6636
rect 20849 6591 20872 6609
rect 20890 6591 20914 6609
rect 20849 6571 20914 6591
rect 19735 6544 20638 6547
rect 19735 6524 19741 6544
rect 19761 6524 20638 6544
rect 19735 6520 20638 6524
rect 20598 6517 20638 6520
rect 20850 6510 20915 6531
rect 19068 6502 19729 6503
rect 19068 6495 20002 6502
rect 19068 6494 19974 6495
rect 19068 6474 19919 6494
rect 19951 6475 19974 6494
rect 19999 6475 20002 6495
rect 19951 6474 20002 6475
rect 19068 6467 20002 6474
rect 18667 6425 18835 6426
rect 19070 6425 19109 6467
rect 19898 6465 20002 6467
rect 19967 6463 20002 6465
rect 20850 6492 20874 6510
rect 20892 6492 20915 6510
rect 20850 6445 20915 6492
rect 18667 6399 19111 6425
rect 18667 6397 18835 6399
rect 18667 6046 18694 6397
rect 19070 6393 19111 6399
rect 18734 6186 18798 6198
rect 19074 6194 19111 6393
rect 19573 6420 19645 6437
rect 19573 6381 19581 6420
rect 19626 6381 19645 6420
rect 19339 6283 19450 6298
rect 19339 6281 19381 6283
rect 19339 6261 19346 6281
rect 19365 6261 19381 6281
rect 19339 6253 19381 6261
rect 19409 6281 19450 6283
rect 19409 6261 19423 6281
rect 19442 6261 19450 6281
rect 19409 6253 19450 6261
rect 19339 6247 19450 6253
rect 19282 6225 19531 6247
rect 19282 6194 19319 6225
rect 19495 6223 19531 6225
rect 19495 6194 19532 6223
rect 18734 6185 18769 6186
rect 18711 6180 18769 6185
rect 18711 6160 18714 6180
rect 18734 6166 18769 6180
rect 18789 6166 18798 6186
rect 18734 6158 18798 6166
rect 18760 6157 18798 6158
rect 18761 6156 18798 6157
rect 18864 6190 18900 6191
rect 18972 6190 19008 6191
rect 18864 6182 19008 6190
rect 18864 6162 18872 6182
rect 18892 6162 18980 6182
rect 19000 6162 19008 6182
rect 18864 6156 19008 6162
rect 19074 6186 19112 6194
rect 19180 6190 19216 6191
rect 19074 6166 19083 6186
rect 19103 6166 19112 6186
rect 19074 6157 19112 6166
rect 19131 6183 19216 6190
rect 19131 6163 19138 6183
rect 19159 6182 19216 6183
rect 19159 6163 19188 6182
rect 19131 6162 19188 6163
rect 19208 6162 19216 6182
rect 19074 6156 19111 6157
rect 19131 6156 19216 6162
rect 19282 6186 19320 6194
rect 19393 6190 19429 6191
rect 19282 6166 19291 6186
rect 19311 6166 19320 6186
rect 19282 6157 19320 6166
rect 19344 6182 19429 6190
rect 19344 6162 19401 6182
rect 19421 6162 19429 6182
rect 19282 6156 19319 6157
rect 19344 6156 19429 6162
rect 19495 6186 19533 6194
rect 19495 6166 19504 6186
rect 19524 6166 19533 6186
rect 19495 6157 19533 6166
rect 19573 6171 19645 6381
rect 19715 6415 20915 6445
rect 19715 6414 20159 6415
rect 19715 6412 19883 6414
rect 19573 6157 19656 6171
rect 19495 6156 19532 6157
rect 18918 6135 18954 6156
rect 19344 6135 19375 6156
rect 19573 6135 19590 6157
rect 18751 6131 18851 6135
rect 18751 6127 18813 6131
rect 18751 6101 18758 6127
rect 18784 6105 18813 6127
rect 18839 6105 18851 6131
rect 18784 6101 18851 6105
rect 18751 6098 18851 6101
rect 18919 6098 18954 6135
rect 19016 6132 19375 6135
rect 19016 6127 19238 6132
rect 19016 6103 19029 6127
rect 19053 6108 19238 6127
rect 19262 6108 19375 6132
rect 19053 6103 19375 6108
rect 19016 6099 19375 6103
rect 19442 6127 19590 6135
rect 19442 6107 19453 6127
rect 19473 6124 19590 6127
rect 19643 6124 19656 6157
rect 19473 6107 19656 6124
rect 19442 6100 19656 6107
rect 19442 6099 19483 6100
rect 19573 6099 19656 6100
rect 18918 6073 18954 6098
rect 18766 6046 18803 6047
rect 18862 6046 18899 6047
rect 18918 6046 18925 6073
rect 18666 6037 18804 6046
rect 18666 6017 18775 6037
rect 18795 6017 18804 6037
rect 18666 6010 18804 6017
rect 18862 6043 18925 6046
rect 18946 6046 18954 6073
rect 18973 6046 19010 6047
rect 18946 6043 19010 6046
rect 18862 6037 19010 6043
rect 18862 6017 18871 6037
rect 18891 6017 18981 6037
rect 19001 6017 19010 6037
rect 18666 6008 18762 6010
rect 18862 6007 19010 6017
rect 19069 6037 19106 6047
rect 19181 6046 19218 6047
rect 19162 6044 19218 6046
rect 19069 6017 19077 6037
rect 19097 6017 19106 6037
rect 18918 6006 18954 6007
rect 18766 5875 18803 5876
rect 19069 5875 19106 6017
rect 19131 6037 19218 6044
rect 19131 6034 19189 6037
rect 19131 6014 19136 6034
rect 19157 6017 19189 6034
rect 19209 6017 19218 6037
rect 19157 6014 19218 6017
rect 19131 6007 19218 6014
rect 19277 6037 19314 6047
rect 19277 6017 19285 6037
rect 19305 6017 19314 6037
rect 19131 6006 19162 6007
rect 19277 5938 19314 6017
rect 19344 6046 19375 6099
rect 19581 6066 19595 6099
rect 19648 6066 19656 6099
rect 19581 6060 19656 6066
rect 19581 6055 19651 6060
rect 19394 6046 19431 6047
rect 19344 6037 19431 6046
rect 19344 6017 19402 6037
rect 19422 6017 19431 6037
rect 19344 6007 19431 6017
rect 19490 6037 19527 6047
rect 19715 6042 19742 6412
rect 19782 6182 19846 6194
rect 20122 6190 20159 6414
rect 20630 6395 20694 6397
rect 20626 6383 20694 6395
rect 20626 6350 20637 6383
rect 20677 6350 20694 6383
rect 20626 6340 20694 6350
rect 20387 6279 20498 6294
rect 20387 6277 20429 6279
rect 20387 6257 20394 6277
rect 20413 6257 20429 6277
rect 20387 6249 20429 6257
rect 20457 6277 20498 6279
rect 20457 6257 20471 6277
rect 20490 6257 20498 6277
rect 20457 6249 20498 6257
rect 20387 6243 20498 6249
rect 20330 6221 20579 6243
rect 20330 6190 20367 6221
rect 20543 6219 20579 6221
rect 20543 6190 20580 6219
rect 19782 6181 19817 6182
rect 19759 6176 19817 6181
rect 19759 6156 19762 6176
rect 19782 6162 19817 6176
rect 19837 6162 19846 6182
rect 19782 6154 19846 6162
rect 19808 6153 19846 6154
rect 19809 6152 19846 6153
rect 19912 6186 19948 6187
rect 20020 6186 20056 6187
rect 19912 6178 20056 6186
rect 19912 6158 19920 6178
rect 19940 6158 20028 6178
rect 20048 6158 20056 6178
rect 19912 6152 20056 6158
rect 20122 6182 20160 6190
rect 20228 6186 20264 6187
rect 20122 6162 20131 6182
rect 20151 6162 20160 6182
rect 20122 6153 20160 6162
rect 20179 6179 20264 6186
rect 20179 6159 20186 6179
rect 20207 6178 20264 6179
rect 20207 6159 20236 6178
rect 20179 6158 20236 6159
rect 20256 6158 20264 6178
rect 20122 6152 20159 6153
rect 20179 6152 20264 6158
rect 20330 6182 20368 6190
rect 20441 6186 20477 6187
rect 20330 6162 20339 6182
rect 20359 6162 20368 6182
rect 20330 6153 20368 6162
rect 20392 6178 20477 6186
rect 20392 6158 20449 6178
rect 20469 6158 20477 6178
rect 20330 6152 20367 6153
rect 20392 6152 20477 6158
rect 20543 6182 20581 6190
rect 20543 6162 20552 6182
rect 20572 6162 20581 6182
rect 20543 6153 20581 6162
rect 20630 6156 20694 6340
rect 20850 6214 20915 6415
rect 20850 6196 20872 6214
rect 20890 6196 20915 6214
rect 20850 6177 20915 6196
rect 20543 6152 20580 6153
rect 19966 6131 20002 6152
rect 20392 6131 20423 6152
rect 20630 6147 20638 6156
rect 20627 6131 20638 6147
rect 19799 6127 19899 6131
rect 19799 6123 19861 6127
rect 19799 6097 19806 6123
rect 19832 6101 19861 6123
rect 19887 6101 19899 6127
rect 19832 6097 19899 6101
rect 19799 6094 19899 6097
rect 19967 6094 20002 6131
rect 20064 6128 20423 6131
rect 20064 6123 20286 6128
rect 20064 6099 20077 6123
rect 20101 6104 20286 6123
rect 20310 6104 20423 6128
rect 20101 6099 20423 6104
rect 20064 6095 20423 6099
rect 20490 6123 20638 6131
rect 20490 6103 20501 6123
rect 20521 6114 20638 6123
rect 20687 6147 20694 6156
rect 20687 6114 20695 6147
rect 20521 6103 20695 6114
rect 20490 6096 20695 6103
rect 20490 6095 20531 6096
rect 19966 6069 20002 6094
rect 19814 6042 19851 6043
rect 19910 6042 19947 6043
rect 19966 6042 19973 6069
rect 19490 6017 19498 6037
rect 19518 6017 19527 6037
rect 19344 6006 19375 6007
rect 19339 5938 19449 5951
rect 19490 5938 19527 6017
rect 19714 6033 19852 6042
rect 19714 6013 19823 6033
rect 19843 6013 19852 6033
rect 19714 6006 19852 6013
rect 19910 6039 19973 6042
rect 19994 6042 20002 6069
rect 20021 6042 20058 6043
rect 19994 6039 20058 6042
rect 19910 6033 20058 6039
rect 19910 6013 19919 6033
rect 19939 6013 20029 6033
rect 20049 6013 20058 6033
rect 19714 6004 19810 6006
rect 19910 6003 20058 6013
rect 20117 6033 20154 6043
rect 20229 6042 20266 6043
rect 20210 6040 20266 6042
rect 20117 6013 20125 6033
rect 20145 6013 20154 6033
rect 19966 6002 20002 6003
rect 19277 5936 19527 5938
rect 19277 5933 19378 5936
rect 19277 5914 19342 5933
rect 19339 5906 19342 5914
rect 19371 5906 19378 5933
rect 19406 5909 19416 5936
rect 19445 5914 19527 5936
rect 19445 5909 19449 5914
rect 19406 5906 19449 5909
rect 19339 5892 19449 5906
rect 18765 5874 19106 5875
rect 18690 5869 19106 5874
rect 19814 5871 19851 5872
rect 20117 5871 20154 6013
rect 20179 6033 20266 6040
rect 20179 6030 20237 6033
rect 20179 6010 20184 6030
rect 20205 6013 20237 6030
rect 20257 6013 20266 6033
rect 20205 6010 20266 6013
rect 20179 6003 20266 6010
rect 20325 6033 20362 6043
rect 20325 6013 20333 6033
rect 20353 6013 20362 6033
rect 20179 6002 20210 6003
rect 20325 5934 20362 6013
rect 20392 6042 20423 6095
rect 20627 6093 20695 6096
rect 20627 6051 20639 6093
rect 20688 6051 20695 6093
rect 20442 6042 20479 6043
rect 20392 6033 20479 6042
rect 20392 6013 20450 6033
rect 20470 6013 20479 6033
rect 20392 6003 20479 6013
rect 20538 6033 20575 6043
rect 20627 6038 20695 6051
rect 20850 6115 20915 6132
rect 20850 6097 20874 6115
rect 20892 6097 20915 6115
rect 20538 6013 20546 6033
rect 20566 6013 20575 6033
rect 20392 6002 20423 6003
rect 20387 5934 20497 5947
rect 20538 5934 20575 6013
rect 20850 5958 20915 6097
rect 20850 5952 20872 5958
rect 20325 5932 20575 5934
rect 20325 5929 20426 5932
rect 20325 5910 20390 5929
rect 20387 5902 20390 5910
rect 20419 5902 20426 5929
rect 20454 5905 20464 5932
rect 20493 5910 20575 5932
rect 20604 5940 20872 5952
rect 20890 5940 20915 5958
rect 20604 5917 20915 5940
rect 20604 5916 20659 5917
rect 20493 5905 20497 5910
rect 20454 5902 20497 5905
rect 20387 5888 20497 5902
rect 19813 5870 20154 5871
rect 18690 5849 18693 5869
rect 18713 5849 19106 5869
rect 19738 5869 20154 5870
rect 20604 5869 20647 5916
rect 19738 5865 20647 5869
rect 19057 5816 19102 5849
rect 19738 5845 19741 5865
rect 19761 5845 20647 5865
rect 20115 5840 20647 5845
rect 20855 5859 20914 5881
rect 20855 5841 20874 5859
rect 20892 5841 20914 5859
rect 19903 5816 20002 5818
rect 19057 5806 20002 5816
rect 19057 5780 19925 5806
rect 19058 5779 19925 5780
rect 19903 5768 19925 5779
rect 19950 5771 19969 5806
rect 19994 5771 20002 5806
rect 19950 5768 20002 5771
rect 20855 5770 20914 5841
rect 19903 5760 20002 5768
rect 19929 5759 20001 5760
rect 19583 5733 19650 5752
rect 19583 5712 19600 5733
rect 19581 5667 19600 5712
rect 19630 5712 19650 5733
rect 19630 5667 19651 5712
rect 20120 5709 20161 5711
rect 20392 5709 20496 5711
rect 20852 5709 20916 5770
rect 19581 5459 19651 5667
rect 19713 5674 20916 5709
rect 19713 5660 19741 5674
rect 19715 5529 19741 5660
rect 20120 5671 20916 5674
rect 18468 5367 18550 5387
rect 18468 5344 18496 5367
rect 18522 5344 18550 5367
rect 18468 5282 18550 5344
rect 18472 5247 18550 5282
rect 19573 5408 19653 5459
rect 19573 5382 19589 5408
rect 19629 5382 19653 5408
rect 19573 5363 19653 5382
rect 19573 5337 19592 5363
rect 19632 5337 19653 5363
rect 19573 5310 19653 5337
rect 19573 5284 19596 5310
rect 19636 5284 19653 5310
rect 19573 5273 19653 5284
rect 19715 5274 19742 5529
rect 20120 5521 20161 5671
rect 20392 5665 20496 5671
rect 20852 5668 20916 5671
rect 20587 5609 20708 5627
rect 20587 5607 20658 5609
rect 20587 5566 20602 5607
rect 20639 5568 20658 5607
rect 20695 5568 20708 5609
rect 20639 5566 20708 5568
rect 20587 5556 20708 5566
rect 19782 5414 19846 5426
rect 20122 5422 20159 5521
rect 20387 5511 20498 5524
rect 20387 5509 20429 5511
rect 20387 5489 20394 5509
rect 20413 5489 20429 5509
rect 20387 5481 20429 5489
rect 20457 5509 20498 5511
rect 20457 5489 20471 5509
rect 20490 5489 20498 5509
rect 20457 5481 20498 5489
rect 20387 5475 20498 5481
rect 20330 5453 20579 5475
rect 20330 5422 20367 5453
rect 20543 5451 20579 5453
rect 20543 5422 20580 5451
rect 19782 5413 19817 5414
rect 19759 5408 19817 5413
rect 19759 5388 19762 5408
rect 19782 5394 19817 5408
rect 19837 5394 19846 5414
rect 19782 5386 19846 5394
rect 19808 5385 19846 5386
rect 19809 5384 19846 5385
rect 19912 5418 19948 5419
rect 20020 5418 20056 5419
rect 19912 5410 20056 5418
rect 19912 5390 19920 5410
rect 19940 5390 20028 5410
rect 20048 5390 20056 5410
rect 19912 5384 20056 5390
rect 20122 5414 20160 5422
rect 20228 5418 20264 5419
rect 20122 5394 20131 5414
rect 20151 5394 20160 5414
rect 20122 5385 20160 5394
rect 20179 5411 20264 5418
rect 20179 5391 20186 5411
rect 20207 5410 20264 5411
rect 20207 5391 20236 5410
rect 20179 5390 20236 5391
rect 20256 5390 20264 5410
rect 20122 5384 20159 5385
rect 20179 5384 20264 5390
rect 20330 5414 20368 5422
rect 20441 5418 20477 5419
rect 20330 5394 20339 5414
rect 20359 5394 20368 5414
rect 20330 5385 20368 5394
rect 20392 5410 20477 5418
rect 20392 5390 20449 5410
rect 20469 5390 20477 5410
rect 20330 5384 20367 5385
rect 20392 5384 20477 5390
rect 20543 5414 20581 5422
rect 20543 5394 20552 5414
rect 20572 5394 20581 5414
rect 20636 5404 20701 5556
rect 20854 5530 20909 5668
rect 20543 5385 20581 5394
rect 20634 5397 20701 5404
rect 20543 5384 20580 5385
rect 19966 5363 20002 5384
rect 20392 5363 20423 5384
rect 20634 5376 20651 5397
rect 20687 5376 20701 5397
rect 20853 5417 20909 5530
rect 20853 5399 20872 5417
rect 20890 5399 20909 5417
rect 20853 5379 20909 5399
rect 20634 5363 20701 5376
rect 19799 5359 19899 5363
rect 19799 5355 19861 5359
rect 19799 5329 19806 5355
rect 19832 5333 19861 5355
rect 19887 5333 19899 5359
rect 19832 5329 19899 5333
rect 19799 5326 19899 5329
rect 19967 5326 20002 5363
rect 20064 5360 20423 5363
rect 20064 5355 20286 5360
rect 20064 5331 20077 5355
rect 20101 5336 20286 5355
rect 20310 5336 20423 5360
rect 20101 5331 20423 5336
rect 20064 5327 20423 5331
rect 20490 5357 20701 5363
rect 20490 5355 20651 5357
rect 20490 5335 20501 5355
rect 20521 5335 20651 5355
rect 20490 5328 20651 5335
rect 20490 5327 20531 5328
rect 19966 5301 20002 5326
rect 19814 5274 19851 5275
rect 19910 5274 19947 5275
rect 19966 5274 19973 5301
rect 19714 5265 19852 5274
rect 18472 4731 18534 5247
rect 19714 5245 19823 5265
rect 19843 5245 19852 5265
rect 19714 5238 19852 5245
rect 19910 5271 19973 5274
rect 19994 5274 20002 5301
rect 20021 5274 20058 5275
rect 19994 5271 20058 5274
rect 19910 5265 20058 5271
rect 19910 5245 19919 5265
rect 19939 5245 20029 5265
rect 20049 5245 20058 5265
rect 19714 5236 19810 5238
rect 19910 5235 20058 5245
rect 20117 5265 20154 5275
rect 20229 5274 20266 5275
rect 20210 5272 20266 5274
rect 20117 5245 20125 5265
rect 20145 5245 20154 5265
rect 19966 5234 20002 5235
rect 19814 5103 19851 5104
rect 20117 5103 20154 5245
rect 20179 5265 20266 5272
rect 20179 5262 20237 5265
rect 20179 5242 20184 5262
rect 20205 5245 20237 5262
rect 20257 5245 20266 5265
rect 20205 5242 20266 5245
rect 20179 5235 20266 5242
rect 20325 5265 20362 5275
rect 20325 5245 20333 5265
rect 20353 5245 20362 5265
rect 20179 5234 20210 5235
rect 20325 5166 20362 5245
rect 20392 5274 20423 5327
rect 20636 5320 20651 5328
rect 20691 5320 20701 5357
rect 20636 5311 20701 5320
rect 20849 5318 20914 5339
rect 20849 5300 20874 5318
rect 20892 5300 20914 5318
rect 20442 5274 20479 5275
rect 20392 5265 20479 5274
rect 20392 5245 20450 5265
rect 20470 5245 20479 5265
rect 20392 5235 20479 5245
rect 20538 5265 20575 5275
rect 20538 5245 20546 5265
rect 20566 5245 20575 5265
rect 20392 5234 20423 5235
rect 20387 5166 20497 5179
rect 20538 5166 20575 5245
rect 20849 5224 20914 5300
rect 20325 5164 20575 5166
rect 20325 5161 20426 5164
rect 20325 5142 20390 5161
rect 20387 5134 20390 5142
rect 20419 5134 20426 5161
rect 20454 5137 20464 5164
rect 20493 5142 20575 5164
rect 20598 5189 20915 5224
rect 20493 5137 20497 5142
rect 20454 5134 20497 5137
rect 20387 5120 20497 5134
rect 19813 5102 20154 5103
rect 19738 5100 20154 5102
rect 20598 5100 20638 5189
rect 20849 5162 20914 5189
rect 20849 5144 20872 5162
rect 20890 5144 20914 5162
rect 20849 5124 20914 5144
rect 19735 5097 20638 5100
rect 19735 5077 19741 5097
rect 19761 5077 20638 5097
rect 19735 5073 20638 5077
rect 20598 5070 20638 5073
rect 20850 5063 20915 5084
rect 19068 5055 19729 5056
rect 19068 5048 20002 5055
rect 19068 5047 19974 5048
rect 19068 5027 19919 5047
rect 19951 5028 19974 5047
rect 19999 5028 20002 5048
rect 19951 5027 20002 5028
rect 19068 5020 20002 5027
rect 18667 4978 18835 4979
rect 19070 4978 19109 5020
rect 19898 5018 20002 5020
rect 19967 5016 20002 5018
rect 20850 5045 20874 5063
rect 20892 5045 20915 5063
rect 20850 4998 20915 5045
rect 18667 4952 19111 4978
rect 18667 4950 18835 4952
rect 18469 4647 18538 4731
rect 18467 4168 18538 4647
rect 18667 4599 18694 4950
rect 19070 4946 19111 4952
rect 18734 4739 18798 4751
rect 19074 4747 19111 4946
rect 19573 4973 19645 4990
rect 19573 4934 19581 4973
rect 19626 4934 19645 4973
rect 19339 4836 19450 4851
rect 19339 4834 19381 4836
rect 19339 4814 19346 4834
rect 19365 4814 19381 4834
rect 19339 4806 19381 4814
rect 19409 4834 19450 4836
rect 19409 4814 19423 4834
rect 19442 4814 19450 4834
rect 19409 4806 19450 4814
rect 19339 4800 19450 4806
rect 19282 4778 19531 4800
rect 19282 4747 19319 4778
rect 19495 4776 19531 4778
rect 19495 4747 19532 4776
rect 18734 4738 18769 4739
rect 18711 4733 18769 4738
rect 18711 4713 18714 4733
rect 18734 4719 18769 4733
rect 18789 4719 18798 4739
rect 18734 4711 18798 4719
rect 18760 4710 18798 4711
rect 18761 4709 18798 4710
rect 18864 4743 18900 4744
rect 18972 4743 19008 4744
rect 18864 4735 19008 4743
rect 18864 4715 18872 4735
rect 18892 4715 18980 4735
rect 19000 4715 19008 4735
rect 18864 4709 19008 4715
rect 19074 4739 19112 4747
rect 19180 4743 19216 4744
rect 19074 4719 19083 4739
rect 19103 4719 19112 4739
rect 19074 4710 19112 4719
rect 19131 4736 19216 4743
rect 19131 4716 19138 4736
rect 19159 4735 19216 4736
rect 19159 4716 19188 4735
rect 19131 4715 19188 4716
rect 19208 4715 19216 4735
rect 19074 4709 19111 4710
rect 19131 4709 19216 4715
rect 19282 4739 19320 4747
rect 19393 4743 19429 4744
rect 19282 4719 19291 4739
rect 19311 4719 19320 4739
rect 19282 4710 19320 4719
rect 19344 4735 19429 4743
rect 19344 4715 19401 4735
rect 19421 4715 19429 4735
rect 19282 4709 19319 4710
rect 19344 4709 19429 4715
rect 19495 4739 19533 4747
rect 19495 4719 19504 4739
rect 19524 4719 19533 4739
rect 19495 4710 19533 4719
rect 19573 4724 19645 4934
rect 19715 4968 20915 4998
rect 19715 4967 20159 4968
rect 19715 4965 19883 4967
rect 19573 4710 19656 4724
rect 19495 4709 19532 4710
rect 18918 4688 18954 4709
rect 19344 4688 19375 4709
rect 19573 4688 19590 4710
rect 18751 4684 18851 4688
rect 18751 4680 18813 4684
rect 18751 4654 18758 4680
rect 18784 4658 18813 4680
rect 18839 4658 18851 4684
rect 18784 4654 18851 4658
rect 18751 4651 18851 4654
rect 18919 4651 18954 4688
rect 19016 4685 19375 4688
rect 19016 4680 19238 4685
rect 19016 4656 19029 4680
rect 19053 4661 19238 4680
rect 19262 4661 19375 4685
rect 19053 4656 19375 4661
rect 19016 4652 19375 4656
rect 19442 4680 19590 4688
rect 19442 4660 19453 4680
rect 19473 4677 19590 4680
rect 19643 4677 19656 4710
rect 19473 4660 19656 4677
rect 19442 4653 19656 4660
rect 19442 4652 19483 4653
rect 19573 4652 19656 4653
rect 18918 4626 18954 4651
rect 18766 4599 18803 4600
rect 18862 4599 18899 4600
rect 18918 4599 18925 4626
rect 18666 4590 18804 4599
rect 18666 4570 18775 4590
rect 18795 4570 18804 4590
rect 18666 4563 18804 4570
rect 18862 4596 18925 4599
rect 18946 4599 18954 4626
rect 18973 4599 19010 4600
rect 18946 4596 19010 4599
rect 18862 4590 19010 4596
rect 18862 4570 18871 4590
rect 18891 4570 18981 4590
rect 19001 4570 19010 4590
rect 18666 4561 18762 4563
rect 18862 4560 19010 4570
rect 19069 4590 19106 4600
rect 19181 4599 19218 4600
rect 19162 4597 19218 4599
rect 19069 4570 19077 4590
rect 19097 4570 19106 4590
rect 18918 4559 18954 4560
rect 18766 4428 18803 4429
rect 19069 4428 19106 4570
rect 19131 4590 19218 4597
rect 19131 4587 19189 4590
rect 19131 4567 19136 4587
rect 19157 4570 19189 4587
rect 19209 4570 19218 4590
rect 19157 4567 19218 4570
rect 19131 4560 19218 4567
rect 19277 4590 19314 4600
rect 19277 4570 19285 4590
rect 19305 4570 19314 4590
rect 19131 4559 19162 4560
rect 19277 4491 19314 4570
rect 19344 4599 19375 4652
rect 19581 4619 19595 4652
rect 19648 4619 19656 4652
rect 19581 4613 19656 4619
rect 19581 4608 19651 4613
rect 19394 4599 19431 4600
rect 19344 4590 19431 4599
rect 19344 4570 19402 4590
rect 19422 4570 19431 4590
rect 19344 4560 19431 4570
rect 19490 4590 19527 4600
rect 19715 4595 19742 4965
rect 19782 4735 19846 4747
rect 20122 4743 20159 4967
rect 20630 4948 20694 4950
rect 20626 4936 20694 4948
rect 20626 4903 20637 4936
rect 20677 4903 20694 4936
rect 20626 4893 20694 4903
rect 20387 4832 20498 4847
rect 20387 4830 20429 4832
rect 20387 4810 20394 4830
rect 20413 4810 20429 4830
rect 20387 4802 20429 4810
rect 20457 4830 20498 4832
rect 20457 4810 20471 4830
rect 20490 4810 20498 4830
rect 20457 4802 20498 4810
rect 20387 4796 20498 4802
rect 20330 4774 20579 4796
rect 20330 4743 20367 4774
rect 20543 4772 20579 4774
rect 20543 4743 20580 4772
rect 19782 4734 19817 4735
rect 19759 4729 19817 4734
rect 19759 4709 19762 4729
rect 19782 4715 19817 4729
rect 19837 4715 19846 4735
rect 19782 4707 19846 4715
rect 19808 4706 19846 4707
rect 19809 4705 19846 4706
rect 19912 4739 19948 4740
rect 20020 4739 20056 4740
rect 19912 4731 20056 4739
rect 19912 4711 19920 4731
rect 19940 4711 20028 4731
rect 20048 4711 20056 4731
rect 19912 4705 20056 4711
rect 20122 4735 20160 4743
rect 20228 4739 20264 4740
rect 20122 4715 20131 4735
rect 20151 4715 20160 4735
rect 20122 4706 20160 4715
rect 20179 4732 20264 4739
rect 20179 4712 20186 4732
rect 20207 4731 20264 4732
rect 20207 4712 20236 4731
rect 20179 4711 20236 4712
rect 20256 4711 20264 4731
rect 20122 4705 20159 4706
rect 20179 4705 20264 4711
rect 20330 4735 20368 4743
rect 20441 4739 20477 4740
rect 20330 4715 20339 4735
rect 20359 4715 20368 4735
rect 20330 4706 20368 4715
rect 20392 4731 20477 4739
rect 20392 4711 20449 4731
rect 20469 4711 20477 4731
rect 20330 4705 20367 4706
rect 20392 4705 20477 4711
rect 20543 4735 20581 4743
rect 20543 4715 20552 4735
rect 20572 4715 20581 4735
rect 20543 4706 20581 4715
rect 20630 4709 20694 4893
rect 20850 4767 20915 4968
rect 20850 4749 20872 4767
rect 20890 4749 20915 4767
rect 20850 4730 20915 4749
rect 20543 4705 20580 4706
rect 19966 4684 20002 4705
rect 20392 4684 20423 4705
rect 20630 4700 20638 4709
rect 20627 4684 20638 4700
rect 19799 4680 19899 4684
rect 19799 4676 19861 4680
rect 19799 4650 19806 4676
rect 19832 4654 19861 4676
rect 19887 4654 19899 4680
rect 19832 4650 19899 4654
rect 19799 4647 19899 4650
rect 19967 4647 20002 4684
rect 20064 4681 20423 4684
rect 20064 4676 20286 4681
rect 20064 4652 20077 4676
rect 20101 4657 20286 4676
rect 20310 4657 20423 4681
rect 20101 4652 20423 4657
rect 20064 4648 20423 4652
rect 20490 4676 20638 4684
rect 20490 4656 20501 4676
rect 20521 4667 20638 4676
rect 20687 4700 20694 4709
rect 20687 4667 20695 4700
rect 20521 4656 20695 4667
rect 20490 4649 20695 4656
rect 20490 4648 20531 4649
rect 19966 4622 20002 4647
rect 19814 4595 19851 4596
rect 19910 4595 19947 4596
rect 19966 4595 19973 4622
rect 19490 4570 19498 4590
rect 19518 4570 19527 4590
rect 19344 4559 19375 4560
rect 19339 4491 19449 4504
rect 19490 4491 19527 4570
rect 19714 4586 19852 4595
rect 19714 4566 19823 4586
rect 19843 4566 19852 4586
rect 19714 4559 19852 4566
rect 19910 4592 19973 4595
rect 19994 4595 20002 4622
rect 20021 4595 20058 4596
rect 19994 4592 20058 4595
rect 19910 4586 20058 4592
rect 19910 4566 19919 4586
rect 19939 4566 20029 4586
rect 20049 4566 20058 4586
rect 19714 4557 19810 4559
rect 19910 4556 20058 4566
rect 20117 4586 20154 4596
rect 20229 4595 20266 4596
rect 20210 4593 20266 4595
rect 20117 4566 20125 4586
rect 20145 4566 20154 4586
rect 19966 4555 20002 4556
rect 19277 4489 19527 4491
rect 19277 4486 19378 4489
rect 19277 4467 19342 4486
rect 19339 4459 19342 4467
rect 19371 4459 19378 4486
rect 19406 4462 19416 4489
rect 19445 4467 19527 4489
rect 19445 4462 19449 4467
rect 19406 4459 19449 4462
rect 19339 4445 19449 4459
rect 18765 4427 19106 4428
rect 18690 4422 19106 4427
rect 19814 4424 19851 4425
rect 20117 4424 20154 4566
rect 20179 4586 20266 4593
rect 20179 4583 20237 4586
rect 20179 4563 20184 4583
rect 20205 4566 20237 4583
rect 20257 4566 20266 4586
rect 20205 4563 20266 4566
rect 20179 4556 20266 4563
rect 20325 4586 20362 4596
rect 20325 4566 20333 4586
rect 20353 4566 20362 4586
rect 20179 4555 20210 4556
rect 20325 4487 20362 4566
rect 20392 4595 20423 4648
rect 20627 4646 20695 4649
rect 20627 4604 20639 4646
rect 20688 4604 20695 4646
rect 20442 4595 20479 4596
rect 20392 4586 20479 4595
rect 20392 4566 20450 4586
rect 20470 4566 20479 4586
rect 20392 4556 20479 4566
rect 20538 4586 20575 4596
rect 20627 4591 20695 4604
rect 20850 4668 20915 4685
rect 20850 4650 20874 4668
rect 20892 4650 20915 4668
rect 20538 4566 20546 4586
rect 20566 4566 20575 4586
rect 20392 4555 20423 4556
rect 20387 4487 20497 4500
rect 20538 4487 20575 4566
rect 20850 4511 20915 4650
rect 20850 4505 20872 4511
rect 20325 4485 20575 4487
rect 20325 4482 20426 4485
rect 20325 4463 20390 4482
rect 20387 4455 20390 4463
rect 20419 4455 20426 4482
rect 20454 4458 20464 4485
rect 20493 4463 20575 4485
rect 20604 4493 20872 4505
rect 20890 4493 20915 4511
rect 20604 4470 20915 4493
rect 20604 4469 20659 4470
rect 20493 4458 20497 4463
rect 20454 4455 20497 4458
rect 20387 4441 20497 4455
rect 19813 4423 20154 4424
rect 18690 4402 18693 4422
rect 18713 4402 19106 4422
rect 19738 4422 20154 4423
rect 20604 4422 20647 4469
rect 19738 4418 20647 4422
rect 19057 4369 19102 4402
rect 19738 4398 19741 4418
rect 19761 4398 20647 4418
rect 20115 4393 20647 4398
rect 20855 4412 20914 4434
rect 20855 4394 20874 4412
rect 20892 4394 20914 4412
rect 19903 4369 20002 4371
rect 19057 4359 20002 4369
rect 19057 4333 19925 4359
rect 19058 4332 19925 4333
rect 19903 4321 19925 4332
rect 19950 4324 19969 4359
rect 19994 4324 20002 4359
rect 19950 4321 20002 4324
rect 19903 4313 20002 4321
rect 19929 4312 20001 4313
rect 20855 4264 20914 4394
rect 19577 4234 19653 4258
rect 19577 4168 19589 4234
rect 19643 4168 19653 4234
rect 20121 4189 20162 4191
rect 20393 4189 20497 4191
rect 20855 4189 20916 4264
rect 18467 4118 18539 4168
rect 18036 3846 18372 3850
rect 17262 3842 17362 3846
rect 17262 3838 17324 3842
rect 17262 3812 17269 3838
rect 17295 3816 17324 3838
rect 17350 3816 17362 3842
rect 17295 3812 17362 3816
rect 17262 3809 17362 3812
rect 17430 3809 17465 3846
rect 17527 3843 17886 3846
rect 17527 3838 17749 3843
rect 17527 3814 17540 3838
rect 17564 3819 17749 3838
rect 17773 3819 17886 3843
rect 17564 3814 17886 3819
rect 17527 3810 17886 3814
rect 17953 3838 18372 3846
rect 17953 3818 17964 3838
rect 17984 3818 18372 3838
rect 17953 3811 18372 3818
rect 17953 3810 17994 3811
rect 18036 3810 18372 3811
rect 17429 3784 17465 3809
rect 17277 3757 17314 3758
rect 17373 3757 17410 3758
rect 17429 3757 17436 3784
rect 17177 3748 17315 3757
rect 17177 3728 17286 3748
rect 17306 3728 17315 3748
rect 17177 3721 17315 3728
rect 17373 3754 17436 3757
rect 17457 3757 17465 3784
rect 17484 3757 17521 3758
rect 17457 3754 17521 3757
rect 17373 3748 17521 3754
rect 17373 3728 17382 3748
rect 17402 3728 17492 3748
rect 17512 3728 17521 3748
rect 17177 3719 17273 3721
rect 17373 3718 17521 3728
rect 17580 3748 17617 3758
rect 17692 3757 17729 3758
rect 17673 3755 17729 3757
rect 17580 3728 17588 3748
rect 17608 3728 17617 3748
rect 17429 3717 17465 3718
rect 17277 3586 17314 3587
rect 17580 3586 17617 3728
rect 17642 3748 17729 3755
rect 17642 3745 17700 3748
rect 17642 3725 17647 3745
rect 17668 3728 17700 3745
rect 17720 3728 17729 3748
rect 17668 3725 17729 3728
rect 17642 3718 17729 3725
rect 17788 3748 17825 3758
rect 17788 3728 17796 3748
rect 17816 3728 17825 3748
rect 17642 3717 17673 3718
rect 17788 3649 17825 3728
rect 17855 3757 17886 3810
rect 18280 3774 18372 3810
rect 17905 3757 17942 3758
rect 17855 3748 17942 3757
rect 17855 3728 17913 3748
rect 17933 3728 17942 3748
rect 17855 3718 17942 3728
rect 18001 3748 18038 3758
rect 18001 3728 18009 3748
rect 18029 3728 18038 3748
rect 17855 3717 17886 3718
rect 17850 3649 17960 3662
rect 18001 3649 18038 3728
rect 17788 3647 18038 3649
rect 17788 3644 17889 3647
rect 17788 3625 17853 3644
rect 17850 3617 17853 3625
rect 17882 3617 17889 3644
rect 17917 3620 17927 3647
rect 17956 3625 18038 3647
rect 17956 3620 17960 3625
rect 17917 3617 17960 3620
rect 17850 3603 17960 3617
rect 17276 3585 17617 3586
rect 17201 3580 17617 3585
rect 17201 3560 17204 3580
rect 17224 3560 17617 3580
rect 17361 3516 17466 3519
rect 17360 3493 17466 3516
rect 16480 3491 16981 3493
rect 17122 3491 17471 3493
rect 14594 3470 14631 3491
rect 14594 3433 14605 3470
rect 14622 3433 14631 3470
rect 16480 3485 17471 3491
rect 16480 3480 17432 3485
rect 16480 3459 17391 3480
rect 17411 3464 17432 3480
rect 17452 3464 17471 3485
rect 17411 3459 17471 3464
rect 16480 3434 17471 3459
rect 16956 3433 17138 3434
rect 14594 3423 14631 3433
rect 14440 3380 14834 3400
rect 14854 3380 14857 3400
rect 14441 3375 14857 3380
rect 14441 3374 14782 3375
rect 14098 3343 14208 3357
rect 14098 3340 14141 3343
rect 14098 3335 14102 3340
rect 14020 3313 14102 3335
rect 14131 3313 14141 3340
rect 14169 3316 14176 3343
rect 14205 3335 14208 3343
rect 14205 3316 14270 3335
rect 14169 3313 14270 3316
rect 14020 3311 14270 3313
rect 14020 3232 14057 3311
rect 14098 3298 14208 3311
rect 14172 3242 14203 3243
rect 14020 3212 14029 3232
rect 14049 3212 14057 3232
rect 14020 3202 14057 3212
rect 14116 3232 14203 3242
rect 14116 3212 14125 3232
rect 14145 3212 14203 3232
rect 14116 3203 14203 3212
rect 14116 3202 14153 3203
rect 14172 3150 14203 3203
rect 14233 3232 14270 3311
rect 14385 3242 14416 3243
rect 14233 3212 14242 3232
rect 14262 3212 14270 3232
rect 14233 3202 14270 3212
rect 14329 3235 14416 3242
rect 14329 3232 14390 3235
rect 14329 3212 14338 3232
rect 14358 3215 14390 3232
rect 14411 3215 14416 3235
rect 14358 3212 14416 3215
rect 14329 3205 14416 3212
rect 14441 3232 14478 3374
rect 14744 3373 14781 3374
rect 14593 3242 14629 3243
rect 14441 3212 14450 3232
rect 14470 3212 14478 3232
rect 14329 3203 14385 3205
rect 14329 3202 14366 3203
rect 14441 3202 14478 3212
rect 14537 3232 14685 3242
rect 14785 3239 14881 3241
rect 14537 3212 14546 3232
rect 14566 3212 14656 3232
rect 14676 3212 14685 3232
rect 14537 3206 14685 3212
rect 14537 3203 14601 3206
rect 14537 3202 14574 3203
rect 14593 3176 14601 3203
rect 14622 3203 14685 3206
rect 14743 3232 14881 3239
rect 14743 3212 14752 3232
rect 14772 3212 14881 3232
rect 14743 3203 14881 3212
rect 17510 3204 17541 3560
rect 14622 3176 14629 3203
rect 14648 3202 14685 3203
rect 14744 3202 14781 3203
rect 14593 3151 14629 3176
rect 14064 3149 14105 3150
rect 13984 3144 14105 3149
rect 13935 3142 14105 3144
rect 13935 3131 14074 3142
rect 13935 3108 13958 3131
rect 13984 3122 14074 3131
rect 14094 3122 14105 3142
rect 13984 3114 14105 3122
rect 14172 3146 14531 3150
rect 14172 3141 14494 3146
rect 14172 3117 14285 3141
rect 14309 3122 14494 3141
rect 14518 3122 14531 3146
rect 14309 3117 14531 3122
rect 14172 3114 14531 3117
rect 14593 3114 14628 3151
rect 14696 3148 14796 3151
rect 14696 3144 14763 3148
rect 14696 3118 14708 3144
rect 14734 3122 14763 3144
rect 14789 3122 14796 3148
rect 14734 3118 14796 3122
rect 14696 3114 14796 3118
rect 13984 3108 13992 3114
rect 13935 3100 13992 3108
rect 14172 3093 14203 3114
rect 14593 3093 14629 3114
rect 14015 3092 14052 3093
rect 14014 3083 14052 3092
rect 14014 3063 14023 3083
rect 14043 3063 14052 3083
rect 14014 3055 14052 3063
rect 14118 3087 14203 3093
rect 14228 3092 14265 3093
rect 14118 3067 14126 3087
rect 14146 3067 14203 3087
rect 14118 3059 14203 3067
rect 14227 3083 14265 3092
rect 14227 3063 14236 3083
rect 14256 3063 14265 3083
rect 14118 3058 14154 3059
rect 14227 3055 14265 3063
rect 14331 3087 14416 3093
rect 14436 3092 14473 3093
rect 14331 3067 14339 3087
rect 14359 3086 14416 3087
rect 14359 3067 14388 3086
rect 14331 3066 14388 3067
rect 14409 3066 14416 3086
rect 14331 3059 14416 3066
rect 14435 3083 14473 3092
rect 14435 3063 14444 3083
rect 14464 3063 14473 3083
rect 14331 3058 14367 3059
rect 14435 3055 14473 3063
rect 14539 3087 14683 3093
rect 14539 3067 14547 3087
rect 14567 3067 14655 3087
rect 14675 3067 14683 3087
rect 14539 3059 14683 3067
rect 14539 3058 14575 3059
rect 14647 3058 14683 3059
rect 14749 3092 14786 3093
rect 14749 3091 14787 3092
rect 14749 3083 14813 3091
rect 14749 3063 14758 3083
rect 14778 3069 14813 3083
rect 14833 3069 14836 3089
rect 14778 3064 14836 3069
rect 14778 3063 14813 3064
rect 14015 3026 14052 3055
rect 14016 3024 14052 3026
rect 14228 3024 14265 3055
rect 14016 3002 14265 3024
rect 14097 2996 14208 3002
rect 14097 2988 14138 2996
rect 14097 2968 14105 2988
rect 14124 2968 14138 2988
rect 14097 2966 14138 2968
rect 14166 2988 14208 2996
rect 14166 2968 14182 2988
rect 14201 2968 14208 2988
rect 14166 2966 14208 2968
rect 14097 2951 14208 2966
rect 14436 2940 14473 3055
rect 14749 3051 14813 3063
rect 14429 2934 14476 2940
rect 14853 2936 14880 3203
rect 17428 3175 17541 3204
rect 14712 2934 14880 2936
rect 14429 2908 14880 2934
rect 14429 2773 14476 2908
rect 14712 2907 14880 2908
rect 17429 2866 17465 3175
rect 18289 3061 18370 3774
rect 18469 3209 18539 4118
rect 19577 4148 19653 4168
rect 19577 4111 19594 4148
rect 19638 4111 19653 4148
rect 19714 4154 20916 4189
rect 19714 4140 19742 4154
rect 19577 4095 19653 4111
rect 19582 3939 19652 4095
rect 19716 4009 19742 4140
rect 20121 4151 20916 4154
rect 19574 3888 19654 3939
rect 19574 3862 19590 3888
rect 19630 3862 19654 3888
rect 19574 3843 19654 3862
rect 19574 3817 19593 3843
rect 19633 3817 19654 3843
rect 19574 3790 19654 3817
rect 19574 3764 19597 3790
rect 19637 3764 19654 3790
rect 19574 3753 19654 3764
rect 19716 3754 19743 4009
rect 20121 4001 20162 4151
rect 20855 4139 20916 4151
rect 20588 4089 20709 4107
rect 20588 4087 20659 4089
rect 20588 4046 20603 4087
rect 20640 4048 20659 4087
rect 20696 4048 20709 4089
rect 20640 4046 20709 4048
rect 20588 4036 20709 4046
rect 20393 4006 20497 4015
rect 19783 3894 19847 3906
rect 20123 3902 20160 4001
rect 20388 3991 20499 4006
rect 20388 3989 20430 3991
rect 20388 3969 20395 3989
rect 20414 3969 20430 3989
rect 20388 3961 20430 3969
rect 20458 3989 20499 3991
rect 20458 3969 20472 3989
rect 20491 3969 20499 3989
rect 20458 3961 20499 3969
rect 20388 3955 20499 3961
rect 20331 3933 20580 3955
rect 20331 3902 20368 3933
rect 20544 3931 20580 3933
rect 20544 3902 20581 3931
rect 19783 3893 19818 3894
rect 19760 3888 19818 3893
rect 19760 3868 19763 3888
rect 19783 3874 19818 3888
rect 19838 3874 19847 3894
rect 19783 3866 19847 3874
rect 19809 3865 19847 3866
rect 19810 3864 19847 3865
rect 19913 3898 19949 3899
rect 20021 3898 20057 3899
rect 19913 3890 20057 3898
rect 19913 3870 19921 3890
rect 19941 3870 20029 3890
rect 20049 3870 20057 3890
rect 19913 3864 20057 3870
rect 20123 3894 20161 3902
rect 20229 3898 20265 3899
rect 20123 3874 20132 3894
rect 20152 3874 20161 3894
rect 20123 3865 20161 3874
rect 20180 3891 20265 3898
rect 20180 3871 20187 3891
rect 20208 3890 20265 3891
rect 20208 3871 20237 3890
rect 20180 3870 20237 3871
rect 20257 3870 20265 3890
rect 20123 3864 20160 3865
rect 20180 3864 20265 3870
rect 20331 3894 20369 3902
rect 20442 3898 20478 3899
rect 20331 3874 20340 3894
rect 20360 3874 20369 3894
rect 20331 3865 20369 3874
rect 20393 3890 20478 3898
rect 20393 3870 20450 3890
rect 20470 3870 20478 3890
rect 20331 3864 20368 3865
rect 20393 3864 20478 3870
rect 20544 3894 20582 3902
rect 20544 3874 20553 3894
rect 20573 3874 20582 3894
rect 20637 3884 20702 4036
rect 20855 4010 20910 4139
rect 20544 3865 20582 3874
rect 20635 3877 20702 3884
rect 20544 3864 20581 3865
rect 19967 3843 20003 3864
rect 20393 3843 20424 3864
rect 20635 3856 20652 3877
rect 20688 3856 20702 3877
rect 20854 3897 20910 4010
rect 20854 3879 20873 3897
rect 20891 3879 20910 3897
rect 20854 3859 20910 3879
rect 20635 3843 20702 3856
rect 19800 3839 19900 3843
rect 19800 3835 19862 3839
rect 19800 3809 19807 3835
rect 19833 3813 19862 3835
rect 19888 3813 19900 3839
rect 19833 3809 19900 3813
rect 19800 3806 19900 3809
rect 19968 3806 20003 3843
rect 20065 3840 20424 3843
rect 20065 3835 20287 3840
rect 20065 3811 20078 3835
rect 20102 3816 20287 3835
rect 20311 3816 20424 3840
rect 20102 3811 20424 3816
rect 20065 3807 20424 3811
rect 20491 3837 20702 3843
rect 20491 3835 20652 3837
rect 20491 3815 20502 3835
rect 20522 3815 20652 3835
rect 20491 3808 20652 3815
rect 20491 3807 20532 3808
rect 19967 3781 20003 3806
rect 19815 3754 19852 3755
rect 19911 3754 19948 3755
rect 19967 3754 19974 3781
rect 19715 3745 19853 3754
rect 19715 3725 19824 3745
rect 19844 3725 19853 3745
rect 19715 3718 19853 3725
rect 19911 3751 19974 3754
rect 19995 3754 20003 3781
rect 20022 3754 20059 3755
rect 19995 3751 20059 3754
rect 19911 3745 20059 3751
rect 19911 3725 19920 3745
rect 19940 3725 20030 3745
rect 20050 3725 20059 3745
rect 19715 3716 19811 3718
rect 19911 3715 20059 3725
rect 20118 3745 20155 3755
rect 20230 3754 20267 3755
rect 20211 3752 20267 3754
rect 20118 3725 20126 3745
rect 20146 3725 20155 3745
rect 19967 3714 20003 3715
rect 19815 3583 19852 3584
rect 20118 3583 20155 3725
rect 20180 3745 20267 3752
rect 20180 3742 20238 3745
rect 20180 3722 20185 3742
rect 20206 3725 20238 3742
rect 20258 3725 20267 3745
rect 20206 3722 20267 3725
rect 20180 3715 20267 3722
rect 20326 3745 20363 3755
rect 20326 3725 20334 3745
rect 20354 3725 20363 3745
rect 20180 3714 20211 3715
rect 20326 3646 20363 3725
rect 20393 3754 20424 3807
rect 20637 3800 20652 3808
rect 20692 3800 20702 3837
rect 20637 3791 20702 3800
rect 20850 3798 20915 3819
rect 20850 3780 20875 3798
rect 20893 3780 20915 3798
rect 20443 3754 20480 3755
rect 20393 3745 20480 3754
rect 20393 3725 20451 3745
rect 20471 3725 20480 3745
rect 20393 3715 20480 3725
rect 20539 3745 20576 3755
rect 20539 3725 20547 3745
rect 20567 3725 20576 3745
rect 20393 3714 20424 3715
rect 20388 3646 20498 3659
rect 20539 3646 20576 3725
rect 20850 3704 20915 3780
rect 20326 3644 20576 3646
rect 20326 3641 20427 3644
rect 20326 3622 20391 3641
rect 20388 3614 20391 3622
rect 20420 3614 20427 3641
rect 20455 3617 20465 3644
rect 20494 3622 20576 3644
rect 20599 3669 20916 3704
rect 20494 3617 20498 3622
rect 20455 3614 20498 3617
rect 20388 3600 20498 3614
rect 19814 3582 20155 3583
rect 19739 3580 20155 3582
rect 20599 3580 20639 3669
rect 20850 3642 20915 3669
rect 20850 3624 20873 3642
rect 20891 3624 20915 3642
rect 20850 3604 20915 3624
rect 19736 3577 20639 3580
rect 19736 3557 19742 3577
rect 19762 3557 20639 3577
rect 19736 3553 20639 3557
rect 20599 3550 20639 3553
rect 20851 3543 20916 3564
rect 19069 3535 19730 3536
rect 19069 3528 20003 3535
rect 19069 3527 19975 3528
rect 19069 3507 19920 3527
rect 19952 3508 19975 3527
rect 20000 3508 20003 3528
rect 19952 3507 20003 3508
rect 19069 3500 20003 3507
rect 18668 3458 18836 3459
rect 19071 3458 19110 3500
rect 19899 3498 20003 3500
rect 19968 3496 20003 3498
rect 20851 3525 20875 3543
rect 20893 3525 20916 3543
rect 20851 3478 20916 3525
rect 18668 3432 19112 3458
rect 18668 3430 18836 3432
rect 17429 2843 17433 2866
rect 17457 2843 17465 2866
rect 17629 2844 17728 2848
rect 17429 2822 17465 2843
rect 17429 2799 17433 2822
rect 17457 2799 17465 2822
rect 17429 2795 17465 2799
rect 17625 2838 17728 2844
rect 17625 2800 17651 2838
rect 17676 2803 17695 2838
rect 17720 2803 17728 2838
rect 17676 2800 17728 2803
rect 17625 2792 17728 2800
rect 17625 2791 17727 2792
rect 14427 2724 14486 2773
rect 14427 2696 14445 2724
rect 14473 2696 14486 2724
rect 14427 2686 14486 2696
rect 17221 2713 17389 2714
rect 17625 2713 17672 2791
rect 17221 2687 17672 2713
rect 17221 2685 17389 2687
rect 17221 2312 17248 2685
rect 17418 2637 17504 2646
rect 17418 2619 17437 2637
rect 17489 2619 17504 2637
rect 17418 2615 17504 2619
rect 17288 2452 17352 2464
rect 17288 2451 17323 2452
rect 17265 2446 17323 2451
rect 17265 2426 17268 2446
rect 17288 2432 17323 2446
rect 17343 2432 17352 2452
rect 17288 2424 17352 2432
rect 17314 2423 17352 2424
rect 17315 2422 17352 2423
rect 17418 2456 17454 2457
rect 17474 2456 17504 2615
rect 17625 2575 17672 2687
rect 17628 2460 17665 2575
rect 17893 2549 18004 2564
rect 17893 2547 17935 2549
rect 17893 2527 17900 2547
rect 17919 2527 17935 2547
rect 17893 2519 17935 2527
rect 17963 2547 18004 2549
rect 17963 2527 17977 2547
rect 17996 2527 18004 2547
rect 17963 2519 18004 2527
rect 17893 2513 18004 2519
rect 17836 2491 18085 2513
rect 17836 2460 17873 2491
rect 18049 2489 18085 2491
rect 18049 2460 18086 2489
rect 18290 2476 18369 3061
rect 18466 2609 18545 3209
rect 18668 3079 18695 3430
rect 19071 3426 19112 3432
rect 18735 3219 18799 3231
rect 19075 3227 19112 3426
rect 19574 3453 19646 3470
rect 19574 3414 19582 3453
rect 19627 3414 19646 3453
rect 19340 3316 19451 3331
rect 19340 3314 19382 3316
rect 19340 3294 19347 3314
rect 19366 3294 19382 3314
rect 19340 3286 19382 3294
rect 19410 3314 19451 3316
rect 19410 3294 19424 3314
rect 19443 3294 19451 3314
rect 19410 3286 19451 3294
rect 19340 3280 19451 3286
rect 19283 3258 19532 3280
rect 19283 3227 19320 3258
rect 19496 3256 19532 3258
rect 19496 3227 19533 3256
rect 18735 3218 18770 3219
rect 18712 3213 18770 3218
rect 18712 3193 18715 3213
rect 18735 3199 18770 3213
rect 18790 3199 18799 3219
rect 18735 3191 18799 3199
rect 18761 3190 18799 3191
rect 18762 3189 18799 3190
rect 18865 3223 18901 3224
rect 18973 3223 19009 3224
rect 18865 3215 19009 3223
rect 18865 3195 18873 3215
rect 18893 3195 18981 3215
rect 19001 3195 19009 3215
rect 18865 3189 19009 3195
rect 19075 3219 19113 3227
rect 19181 3223 19217 3224
rect 19075 3199 19084 3219
rect 19104 3199 19113 3219
rect 19075 3190 19113 3199
rect 19132 3216 19217 3223
rect 19132 3196 19139 3216
rect 19160 3215 19217 3216
rect 19160 3196 19189 3215
rect 19132 3195 19189 3196
rect 19209 3195 19217 3215
rect 19075 3189 19112 3190
rect 19132 3189 19217 3195
rect 19283 3219 19321 3227
rect 19394 3223 19430 3224
rect 19283 3199 19292 3219
rect 19312 3199 19321 3219
rect 19283 3190 19321 3199
rect 19345 3215 19430 3223
rect 19345 3195 19402 3215
rect 19422 3195 19430 3215
rect 19283 3189 19320 3190
rect 19345 3189 19430 3195
rect 19496 3219 19534 3227
rect 19496 3199 19505 3219
rect 19525 3199 19534 3219
rect 19496 3190 19534 3199
rect 19574 3204 19646 3414
rect 19716 3448 20916 3478
rect 19716 3447 20160 3448
rect 19716 3445 19884 3447
rect 19574 3190 19657 3204
rect 19496 3189 19533 3190
rect 18919 3168 18955 3189
rect 19345 3168 19376 3189
rect 19574 3168 19591 3190
rect 18752 3164 18852 3168
rect 18752 3160 18814 3164
rect 18752 3134 18759 3160
rect 18785 3138 18814 3160
rect 18840 3138 18852 3164
rect 18785 3134 18852 3138
rect 18752 3131 18852 3134
rect 18920 3131 18955 3168
rect 19017 3165 19376 3168
rect 19017 3160 19239 3165
rect 19017 3136 19030 3160
rect 19054 3141 19239 3160
rect 19263 3141 19376 3165
rect 19054 3136 19376 3141
rect 19017 3132 19376 3136
rect 19443 3160 19591 3168
rect 19443 3140 19454 3160
rect 19474 3157 19591 3160
rect 19644 3157 19657 3190
rect 19474 3140 19657 3157
rect 19443 3133 19657 3140
rect 19443 3132 19484 3133
rect 19574 3132 19657 3133
rect 18919 3106 18955 3131
rect 18767 3079 18804 3080
rect 18863 3079 18900 3080
rect 18919 3079 18926 3106
rect 18667 3070 18805 3079
rect 18667 3050 18776 3070
rect 18796 3050 18805 3070
rect 18667 3043 18805 3050
rect 18863 3076 18926 3079
rect 18947 3079 18955 3106
rect 18974 3079 19011 3080
rect 18947 3076 19011 3079
rect 18863 3070 19011 3076
rect 18863 3050 18872 3070
rect 18892 3050 18982 3070
rect 19002 3050 19011 3070
rect 18667 3041 18763 3043
rect 18863 3040 19011 3050
rect 19070 3070 19107 3080
rect 19182 3079 19219 3080
rect 19163 3077 19219 3079
rect 19070 3050 19078 3070
rect 19098 3050 19107 3070
rect 18919 3039 18955 3040
rect 18767 2908 18804 2909
rect 19070 2908 19107 3050
rect 19132 3070 19219 3077
rect 19132 3067 19190 3070
rect 19132 3047 19137 3067
rect 19158 3050 19190 3067
rect 19210 3050 19219 3070
rect 19158 3047 19219 3050
rect 19132 3040 19219 3047
rect 19278 3070 19315 3080
rect 19278 3050 19286 3070
rect 19306 3050 19315 3070
rect 19132 3039 19163 3040
rect 19278 2971 19315 3050
rect 19345 3079 19376 3132
rect 19582 3099 19596 3132
rect 19649 3099 19657 3132
rect 19582 3093 19657 3099
rect 19582 3088 19652 3093
rect 19395 3079 19432 3080
rect 19345 3070 19432 3079
rect 19345 3050 19403 3070
rect 19423 3050 19432 3070
rect 19345 3040 19432 3050
rect 19491 3070 19528 3080
rect 19716 3075 19743 3445
rect 19783 3215 19847 3227
rect 20123 3223 20160 3447
rect 20631 3428 20695 3430
rect 20627 3416 20695 3428
rect 20627 3383 20638 3416
rect 20678 3383 20695 3416
rect 20627 3373 20695 3383
rect 20388 3312 20499 3327
rect 20388 3310 20430 3312
rect 20388 3290 20395 3310
rect 20414 3290 20430 3310
rect 20388 3282 20430 3290
rect 20458 3310 20499 3312
rect 20458 3290 20472 3310
rect 20491 3290 20499 3310
rect 20458 3282 20499 3290
rect 20388 3276 20499 3282
rect 20331 3254 20580 3276
rect 20331 3223 20368 3254
rect 20544 3252 20580 3254
rect 20544 3223 20581 3252
rect 19783 3214 19818 3215
rect 19760 3209 19818 3214
rect 19760 3189 19763 3209
rect 19783 3195 19818 3209
rect 19838 3195 19847 3215
rect 19783 3187 19847 3195
rect 19809 3186 19847 3187
rect 19810 3185 19847 3186
rect 19913 3219 19949 3220
rect 20021 3219 20057 3220
rect 19913 3211 20057 3219
rect 19913 3191 19921 3211
rect 19941 3191 20029 3211
rect 20049 3191 20057 3211
rect 19913 3185 20057 3191
rect 20123 3215 20161 3223
rect 20229 3219 20265 3220
rect 20123 3195 20132 3215
rect 20152 3195 20161 3215
rect 20123 3186 20161 3195
rect 20180 3212 20265 3219
rect 20180 3192 20187 3212
rect 20208 3211 20265 3212
rect 20208 3192 20237 3211
rect 20180 3191 20237 3192
rect 20257 3191 20265 3211
rect 20123 3185 20160 3186
rect 20180 3185 20265 3191
rect 20331 3215 20369 3223
rect 20442 3219 20478 3220
rect 20331 3195 20340 3215
rect 20360 3195 20369 3215
rect 20331 3186 20369 3195
rect 20393 3211 20478 3219
rect 20393 3191 20450 3211
rect 20470 3191 20478 3211
rect 20331 3185 20368 3186
rect 20393 3185 20478 3191
rect 20544 3215 20582 3223
rect 20544 3195 20553 3215
rect 20573 3195 20582 3215
rect 20544 3186 20582 3195
rect 20631 3189 20695 3373
rect 20851 3247 20916 3448
rect 20851 3229 20873 3247
rect 20891 3229 20916 3247
rect 20851 3210 20916 3229
rect 20544 3185 20581 3186
rect 19967 3164 20003 3185
rect 20393 3164 20424 3185
rect 20631 3180 20639 3189
rect 20628 3164 20639 3180
rect 19800 3160 19900 3164
rect 19800 3156 19862 3160
rect 19800 3130 19807 3156
rect 19833 3134 19862 3156
rect 19888 3134 19900 3160
rect 19833 3130 19900 3134
rect 19800 3127 19900 3130
rect 19968 3127 20003 3164
rect 20065 3161 20424 3164
rect 20065 3156 20287 3161
rect 20065 3132 20078 3156
rect 20102 3137 20287 3156
rect 20311 3137 20424 3161
rect 20102 3132 20424 3137
rect 20065 3128 20424 3132
rect 20491 3156 20639 3164
rect 20491 3136 20502 3156
rect 20522 3147 20639 3156
rect 20688 3180 20695 3189
rect 20688 3147 20696 3180
rect 20522 3136 20696 3147
rect 20491 3129 20696 3136
rect 20491 3128 20532 3129
rect 19967 3102 20003 3127
rect 19815 3075 19852 3076
rect 19911 3075 19948 3076
rect 19967 3075 19974 3102
rect 19491 3050 19499 3070
rect 19519 3050 19528 3070
rect 19345 3039 19376 3040
rect 19340 2971 19450 2984
rect 19491 2971 19528 3050
rect 19715 3066 19853 3075
rect 19715 3046 19824 3066
rect 19844 3046 19853 3066
rect 19715 3039 19853 3046
rect 19911 3072 19974 3075
rect 19995 3075 20003 3102
rect 20022 3075 20059 3076
rect 19995 3072 20059 3075
rect 19911 3066 20059 3072
rect 19911 3046 19920 3066
rect 19940 3046 20030 3066
rect 20050 3046 20059 3066
rect 19715 3037 19811 3039
rect 19911 3036 20059 3046
rect 20118 3066 20155 3076
rect 20230 3075 20267 3076
rect 20211 3073 20267 3075
rect 20118 3046 20126 3066
rect 20146 3046 20155 3066
rect 19967 3035 20003 3036
rect 19278 2969 19528 2971
rect 19278 2966 19379 2969
rect 19278 2947 19343 2966
rect 19340 2939 19343 2947
rect 19372 2939 19379 2966
rect 19407 2942 19417 2969
rect 19446 2947 19528 2969
rect 19446 2942 19450 2947
rect 19407 2939 19450 2942
rect 19340 2925 19450 2939
rect 18766 2907 19107 2908
rect 18691 2902 19107 2907
rect 19815 2904 19852 2905
rect 20118 2904 20155 3046
rect 20180 3066 20267 3073
rect 20180 3063 20238 3066
rect 20180 3043 20185 3063
rect 20206 3046 20238 3063
rect 20258 3046 20267 3066
rect 20206 3043 20267 3046
rect 20180 3036 20267 3043
rect 20326 3066 20363 3076
rect 20326 3046 20334 3066
rect 20354 3046 20363 3066
rect 20180 3035 20211 3036
rect 20326 2967 20363 3046
rect 20393 3075 20424 3128
rect 20628 3126 20696 3129
rect 20628 3084 20640 3126
rect 20689 3084 20696 3126
rect 20443 3075 20480 3076
rect 20393 3066 20480 3075
rect 20393 3046 20451 3066
rect 20471 3046 20480 3066
rect 20393 3036 20480 3046
rect 20539 3066 20576 3076
rect 20628 3071 20696 3084
rect 20851 3148 20916 3165
rect 20851 3130 20875 3148
rect 20893 3130 20916 3148
rect 20539 3046 20547 3066
rect 20567 3046 20576 3066
rect 20393 3035 20424 3036
rect 20388 2967 20498 2980
rect 20539 2967 20576 3046
rect 20851 2991 20916 3130
rect 20851 2985 20873 2991
rect 20326 2965 20576 2967
rect 20326 2962 20427 2965
rect 20326 2943 20391 2962
rect 20388 2935 20391 2943
rect 20420 2935 20427 2962
rect 20455 2938 20465 2965
rect 20494 2943 20576 2965
rect 20605 2973 20873 2985
rect 20891 2973 20916 2991
rect 20605 2950 20916 2973
rect 20605 2949 20660 2950
rect 20494 2938 20498 2943
rect 20455 2935 20498 2938
rect 20388 2921 20498 2935
rect 19814 2903 20155 2904
rect 18691 2882 18694 2902
rect 18714 2882 19107 2902
rect 19739 2902 20155 2903
rect 20605 2902 20648 2949
rect 19739 2898 20648 2902
rect 19058 2849 19103 2882
rect 19739 2878 19742 2898
rect 19762 2878 20648 2898
rect 20116 2873 20648 2878
rect 20856 2892 20915 2914
rect 20856 2874 20875 2892
rect 20893 2874 20915 2892
rect 19904 2849 20003 2851
rect 19058 2839 20003 2849
rect 19058 2813 19926 2839
rect 19059 2812 19926 2813
rect 19904 2801 19926 2812
rect 19951 2804 19970 2839
rect 19995 2804 20003 2839
rect 19951 2801 20003 2804
rect 20856 2803 20915 2874
rect 19904 2793 20003 2801
rect 19930 2792 20002 2793
rect 19584 2766 19651 2785
rect 19584 2745 19601 2766
rect 18465 2567 18545 2609
rect 19582 2700 19601 2745
rect 19631 2745 19651 2766
rect 19631 2700 19652 2745
rect 20121 2742 20162 2744
rect 20393 2742 20497 2744
rect 20853 2742 20917 2803
rect 17526 2456 17562 2457
rect 17418 2448 17562 2456
rect 17418 2428 17426 2448
rect 17446 2428 17534 2448
rect 17554 2428 17562 2448
rect 17418 2422 17562 2428
rect 17628 2452 17666 2460
rect 17734 2456 17770 2457
rect 17628 2432 17637 2452
rect 17657 2432 17666 2452
rect 17628 2423 17666 2432
rect 17685 2449 17770 2456
rect 17685 2429 17692 2449
rect 17713 2448 17770 2449
rect 17713 2429 17742 2448
rect 17685 2428 17742 2429
rect 17762 2428 17770 2448
rect 17628 2422 17665 2423
rect 17685 2422 17770 2428
rect 17836 2452 17874 2460
rect 17947 2456 17983 2457
rect 17836 2432 17845 2452
rect 17865 2432 17874 2452
rect 17836 2423 17874 2432
rect 17898 2448 17983 2456
rect 17898 2428 17955 2448
rect 17975 2428 17983 2448
rect 17836 2422 17873 2423
rect 17898 2422 17983 2428
rect 18049 2452 18087 2460
rect 18049 2432 18058 2452
rect 18078 2432 18087 2452
rect 18049 2423 18087 2432
rect 18287 2440 18373 2476
rect 18049 2422 18086 2423
rect 17472 2401 17508 2422
rect 17898 2401 17929 2422
rect 18125 2401 18171 2405
rect 17305 2397 17405 2401
rect 17305 2393 17367 2397
rect 17305 2367 17312 2393
rect 17338 2371 17367 2393
rect 17393 2371 17405 2397
rect 17338 2367 17405 2371
rect 17305 2364 17405 2367
rect 17473 2364 17508 2401
rect 17570 2398 17929 2401
rect 17570 2393 17792 2398
rect 17570 2369 17583 2393
rect 17607 2374 17792 2393
rect 17816 2374 17929 2398
rect 17607 2369 17929 2374
rect 17570 2365 17929 2369
rect 17996 2393 18171 2401
rect 17996 2373 18007 2393
rect 18027 2373 18171 2393
rect 18287 2399 18304 2440
rect 18358 2399 18373 2440
rect 18287 2380 18373 2399
rect 17996 2366 18171 2373
rect 17996 2365 18037 2366
rect 17472 2339 17508 2364
rect 17320 2312 17357 2313
rect 17416 2312 17453 2313
rect 17472 2312 17479 2339
rect 17220 2303 17358 2312
rect 17220 2283 17329 2303
rect 17349 2283 17358 2303
rect 17220 2276 17358 2283
rect 17416 2309 17479 2312
rect 17500 2312 17508 2339
rect 17527 2312 17564 2313
rect 17500 2309 17564 2312
rect 17416 2303 17564 2309
rect 17416 2283 17425 2303
rect 17445 2283 17535 2303
rect 17555 2283 17564 2303
rect 17220 2274 17316 2276
rect 17416 2273 17564 2283
rect 17623 2303 17660 2313
rect 17735 2312 17772 2313
rect 17716 2310 17772 2312
rect 17623 2283 17631 2303
rect 17651 2283 17660 2303
rect 17472 2272 17508 2273
rect 17320 2141 17357 2142
rect 17623 2141 17660 2283
rect 17685 2303 17772 2310
rect 17685 2300 17743 2303
rect 17685 2280 17690 2300
rect 17711 2283 17743 2300
rect 17763 2283 17772 2303
rect 17711 2280 17772 2283
rect 17685 2273 17772 2280
rect 17831 2303 17868 2313
rect 17831 2283 17839 2303
rect 17859 2283 17868 2303
rect 17685 2272 17716 2273
rect 17831 2204 17868 2283
rect 17898 2312 17929 2365
rect 17948 2312 17985 2313
rect 17898 2303 17985 2312
rect 17898 2283 17956 2303
rect 17976 2283 17985 2303
rect 17898 2273 17985 2283
rect 18044 2303 18081 2313
rect 18044 2283 18052 2303
rect 18072 2283 18081 2303
rect 17898 2272 17929 2273
rect 17893 2204 18003 2217
rect 18044 2204 18081 2283
rect 18125 2283 18171 2366
rect 18465 2283 18540 2567
rect 19582 2492 19652 2700
rect 19714 2707 20917 2742
rect 19714 2693 19742 2707
rect 19716 2562 19742 2693
rect 20121 2704 20917 2707
rect 19574 2441 19654 2492
rect 19574 2415 19590 2441
rect 19630 2415 19654 2441
rect 19574 2396 19654 2415
rect 19574 2370 19593 2396
rect 19633 2370 19654 2396
rect 19574 2343 19654 2370
rect 19574 2317 19597 2343
rect 19637 2317 19654 2343
rect 19574 2306 19654 2317
rect 19716 2307 19743 2562
rect 20121 2554 20162 2704
rect 20393 2698 20497 2704
rect 20853 2701 20917 2704
rect 20588 2642 20709 2660
rect 20588 2640 20659 2642
rect 20588 2599 20603 2640
rect 20640 2601 20659 2640
rect 20696 2601 20709 2642
rect 20640 2599 20709 2601
rect 20588 2589 20709 2599
rect 19783 2447 19847 2459
rect 20123 2455 20160 2554
rect 20388 2544 20499 2557
rect 20388 2542 20430 2544
rect 20388 2522 20395 2542
rect 20414 2522 20430 2542
rect 20388 2514 20430 2522
rect 20458 2542 20499 2544
rect 20458 2522 20472 2542
rect 20491 2522 20499 2542
rect 20458 2514 20499 2522
rect 20388 2508 20499 2514
rect 20331 2486 20580 2508
rect 20331 2455 20368 2486
rect 20544 2484 20580 2486
rect 20544 2455 20581 2484
rect 19783 2446 19818 2447
rect 19760 2441 19818 2446
rect 19760 2421 19763 2441
rect 19783 2427 19818 2441
rect 19838 2427 19847 2447
rect 19783 2419 19847 2427
rect 19809 2418 19847 2419
rect 19810 2417 19847 2418
rect 19913 2451 19949 2452
rect 20021 2451 20057 2452
rect 19913 2443 20057 2451
rect 19913 2423 19921 2443
rect 19941 2423 20029 2443
rect 20049 2423 20057 2443
rect 19913 2417 20057 2423
rect 20123 2447 20161 2455
rect 20229 2451 20265 2452
rect 20123 2427 20132 2447
rect 20152 2427 20161 2447
rect 20123 2418 20161 2427
rect 20180 2444 20265 2451
rect 20180 2424 20187 2444
rect 20208 2443 20265 2444
rect 20208 2424 20237 2443
rect 20180 2423 20237 2424
rect 20257 2423 20265 2443
rect 20123 2417 20160 2418
rect 20180 2417 20265 2423
rect 20331 2447 20369 2455
rect 20442 2451 20478 2452
rect 20331 2427 20340 2447
rect 20360 2427 20369 2447
rect 20331 2418 20369 2427
rect 20393 2443 20478 2451
rect 20393 2423 20450 2443
rect 20470 2423 20478 2443
rect 20331 2417 20368 2418
rect 20393 2417 20478 2423
rect 20544 2447 20582 2455
rect 20544 2427 20553 2447
rect 20573 2427 20582 2447
rect 20637 2437 20702 2589
rect 20855 2563 20910 2701
rect 20544 2418 20582 2427
rect 20635 2430 20702 2437
rect 20544 2417 20581 2418
rect 19967 2396 20003 2417
rect 20393 2396 20424 2417
rect 20635 2409 20652 2430
rect 20688 2409 20702 2430
rect 20854 2450 20910 2563
rect 20854 2432 20873 2450
rect 20891 2432 20910 2450
rect 20854 2412 20910 2432
rect 20635 2396 20702 2409
rect 19800 2392 19900 2396
rect 19800 2388 19862 2392
rect 19800 2362 19807 2388
rect 19833 2366 19862 2388
rect 19888 2366 19900 2392
rect 19833 2362 19900 2366
rect 19800 2359 19900 2362
rect 19968 2359 20003 2396
rect 20065 2393 20424 2396
rect 20065 2388 20287 2393
rect 20065 2364 20078 2388
rect 20102 2369 20287 2388
rect 20311 2369 20424 2393
rect 20102 2364 20424 2369
rect 20065 2360 20424 2364
rect 20491 2390 20702 2396
rect 20491 2388 20652 2390
rect 20491 2368 20502 2388
rect 20522 2368 20652 2388
rect 20491 2361 20652 2368
rect 20491 2360 20532 2361
rect 19967 2334 20003 2359
rect 19815 2307 19852 2308
rect 19911 2307 19948 2308
rect 19967 2307 19974 2334
rect 18125 2248 18540 2283
rect 19715 2298 19853 2307
rect 19715 2278 19824 2298
rect 19844 2278 19853 2298
rect 19715 2271 19853 2278
rect 19911 2304 19974 2307
rect 19995 2307 20003 2334
rect 20022 2307 20059 2308
rect 19995 2304 20059 2307
rect 19911 2298 20059 2304
rect 19911 2278 19920 2298
rect 19940 2278 20030 2298
rect 20050 2278 20059 2298
rect 19715 2269 19811 2271
rect 19911 2268 20059 2278
rect 20118 2298 20155 2308
rect 20230 2307 20267 2308
rect 20211 2305 20267 2307
rect 20118 2278 20126 2298
rect 20146 2278 20155 2298
rect 19967 2267 20003 2268
rect 18125 2247 18171 2248
rect 17831 2202 18081 2204
rect 17831 2199 17932 2202
rect 17831 2180 17896 2199
rect 17893 2172 17896 2180
rect 17925 2172 17932 2199
rect 17960 2175 17970 2202
rect 17999 2180 18081 2202
rect 18465 2196 18540 2248
rect 17999 2175 18003 2180
rect 17960 2172 18003 2175
rect 17893 2158 18003 2172
rect 17319 2140 17660 2141
rect 17244 2135 17660 2140
rect 17244 2115 17247 2135
rect 17267 2115 17661 2135
rect 13724 1706 16792 1731
rect 13724 1641 16587 1706
rect 16718 1641 16792 1706
rect 13724 1624 16792 1641
rect 17618 1611 17661 2115
rect 18278 2026 18373 2046
rect 18278 1982 18298 2026
rect 18358 1982 18373 2026
rect 18278 1686 18373 1982
rect 18278 1645 18311 1686
rect 18347 1645 18373 1686
rect 18473 1725 18535 2196
rect 19815 2136 19852 2137
rect 20118 2136 20155 2278
rect 20180 2298 20267 2305
rect 20180 2295 20238 2298
rect 20180 2275 20185 2295
rect 20206 2278 20238 2295
rect 20258 2278 20267 2298
rect 20206 2275 20267 2278
rect 20180 2268 20267 2275
rect 20326 2298 20363 2308
rect 20326 2278 20334 2298
rect 20354 2278 20363 2298
rect 20180 2267 20211 2268
rect 20326 2199 20363 2278
rect 20393 2307 20424 2360
rect 20637 2353 20652 2361
rect 20692 2353 20702 2390
rect 20637 2344 20702 2353
rect 20850 2351 20915 2372
rect 20850 2333 20875 2351
rect 20893 2333 20915 2351
rect 20443 2307 20480 2308
rect 20393 2298 20480 2307
rect 20393 2278 20451 2298
rect 20471 2278 20480 2298
rect 20393 2268 20480 2278
rect 20539 2298 20576 2308
rect 20539 2278 20547 2298
rect 20567 2278 20576 2298
rect 20393 2267 20424 2268
rect 20388 2199 20498 2212
rect 20539 2199 20576 2278
rect 20850 2257 20915 2333
rect 20326 2197 20576 2199
rect 20326 2194 20427 2197
rect 20326 2175 20391 2194
rect 20388 2167 20391 2175
rect 20420 2167 20427 2194
rect 20455 2170 20465 2197
rect 20494 2175 20576 2197
rect 20599 2222 20916 2257
rect 20494 2170 20498 2175
rect 20455 2167 20498 2170
rect 20388 2153 20498 2167
rect 19814 2135 20155 2136
rect 19739 2133 20155 2135
rect 20599 2133 20639 2222
rect 20850 2195 20915 2222
rect 20850 2177 20873 2195
rect 20891 2177 20915 2195
rect 20850 2157 20915 2177
rect 19736 2130 20639 2133
rect 19736 2110 19742 2130
rect 19762 2110 20639 2130
rect 19736 2106 20639 2110
rect 20599 2103 20639 2106
rect 20851 2096 20916 2117
rect 19069 2088 19730 2089
rect 19069 2081 20003 2088
rect 19069 2080 19975 2081
rect 19069 2060 19920 2080
rect 19952 2061 19975 2080
rect 20000 2061 20003 2081
rect 19952 2060 20003 2061
rect 19069 2053 20003 2060
rect 18668 2011 18836 2012
rect 19071 2011 19110 2053
rect 19899 2051 20003 2053
rect 19968 2049 20003 2051
rect 20851 2078 20875 2096
rect 20893 2078 20916 2096
rect 20851 2031 20916 2078
rect 18668 1985 19112 2011
rect 18668 1983 18836 1985
rect 18473 1706 18537 1725
rect 18473 1667 18490 1706
rect 18524 1667 18537 1706
rect 18473 1648 18537 1667
rect 18278 1619 18373 1645
rect 18668 1632 18695 1983
rect 19071 1979 19112 1985
rect 18735 1772 18799 1784
rect 19075 1780 19112 1979
rect 19574 2006 19646 2023
rect 19574 1967 19582 2006
rect 19627 1967 19646 2006
rect 19340 1869 19451 1884
rect 19340 1867 19382 1869
rect 19340 1847 19347 1867
rect 19366 1847 19382 1867
rect 19340 1839 19382 1847
rect 19410 1867 19451 1869
rect 19410 1847 19424 1867
rect 19443 1847 19451 1867
rect 19410 1839 19451 1847
rect 19340 1833 19451 1839
rect 19283 1811 19532 1833
rect 19283 1780 19320 1811
rect 19496 1809 19532 1811
rect 19496 1780 19533 1809
rect 18735 1771 18770 1772
rect 18712 1766 18770 1771
rect 18712 1746 18715 1766
rect 18735 1752 18770 1766
rect 18790 1752 18799 1772
rect 18735 1744 18799 1752
rect 18761 1743 18799 1744
rect 18762 1742 18799 1743
rect 18865 1776 18901 1777
rect 18973 1776 19009 1777
rect 18865 1768 19009 1776
rect 18865 1748 18873 1768
rect 18893 1748 18981 1768
rect 19001 1748 19009 1768
rect 18865 1742 19009 1748
rect 19075 1772 19113 1780
rect 19181 1776 19217 1777
rect 19075 1752 19084 1772
rect 19104 1752 19113 1772
rect 19075 1743 19113 1752
rect 19132 1769 19217 1776
rect 19132 1749 19139 1769
rect 19160 1768 19217 1769
rect 19160 1749 19189 1768
rect 19132 1748 19189 1749
rect 19209 1748 19217 1768
rect 19075 1742 19112 1743
rect 19132 1742 19217 1748
rect 19283 1772 19321 1780
rect 19394 1776 19430 1777
rect 19283 1752 19292 1772
rect 19312 1752 19321 1772
rect 19283 1743 19321 1752
rect 19345 1768 19430 1776
rect 19345 1748 19402 1768
rect 19422 1748 19430 1768
rect 19283 1742 19320 1743
rect 19345 1742 19430 1748
rect 19496 1772 19534 1780
rect 19496 1752 19505 1772
rect 19525 1752 19534 1772
rect 19496 1743 19534 1752
rect 19574 1757 19646 1967
rect 19716 2001 20916 2031
rect 19716 2000 20160 2001
rect 19716 1998 19884 2000
rect 19574 1743 19657 1757
rect 19496 1742 19533 1743
rect 18919 1721 18955 1742
rect 19345 1721 19376 1742
rect 19574 1721 19591 1743
rect 18752 1717 18852 1721
rect 18752 1713 18814 1717
rect 18752 1687 18759 1713
rect 18785 1691 18814 1713
rect 18840 1691 18852 1717
rect 18785 1687 18852 1691
rect 18752 1684 18852 1687
rect 18920 1684 18955 1721
rect 19017 1718 19376 1721
rect 19017 1713 19239 1718
rect 19017 1689 19030 1713
rect 19054 1694 19239 1713
rect 19263 1694 19376 1718
rect 19054 1689 19376 1694
rect 19017 1685 19376 1689
rect 19443 1713 19591 1721
rect 19443 1693 19454 1713
rect 19474 1710 19591 1713
rect 19644 1710 19657 1743
rect 19474 1693 19657 1710
rect 19443 1686 19657 1693
rect 19443 1685 19484 1686
rect 19574 1685 19657 1686
rect 18919 1659 18955 1684
rect 18767 1632 18804 1633
rect 18863 1632 18900 1633
rect 18919 1632 18926 1659
rect 18667 1623 18805 1632
rect 13479 1525 13636 1538
rect 13479 1521 13640 1525
rect 12359 1375 12385 1480
rect 13479 1414 13520 1521
rect 13620 1414 13640 1521
rect 13479 1385 13640 1414
rect 17616 1402 17665 1611
rect 18667 1603 18776 1623
rect 18796 1603 18805 1623
rect 18667 1596 18805 1603
rect 18863 1629 18926 1632
rect 18947 1632 18955 1659
rect 18974 1632 19011 1633
rect 18947 1629 19011 1632
rect 18863 1623 19011 1629
rect 18863 1603 18872 1623
rect 18892 1603 18982 1623
rect 19002 1603 19011 1623
rect 18667 1594 18763 1596
rect 18863 1593 19011 1603
rect 19070 1623 19107 1633
rect 19182 1632 19219 1633
rect 19163 1630 19219 1632
rect 19070 1603 19078 1623
rect 19098 1603 19107 1623
rect 18919 1592 18955 1593
rect 18767 1461 18804 1462
rect 19070 1461 19107 1603
rect 19132 1623 19219 1630
rect 19132 1620 19190 1623
rect 19132 1600 19137 1620
rect 19158 1603 19190 1620
rect 19210 1603 19219 1623
rect 19158 1600 19219 1603
rect 19132 1593 19219 1600
rect 19278 1623 19315 1633
rect 19278 1603 19286 1623
rect 19306 1603 19315 1623
rect 19132 1592 19163 1593
rect 19278 1524 19315 1603
rect 19345 1632 19376 1685
rect 19582 1652 19596 1685
rect 19649 1652 19657 1685
rect 19582 1646 19657 1652
rect 19582 1641 19652 1646
rect 19395 1632 19432 1633
rect 19345 1623 19432 1632
rect 19345 1603 19403 1623
rect 19423 1603 19432 1623
rect 19345 1593 19432 1603
rect 19491 1623 19528 1633
rect 19716 1628 19743 1998
rect 19783 1768 19847 1780
rect 20123 1776 20160 2000
rect 20631 1981 20695 1983
rect 20627 1969 20695 1981
rect 20627 1936 20638 1969
rect 20678 1936 20695 1969
rect 20627 1926 20695 1936
rect 20388 1865 20499 1880
rect 20388 1863 20430 1865
rect 20388 1843 20395 1863
rect 20414 1843 20430 1863
rect 20388 1835 20430 1843
rect 20458 1863 20499 1865
rect 20458 1843 20472 1863
rect 20491 1843 20499 1863
rect 20458 1835 20499 1843
rect 20388 1829 20499 1835
rect 20331 1807 20580 1829
rect 20331 1776 20368 1807
rect 20544 1805 20580 1807
rect 20544 1776 20581 1805
rect 19783 1767 19818 1768
rect 19760 1762 19818 1767
rect 19760 1742 19763 1762
rect 19783 1748 19818 1762
rect 19838 1748 19847 1768
rect 19783 1740 19847 1748
rect 19809 1739 19847 1740
rect 19810 1738 19847 1739
rect 19913 1772 19949 1773
rect 20021 1772 20057 1773
rect 19913 1764 20057 1772
rect 19913 1744 19921 1764
rect 19941 1744 20029 1764
rect 20049 1744 20057 1764
rect 19913 1738 20057 1744
rect 20123 1768 20161 1776
rect 20229 1772 20265 1773
rect 20123 1748 20132 1768
rect 20152 1748 20161 1768
rect 20123 1739 20161 1748
rect 20180 1765 20265 1772
rect 20180 1745 20187 1765
rect 20208 1764 20265 1765
rect 20208 1745 20237 1764
rect 20180 1744 20237 1745
rect 20257 1744 20265 1764
rect 20123 1738 20160 1739
rect 20180 1738 20265 1744
rect 20331 1768 20369 1776
rect 20442 1772 20478 1773
rect 20331 1748 20340 1768
rect 20360 1748 20369 1768
rect 20331 1739 20369 1748
rect 20393 1764 20478 1772
rect 20393 1744 20450 1764
rect 20470 1744 20478 1764
rect 20331 1738 20368 1739
rect 20393 1738 20478 1744
rect 20544 1768 20582 1776
rect 20544 1748 20553 1768
rect 20573 1748 20582 1768
rect 20544 1739 20582 1748
rect 20631 1742 20695 1926
rect 20851 1800 20916 2001
rect 20851 1782 20873 1800
rect 20891 1782 20916 1800
rect 20851 1763 20916 1782
rect 20544 1738 20581 1739
rect 19967 1717 20003 1738
rect 20393 1717 20424 1738
rect 20631 1733 20639 1742
rect 20628 1717 20639 1733
rect 19800 1713 19900 1717
rect 19800 1709 19862 1713
rect 19800 1683 19807 1709
rect 19833 1687 19862 1709
rect 19888 1687 19900 1713
rect 19833 1683 19900 1687
rect 19800 1680 19900 1683
rect 19968 1680 20003 1717
rect 20065 1714 20424 1717
rect 20065 1709 20287 1714
rect 20065 1685 20078 1709
rect 20102 1690 20287 1709
rect 20311 1690 20424 1714
rect 20102 1685 20424 1690
rect 20065 1681 20424 1685
rect 20491 1709 20639 1717
rect 20491 1689 20502 1709
rect 20522 1700 20639 1709
rect 20688 1733 20695 1742
rect 20688 1700 20696 1733
rect 20522 1689 20696 1700
rect 20491 1682 20696 1689
rect 20491 1681 20532 1682
rect 19967 1655 20003 1680
rect 19815 1628 19852 1629
rect 19911 1628 19948 1629
rect 19967 1628 19974 1655
rect 19491 1603 19499 1623
rect 19519 1603 19528 1623
rect 19345 1592 19376 1593
rect 19340 1524 19450 1537
rect 19491 1524 19528 1603
rect 19715 1619 19853 1628
rect 19715 1599 19824 1619
rect 19844 1599 19853 1619
rect 19715 1592 19853 1599
rect 19911 1625 19974 1628
rect 19995 1628 20003 1655
rect 20022 1628 20059 1629
rect 19995 1625 20059 1628
rect 19911 1619 20059 1625
rect 19911 1599 19920 1619
rect 19940 1599 20030 1619
rect 20050 1599 20059 1619
rect 19715 1590 19811 1592
rect 19911 1589 20059 1599
rect 20118 1619 20155 1629
rect 20230 1628 20267 1629
rect 20211 1626 20267 1628
rect 20118 1599 20126 1619
rect 20146 1599 20155 1619
rect 19967 1588 20003 1589
rect 19278 1522 19528 1524
rect 19278 1519 19379 1522
rect 19278 1500 19343 1519
rect 19340 1492 19343 1500
rect 19372 1492 19379 1519
rect 19407 1495 19417 1522
rect 19446 1500 19528 1522
rect 19446 1495 19450 1500
rect 19407 1492 19450 1495
rect 19340 1478 19450 1492
rect 18766 1460 19107 1461
rect 18691 1455 19107 1460
rect 19815 1457 19852 1458
rect 20118 1457 20155 1599
rect 20180 1619 20267 1626
rect 20180 1616 20238 1619
rect 20180 1596 20185 1616
rect 20206 1599 20238 1616
rect 20258 1599 20267 1619
rect 20206 1596 20267 1599
rect 20180 1589 20267 1596
rect 20326 1619 20363 1629
rect 20326 1599 20334 1619
rect 20354 1599 20363 1619
rect 20180 1588 20211 1589
rect 20326 1520 20363 1599
rect 20393 1628 20424 1681
rect 20628 1679 20696 1682
rect 20628 1637 20640 1679
rect 20689 1637 20696 1679
rect 20443 1628 20480 1629
rect 20393 1619 20480 1628
rect 20393 1599 20451 1619
rect 20471 1599 20480 1619
rect 20393 1589 20480 1599
rect 20539 1619 20576 1629
rect 20628 1624 20696 1637
rect 20851 1701 20916 1718
rect 20851 1683 20875 1701
rect 20893 1683 20916 1701
rect 20539 1599 20547 1619
rect 20567 1599 20576 1619
rect 20393 1588 20424 1589
rect 20388 1520 20498 1533
rect 20539 1520 20576 1599
rect 20851 1544 20916 1683
rect 20851 1538 20873 1544
rect 20326 1518 20576 1520
rect 20326 1515 20427 1518
rect 20326 1496 20391 1515
rect 20388 1488 20391 1496
rect 20420 1488 20427 1515
rect 20455 1491 20465 1518
rect 20494 1496 20576 1518
rect 20605 1526 20873 1538
rect 20891 1526 20916 1544
rect 20605 1503 20916 1526
rect 20605 1502 20660 1503
rect 20494 1491 20498 1496
rect 20455 1488 20498 1491
rect 20388 1474 20498 1488
rect 19814 1456 20155 1457
rect 18691 1435 18694 1455
rect 18714 1435 19107 1455
rect 19739 1455 20155 1456
rect 20605 1455 20648 1502
rect 19739 1451 20648 1455
rect 12359 1361 12387 1375
rect 13483 1372 13640 1385
rect 17614 1400 18431 1402
rect 18864 1400 18953 1403
rect 17614 1391 18953 1400
rect 11161 1326 12387 1361
rect 17614 1353 18876 1391
rect 18901 1356 18920 1391
rect 18945 1356 18953 1391
rect 19058 1402 19103 1435
rect 19739 1431 19742 1451
rect 19762 1431 20648 1451
rect 20116 1426 20648 1431
rect 20856 1445 20915 1467
rect 20856 1427 20875 1445
rect 20893 1427 20915 1445
rect 19904 1402 20003 1404
rect 19058 1392 20003 1402
rect 19058 1366 19926 1392
rect 19059 1365 19926 1366
rect 18901 1353 18953 1356
rect 17614 1345 18953 1353
rect 19904 1354 19926 1365
rect 19951 1357 19970 1392
rect 19995 1357 20003 1392
rect 19951 1354 20003 1357
rect 19904 1346 20003 1354
rect 19930 1345 20002 1346
rect 17614 1344 18952 1345
rect 17614 1342 18431 1344
rect 18205 1338 18431 1342
rect 453 1183 10221 1256
rect 467 1168 10221 1183
rect 11161 1250 11246 1326
rect 11604 1324 11708 1326
rect 11939 1324 11980 1326
rect 20856 1250 20915 1427
rect 11161 1177 20929 1250
rect 7536 1163 7690 1168
rect 11175 1162 20929 1177
rect 18244 1157 18398 1162
rect 10117 23 11004 25
rect 10117 12 11011 23
rect 10117 -34 10139 12
rect 10215 -34 11011 12
rect 10117 -47 11011 -34
rect 10945 -195 11011 -47
rect 11586 -64 11651 -58
rect 11586 -112 11601 -64
rect 11642 -112 11651 -64
rect 11586 -132 11651 -112
rect 10945 -215 11342 -195
rect 11362 -215 11365 -195
rect 10945 -220 11365 -215
rect 10945 -221 11290 -220
rect 10945 -233 11011 -221
rect 11252 -222 11289 -221
rect 10606 -252 10716 -238
rect 10606 -255 10649 -252
rect 10606 -260 10610 -255
rect 10528 -282 10610 -260
rect 10639 -282 10649 -255
rect 10677 -279 10684 -252
rect 10713 -260 10716 -252
rect 10713 -279 10778 -260
rect 10677 -282 10778 -279
rect 10528 -284 10778 -282
rect 10528 -363 10565 -284
rect 10606 -297 10716 -284
rect 10680 -353 10711 -352
rect 10528 -383 10537 -363
rect 10557 -383 10565 -363
rect 10528 -393 10565 -383
rect 10624 -363 10711 -353
rect 10624 -383 10633 -363
rect 10653 -383 10711 -363
rect 10624 -392 10711 -383
rect 10624 -393 10661 -392
rect 10089 -430 10218 -423
rect 10089 -489 10113 -430
rect 10144 -489 10175 -430
rect 10206 -445 10218 -430
rect 10680 -445 10711 -392
rect 10741 -363 10778 -284
rect 10893 -353 10924 -352
rect 10741 -383 10750 -363
rect 10770 -383 10778 -363
rect 10741 -393 10778 -383
rect 10837 -360 10924 -353
rect 10837 -363 10898 -360
rect 10837 -383 10846 -363
rect 10866 -380 10898 -363
rect 10919 -380 10924 -360
rect 10866 -383 10924 -380
rect 10837 -390 10924 -383
rect 10949 -363 10986 -233
rect 11101 -353 11137 -352
rect 10949 -383 10958 -363
rect 10978 -383 10986 -363
rect 10837 -392 10893 -390
rect 10837 -393 10874 -392
rect 10949 -393 10986 -383
rect 11045 -363 11193 -353
rect 11293 -356 11389 -354
rect 11045 -383 11054 -363
rect 11074 -383 11164 -363
rect 11184 -383 11193 -363
rect 11045 -389 11193 -383
rect 11045 -392 11109 -389
rect 11045 -393 11082 -392
rect 11101 -419 11109 -392
rect 11130 -392 11193 -389
rect 11251 -363 11389 -356
rect 11251 -383 11260 -363
rect 11280 -383 11389 -363
rect 11251 -392 11389 -383
rect 11130 -419 11137 -392
rect 11156 -393 11193 -392
rect 11252 -393 11289 -392
rect 11101 -444 11137 -419
rect 10206 -446 10503 -445
rect 10572 -446 10613 -445
rect 10206 -453 10613 -446
rect 10206 -473 10582 -453
rect 10602 -473 10613 -453
rect 10206 -481 10613 -473
rect 10680 -449 11039 -445
rect 10680 -454 11002 -449
rect 10680 -478 10793 -454
rect 10817 -473 11002 -454
rect 11026 -473 11039 -449
rect 10817 -478 11039 -473
rect 10680 -481 11039 -478
rect 11101 -481 11136 -444
rect 11204 -447 11304 -444
rect 11204 -451 11271 -447
rect 11204 -477 11216 -451
rect 11242 -473 11271 -451
rect 11297 -473 11304 -447
rect 11242 -477 11304 -473
rect 11204 -481 11304 -477
rect 10206 -489 10503 -481
rect 10089 -502 10218 -489
rect 10680 -502 10711 -481
rect 11101 -502 11137 -481
rect 10523 -503 10560 -502
rect 10522 -512 10560 -503
rect 10522 -532 10531 -512
rect 10551 -532 10560 -512
rect 10522 -540 10560 -532
rect 10626 -508 10711 -502
rect 10736 -503 10773 -502
rect 10626 -528 10634 -508
rect 10654 -528 10711 -508
rect 10626 -536 10711 -528
rect 10735 -512 10773 -503
rect 10735 -532 10744 -512
rect 10764 -532 10773 -512
rect 10626 -537 10662 -536
rect 10735 -540 10773 -532
rect 10839 -508 10924 -502
rect 10944 -503 10981 -502
rect 10839 -528 10847 -508
rect 10867 -509 10924 -508
rect 10867 -528 10896 -509
rect 10839 -529 10896 -528
rect 10917 -529 10924 -509
rect 10839 -536 10924 -529
rect 10943 -512 10981 -503
rect 10943 -532 10952 -512
rect 10972 -532 10981 -512
rect 10839 -537 10875 -536
rect 10943 -540 10981 -532
rect 11047 -508 11191 -502
rect 11047 -528 11055 -508
rect 11075 -528 11110 -508
rect 11047 -531 11110 -528
rect 11130 -528 11163 -508
rect 11183 -528 11191 -508
rect 11130 -531 11191 -528
rect 11047 -536 11191 -531
rect 11047 -537 11083 -536
rect 11155 -537 11191 -536
rect 11257 -503 11294 -502
rect 11257 -504 11295 -503
rect 11257 -512 11321 -504
rect 11257 -532 11266 -512
rect 11286 -526 11321 -512
rect 11341 -526 11344 -506
rect 11286 -531 11344 -526
rect 11286 -532 11321 -531
rect 10523 -569 10560 -540
rect 10524 -571 10560 -569
rect 10736 -571 10773 -540
rect 10524 -593 10773 -571
rect 10605 -599 10716 -593
rect 10605 -607 10646 -599
rect 10605 -627 10613 -607
rect 10632 -627 10646 -607
rect 10605 -629 10646 -627
rect 10674 -607 10716 -599
rect 10674 -627 10690 -607
rect 10709 -627 10716 -607
rect 10674 -629 10716 -627
rect 10605 -644 10716 -629
rect 10944 -661 10981 -540
rect 11257 -544 11321 -532
rect 11361 -654 11388 -392
rect 11586 -654 11634 -132
rect 11339 -659 11634 -654
rect 11220 -661 11634 -659
rect 10944 -687 11634 -661
rect 11220 -688 11634 -687
rect 11339 -689 11634 -688
rect 11586 -694 11634 -689
<< viali >>
rect 2869 13645 2906 13693
rect 1399 13104 1424 13139
rect 1443 13104 1468 13142
rect 1632 13045 1652 13065
rect 2449 13105 2474 13140
rect 2493 13105 2518 13143
rect 2680 13041 2700 13061
rect 900 12978 929 13005
rect 974 12981 1003 13008
rect 705 12817 754 12859
rect 1188 12880 1209 12900
rect 1948 12974 1977 13001
rect 2022 12977 2051 13004
rect 1399 12841 1420 12871
rect 706 12754 755 12796
rect 1561 12787 1587 12813
rect 1186 12731 1207 12751
rect 1611 12734 1631 12754
rect 903 12633 922 12653
rect 980 12633 999 12653
rect 716 12527 756 12560
rect 1745 12811 1798 12844
rect 2236 12876 2257 12896
rect 2447 12837 2468 12867
rect 1750 12753 1803 12786
rect 2609 12783 2635 12809
rect 2234 12727 2255 12747
rect 2659 12730 2679 12750
rect 1951 12629 1970 12649
rect 2028 12629 2047 12649
rect 1767 12490 1812 12529
rect 2870 12790 2904 12829
rect 1394 12415 1419 12435
rect 1442 12416 1474 12436
rect 1632 12366 1652 12386
rect 900 12299 929 12326
rect 974 12302 1003 12329
rect 702 12106 742 12143
rect 1188 12201 1209 12221
rect 3047 12810 3083 12851
rect 3036 12470 3096 12514
rect 4842 12917 4928 12984
rect 8883 12843 8923 12869
rect 8886 12798 8926 12824
rect 4127 12361 4147 12381
rect 3395 12294 3424 12321
rect 3469 12297 3498 12324
rect 1399 12162 1420 12192
rect 1561 12108 1587 12134
rect 706 12066 742 12087
rect 1186 12052 1207 12072
rect 1611 12055 1631 12075
rect 903 11954 922 11974
rect 980 11954 999 11974
rect 698 11854 735 11895
rect 754 11856 791 11897
rect 1757 12153 1797 12179
rect 1761 12100 1801 12126
rect 1764 12055 1804 12081
rect 3683 12196 3704 12216
rect 3894 12157 3915 12187
rect 3036 12056 3090 12097
rect 4056 12103 4082 12129
rect 3681 12047 3702 12067
rect 1763 11730 1793 11796
rect 1399 11657 1424 11692
rect 1443 11657 1468 11695
rect 1632 11598 1652 11618
rect 2680 11594 2700 11614
rect 900 11531 929 11558
rect 974 11534 1003 11561
rect 705 11370 754 11412
rect 1188 11433 1209 11453
rect 1948 11527 1977 11554
rect 2022 11530 2051 11557
rect 1399 11394 1420 11424
rect 706 11307 755 11349
rect 1561 11340 1587 11366
rect 1186 11284 1207 11304
rect 1611 11287 1631 11307
rect 903 11186 922 11206
rect 980 11186 999 11206
rect 716 11080 756 11113
rect 1745 11364 1798 11397
rect 2236 11429 2257 11449
rect 2447 11390 2468 11420
rect 1750 11306 1803 11339
rect 2609 11336 2635 11362
rect 2234 11280 2255 11300
rect 2659 11283 2679 11303
rect 1951 11182 1970 11202
rect 2028 11182 2047 11202
rect 1767 11043 1812 11082
rect 3398 11949 3417 11969
rect 3475 11949 3494 11969
rect 4106 12050 4126 12070
rect 3905 11859 3957 11877
rect 3674 11658 3699 11693
rect 3718 11658 3743 11696
rect 3937 11674 3961 11697
rect 3937 11630 3961 11653
rect 1394 10968 1419 10988
rect 1442 10969 1474 10989
rect 1632 10919 1652 10939
rect 900 10852 929 10879
rect 974 10855 1003 10882
rect 702 10659 742 10696
rect 1188 10754 1209 10774
rect 1399 10715 1420 10745
rect 1561 10661 1587 10687
rect 706 10619 742 10640
rect 1186 10605 1207 10625
rect 1611 10608 1631 10628
rect 903 10507 922 10527
rect 980 10507 999 10527
rect 698 10407 735 10448
rect 754 10409 791 10450
rect 1757 10706 1797 10732
rect 1761 10653 1801 10679
rect 1764 10608 1804 10634
rect 1756 10348 1800 10385
rect 3942 11011 3962 11032
rect 3983 11016 4003 11037
rect 4170 10916 4190 10936
rect 3438 10849 3467 10876
rect 3512 10852 3541 10879
rect 3726 10751 3747 10771
rect 3937 10712 3958 10742
rect 4099 10658 4125 10684
rect 1751 10262 1805 10328
rect 1400 10137 1425 10172
rect 1444 10137 1469 10175
rect 1633 10078 1653 10098
rect 2681 10074 2701 10094
rect 901 10011 930 10038
rect 975 10014 1004 10041
rect 706 9850 755 9892
rect 1189 9913 1210 9933
rect 1949 10007 1978 10034
rect 2023 10010 2052 10037
rect 1400 9874 1421 9904
rect 707 9787 756 9829
rect 1562 9820 1588 9846
rect 1187 9764 1208 9784
rect 1612 9767 1632 9787
rect 904 9666 923 9686
rect 981 9666 1000 9686
rect 717 9560 757 9593
rect 1746 9844 1799 9877
rect 2237 9909 2258 9929
rect 2448 9870 2469 9900
rect 1751 9786 1804 9819
rect 2610 9816 2636 9842
rect 2235 9760 2256 9780
rect 2660 9763 2680 9783
rect 1952 9662 1971 9682
rect 2029 9662 2048 9682
rect 1768 9523 1813 9562
rect 1395 9448 1420 9468
rect 1443 9449 1475 9469
rect 1633 9399 1653 9419
rect 901 9332 930 9359
rect 975 9335 1004 9362
rect 703 9139 743 9176
rect 1189 9234 1210 9254
rect 1400 9195 1421 9225
rect 1562 9141 1588 9167
rect 707 9099 743 9120
rect 1187 9085 1208 9105
rect 1612 9088 1632 9108
rect 904 8987 923 9007
rect 981 8987 1000 9007
rect 699 8887 736 8928
rect 755 8889 792 8930
rect 1758 9186 1798 9212
rect 1762 9133 1802 9159
rect 1765 9088 1805 9114
rect 2872 9129 2898 9152
rect 1764 8763 1794 8829
rect 1400 8690 1425 8725
rect 1444 8690 1469 8728
rect 1633 8631 1653 8651
rect 2681 8627 2701 8647
rect 901 8564 930 8591
rect 975 8567 1004 8594
rect 706 8403 755 8445
rect 1189 8466 1210 8486
rect 1949 8560 1978 8587
rect 2023 8563 2052 8590
rect 1400 8427 1421 8457
rect 707 8340 756 8382
rect 1562 8373 1588 8399
rect 1187 8317 1208 8337
rect 1612 8320 1632 8340
rect 904 8219 923 8239
rect 981 8219 1000 8239
rect 717 8113 757 8146
rect 1746 8397 1799 8430
rect 2237 8462 2258 8482
rect 2448 8423 2469 8453
rect 1751 8339 1804 8372
rect 2610 8369 2636 8395
rect 2235 8313 2256 8333
rect 2660 8316 2680 8336
rect 1952 8215 1971 8235
rect 2029 8215 2048 8235
rect 1768 8076 1813 8115
rect 1395 8001 1420 8021
rect 1443 8002 1475 8022
rect 1633 7952 1653 7972
rect 901 7885 930 7912
rect 975 7888 1004 7915
rect 703 7692 743 7729
rect 1189 7787 1210 7807
rect 1400 7748 1421 7778
rect 1562 7694 1588 7720
rect 707 7652 743 7673
rect 1187 7638 1208 7658
rect 1612 7641 1632 7661
rect 904 7540 923 7560
rect 981 7540 1000 7560
rect 699 7440 736 7481
rect 755 7442 792 7483
rect 1758 7739 1798 7765
rect 1762 7686 1802 7712
rect 1765 7641 1805 7667
rect 1756 7320 1802 7368
rect 3724 10602 3745 10622
rect 4149 10605 4169 10625
rect 3441 10504 3460 10524
rect 3518 10504 3537 10524
rect 3741 10138 3766 10176
rect 3899 9447 3916 9484
rect 4128 9394 4148 9414
rect 3396 9327 3425 9354
rect 3470 9330 3499 9357
rect 3684 9229 3705 9249
rect 3895 9190 3916 9220
rect 3252 9122 3278 9145
rect 4057 9136 4083 9162
rect 3682 9080 3703 9100
rect 4107 9083 4127 9103
rect 3399 8982 3418 9002
rect 3476 8982 3495 9002
rect 3739 8710 3767 8738
rect 5236 7943 5256 7963
rect 4504 7876 4533 7903
rect 4578 7879 4607 7906
rect 4792 7778 4813 7798
rect 5003 7739 5024 7769
rect 4300 7680 4324 7704
rect 4357 7681 4381 7705
rect 5165 7685 5191 7711
rect 4790 7629 4811 7649
rect 5003 7627 5027 7649
rect 5215 7632 5235 7652
rect 4507 7531 4526 7551
rect 4584 7531 4603 7551
rect 8890 12745 8930 12771
rect 9896 13027 9933 13068
rect 9952 13029 9989 13070
rect 9688 12950 9707 12970
rect 9765 12950 9784 12970
rect 9056 12849 9076 12869
rect 9480 12852 9501 12872
rect 12107 13098 12132 13133
rect 12151 13098 12176 13136
rect 12340 13039 12360 13059
rect 13157 13099 13182 13134
rect 13201 13099 13226 13137
rect 9945 12837 9981 12858
rect 13388 13035 13408 13055
rect 11608 12972 11637 12999
rect 11682 12975 11711 13002
rect 9100 12790 9126 12816
rect 9267 12732 9288 12762
rect 9478 12703 9499 12723
rect 9945 12781 9985 12818
rect 11413 12811 11462 12853
rect 11896 12874 11917 12894
rect 12656 12968 12685 12995
rect 12730 12971 12759 12998
rect 12107 12835 12128 12865
rect 11414 12748 11463 12790
rect 12269 12781 12295 12807
rect 9684 12595 9713 12622
rect 9758 12598 9787 12625
rect 9035 12538 9055 12558
rect 9213 12488 9245 12508
rect 9268 12489 9293 12509
rect 8875 12395 8920 12434
rect 8640 12275 8659 12295
rect 8717 12275 8736 12295
rect 8008 12174 8028 12194
rect 8432 12177 8453 12197
rect 8052 12115 8078 12141
rect 8884 12138 8937 12171
rect 8219 12057 8240 12087
rect 8430 12028 8451 12048
rect 8889 12080 8942 12113
rect 9931 12364 9971 12397
rect 9688 12271 9707 12291
rect 9765 12271 9784 12291
rect 9056 12170 9076 12190
rect 9480 12173 9501 12193
rect 11894 12725 11915 12745
rect 12319 12728 12339 12748
rect 11611 12627 11630 12647
rect 11688 12627 11707 12647
rect 11424 12521 11464 12554
rect 12453 12805 12506 12838
rect 12944 12870 12965 12890
rect 13155 12831 13176 12861
rect 12458 12747 12511 12780
rect 13317 12777 13343 12803
rect 12942 12721 12963 12741
rect 13367 12724 13387 12744
rect 12659 12623 12678 12643
rect 12736 12623 12755 12643
rect 12475 12484 12520 12523
rect 13578 12784 13612 12823
rect 12102 12409 12127 12429
rect 12150 12410 12182 12430
rect 12340 12360 12360 12380
rect 11608 12293 11637 12320
rect 11682 12296 11711 12323
rect 9100 12111 9126 12137
rect 9932 12128 9981 12170
rect 9267 12053 9288 12083
rect 8636 11920 8665 11947
rect 8710 11923 8739 11950
rect 9478 12024 9499 12044
rect 9933 12065 9982 12107
rect 11410 12100 11450 12137
rect 11896 12195 11917 12215
rect 13755 12804 13791 12845
rect 13744 12464 13804 12508
rect 15056 12906 15094 13003
rect 15116 12912 15154 13009
rect 19591 12837 19631 12863
rect 14835 12355 14855 12375
rect 14103 12288 14132 12315
rect 14177 12291 14206 12318
rect 12107 12156 12128 12186
rect 12269 12102 12295 12128
rect 9684 11916 9713 11943
rect 9758 11919 9787 11946
rect 7987 11863 8007 11883
rect 11414 12060 11450 12081
rect 9035 11859 9055 11879
rect 6921 11772 6949 11800
rect 9219 11782 9244 11820
rect 9263 11785 9288 11820
rect 11894 12046 11915 12066
rect 12319 12049 12339 12069
rect 11611 11948 11630 11968
rect 11688 11948 11707 11968
rect 11406 11848 11443 11889
rect 11462 11850 11499 11891
rect 12465 12147 12505 12173
rect 12469 12094 12509 12120
rect 12472 12049 12512 12075
rect 8894 11681 8924 11747
rect 7193 11508 7212 11528
rect 7270 11508 7289 11528
rect 14391 12190 14412 12210
rect 14602 12151 14623 12181
rect 13744 12050 13798 12091
rect 14764 12097 14790 12123
rect 14389 12041 14410 12061
rect 12471 11724 12501 11790
rect 6561 11407 6581 11427
rect 6985 11410 7006 11430
rect 6605 11348 6631 11374
rect 7410 11365 7436 11388
rect 7790 11358 7816 11381
rect 6772 11290 6793 11320
rect 6983 11261 7004 11281
rect 8883 11396 8923 11422
rect 8886 11351 8926 11377
rect 8890 11298 8930 11324
rect 7189 11153 7218 11180
rect 7263 11156 7292 11183
rect 6540 11096 6560 11116
rect 6772 11026 6789 11063
rect 9896 11580 9933 11621
rect 9952 11582 9989 11623
rect 9688 11503 9707 11523
rect 9765 11503 9784 11523
rect 9056 11402 9076 11422
rect 9480 11405 9501 11425
rect 12107 11651 12132 11686
rect 12151 11651 12176 11689
rect 12340 11592 12360 11612
rect 9945 11390 9981 11411
rect 13388 11588 13408 11608
rect 11608 11525 11637 11552
rect 11682 11528 11711 11555
rect 9100 11343 9126 11369
rect 9267 11285 9288 11315
rect 9478 11256 9499 11276
rect 9945 11334 9985 11371
rect 11413 11364 11462 11406
rect 11896 11427 11917 11447
rect 12656 11521 12685 11548
rect 12730 11524 12759 11551
rect 12107 11388 12128 11418
rect 11414 11301 11463 11343
rect 12269 11334 12295 11360
rect 9684 11148 9713 11175
rect 9758 11151 9787 11178
rect 9035 11091 9055 11111
rect 9213 11041 9245 11061
rect 9268 11042 9293 11062
rect 6922 10334 6947 10372
rect 8875 10948 8920 10987
rect 8640 10828 8659 10848
rect 8717 10828 8736 10848
rect 8008 10727 8028 10747
rect 8432 10730 8453 10750
rect 8052 10668 8078 10694
rect 8884 10691 8937 10724
rect 8219 10610 8240 10640
rect 8430 10581 8451 10601
rect 8889 10633 8942 10666
rect 9931 10917 9971 10950
rect 9688 10824 9707 10844
rect 9765 10824 9784 10844
rect 9056 10723 9076 10743
rect 9480 10726 9501 10746
rect 11894 11278 11915 11298
rect 12319 11281 12339 11301
rect 11611 11180 11630 11200
rect 11688 11180 11707 11200
rect 11424 11074 11464 11107
rect 12453 11358 12506 11391
rect 12944 11423 12965 11443
rect 13155 11384 13176 11414
rect 12458 11300 12511 11333
rect 13317 11330 13343 11356
rect 12942 11274 12963 11294
rect 13367 11277 13387 11297
rect 12659 11176 12678 11196
rect 12736 11176 12755 11196
rect 12475 11037 12520 11076
rect 14106 11943 14125 11963
rect 14183 11943 14202 11963
rect 14814 12044 14834 12064
rect 14613 11853 14665 11871
rect 14382 11652 14407 11687
rect 14426 11652 14451 11690
rect 14645 11668 14669 11691
rect 14645 11624 14669 11647
rect 12102 10962 12127 10982
rect 12150 10963 12182 10983
rect 12340 10913 12360 10933
rect 11608 10846 11637 10873
rect 11682 10849 11711 10876
rect 9100 10664 9126 10690
rect 9932 10681 9981 10723
rect 9267 10606 9288 10636
rect 8636 10473 8665 10500
rect 8710 10476 8739 10503
rect 9478 10577 9499 10597
rect 9933 10618 9982 10660
rect 11410 10653 11450 10690
rect 11896 10748 11917 10768
rect 12107 10709 12128 10739
rect 12269 10655 12295 10681
rect 9684 10469 9713 10496
rect 9758 10472 9787 10499
rect 7987 10416 8007 10436
rect 11414 10613 11450 10634
rect 9035 10412 9055 10432
rect 9219 10335 9244 10373
rect 9263 10338 9288 10373
rect 11894 10599 11915 10619
rect 12319 10602 12339 10622
rect 11611 10501 11630 10521
rect 11688 10501 11707 10521
rect 11406 10401 11443 10442
rect 11462 10403 11499 10444
rect 12465 10700 12505 10726
rect 12469 10647 12509 10673
rect 12472 10602 12512 10628
rect 12464 10342 12508 10379
rect 14650 11005 14670 11026
rect 14691 11010 14711 11031
rect 14878 10910 14898 10930
rect 14146 10843 14175 10870
rect 14220 10846 14249 10873
rect 14434 10745 14455 10765
rect 14645 10706 14666 10736
rect 14807 10652 14833 10678
rect 8883 10182 8937 10248
rect 12459 10256 12513 10322
rect 7151 9986 7170 10006
rect 7228 9986 7247 10006
rect 6519 9885 6539 9905
rect 6943 9888 6964 9908
rect 6563 9826 6589 9852
rect 6730 9768 6751 9798
rect 6941 9739 6962 9759
rect 7147 9631 7176 9658
rect 7221 9634 7250 9661
rect 6498 9574 6518 9594
rect 8888 10125 8932 10162
rect 8884 9876 8924 9902
rect 8887 9831 8927 9857
rect 8891 9778 8931 9804
rect 9897 10060 9934 10101
rect 9953 10062 9990 10103
rect 9689 9983 9708 10003
rect 9766 9983 9785 10003
rect 9057 9882 9077 9902
rect 9481 9885 9502 9905
rect 12108 10131 12133 10166
rect 12152 10131 12177 10169
rect 12341 10072 12361 10092
rect 9946 9870 9982 9891
rect 13389 10068 13409 10088
rect 11609 10005 11638 10032
rect 11683 10008 11712 10035
rect 9101 9823 9127 9849
rect 9268 9765 9289 9795
rect 9479 9736 9500 9756
rect 9946 9814 9986 9851
rect 11414 9844 11463 9886
rect 11897 9907 11918 9927
rect 12657 10001 12686 10028
rect 12731 10004 12760 10031
rect 12108 9868 12129 9898
rect 11415 9781 11464 9823
rect 12270 9814 12296 9840
rect 9685 9628 9714 9655
rect 9759 9631 9788 9658
rect 9036 9571 9056 9591
rect 9214 9521 9246 9541
rect 9269 9522 9294 9542
rect 6727 8857 6751 8880
rect 6727 8813 6751 8836
rect 6945 8814 6970 8852
rect 6989 8817 7014 8852
rect 6731 8633 6783 8651
rect 6562 8440 6582 8460
rect 7194 8541 7213 8561
rect 7271 8541 7290 8561
rect 8876 9428 8921 9467
rect 8641 9308 8660 9328
rect 8718 9308 8737 9328
rect 8009 9207 8029 9227
rect 8433 9210 8454 9230
rect 8053 9148 8079 9174
rect 8885 9171 8938 9204
rect 8220 9090 8241 9120
rect 8431 9061 8452 9081
rect 8890 9113 8943 9146
rect 9932 9397 9972 9430
rect 9689 9304 9708 9324
rect 9766 9304 9785 9324
rect 9057 9203 9077 9223
rect 9481 9206 9502 9226
rect 11895 9758 11916 9778
rect 12320 9761 12340 9781
rect 11612 9660 11631 9680
rect 11689 9660 11708 9680
rect 11425 9554 11465 9587
rect 12454 9838 12507 9871
rect 12945 9903 12966 9923
rect 13156 9864 13177 9894
rect 12459 9780 12512 9813
rect 13318 9810 13344 9836
rect 12943 9754 12964 9774
rect 13368 9757 13388 9777
rect 12660 9656 12679 9676
rect 12737 9656 12756 9676
rect 12476 9517 12521 9556
rect 12103 9442 12128 9462
rect 12151 9443 12183 9463
rect 12341 9393 12361 9413
rect 11609 9326 11638 9353
rect 11683 9329 11712 9356
rect 9101 9144 9127 9170
rect 9933 9161 9982 9203
rect 9268 9086 9289 9116
rect 8637 8953 8666 8980
rect 8711 8956 8740 8983
rect 9479 9057 9500 9077
rect 9934 9098 9983 9140
rect 11411 9133 11451 9170
rect 11897 9228 11918 9248
rect 12108 9189 12129 9219
rect 12270 9135 12296 9161
rect 9685 8949 9714 8976
rect 9759 8952 9788 8979
rect 7988 8896 8008 8916
rect 11415 9093 11451 9114
rect 9036 8892 9056 8912
rect 9220 8815 9245 8853
rect 9264 8818 9289 8853
rect 11895 9079 11916 9099
rect 12320 9082 12340 9102
rect 11612 8981 11631 9001
rect 11689 8981 11708 9001
rect 11407 8881 11444 8922
rect 11463 8883 11500 8924
rect 12466 9180 12506 9206
rect 12470 9127 12510 9153
rect 12473 9082 12513 9108
rect 13580 9123 13606 9146
rect 8895 8714 8925 8780
rect 6986 8443 7007 8463
rect 6606 8381 6632 8407
rect 7598 8413 7652 8454
rect 6773 8323 6794 8353
rect 6984 8294 7005 8314
rect 12472 8757 12502 8823
rect 8884 8429 8924 8455
rect 8887 8384 8927 8410
rect 8891 8331 8931 8357
rect 9897 8613 9934 8654
rect 9953 8615 9990 8656
rect 9689 8536 9708 8556
rect 9766 8536 9785 8556
rect 9057 8435 9077 8455
rect 9481 8438 9502 8458
rect 12108 8684 12133 8719
rect 12152 8684 12177 8722
rect 12341 8625 12361 8645
rect 9946 8423 9982 8444
rect 13389 8621 13409 8641
rect 11609 8558 11638 8585
rect 11683 8561 11712 8588
rect 9101 8376 9127 8402
rect 9268 8318 9289 8348
rect 7190 8186 7219 8213
rect 7264 8189 7293 8216
rect 6541 8129 6561 8149
rect 4843 7438 4872 7472
rect 4842 7378 4871 7412
rect 3058 7293 3102 7321
rect 2867 7194 2904 7242
rect 3055 7236 3099 7264
rect 5350 7154 5413 7208
rect 1397 7096 1422 7131
rect 1441 7096 1466 7134
rect 1630 7037 1650 7057
rect 2447 7097 2472 7132
rect 2491 7097 2516 7135
rect 2678 7033 2698 7053
rect 898 6970 927 6997
rect 972 6973 1001 7000
rect 703 6809 752 6851
rect 1186 6872 1207 6892
rect 1946 6966 1975 6993
rect 2020 6969 2049 6996
rect 1397 6833 1418 6863
rect 704 6746 753 6788
rect 1559 6779 1585 6805
rect 1184 6723 1205 6743
rect 1609 6726 1629 6746
rect 901 6625 920 6645
rect 978 6625 997 6645
rect 714 6519 754 6552
rect 1743 6803 1796 6836
rect 2234 6868 2255 6888
rect 2445 6829 2466 6859
rect 1748 6745 1801 6778
rect 2607 6775 2633 6801
rect 2232 6719 2253 6739
rect 2657 6722 2677 6742
rect 1949 6621 1968 6641
rect 2026 6621 2045 6641
rect 1765 6482 1810 6521
rect 2868 6782 2902 6821
rect 1392 6407 1417 6427
rect 1440 6408 1472 6428
rect 1630 6358 1650 6378
rect 898 6291 927 6318
rect 972 6294 1001 6321
rect 700 6098 740 6135
rect 1186 6193 1207 6213
rect 3045 6802 3081 6843
rect 3034 6462 3094 6506
rect 4125 6353 4145 6373
rect 3393 6286 3422 6313
rect 3467 6289 3496 6316
rect 1397 6154 1418 6184
rect 1559 6100 1585 6126
rect 704 6058 740 6079
rect 1184 6044 1205 6064
rect 1609 6047 1629 6067
rect 901 5946 920 5966
rect 978 5946 997 5966
rect 696 5846 733 5887
rect 752 5848 789 5889
rect 1755 6145 1795 6171
rect 1759 6092 1799 6118
rect 1762 6047 1802 6073
rect 3681 6188 3702 6208
rect 3892 6149 3913 6179
rect 3034 6048 3088 6089
rect 4054 6095 4080 6121
rect 3679 6039 3700 6059
rect 1761 5722 1791 5788
rect 1397 5649 1422 5684
rect 1441 5649 1466 5687
rect 1630 5590 1650 5610
rect 2678 5586 2698 5606
rect 898 5523 927 5550
rect 972 5526 1001 5553
rect 703 5362 752 5404
rect 1186 5425 1207 5445
rect 1946 5519 1975 5546
rect 2020 5522 2049 5549
rect 1397 5386 1418 5416
rect 704 5299 753 5341
rect 1559 5332 1585 5358
rect 1184 5276 1205 5296
rect 1609 5279 1629 5299
rect 901 5178 920 5198
rect 978 5178 997 5198
rect 714 5072 754 5105
rect 1743 5356 1796 5389
rect 2234 5421 2255 5441
rect 2445 5382 2466 5412
rect 1748 5298 1801 5331
rect 2607 5328 2633 5354
rect 2232 5272 2253 5292
rect 2657 5275 2677 5295
rect 1949 5174 1968 5194
rect 2026 5174 2045 5194
rect 1765 5035 1810 5074
rect 3396 5941 3415 5961
rect 3473 5941 3492 5961
rect 4104 6042 4124 6062
rect 3903 5851 3955 5869
rect 3672 5650 3697 5685
rect 3716 5650 3741 5688
rect 3935 5666 3959 5689
rect 3935 5622 3959 5645
rect 1392 4960 1417 4980
rect 1440 4961 1472 4981
rect 1630 4911 1650 4931
rect 898 4844 927 4871
rect 972 4847 1001 4874
rect 700 4651 740 4688
rect 1186 4746 1207 4766
rect 1397 4707 1418 4737
rect 1559 4653 1585 4679
rect 704 4611 740 4632
rect 1184 4597 1205 4617
rect 1609 4600 1629 4620
rect 901 4499 920 4519
rect 978 4499 997 4519
rect 696 4399 733 4440
rect 752 4401 789 4442
rect 1755 4698 1795 4724
rect 1759 4645 1799 4671
rect 1762 4600 1802 4626
rect 1754 4340 1798 4377
rect 4168 4908 4188 4928
rect 3436 4841 3465 4868
rect 3510 4844 3539 4871
rect 3724 4743 3745 4763
rect 3935 4704 3956 4734
rect 4097 4650 4123 4676
rect 1749 4254 1803 4320
rect 1398 4129 1423 4164
rect 1442 4129 1467 4167
rect 1631 4070 1651 4090
rect 2679 4066 2699 4086
rect 899 4003 928 4030
rect 973 4006 1002 4033
rect 704 3842 753 3884
rect 1187 3905 1208 3925
rect 1947 3999 1976 4026
rect 2021 4002 2050 4029
rect 1398 3866 1419 3896
rect 705 3779 754 3821
rect 1560 3812 1586 3838
rect 1185 3756 1206 3776
rect 1610 3759 1630 3779
rect 902 3658 921 3678
rect 979 3658 998 3678
rect 715 3552 755 3585
rect 1744 3836 1797 3869
rect 2235 3901 2256 3921
rect 2446 3862 2467 3892
rect 1749 3778 1802 3811
rect 2608 3808 2634 3834
rect 2233 3752 2254 3772
rect 2658 3755 2678 3775
rect 1950 3654 1969 3674
rect 2027 3654 2046 3674
rect 1766 3515 1811 3554
rect 1393 3440 1418 3460
rect 1441 3441 1473 3461
rect 1631 3391 1651 3411
rect 899 3324 928 3351
rect 973 3327 1002 3354
rect 701 3131 741 3168
rect 1187 3226 1208 3246
rect 1398 3187 1419 3217
rect 1560 3133 1586 3159
rect 705 3091 741 3112
rect 1185 3077 1206 3097
rect 1610 3080 1630 3100
rect 902 2979 921 2999
rect 979 2979 998 2999
rect 697 2879 734 2920
rect 753 2881 790 2922
rect 1756 3178 1796 3204
rect 1760 3125 1800 3151
rect 1763 3080 1803 3106
rect 2825 3111 2850 3142
rect 2870 3121 2896 3144
rect 1762 2755 1792 2821
rect 1398 2682 1423 2717
rect 1442 2682 1467 2720
rect 1631 2623 1651 2643
rect 2679 2619 2699 2639
rect 899 2556 928 2583
rect 973 2559 1002 2586
rect 704 2395 753 2437
rect 1187 2458 1208 2478
rect 1947 2552 1976 2579
rect 2021 2555 2050 2582
rect 1398 2419 1419 2449
rect 705 2332 754 2374
rect 1560 2365 1586 2391
rect 1185 2309 1206 2329
rect 1610 2312 1630 2332
rect 902 2211 921 2231
rect 979 2211 998 2231
rect 715 2105 755 2138
rect 1744 2389 1797 2422
rect 2235 2454 2256 2474
rect 2446 2415 2467 2445
rect 1749 2331 1802 2364
rect 2608 2361 2634 2387
rect 2233 2305 2254 2325
rect 2658 2308 2678 2328
rect 1950 2207 1969 2227
rect 2027 2207 2046 2227
rect 1766 2068 1811 2107
rect 1393 1993 1418 2013
rect 1441 1994 1473 2014
rect 1631 1944 1651 1964
rect 899 1877 928 1904
rect 973 1880 1002 1907
rect 701 1684 741 1721
rect 1187 1779 1208 1799
rect 1398 1740 1419 1770
rect 1560 1686 1586 1712
rect 705 1644 741 1665
rect 1185 1630 1206 1650
rect 1610 1633 1630 1653
rect 902 1532 921 1552
rect 979 1532 998 1552
rect 697 1432 734 1473
rect 753 1434 790 1475
rect 3722 4594 3743 4614
rect 4147 4597 4167 4617
rect 3439 4496 3458 4516
rect 3516 4496 3535 4516
rect 3739 4130 3764 4168
rect 5815 7090 5844 7124
rect 5814 7030 5843 7064
rect 6083 6951 6102 6971
rect 6160 6951 6179 6971
rect 5451 6850 5471 6870
rect 5875 6853 5896 6873
rect 7592 7996 7652 8040
rect 7605 7659 7641 7700
rect 9479 8289 9500 8309
rect 9946 8367 9986 8404
rect 11414 8397 11463 8439
rect 11897 8460 11918 8480
rect 12657 8554 12686 8581
rect 12731 8557 12760 8584
rect 12108 8421 12129 8451
rect 11415 8334 11464 8376
rect 12270 8367 12296 8393
rect 9685 8181 9714 8208
rect 9759 8184 9788 8211
rect 9036 8124 9056 8144
rect 9214 8074 9246 8094
rect 9269 8075 9294 8095
rect 7784 7681 7818 7720
rect 8876 7981 8921 8020
rect 8641 7861 8660 7881
rect 8718 7861 8737 7881
rect 8009 7760 8029 7780
rect 8433 7763 8454 7783
rect 8053 7701 8079 7727
rect 8885 7724 8938 7757
rect 8220 7643 8241 7673
rect 8431 7614 8452 7634
rect 8890 7666 8943 7699
rect 9932 7950 9972 7983
rect 9689 7857 9708 7877
rect 9766 7857 9785 7877
rect 9057 7756 9077 7776
rect 9481 7759 9502 7779
rect 11895 8311 11916 8331
rect 12320 8314 12340 8334
rect 11612 8213 11631 8233
rect 11689 8213 11708 8233
rect 11425 8107 11465 8140
rect 12454 8391 12507 8424
rect 12945 8456 12966 8476
rect 13156 8417 13177 8447
rect 12459 8333 12512 8366
rect 13318 8363 13344 8389
rect 12943 8307 12964 8327
rect 13368 8310 13388 8330
rect 12660 8209 12679 8229
rect 12737 8209 12756 8229
rect 12476 8070 12521 8109
rect 12103 7995 12128 8015
rect 12151 7996 12183 8016
rect 12341 7946 12361 7966
rect 11609 7879 11638 7906
rect 11683 7882 11712 7909
rect 9101 7697 9127 7723
rect 9933 7714 9982 7756
rect 9268 7639 9289 7669
rect 8637 7506 8666 7533
rect 8711 7509 8740 7536
rect 9479 7610 9500 7630
rect 9934 7651 9983 7693
rect 11411 7686 11451 7723
rect 11897 7781 11918 7801
rect 12108 7742 12129 7772
rect 12270 7688 12296 7714
rect 9685 7502 9714 7529
rect 9759 7505 9788 7532
rect 7988 7449 8008 7469
rect 11415 7646 11451 7667
rect 8170 7367 8195 7405
rect 8214 7370 8239 7405
rect 9036 7445 9056 7465
rect 9220 7368 9245 7406
rect 9264 7371 9289 7406
rect 11895 7632 11916 7652
rect 12320 7635 12340 7655
rect 11612 7534 11631 7554
rect 11689 7534 11708 7554
rect 11407 7434 11444 7475
rect 11463 7436 11500 7477
rect 12466 7733 12506 7759
rect 12470 7680 12510 7706
rect 12473 7635 12513 7661
rect 5495 6791 5521 6817
rect 6305 6797 6329 6821
rect 6362 6798 6386 6822
rect 5662 6733 5683 6763
rect 5873 6704 5894 6724
rect 7587 7238 7631 7266
rect 7782 7260 7819 7308
rect 7584 7181 7628 7209
rect 6079 6596 6108 6623
rect 6153 6599 6182 6626
rect 5430 6539 5450 6559
rect 5192 4141 5217 4167
rect 5581 4072 5601 4092
rect 4849 4005 4878 4032
rect 4923 4008 4952 4035
rect 5137 3907 5158 3927
rect 5348 3868 5369 3898
rect 5510 3814 5536 3840
rect 5135 3758 5156 3778
rect 5339 3760 5372 3780
rect 5560 3761 5580 3781
rect 4852 3660 4871 3680
rect 4929 3660 4948 3680
rect 5660 3603 5683 3641
rect 6919 5764 6947 5792
rect 7191 5500 7210 5520
rect 7268 5500 7287 5520
rect 6559 5399 6579 5419
rect 6983 5402 7004 5422
rect 6603 5340 6629 5366
rect 7408 5357 7434 5380
rect 6770 5282 6791 5312
rect 6981 5253 7002 5273
rect 7187 5145 7216 5172
rect 7261 5148 7290 5175
rect 6538 5088 6558 5108
rect 6770 5018 6787 5055
rect 6920 4326 6945 4364
rect 7149 3978 7168 3998
rect 7226 3978 7245 3998
rect 6517 3877 6537 3897
rect 6941 3880 6962 3900
rect 8884 7134 8930 7182
rect 12464 7314 12510 7362
rect 14432 10596 14453 10616
rect 14857 10599 14877 10619
rect 14149 10498 14168 10518
rect 14226 10498 14245 10518
rect 14449 10132 14474 10170
rect 14607 9441 14624 9478
rect 14836 9388 14856 9408
rect 14104 9321 14133 9348
rect 14178 9324 14207 9351
rect 14392 9223 14413 9243
rect 14603 9184 14624 9214
rect 13960 9116 13986 9139
rect 14765 9130 14791 9156
rect 14390 9074 14411 9094
rect 14815 9077 14835 9097
rect 14107 8976 14126 8996
rect 14184 8976 14203 8996
rect 14447 8704 14475 8732
rect 15944 7937 15964 7957
rect 15212 7870 15241 7897
rect 15286 7873 15315 7900
rect 15500 7772 15521 7792
rect 15711 7733 15732 7763
rect 15008 7674 15032 7698
rect 15065 7675 15089 7699
rect 15873 7679 15899 7705
rect 15498 7623 15519 7643
rect 15711 7621 15735 7643
rect 15923 7626 15943 7646
rect 15215 7525 15234 7545
rect 15292 7525 15311 7545
rect 19594 12792 19634 12818
rect 19598 12739 19638 12765
rect 20604 13021 20641 13062
rect 20660 13023 20697 13064
rect 20396 12944 20415 12964
rect 20473 12944 20492 12964
rect 19764 12843 19784 12863
rect 20188 12846 20209 12866
rect 20653 12831 20689 12852
rect 19808 12784 19834 12810
rect 19975 12726 19996 12756
rect 20186 12697 20207 12717
rect 20653 12775 20693 12812
rect 20392 12589 20421 12616
rect 20466 12592 20495 12619
rect 19743 12532 19763 12552
rect 19921 12482 19953 12502
rect 19976 12483 20001 12503
rect 19583 12389 19628 12428
rect 19348 12269 19367 12289
rect 19425 12269 19444 12289
rect 18716 12168 18736 12188
rect 19140 12171 19161 12191
rect 18760 12109 18786 12135
rect 19592 12132 19645 12165
rect 18927 12051 18948 12081
rect 19138 12022 19159 12042
rect 19597 12074 19650 12107
rect 20639 12358 20679 12391
rect 20396 12265 20415 12285
rect 20473 12265 20492 12285
rect 19764 12164 19784 12184
rect 20188 12167 20209 12187
rect 19808 12105 19834 12131
rect 20640 12122 20689 12164
rect 19975 12047 19996 12077
rect 19344 11914 19373 11941
rect 19418 11917 19447 11944
rect 20186 12018 20207 12038
rect 20641 12059 20690 12101
rect 20392 11910 20421 11937
rect 20466 11913 20495 11940
rect 18695 11857 18715 11877
rect 19743 11853 19763 11873
rect 17629 11766 17657 11794
rect 19927 11776 19952 11814
rect 19971 11779 19996 11814
rect 19602 11675 19632 11741
rect 17901 11502 17920 11522
rect 17978 11502 17997 11522
rect 17269 11401 17289 11421
rect 17693 11404 17714 11424
rect 17313 11342 17339 11368
rect 18118 11359 18144 11382
rect 18498 11352 18524 11375
rect 17480 11284 17501 11314
rect 17691 11255 17712 11275
rect 19591 11390 19631 11416
rect 19594 11345 19634 11371
rect 19598 11292 19638 11318
rect 17897 11147 17926 11174
rect 17971 11150 18000 11177
rect 17248 11090 17268 11110
rect 17480 11020 17497 11057
rect 20604 11574 20641 11615
rect 20660 11576 20697 11617
rect 20396 11497 20415 11517
rect 20473 11497 20492 11517
rect 19764 11396 19784 11416
rect 20188 11399 20209 11419
rect 20653 11384 20689 11405
rect 19808 11337 19834 11363
rect 19975 11279 19996 11309
rect 20186 11250 20207 11270
rect 20653 11328 20693 11365
rect 20392 11142 20421 11169
rect 20466 11145 20495 11172
rect 19743 11085 19763 11105
rect 19921 11035 19953 11055
rect 19976 11036 20001 11056
rect 17630 10328 17655 10366
rect 19583 10942 19628 10981
rect 19348 10822 19367 10842
rect 19425 10822 19444 10842
rect 18716 10721 18736 10741
rect 19140 10724 19161 10744
rect 18760 10662 18786 10688
rect 19592 10685 19645 10718
rect 18927 10604 18948 10634
rect 19138 10575 19159 10595
rect 19597 10627 19650 10660
rect 20639 10911 20679 10944
rect 20396 10818 20415 10838
rect 20473 10818 20492 10838
rect 19764 10717 19784 10737
rect 20188 10720 20209 10740
rect 19808 10658 19834 10684
rect 20640 10675 20689 10717
rect 19975 10600 19996 10630
rect 19344 10467 19373 10494
rect 19418 10470 19447 10497
rect 20186 10571 20207 10591
rect 20641 10612 20690 10654
rect 20392 10463 20421 10490
rect 20466 10466 20495 10493
rect 18695 10410 18715 10430
rect 19743 10406 19763 10426
rect 19927 10329 19952 10367
rect 19971 10332 19996 10367
rect 19591 10176 19645 10242
rect 17859 9980 17878 10000
rect 17936 9980 17955 10000
rect 17227 9879 17247 9899
rect 17651 9882 17672 9902
rect 17271 9820 17297 9846
rect 17438 9762 17459 9792
rect 17649 9733 17670 9753
rect 17855 9625 17884 9652
rect 17929 9628 17958 9655
rect 17206 9568 17226 9588
rect 19596 10119 19640 10156
rect 19592 9870 19632 9896
rect 19595 9825 19635 9851
rect 19599 9772 19639 9798
rect 20605 10054 20642 10095
rect 20661 10056 20698 10097
rect 20397 9977 20416 9997
rect 20474 9977 20493 9997
rect 19765 9876 19785 9896
rect 20189 9879 20210 9899
rect 20654 9864 20690 9885
rect 19809 9817 19835 9843
rect 19976 9759 19997 9789
rect 20187 9730 20208 9750
rect 20654 9808 20694 9845
rect 20393 9622 20422 9649
rect 20467 9625 20496 9652
rect 19744 9565 19764 9585
rect 19922 9515 19954 9535
rect 19977 9516 20002 9536
rect 17435 8851 17459 8874
rect 17435 8807 17459 8830
rect 17653 8808 17678 8846
rect 17697 8811 17722 8846
rect 17439 8627 17491 8645
rect 17270 8434 17290 8454
rect 17902 8535 17921 8555
rect 17979 8535 17998 8555
rect 19584 9422 19629 9461
rect 19349 9302 19368 9322
rect 19426 9302 19445 9322
rect 18717 9201 18737 9221
rect 19141 9204 19162 9224
rect 18761 9142 18787 9168
rect 19593 9165 19646 9198
rect 18928 9084 18949 9114
rect 19139 9055 19160 9075
rect 19598 9107 19651 9140
rect 20640 9391 20680 9424
rect 20397 9298 20416 9318
rect 20474 9298 20493 9318
rect 19765 9197 19785 9217
rect 20189 9200 20210 9220
rect 19809 9138 19835 9164
rect 20641 9155 20690 9197
rect 19976 9080 19997 9110
rect 19345 8947 19374 8974
rect 19419 8950 19448 8977
rect 20187 9051 20208 9071
rect 20642 9092 20691 9134
rect 20393 8943 20422 8970
rect 20467 8946 20496 8973
rect 18696 8890 18716 8910
rect 19744 8886 19764 8906
rect 19928 8809 19953 8847
rect 19972 8812 19997 8847
rect 19603 8708 19633 8774
rect 17694 8437 17715 8457
rect 17314 8375 17340 8401
rect 18306 8407 18360 8448
rect 17481 8317 17502 8347
rect 17692 8288 17713 8308
rect 19592 8423 19632 8449
rect 19595 8378 19635 8404
rect 19599 8325 19639 8351
rect 20605 8607 20642 8648
rect 20661 8609 20698 8650
rect 20397 8530 20416 8550
rect 20474 8530 20493 8550
rect 19765 8429 19785 8449
rect 20189 8432 20210 8452
rect 20654 8417 20690 8438
rect 19809 8370 19835 8396
rect 19976 8312 19997 8342
rect 17898 8180 17927 8207
rect 17972 8183 18001 8210
rect 17249 8123 17269 8143
rect 15551 7432 15580 7466
rect 15550 7372 15579 7406
rect 13766 7287 13810 7315
rect 13575 7188 13612 7236
rect 13763 7230 13807 7258
rect 8881 6835 8921 6861
rect 8884 6790 8924 6816
rect 8888 6737 8928 6763
rect 16058 7148 16121 7202
rect 9894 7019 9931 7060
rect 9950 7021 9987 7062
rect 9686 6942 9705 6962
rect 9763 6942 9782 6962
rect 9054 6841 9074 6861
rect 9478 6844 9499 6864
rect 12105 7090 12130 7125
rect 12149 7090 12174 7128
rect 12338 7031 12358 7051
rect 13155 7091 13180 7126
rect 13199 7091 13224 7129
rect 9943 6829 9979 6850
rect 13386 7027 13406 7047
rect 11606 6964 11635 6991
rect 11680 6967 11709 6994
rect 9098 6782 9124 6808
rect 9265 6724 9286 6754
rect 9476 6695 9497 6715
rect 9943 6773 9983 6810
rect 11411 6803 11460 6845
rect 11894 6866 11915 6886
rect 12654 6960 12683 6987
rect 12728 6963 12757 6990
rect 12105 6827 12126 6857
rect 11412 6740 11461 6782
rect 12267 6773 12293 6799
rect 9682 6587 9711 6614
rect 9756 6590 9785 6617
rect 9033 6530 9053 6550
rect 9211 6480 9243 6500
rect 9266 6481 9291 6501
rect 8873 6387 8918 6426
rect 8638 6267 8657 6287
rect 8715 6267 8734 6287
rect 8006 6166 8026 6186
rect 8430 6169 8451 6189
rect 8050 6107 8076 6133
rect 8882 6130 8935 6163
rect 8217 6049 8238 6079
rect 8428 6020 8449 6040
rect 8887 6072 8940 6105
rect 9929 6356 9969 6389
rect 9686 6263 9705 6283
rect 9763 6263 9782 6283
rect 9054 6162 9074 6182
rect 9478 6165 9499 6185
rect 11892 6717 11913 6737
rect 12317 6720 12337 6740
rect 11609 6619 11628 6639
rect 11686 6619 11705 6639
rect 11422 6513 11462 6546
rect 12451 6797 12504 6830
rect 12942 6862 12963 6882
rect 13153 6823 13174 6853
rect 12456 6739 12509 6772
rect 13315 6769 13341 6795
rect 12940 6713 12961 6733
rect 13365 6716 13385 6736
rect 12657 6615 12676 6635
rect 12734 6615 12753 6635
rect 12473 6476 12518 6515
rect 13576 6776 13610 6815
rect 12100 6401 12125 6421
rect 12148 6402 12180 6422
rect 12338 6352 12358 6372
rect 11606 6285 11635 6312
rect 11680 6288 11709 6315
rect 9098 6103 9124 6129
rect 9930 6120 9979 6162
rect 9265 6045 9286 6075
rect 8634 5912 8663 5939
rect 8708 5915 8737 5942
rect 9476 6016 9497 6036
rect 9931 6057 9980 6099
rect 11408 6092 11448 6129
rect 11894 6187 11915 6207
rect 13753 6796 13789 6837
rect 13742 6456 13802 6500
rect 14833 6347 14853 6367
rect 14101 6280 14130 6307
rect 14175 6283 14204 6310
rect 12105 6148 12126 6178
rect 12267 6094 12293 6120
rect 9682 5908 9711 5935
rect 9756 5911 9785 5938
rect 7985 5855 8005 5875
rect 11412 6052 11448 6073
rect 9033 5851 9053 5871
rect 9217 5774 9242 5812
rect 9261 5777 9286 5812
rect 11892 6038 11913 6058
rect 12317 6041 12337 6061
rect 11609 5940 11628 5960
rect 11686 5940 11705 5960
rect 11404 5840 11441 5881
rect 11460 5842 11497 5883
rect 12463 6139 12503 6165
rect 12467 6086 12507 6112
rect 12470 6041 12510 6067
rect 8892 5673 8922 5739
rect 14389 6182 14410 6202
rect 14600 6143 14621 6173
rect 13742 6042 13796 6083
rect 14762 6089 14788 6115
rect 14387 6033 14408 6053
rect 12469 5716 12499 5782
rect 7788 5350 7814 5373
rect 8881 5388 8921 5414
rect 8884 5343 8924 5369
rect 8888 5290 8928 5316
rect 9894 5572 9931 5613
rect 9950 5574 9987 5615
rect 9686 5495 9705 5515
rect 9763 5495 9782 5515
rect 9054 5394 9074 5414
rect 9478 5397 9499 5417
rect 12105 5643 12130 5678
rect 12149 5643 12174 5681
rect 12338 5584 12358 5604
rect 9943 5382 9979 5403
rect 13386 5580 13406 5600
rect 11606 5517 11635 5544
rect 11680 5520 11709 5547
rect 9098 5335 9124 5361
rect 9265 5277 9286 5307
rect 9476 5248 9497 5268
rect 9943 5326 9983 5363
rect 11411 5356 11460 5398
rect 11894 5419 11915 5439
rect 12654 5513 12683 5540
rect 12728 5516 12757 5543
rect 12105 5380 12126 5410
rect 11412 5293 11461 5335
rect 12267 5326 12293 5352
rect 9682 5140 9711 5167
rect 9756 5143 9785 5170
rect 9033 5083 9053 5103
rect 9211 5033 9243 5053
rect 9266 5034 9291 5054
rect 8873 4940 8918 4979
rect 8638 4820 8657 4840
rect 8715 4820 8734 4840
rect 8006 4719 8026 4739
rect 8430 4722 8451 4742
rect 8050 4660 8076 4686
rect 8882 4683 8935 4716
rect 8217 4602 8238 4632
rect 8428 4573 8449 4593
rect 8887 4625 8940 4658
rect 9929 4909 9969 4942
rect 9686 4816 9705 4836
rect 9763 4816 9782 4836
rect 9054 4715 9074 4735
rect 9478 4718 9499 4738
rect 11892 5270 11913 5290
rect 12317 5273 12337 5293
rect 11609 5172 11628 5192
rect 11686 5172 11705 5192
rect 11422 5066 11462 5099
rect 12451 5350 12504 5383
rect 12942 5415 12963 5435
rect 13153 5376 13174 5406
rect 12456 5292 12509 5325
rect 13315 5322 13341 5348
rect 12940 5266 12961 5286
rect 13365 5269 13385 5289
rect 12657 5168 12676 5188
rect 12734 5168 12753 5188
rect 12473 5029 12518 5068
rect 14104 5935 14123 5955
rect 14181 5935 14200 5955
rect 14812 6036 14832 6056
rect 14611 5845 14663 5863
rect 14380 5644 14405 5679
rect 14424 5644 14449 5682
rect 14643 5660 14667 5683
rect 14643 5616 14667 5639
rect 12100 4954 12125 4974
rect 12148 4955 12180 4975
rect 12338 4905 12358 4925
rect 11606 4838 11635 4865
rect 11680 4841 11709 4868
rect 9098 4656 9124 4682
rect 9930 4673 9979 4715
rect 9265 4598 9286 4628
rect 8634 4465 8663 4492
rect 8708 4468 8737 4495
rect 9476 4569 9497 4589
rect 9931 4610 9980 4652
rect 11408 4645 11448 4682
rect 11894 4740 11915 4760
rect 12105 4701 12126 4731
rect 12267 4647 12293 4673
rect 9682 4461 9711 4488
rect 9756 4464 9785 4491
rect 7985 4408 8005 4428
rect 11412 4605 11448 4626
rect 9033 4404 9053 4424
rect 9217 4327 9242 4365
rect 9261 4330 9286 4365
rect 11892 4591 11913 4611
rect 12317 4594 12337 4614
rect 11609 4493 11628 4513
rect 11686 4493 11705 4513
rect 11404 4393 11441 4434
rect 11460 4395 11497 4436
rect 12463 4692 12503 4718
rect 12467 4639 12507 4665
rect 12470 4594 12510 4620
rect 12462 4334 12506 4371
rect 14876 4902 14896 4922
rect 14144 4835 14173 4862
rect 14218 4838 14247 4865
rect 14432 4737 14453 4757
rect 14643 4698 14664 4728
rect 14805 4644 14831 4670
rect 8881 4174 8935 4240
rect 12457 4248 12511 4314
rect 6561 3818 6587 3844
rect 6728 3760 6749 3790
rect 6939 3731 6960 3751
rect 7145 3623 7174 3650
rect 7219 3626 7248 3653
rect 6496 3566 6516 3586
rect 3897 3439 3914 3476
rect 6683 3465 6703 3486
rect 6724 3470 6744 3491
rect 4126 3386 4146 3406
rect 3394 3319 3423 3346
rect 3468 3322 3497 3349
rect 3682 3221 3703 3241
rect 3893 3182 3914 3212
rect 3250 3114 3276 3137
rect 4055 3128 4081 3154
rect 3680 3072 3701 3092
rect 4105 3075 4125 3095
rect 3397 2974 3416 2994
rect 3474 2974 3493 2994
rect 8886 4117 8930 4154
rect 8882 3868 8922 3894
rect 8885 3823 8925 3849
rect 8889 3770 8929 3796
rect 9895 4052 9932 4093
rect 9951 4054 9988 4095
rect 9687 3975 9706 3995
rect 9764 3975 9783 3995
rect 9055 3874 9075 3894
rect 9479 3877 9500 3897
rect 12106 4123 12131 4158
rect 12150 4123 12175 4161
rect 12339 4064 12359 4084
rect 9944 3862 9980 3883
rect 13387 4060 13407 4080
rect 11607 3997 11636 4024
rect 11681 4000 11710 4027
rect 9099 3815 9125 3841
rect 9266 3757 9287 3787
rect 9477 3728 9498 3748
rect 9944 3806 9984 3843
rect 11412 3836 11461 3878
rect 11895 3899 11916 3919
rect 12655 3993 12684 4020
rect 12729 3996 12758 4023
rect 12106 3860 12127 3890
rect 11413 3773 11462 3815
rect 12268 3806 12294 3832
rect 9683 3620 9712 3647
rect 9757 3623 9786 3650
rect 9034 3563 9054 3583
rect 9212 3513 9244 3533
rect 9267 3514 9292 3534
rect 6725 2849 6749 2872
rect 6725 2805 6749 2828
rect 6943 2806 6968 2844
rect 6987 2809 7012 2844
rect 3737 2702 3765 2730
rect 6729 2625 6781 2643
rect 6560 2432 6580 2452
rect 7192 2533 7211 2553
rect 7269 2533 7288 2553
rect 8874 3420 8919 3459
rect 8639 3300 8658 3320
rect 8716 3300 8735 3320
rect 8007 3199 8027 3219
rect 8431 3202 8452 3222
rect 8051 3140 8077 3166
rect 8883 3163 8936 3196
rect 8218 3082 8239 3112
rect 8429 3053 8450 3073
rect 8888 3105 8941 3138
rect 9930 3389 9970 3422
rect 9687 3296 9706 3316
rect 9764 3296 9783 3316
rect 9055 3195 9075 3215
rect 9479 3198 9500 3218
rect 11893 3750 11914 3770
rect 12318 3753 12338 3773
rect 11610 3652 11629 3672
rect 11687 3652 11706 3672
rect 11423 3546 11463 3579
rect 12452 3830 12505 3863
rect 12943 3895 12964 3915
rect 13154 3856 13175 3886
rect 12457 3772 12510 3805
rect 13316 3802 13342 3828
rect 12941 3746 12962 3766
rect 13366 3749 13386 3769
rect 12658 3648 12677 3668
rect 12735 3648 12754 3668
rect 12474 3509 12519 3548
rect 12101 3434 12126 3454
rect 12149 3435 12181 3455
rect 12339 3385 12359 3405
rect 11607 3318 11636 3345
rect 11681 3321 11710 3348
rect 9099 3136 9125 3162
rect 9931 3153 9980 3195
rect 9266 3078 9287 3108
rect 8635 2945 8664 2972
rect 8709 2948 8738 2975
rect 9477 3049 9498 3069
rect 9932 3090 9981 3132
rect 11409 3125 11449 3162
rect 11895 3220 11916 3240
rect 12106 3181 12127 3211
rect 12268 3127 12294 3153
rect 9683 2941 9712 2968
rect 9757 2944 9786 2971
rect 7986 2888 8006 2908
rect 11413 3085 11449 3106
rect 9034 2884 9054 2904
rect 9218 2807 9243 2845
rect 9262 2810 9287 2845
rect 11893 3071 11914 3091
rect 12318 3074 12338 3094
rect 11610 2973 11629 2993
rect 11687 2973 11706 2993
rect 11405 2873 11442 2914
rect 11461 2875 11498 2916
rect 12464 3172 12504 3198
rect 12468 3119 12508 3145
rect 12471 3074 12511 3100
rect 13533 3105 13558 3136
rect 13578 3115 13604 3138
rect 8893 2706 8923 2772
rect 6984 2435 7005 2455
rect 6604 2373 6630 2399
rect 7596 2405 7650 2446
rect 6771 2315 6792 2345
rect 6982 2286 7003 2306
rect 12470 2749 12500 2815
rect 8882 2421 8922 2447
rect 8885 2376 8925 2402
rect 8889 2323 8929 2349
rect 9895 2605 9932 2646
rect 9951 2607 9988 2648
rect 9687 2528 9706 2548
rect 9764 2528 9783 2548
rect 9055 2427 9075 2447
rect 9479 2430 9500 2450
rect 12106 2676 12131 2711
rect 12150 2676 12175 2714
rect 12339 2617 12359 2637
rect 9944 2415 9980 2436
rect 13387 2613 13407 2633
rect 11607 2550 11636 2577
rect 11681 2553 11710 2580
rect 9099 2368 9125 2394
rect 9266 2310 9287 2340
rect 7188 2178 7217 2205
rect 7262 2181 7291 2208
rect 6539 2121 6559 2141
rect 5879 1647 6010 1712
rect 7590 1988 7650 2032
rect 7603 1651 7639 1692
rect 9477 2281 9498 2301
rect 9944 2359 9984 2396
rect 11412 2389 11461 2431
rect 11895 2452 11916 2472
rect 12655 2546 12684 2573
rect 12729 2549 12758 2576
rect 12106 2413 12127 2443
rect 11413 2326 11462 2368
rect 12268 2359 12294 2385
rect 9683 2173 9712 2200
rect 9757 2176 9786 2203
rect 9034 2116 9054 2136
rect 9212 2066 9244 2086
rect 9267 2067 9292 2087
rect 7782 1673 7816 1712
rect 8874 1973 8919 2012
rect 8639 1853 8658 1873
rect 8716 1853 8735 1873
rect 8007 1752 8027 1772
rect 8431 1755 8452 1775
rect 8051 1693 8077 1719
rect 8883 1716 8936 1749
rect 2812 1420 2912 1527
rect 8218 1635 8239 1665
rect 8429 1606 8450 1626
rect 8888 1658 8941 1691
rect 9930 1942 9970 1975
rect 9687 1849 9706 1869
rect 9764 1849 9783 1869
rect 9055 1748 9075 1768
rect 9479 1751 9500 1771
rect 11893 2303 11914 2323
rect 12318 2306 12338 2326
rect 11610 2205 11629 2225
rect 11687 2205 11706 2225
rect 11423 2099 11463 2132
rect 12452 2383 12505 2416
rect 12943 2448 12964 2468
rect 13154 2409 13175 2439
rect 12457 2325 12510 2358
rect 13316 2355 13342 2381
rect 12941 2299 12962 2319
rect 13366 2302 13386 2322
rect 12658 2201 12677 2221
rect 12735 2201 12754 2221
rect 12474 2062 12519 2101
rect 12101 1987 12126 2007
rect 12149 1988 12181 2008
rect 12339 1938 12359 1958
rect 11607 1871 11636 1898
rect 11681 1874 11710 1901
rect 9099 1689 9125 1715
rect 9931 1706 9980 1748
rect 9266 1631 9287 1661
rect 8635 1498 8664 1525
rect 8709 1501 8738 1528
rect 9477 1602 9498 1622
rect 9932 1643 9981 1685
rect 11409 1678 11449 1715
rect 11895 1773 11916 1793
rect 12106 1734 12127 1764
rect 12268 1680 12294 1706
rect 9683 1494 9712 1521
rect 9757 1497 9786 1524
rect 7986 1441 8006 1461
rect 11413 1638 11449 1659
rect 8168 1359 8193 1397
rect 8212 1362 8237 1397
rect 9034 1437 9054 1457
rect 9218 1360 9243 1398
rect 9262 1363 9287 1398
rect 11893 1624 11914 1644
rect 12318 1627 12338 1647
rect 11610 1526 11629 1546
rect 11687 1526 11706 1546
rect 11405 1426 11442 1467
rect 11461 1428 11498 1469
rect 14430 4588 14451 4608
rect 14855 4591 14875 4611
rect 14147 4490 14166 4510
rect 14224 4490 14243 4510
rect 14447 4124 14472 4162
rect 16523 7084 16552 7118
rect 16522 7024 16551 7058
rect 16791 6945 16810 6965
rect 16868 6945 16887 6965
rect 16159 6844 16179 6864
rect 16583 6847 16604 6867
rect 18300 7990 18360 8034
rect 18313 7653 18349 7694
rect 20187 8283 20208 8303
rect 20654 8361 20694 8398
rect 20393 8175 20422 8202
rect 20467 8178 20496 8205
rect 19744 8118 19764 8138
rect 19922 8068 19954 8088
rect 19977 8069 20002 8089
rect 18492 7675 18526 7714
rect 19584 7975 19629 8014
rect 19349 7855 19368 7875
rect 19426 7855 19445 7875
rect 18717 7754 18737 7774
rect 19141 7757 19162 7777
rect 18761 7695 18787 7721
rect 19593 7718 19646 7751
rect 18928 7637 18949 7667
rect 19139 7608 19160 7628
rect 19598 7660 19651 7693
rect 20640 7944 20680 7977
rect 20397 7851 20416 7871
rect 20474 7851 20493 7871
rect 19765 7750 19785 7770
rect 20189 7753 20210 7773
rect 19809 7691 19835 7717
rect 20641 7708 20690 7750
rect 19976 7633 19997 7663
rect 19345 7500 19374 7527
rect 19419 7503 19448 7530
rect 20187 7604 20208 7624
rect 20642 7645 20691 7687
rect 20393 7496 20422 7523
rect 20467 7499 20496 7526
rect 18696 7443 18716 7463
rect 18878 7361 18903 7399
rect 18922 7364 18947 7399
rect 19744 7439 19764 7459
rect 19928 7362 19953 7400
rect 19972 7365 19997 7400
rect 16203 6785 16229 6811
rect 17013 6791 17037 6815
rect 17070 6792 17094 6816
rect 16370 6727 16391 6757
rect 16581 6698 16602 6718
rect 18295 7232 18339 7260
rect 18490 7254 18527 7302
rect 18292 7175 18336 7203
rect 16787 6590 16816 6617
rect 16861 6593 16890 6620
rect 16138 6533 16158 6553
rect 15900 4135 15925 4161
rect 16289 4066 16309 4086
rect 15557 3999 15586 4026
rect 15631 4002 15660 4029
rect 15845 3901 15866 3921
rect 16056 3862 16077 3892
rect 16218 3808 16244 3834
rect 15843 3752 15864 3772
rect 16047 3754 16080 3774
rect 16268 3755 16288 3775
rect 15560 3654 15579 3674
rect 15637 3654 15656 3674
rect 16368 3597 16391 3635
rect 17627 5758 17655 5786
rect 17899 5494 17918 5514
rect 17976 5494 17995 5514
rect 17267 5393 17287 5413
rect 17691 5396 17712 5416
rect 17311 5334 17337 5360
rect 18116 5351 18142 5374
rect 17478 5276 17499 5306
rect 17689 5247 17710 5267
rect 17895 5139 17924 5166
rect 17969 5142 17998 5169
rect 17246 5082 17266 5102
rect 17478 5012 17495 5049
rect 17628 4320 17653 4358
rect 17857 3972 17876 3992
rect 17934 3972 17953 3992
rect 17225 3871 17245 3891
rect 17649 3874 17670 3894
rect 19592 7128 19638 7176
rect 19589 6829 19629 6855
rect 19592 6784 19632 6810
rect 19596 6731 19636 6757
rect 20602 7013 20639 7054
rect 20658 7015 20695 7056
rect 20394 6936 20413 6956
rect 20471 6936 20490 6956
rect 19762 6835 19782 6855
rect 20186 6838 20207 6858
rect 20651 6823 20687 6844
rect 19806 6776 19832 6802
rect 19973 6718 19994 6748
rect 20184 6689 20205 6709
rect 20651 6767 20691 6804
rect 20390 6581 20419 6608
rect 20464 6584 20493 6611
rect 19741 6524 19761 6544
rect 19919 6474 19951 6494
rect 19974 6475 19999 6495
rect 19581 6381 19626 6420
rect 19346 6261 19365 6281
rect 19423 6261 19442 6281
rect 18714 6160 18734 6180
rect 19138 6163 19159 6183
rect 18758 6101 18784 6127
rect 19590 6124 19643 6157
rect 18925 6043 18946 6073
rect 19136 6014 19157 6034
rect 19595 6066 19648 6099
rect 20637 6350 20677 6383
rect 20394 6257 20413 6277
rect 20471 6257 20490 6277
rect 19762 6156 19782 6176
rect 20186 6159 20207 6179
rect 19806 6097 19832 6123
rect 20638 6114 20687 6156
rect 19973 6039 19994 6069
rect 19342 5906 19371 5933
rect 19416 5909 19445 5936
rect 20184 6010 20205 6030
rect 20639 6051 20688 6093
rect 20390 5902 20419 5929
rect 20464 5905 20493 5932
rect 18693 5849 18713 5869
rect 19741 5845 19761 5865
rect 19925 5768 19950 5806
rect 19969 5771 19994 5806
rect 19600 5667 19630 5733
rect 18496 5344 18522 5367
rect 19589 5382 19629 5408
rect 19592 5337 19632 5363
rect 19596 5284 19636 5310
rect 20602 5566 20639 5607
rect 20658 5568 20695 5609
rect 20394 5489 20413 5509
rect 20471 5489 20490 5509
rect 19762 5388 19782 5408
rect 20186 5391 20207 5411
rect 20651 5376 20687 5397
rect 19806 5329 19832 5355
rect 19973 5271 19994 5301
rect 20184 5242 20205 5262
rect 20651 5320 20691 5357
rect 20390 5134 20419 5161
rect 20464 5137 20493 5164
rect 19741 5077 19761 5097
rect 19919 5027 19951 5047
rect 19974 5028 19999 5048
rect 19581 4934 19626 4973
rect 19346 4814 19365 4834
rect 19423 4814 19442 4834
rect 18714 4713 18734 4733
rect 19138 4716 19159 4736
rect 18758 4654 18784 4680
rect 19590 4677 19643 4710
rect 18925 4596 18946 4626
rect 19136 4567 19157 4587
rect 19595 4619 19648 4652
rect 20637 4903 20677 4936
rect 20394 4810 20413 4830
rect 20471 4810 20490 4830
rect 19762 4709 19782 4729
rect 20186 4712 20207 4732
rect 19806 4650 19832 4676
rect 20638 4667 20687 4709
rect 19973 4592 19994 4622
rect 19342 4459 19371 4486
rect 19416 4462 19445 4489
rect 20184 4563 20205 4583
rect 20639 4604 20688 4646
rect 20390 4455 20419 4482
rect 20464 4458 20493 4485
rect 18693 4402 18713 4422
rect 19741 4398 19761 4418
rect 19925 4321 19950 4359
rect 19969 4324 19994 4359
rect 19589 4168 19643 4234
rect 17269 3812 17295 3838
rect 17436 3754 17457 3784
rect 17647 3725 17668 3745
rect 17853 3617 17882 3644
rect 17927 3620 17956 3647
rect 17204 3560 17224 3580
rect 14605 3433 14622 3470
rect 17391 3459 17411 3480
rect 17432 3464 17452 3485
rect 14834 3380 14854 3400
rect 14102 3313 14131 3340
rect 14176 3316 14205 3343
rect 14390 3215 14411 3235
rect 14601 3176 14622 3206
rect 13958 3108 13984 3131
rect 14763 3122 14789 3148
rect 14388 3066 14409 3086
rect 14813 3069 14833 3089
rect 14105 2968 14124 2988
rect 14182 2968 14201 2988
rect 19594 4111 19638 4148
rect 19590 3862 19630 3888
rect 19593 3817 19633 3843
rect 19597 3764 19637 3790
rect 20603 4046 20640 4087
rect 20659 4048 20696 4089
rect 20395 3969 20414 3989
rect 20472 3969 20491 3989
rect 19763 3868 19783 3888
rect 20187 3871 20208 3891
rect 20652 3856 20688 3877
rect 19807 3809 19833 3835
rect 19974 3751 19995 3781
rect 20185 3722 20206 3742
rect 20652 3800 20692 3837
rect 20391 3614 20420 3641
rect 20465 3617 20494 3644
rect 19742 3557 19762 3577
rect 19920 3507 19952 3527
rect 19975 3508 20000 3528
rect 17433 2843 17457 2866
rect 17433 2799 17457 2822
rect 17651 2800 17676 2838
rect 17695 2803 17720 2838
rect 14445 2696 14473 2724
rect 17437 2619 17489 2637
rect 17268 2426 17288 2446
rect 17900 2527 17919 2547
rect 17977 2527 17996 2547
rect 19582 3414 19627 3453
rect 19347 3294 19366 3314
rect 19424 3294 19443 3314
rect 18715 3193 18735 3213
rect 19139 3196 19160 3216
rect 18759 3134 18785 3160
rect 19591 3157 19644 3190
rect 18926 3076 18947 3106
rect 19137 3047 19158 3067
rect 19596 3099 19649 3132
rect 20638 3383 20678 3416
rect 20395 3290 20414 3310
rect 20472 3290 20491 3310
rect 19763 3189 19783 3209
rect 20187 3192 20208 3212
rect 19807 3130 19833 3156
rect 20639 3147 20688 3189
rect 19974 3072 19995 3102
rect 19343 2939 19372 2966
rect 19417 2942 19446 2969
rect 20185 3043 20206 3063
rect 20640 3084 20689 3126
rect 20391 2935 20420 2962
rect 20465 2938 20494 2965
rect 18694 2882 18714 2902
rect 19742 2878 19762 2898
rect 19926 2801 19951 2839
rect 19970 2804 19995 2839
rect 19601 2700 19631 2766
rect 17692 2429 17713 2449
rect 17312 2367 17338 2393
rect 18304 2399 18358 2440
rect 17479 2309 17500 2339
rect 17690 2280 17711 2300
rect 19590 2415 19630 2441
rect 19593 2370 19633 2396
rect 19597 2317 19637 2343
rect 20603 2599 20640 2640
rect 20659 2601 20696 2642
rect 20395 2522 20414 2542
rect 20472 2522 20491 2542
rect 19763 2421 19783 2441
rect 20187 2424 20208 2444
rect 20652 2409 20688 2430
rect 19807 2362 19833 2388
rect 19974 2304 19995 2334
rect 17896 2172 17925 2199
rect 17970 2175 17999 2202
rect 17247 2115 17267 2135
rect 16587 1641 16718 1706
rect 18298 1982 18358 2026
rect 18311 1645 18347 1686
rect 20185 2275 20206 2295
rect 20652 2353 20692 2390
rect 20391 2167 20420 2194
rect 20465 2170 20494 2197
rect 19742 2110 19762 2130
rect 19920 2060 19952 2080
rect 19975 2061 20000 2081
rect 18490 1667 18524 1706
rect 19582 1967 19627 2006
rect 19347 1847 19366 1867
rect 19424 1847 19443 1867
rect 18715 1746 18735 1766
rect 19139 1749 19160 1769
rect 18759 1687 18785 1713
rect 19591 1710 19644 1743
rect 13520 1414 13620 1521
rect 18926 1629 18947 1659
rect 19137 1600 19158 1620
rect 19596 1652 19649 1685
rect 20638 1936 20678 1969
rect 20395 1843 20414 1863
rect 20472 1843 20491 1863
rect 19763 1742 19783 1762
rect 20187 1745 20208 1765
rect 19807 1683 19833 1709
rect 20639 1700 20688 1742
rect 19974 1625 19995 1655
rect 19343 1492 19372 1519
rect 19417 1495 19446 1522
rect 20185 1596 20206 1616
rect 20640 1637 20689 1679
rect 20391 1488 20420 1515
rect 20465 1491 20494 1518
rect 18694 1435 18714 1455
rect 18876 1353 18901 1391
rect 18920 1356 18945 1391
rect 19742 1431 19762 1451
rect 19926 1354 19951 1392
rect 19970 1357 19995 1392
rect 10139 -34 10215 12
rect 11601 -112 11642 -64
rect 11342 -215 11362 -195
rect 10610 -282 10639 -255
rect 10684 -279 10713 -252
rect 10113 -489 10144 -430
rect 10175 -489 10206 -430
rect 10898 -380 10919 -360
rect 11109 -419 11130 -389
rect 11271 -473 11297 -447
rect 10896 -529 10917 -509
rect 11110 -531 11130 -508
rect 11321 -526 11341 -506
rect 10613 -627 10632 -607
rect 10690 -627 10709 -607
<< metal1 >>
rect 2856 13693 2921 13728
rect 2856 13689 2869 13693
rect 2857 13645 2869 13689
rect 2906 13689 2921 13693
rect 2906 13645 2919 13689
rect 217 12671 324 13461
rect 696 12859 768 13452
rect 1392 13150 1464 13151
rect 1391 13142 1490 13150
rect 1391 13139 1443 13142
rect 1391 13104 1399 13139
rect 1424 13104 1443 13139
rect 1468 13104 1490 13142
rect 1391 13092 1490 13104
rect 1392 13073 1460 13092
rect 1393 13070 1426 13073
rect 1628 13070 1660 13071
rect 803 13009 1006 13022
rect 803 12976 827 13009
rect 863 13008 1006 13009
rect 863 13005 974 13008
rect 863 12978 900 13005
rect 929 12981 974 13005
rect 1003 12981 1006 13008
rect 929 12978 1006 12981
rect 863 12976 1006 12978
rect 803 12963 1006 12976
rect 803 12962 904 12963
rect 696 12817 705 12859
rect 754 12817 768 12859
rect 696 12796 768 12817
rect 696 12754 706 12796
rect 755 12754 768 12796
rect 696 12736 768 12754
rect 1181 12900 1213 12907
rect 1181 12880 1188 12900
rect 1209 12880 1213 12900
rect 1181 12815 1213 12880
rect 1393 12871 1424 13070
rect 1625 13065 1660 13070
rect 1625 13045 1632 13065
rect 1652 13045 1660 13065
rect 1625 13037 1660 13045
rect 1393 12841 1399 12871
rect 1420 12841 1424 12871
rect 1393 12833 1424 12841
rect 1551 12815 1591 12816
rect 1181 12813 1593 12815
rect 1181 12787 1561 12813
rect 1587 12787 1593 12813
rect 1181 12779 1593 12787
rect 1181 12751 1213 12779
rect 1626 12759 1660 13037
rect 1742 12850 1812 13453
rect 2442 13151 2514 13152
rect 2441 13143 2530 13151
rect 2441 13140 2493 13143
rect 2441 13105 2449 13140
rect 2474 13105 2493 13140
rect 2518 13105 2530 13143
rect 2441 13093 2530 13105
rect 2441 13092 2510 13093
rect 2441 13074 2477 13092
rect 1851 13005 2054 13018
rect 1851 12972 1875 13005
rect 1911 13004 2054 13005
rect 1911 13001 2022 13004
rect 1911 12974 1948 13001
rect 1977 12977 2022 13001
rect 2051 12977 2054 13004
rect 1977 12974 2054 12977
rect 1911 12972 2054 12974
rect 1851 12959 2054 12972
rect 1851 12958 1952 12959
rect 1181 12731 1186 12751
rect 1207 12731 1213 12751
rect 1181 12724 1213 12731
rect 1604 12754 1660 12759
rect 1604 12734 1611 12754
rect 1631 12734 1660 12754
rect 1737 12844 1812 12850
rect 1737 12811 1745 12844
rect 1798 12811 1812 12844
rect 1737 12786 1812 12811
rect 1737 12753 1750 12786
rect 1803 12753 1812 12786
rect 1737 12744 1812 12753
rect 2229 12896 2261 12903
rect 2229 12876 2236 12896
rect 2257 12876 2261 12896
rect 2229 12811 2261 12876
rect 2441 12867 2472 13074
rect 2676 13066 2708 13067
rect 2673 13061 2708 13066
rect 2673 13041 2680 13061
rect 2700 13041 2708 13061
rect 2673 13033 2708 13041
rect 2441 12837 2447 12867
rect 2468 12837 2472 12867
rect 2441 12829 2472 12837
rect 2599 12811 2639 12812
rect 2229 12809 2641 12811
rect 2229 12783 2609 12809
rect 2635 12783 2641 12809
rect 2229 12775 2641 12783
rect 2229 12747 2261 12775
rect 2674 12755 2708 13033
rect 2857 12848 2919 13645
rect 3026 13316 3108 13723
rect 4293 13417 4342 13763
rect 5330 13756 5432 13772
rect 5330 13531 5438 13756
rect 5330 13473 5350 13531
rect 5428 13473 5438 13531
rect 16052 13528 16160 13548
rect 16052 13522 16069 13528
rect 4271 13406 4370 13417
rect 4271 13351 4287 13406
rect 4353 13351 4370 13406
rect 4271 13337 4370 13351
rect 3011 13295 3132 13316
rect 3011 13222 3025 13295
rect 3095 13222 3132 13295
rect 3011 13206 3132 13222
rect 3026 12851 3108 13206
rect 4293 13000 4342 13337
rect 4810 13012 4948 13016
rect 4790 13000 4948 13012
rect 4283 12984 4948 13000
rect 4283 12917 4842 12984
rect 4928 12917 4948 12984
rect 4283 12901 4948 12917
rect 2857 12829 2921 12848
rect 2857 12790 2870 12829
rect 2904 12790 2921 12829
rect 2857 12771 2921 12790
rect 3026 12810 3047 12851
rect 3083 12810 3108 12851
rect 3026 12781 3108 12810
rect 1737 12739 1795 12744
rect 1604 12727 1660 12734
rect 2229 12727 2234 12747
rect 2255 12727 2261 12747
rect 1604 12726 1639 12727
rect 2229 12720 2261 12727
rect 2652 12750 2708 12755
rect 2652 12730 2659 12750
rect 2679 12730 2708 12750
rect 2652 12723 2708 12730
rect 2652 12722 2687 12723
rect 895 12671 1006 12675
rect 2678 12671 3791 12672
rect 217 12653 3791 12671
rect 217 12633 903 12653
rect 922 12633 980 12653
rect 999 12649 3791 12653
rect 999 12633 1951 12649
rect 217 12629 1951 12633
rect 1970 12629 2028 12649
rect 2047 12629 3791 12649
rect 217 12615 3791 12629
rect 217 11992 324 12615
rect 1943 12612 2054 12615
rect 703 12566 767 12570
rect 699 12560 767 12566
rect 699 12527 716 12560
rect 756 12527 767 12560
rect 699 12515 767 12527
rect 1750 12529 1815 12551
rect 699 12513 756 12515
rect 703 12152 754 12513
rect 1750 12490 1767 12529
rect 1812 12490 1815 12529
rect 1391 12445 1426 12447
rect 1391 12436 1495 12445
rect 1391 12435 1442 12436
rect 1391 12415 1394 12435
rect 1419 12416 1442 12435
rect 1474 12416 1495 12436
rect 1419 12415 1495 12416
rect 1391 12408 1495 12415
rect 1391 12396 1426 12408
rect 803 12330 1006 12343
rect 803 12297 827 12330
rect 863 12329 1006 12330
rect 863 12326 974 12329
rect 863 12299 900 12326
rect 929 12302 974 12326
rect 1003 12302 1006 12329
rect 929 12299 1006 12302
rect 863 12297 1006 12299
rect 803 12284 1006 12297
rect 803 12283 904 12284
rect 1181 12221 1213 12228
rect 1181 12201 1188 12221
rect 1209 12201 1213 12221
rect 692 12143 757 12152
rect 692 12106 702 12143
rect 742 12109 757 12143
rect 1181 12136 1213 12201
rect 1393 12192 1424 12396
rect 1628 12391 1660 12392
rect 1625 12386 1660 12391
rect 1625 12366 1632 12386
rect 1652 12366 1660 12386
rect 1625 12358 1660 12366
rect 1393 12162 1399 12192
rect 1420 12162 1424 12192
rect 1393 12154 1424 12162
rect 1551 12136 1591 12137
rect 1181 12134 1593 12136
rect 742 12106 759 12109
rect 692 12087 759 12106
rect 692 12066 706 12087
rect 742 12066 759 12087
rect 692 12059 759 12066
rect 1181 12108 1561 12134
rect 1587 12108 1593 12134
rect 1181 12100 1593 12108
rect 1181 12072 1213 12100
rect 1626 12080 1660 12358
rect 1750 12190 1815 12490
rect 3021 12514 3114 12529
rect 3021 12470 3036 12514
rect 3096 12470 3114 12514
rect 1181 12052 1186 12072
rect 1207 12052 1213 12072
rect 1181 12045 1213 12052
rect 1604 12075 1660 12080
rect 1604 12055 1611 12075
rect 1631 12055 1660 12075
rect 1604 12048 1660 12055
rect 1740 12179 1820 12190
rect 1740 12153 1757 12179
rect 1797 12153 1820 12179
rect 1740 12126 1820 12153
rect 1740 12100 1761 12126
rect 1801 12100 1820 12126
rect 1740 12081 1820 12100
rect 1740 12055 1764 12081
rect 1804 12055 1820 12081
rect 1604 12047 1639 12048
rect 1740 12043 1820 12055
rect 3021 12097 3114 12470
rect 3298 12325 3501 12338
rect 3298 12292 3322 12325
rect 3358 12324 3501 12325
rect 3358 12321 3469 12324
rect 3358 12294 3395 12321
rect 3424 12297 3469 12321
rect 3498 12297 3501 12324
rect 3424 12294 3501 12297
rect 3358 12292 3501 12294
rect 3298 12279 3501 12292
rect 3298 12278 3399 12279
rect 3021 12056 3036 12097
rect 3090 12056 3114 12097
rect 3021 12049 3114 12056
rect 3676 12216 3708 12223
rect 3676 12196 3683 12216
rect 3704 12196 3708 12216
rect 3676 12131 3708 12196
rect 3888 12187 3919 12388
rect 4123 12386 4155 12387
rect 4120 12381 4155 12386
rect 4120 12361 4127 12381
rect 4147 12361 4155 12381
rect 4120 12353 4155 12361
rect 3888 12157 3894 12187
rect 3915 12157 3919 12187
rect 3888 12149 3919 12157
rect 4046 12131 4086 12132
rect 3676 12129 4088 12131
rect 3676 12103 4056 12129
rect 4082 12103 4088 12129
rect 3676 12095 4088 12103
rect 3676 12067 3708 12095
rect 4121 12075 4155 12353
rect 3676 12047 3681 12067
rect 3702 12047 3708 12067
rect 3676 12040 3708 12047
rect 4099 12070 4155 12075
rect 4099 12050 4106 12070
rect 4126 12050 4155 12070
rect 4099 12043 4155 12050
rect 4099 12042 4134 12043
rect 895 11992 1006 11996
rect 2637 11992 4186 11995
rect 215 11974 4186 11992
rect 215 11954 903 11974
rect 922 11954 980 11974
rect 999 11969 4186 11974
rect 999 11954 3398 11969
rect 215 11949 3398 11954
rect 3417 11949 3475 11969
rect 3494 11949 4186 11969
rect 215 11939 4186 11949
rect 215 11936 840 11939
rect 1027 11936 4186 11939
rect 217 11708 324 11936
rect 2637 11935 4186 11936
rect 3390 11932 3501 11935
rect 685 11897 806 11907
rect 685 11895 754 11897
rect 685 11854 698 11895
rect 735 11856 754 11895
rect 791 11856 806 11897
rect 735 11854 806 11856
rect 685 11836 806 11854
rect 3890 11877 3976 11881
rect 3890 11859 3905 11877
rect 3957 11859 3976 11877
rect 3890 11850 3976 11859
rect 691 11734 770 11836
rect 1743 11796 1810 11815
rect 1743 11776 1763 11796
rect 217 11653 325 11708
rect 692 11653 770 11734
rect 1742 11730 1763 11776
rect 1793 11776 1810 11796
rect 1793 11746 1812 11776
rect 1793 11730 1813 11746
rect 1742 11714 1813 11730
rect 1392 11703 1464 11704
rect 1391 11695 1490 11703
rect 1391 11692 1443 11695
rect 1391 11657 1399 11692
rect 1424 11657 1443 11692
rect 1468 11657 1490 11695
rect 217 11224 324 11653
rect 696 11412 768 11653
rect 1391 11645 1490 11657
rect 1392 11626 1460 11645
rect 1393 11623 1426 11626
rect 1628 11623 1660 11624
rect 803 11562 1006 11575
rect 803 11529 827 11562
rect 863 11561 1006 11562
rect 863 11558 974 11561
rect 863 11531 900 11558
rect 929 11534 974 11558
rect 1003 11534 1006 11561
rect 929 11531 1006 11534
rect 863 11529 1006 11531
rect 803 11516 1006 11529
rect 803 11515 904 11516
rect 696 11370 705 11412
rect 754 11370 768 11412
rect 696 11349 768 11370
rect 696 11307 706 11349
rect 755 11307 768 11349
rect 696 11289 768 11307
rect 1181 11453 1213 11460
rect 1181 11433 1188 11453
rect 1209 11433 1213 11453
rect 1181 11368 1213 11433
rect 1393 11424 1424 11623
rect 1625 11618 1660 11623
rect 1625 11598 1632 11618
rect 1652 11598 1660 11618
rect 1625 11590 1660 11598
rect 1393 11394 1399 11424
rect 1420 11394 1424 11424
rect 1393 11386 1424 11394
rect 1551 11368 1591 11369
rect 1181 11366 1593 11368
rect 1181 11340 1561 11366
rect 1587 11340 1593 11366
rect 1181 11332 1593 11340
rect 1181 11304 1213 11332
rect 1626 11312 1660 11590
rect 1742 11403 1812 11714
rect 3667 11704 3739 11705
rect 3666 11701 3755 11704
rect 2438 11699 3755 11701
rect 2435 11696 3755 11699
rect 2435 11693 3718 11696
rect 2435 11658 3674 11693
rect 3699 11658 3718 11693
rect 3743 11658 3755 11696
rect 2435 11648 3755 11658
rect 3931 11697 3967 11850
rect 3931 11674 3937 11697
rect 3961 11674 3967 11697
rect 3931 11653 3967 11674
rect 2435 11646 3720 11648
rect 2435 11636 2532 11646
rect 2441 11627 2477 11636
rect 3931 11630 3937 11653
rect 3961 11630 3967 11653
rect 1851 11558 2054 11571
rect 1851 11525 1875 11558
rect 1911 11557 2054 11558
rect 1911 11554 2022 11557
rect 1911 11527 1948 11554
rect 1977 11530 2022 11554
rect 2051 11530 2054 11557
rect 1977 11527 2054 11530
rect 1911 11525 2054 11527
rect 1851 11512 2054 11525
rect 1851 11511 1952 11512
rect 1181 11284 1186 11304
rect 1207 11284 1213 11304
rect 1181 11277 1213 11284
rect 1604 11307 1660 11312
rect 1604 11287 1611 11307
rect 1631 11287 1660 11307
rect 1737 11397 1812 11403
rect 1737 11364 1745 11397
rect 1798 11364 1812 11397
rect 1737 11339 1812 11364
rect 1737 11306 1750 11339
rect 1803 11306 1812 11339
rect 1737 11297 1812 11306
rect 2229 11449 2261 11456
rect 2229 11429 2236 11449
rect 2257 11429 2261 11449
rect 2229 11364 2261 11429
rect 2441 11420 2472 11627
rect 2676 11619 2708 11620
rect 3931 11619 3967 11630
rect 2673 11614 2708 11619
rect 2673 11594 2680 11614
rect 2700 11594 2708 11614
rect 2673 11586 2708 11594
rect 2441 11390 2447 11420
rect 2468 11390 2472 11420
rect 2441 11382 2472 11390
rect 2599 11364 2639 11365
rect 2229 11362 2641 11364
rect 2229 11336 2609 11362
rect 2635 11336 2641 11362
rect 2229 11328 2641 11336
rect 2229 11300 2261 11328
rect 2674 11308 2708 11586
rect 1737 11292 1795 11297
rect 1604 11280 1660 11287
rect 2229 11280 2234 11300
rect 2255 11280 2261 11300
rect 1604 11279 1639 11280
rect 2229 11273 2261 11280
rect 2652 11303 2708 11308
rect 2652 11283 2659 11303
rect 2679 11283 2708 11303
rect 2652 11276 2708 11283
rect 2652 11275 2687 11276
rect 895 11224 1006 11228
rect 2770 11224 4011 11225
rect 217 11206 4011 11224
rect 217 11186 903 11206
rect 922 11186 980 11206
rect 999 11202 4011 11206
rect 999 11186 1951 11202
rect 217 11182 1951 11186
rect 1970 11182 2028 11202
rect 2047 11182 4011 11202
rect 217 11168 4011 11182
rect 217 10545 324 11168
rect 1943 11165 2054 11168
rect 703 11119 767 11123
rect 699 11113 767 11119
rect 699 11080 716 11113
rect 756 11080 767 11113
rect 699 11068 767 11080
rect 1750 11082 1815 11104
rect 699 11066 756 11068
rect 703 10705 754 11066
rect 1750 11043 1767 11082
rect 1812 11043 1815 11082
rect 1391 10998 1426 11000
rect 1391 10989 1495 10998
rect 1391 10988 1442 10989
rect 1391 10968 1394 10988
rect 1419 10969 1442 10988
rect 1474 10969 1495 10989
rect 1419 10968 1495 10969
rect 1391 10961 1495 10968
rect 1391 10949 1426 10961
rect 803 10883 1006 10896
rect 803 10850 827 10883
rect 863 10882 1006 10883
rect 863 10879 974 10882
rect 863 10852 900 10879
rect 929 10855 974 10879
rect 1003 10855 1006 10882
rect 929 10852 1006 10855
rect 863 10850 1006 10852
rect 803 10837 1006 10850
rect 803 10836 904 10837
rect 1181 10774 1213 10781
rect 1181 10754 1188 10774
rect 1209 10754 1213 10774
rect 692 10696 757 10705
rect 692 10659 702 10696
rect 742 10662 757 10696
rect 1181 10689 1213 10754
rect 1393 10745 1424 10949
rect 1628 10944 1660 10945
rect 1625 10939 1660 10944
rect 1625 10919 1632 10939
rect 1652 10919 1660 10939
rect 1625 10911 1660 10919
rect 1393 10715 1399 10745
rect 1420 10715 1424 10745
rect 1393 10707 1424 10715
rect 1551 10689 1591 10690
rect 1181 10687 1593 10689
rect 742 10659 759 10662
rect 692 10640 759 10659
rect 692 10619 706 10640
rect 742 10619 759 10640
rect 692 10612 759 10619
rect 1181 10661 1561 10687
rect 1587 10661 1593 10687
rect 1181 10653 1593 10661
rect 1181 10625 1213 10653
rect 1626 10633 1660 10911
rect 1750 10743 1815 11043
rect 3929 11037 4034 11046
rect 3929 11032 3983 11037
rect 3929 11011 3942 11032
rect 3962 11016 3983 11032
rect 4003 11016 4034 11037
rect 3962 11011 4034 11016
rect 3929 10980 4034 11011
rect 3932 10963 3967 10980
rect 3931 10945 3967 10963
rect 3341 10880 3544 10893
rect 3341 10847 3365 10880
rect 3401 10879 3544 10880
rect 3401 10876 3512 10879
rect 3401 10849 3438 10876
rect 3467 10852 3512 10876
rect 3541 10852 3544 10879
rect 3467 10849 3544 10852
rect 3401 10847 3544 10849
rect 3341 10834 3544 10847
rect 3341 10833 3442 10834
rect 3719 10771 3751 10778
rect 3719 10751 3726 10771
rect 3747 10751 3751 10771
rect 1181 10605 1186 10625
rect 1207 10605 1213 10625
rect 1181 10598 1213 10605
rect 1604 10628 1660 10633
rect 1604 10608 1611 10628
rect 1631 10608 1660 10628
rect 1604 10601 1660 10608
rect 1740 10732 1820 10743
rect 1740 10706 1757 10732
rect 1797 10706 1820 10732
rect 1740 10679 1820 10706
rect 1740 10653 1761 10679
rect 1801 10653 1820 10679
rect 1740 10634 1820 10653
rect 1740 10608 1764 10634
rect 1804 10608 1820 10634
rect 1604 10600 1639 10601
rect 1740 10596 1820 10608
rect 3719 10686 3751 10751
rect 3931 10742 3962 10945
rect 4166 10941 4198 10942
rect 4163 10936 4198 10941
rect 4163 10916 4170 10936
rect 4190 10916 4198 10936
rect 4163 10908 4198 10916
rect 3931 10712 3937 10742
rect 3958 10712 3962 10742
rect 3931 10704 3962 10712
rect 4089 10686 4129 10687
rect 3719 10684 4131 10686
rect 3719 10658 4099 10684
rect 4125 10658 4131 10684
rect 3719 10650 4131 10658
rect 3719 10622 3751 10650
rect 4164 10630 4198 10908
rect 3719 10602 3724 10622
rect 3745 10602 3751 10622
rect 3719 10595 3751 10602
rect 4142 10625 4198 10630
rect 4142 10605 4149 10625
rect 4169 10605 4198 10625
rect 4142 10598 4198 10605
rect 4142 10597 4177 10598
rect 895 10545 1006 10549
rect 2650 10545 2857 10546
rect 3433 10545 3544 10546
rect 215 10527 4235 10545
rect 215 10507 903 10527
rect 922 10507 980 10527
rect 999 10524 4235 10527
rect 999 10507 3441 10524
rect 215 10504 3441 10507
rect 3460 10504 3518 10524
rect 3537 10504 4235 10524
rect 215 10489 4235 10504
rect 217 10301 324 10489
rect 2812 10487 4235 10489
rect 685 10450 806 10460
rect 685 10448 754 10450
rect 685 10407 698 10448
rect 735 10409 754 10448
rect 791 10409 806 10450
rect 735 10407 806 10409
rect 685 10389 806 10407
rect 217 10297 325 10301
rect 691 10297 768 10389
rect 1741 10385 1817 10401
rect 1741 10362 1756 10385
rect 218 9704 325 10297
rect 693 10246 768 10297
rect 1734 10348 1756 10362
rect 1800 10348 1817 10385
rect 1734 10328 1817 10348
rect 1734 10262 1751 10328
rect 1805 10262 1817 10328
rect 693 10203 769 10246
rect 697 9892 769 10203
rect 1734 10238 1817 10262
rect 1734 10218 1810 10238
rect 1734 10199 1813 10218
rect 1393 10183 1465 10184
rect 1392 10175 1491 10183
rect 1392 10172 1444 10175
rect 1392 10137 1400 10172
rect 1425 10137 1444 10172
rect 1469 10137 1491 10175
rect 1392 10125 1491 10137
rect 1393 10106 1461 10125
rect 1394 10103 1427 10106
rect 1629 10103 1661 10104
rect 804 10042 1007 10055
rect 804 10009 828 10042
rect 864 10041 1007 10042
rect 864 10038 975 10041
rect 864 10011 901 10038
rect 930 10014 975 10038
rect 1004 10014 1007 10041
rect 930 10011 1007 10014
rect 864 10009 1007 10011
rect 804 9996 1007 10009
rect 804 9995 905 9996
rect 697 9850 706 9892
rect 755 9850 769 9892
rect 697 9829 769 9850
rect 697 9787 707 9829
rect 756 9787 769 9829
rect 697 9769 769 9787
rect 1182 9933 1214 9940
rect 1182 9913 1189 9933
rect 1210 9913 1214 9933
rect 1182 9848 1214 9913
rect 1394 9904 1425 10103
rect 1626 10098 1661 10103
rect 1626 10078 1633 10098
rect 1653 10078 1661 10098
rect 1626 10070 1661 10078
rect 1394 9874 1400 9904
rect 1421 9874 1425 9904
rect 1394 9866 1425 9874
rect 1552 9848 1592 9849
rect 1182 9846 1594 9848
rect 1182 9820 1562 9846
rect 1588 9820 1594 9846
rect 1182 9812 1594 9820
rect 1182 9784 1214 9812
rect 1627 9792 1661 10070
rect 1743 9883 1813 10199
rect 3731 10184 3762 10185
rect 3731 10176 3776 10184
rect 2811 10153 2975 10160
rect 3731 10153 3741 10176
rect 2437 10138 3741 10153
rect 3766 10138 3776 10176
rect 2437 10120 3776 10138
rect 2442 10107 2478 10120
rect 2811 10117 2975 10120
rect 1852 10038 2055 10051
rect 1852 10005 1876 10038
rect 1912 10037 2055 10038
rect 1912 10034 2023 10037
rect 1912 10007 1949 10034
rect 1978 10010 2023 10034
rect 2052 10010 2055 10037
rect 1978 10007 2055 10010
rect 1912 10005 2055 10007
rect 1852 9992 2055 10005
rect 1852 9991 1953 9992
rect 1182 9764 1187 9784
rect 1208 9764 1214 9784
rect 1182 9757 1214 9764
rect 1605 9787 1661 9792
rect 1605 9767 1612 9787
rect 1632 9767 1661 9787
rect 1738 9877 1813 9883
rect 1738 9844 1746 9877
rect 1799 9844 1813 9877
rect 1738 9819 1813 9844
rect 1738 9786 1751 9819
rect 1804 9786 1813 9819
rect 1738 9777 1813 9786
rect 2230 9929 2262 9936
rect 2230 9909 2237 9929
rect 2258 9909 2262 9929
rect 2230 9844 2262 9909
rect 2442 9900 2473 10107
rect 2677 10099 2709 10100
rect 2674 10094 2709 10099
rect 2674 10074 2681 10094
rect 2701 10074 2709 10094
rect 2674 10066 2709 10074
rect 2442 9870 2448 9900
rect 2469 9870 2473 9900
rect 2442 9862 2473 9870
rect 2600 9844 2640 9845
rect 2230 9842 2642 9844
rect 2230 9816 2610 9842
rect 2636 9816 2642 9842
rect 2230 9808 2642 9816
rect 2230 9780 2262 9808
rect 2675 9788 2709 10066
rect 1738 9772 1796 9777
rect 1605 9760 1661 9767
rect 2230 9760 2235 9780
rect 2256 9760 2262 9780
rect 1605 9759 1640 9760
rect 2230 9753 2262 9760
rect 2653 9783 2709 9788
rect 2653 9763 2660 9783
rect 2680 9763 2709 9783
rect 2653 9756 2709 9763
rect 2653 9755 2688 9756
rect 896 9704 1007 9708
rect 2679 9704 3979 9705
rect 218 9686 3979 9704
rect 218 9666 904 9686
rect 923 9666 981 9686
rect 1000 9682 3979 9686
rect 1000 9666 1952 9682
rect 218 9662 1952 9666
rect 1971 9662 2029 9682
rect 2048 9662 3979 9682
rect 218 9648 3979 9662
rect 218 9025 325 9648
rect 1944 9645 2055 9648
rect 704 9599 768 9603
rect 700 9593 768 9599
rect 700 9560 717 9593
rect 757 9560 768 9593
rect 700 9548 768 9560
rect 1751 9562 1816 9584
rect 700 9546 757 9548
rect 704 9185 755 9546
rect 1751 9523 1768 9562
rect 1813 9523 1816 9562
rect 1392 9478 1427 9480
rect 1392 9469 1496 9478
rect 1392 9468 1443 9469
rect 1392 9448 1395 9468
rect 1420 9449 1443 9468
rect 1475 9449 1496 9469
rect 1420 9448 1496 9449
rect 1392 9441 1496 9448
rect 1392 9429 1427 9441
rect 804 9363 1007 9376
rect 804 9330 828 9363
rect 864 9362 1007 9363
rect 864 9359 975 9362
rect 864 9332 901 9359
rect 930 9335 975 9359
rect 1004 9335 1007 9362
rect 930 9332 1007 9335
rect 864 9330 1007 9332
rect 804 9317 1007 9330
rect 804 9316 905 9317
rect 1182 9254 1214 9261
rect 1182 9234 1189 9254
rect 1210 9234 1214 9254
rect 693 9176 758 9185
rect 693 9139 703 9176
rect 743 9142 758 9176
rect 1182 9169 1214 9234
rect 1394 9225 1425 9429
rect 1629 9424 1661 9425
rect 1626 9419 1661 9424
rect 1626 9399 1633 9419
rect 1653 9399 1661 9419
rect 1626 9391 1661 9399
rect 1394 9195 1400 9225
rect 1421 9195 1425 9225
rect 1394 9187 1425 9195
rect 1552 9169 1592 9170
rect 1182 9167 1594 9169
rect 743 9139 760 9142
rect 693 9120 760 9139
rect 693 9099 707 9120
rect 743 9099 760 9120
rect 693 9092 760 9099
rect 1182 9141 1562 9167
rect 1588 9141 1594 9167
rect 1182 9133 1594 9141
rect 1182 9105 1214 9133
rect 1627 9113 1661 9391
rect 1751 9223 1816 9523
rect 3888 9484 3925 9505
rect 3888 9447 3899 9484
rect 3916 9460 3925 9484
rect 3916 9447 3926 9460
rect 3888 9437 3926 9447
rect 3889 9433 3926 9437
rect 3889 9427 3922 9433
rect 3299 9358 3502 9371
rect 3299 9325 3323 9358
rect 3359 9357 3502 9358
rect 3359 9354 3470 9357
rect 3359 9327 3396 9354
rect 3425 9330 3470 9354
rect 3499 9330 3502 9357
rect 3425 9327 3502 9330
rect 3359 9325 3502 9327
rect 3299 9312 3502 9325
rect 3299 9311 3400 9312
rect 3677 9249 3709 9256
rect 3677 9229 3684 9249
rect 3705 9229 3709 9249
rect 1182 9085 1187 9105
rect 1208 9085 1214 9105
rect 1182 9078 1214 9085
rect 1605 9108 1661 9113
rect 1605 9088 1612 9108
rect 1632 9088 1661 9108
rect 1605 9081 1661 9088
rect 1741 9212 1821 9223
rect 1741 9186 1758 9212
rect 1798 9186 1821 9212
rect 1741 9159 1821 9186
rect 1741 9133 1762 9159
rect 1802 9133 1821 9159
rect 3677 9164 3709 9229
rect 3889 9220 3920 9427
rect 4124 9419 4156 9420
rect 4121 9414 4156 9419
rect 4121 9394 4128 9414
rect 4148 9394 4156 9414
rect 4121 9386 4156 9394
rect 3889 9190 3895 9220
rect 3916 9190 3920 9220
rect 3889 9182 3920 9190
rect 4047 9164 4087 9165
rect 3677 9162 4089 9164
rect 1741 9114 1821 9133
rect 1741 9088 1765 9114
rect 1805 9088 1821 9114
rect 2854 9152 3291 9158
rect 2854 9129 2872 9152
rect 2898 9145 3291 9152
rect 2898 9129 3252 9145
rect 2854 9122 3252 9129
rect 3278 9122 3291 9145
rect 2854 9109 3291 9122
rect 3677 9136 4057 9162
rect 4083 9136 4089 9162
rect 3677 9128 4089 9136
rect 1605 9080 1640 9081
rect 1741 9076 1821 9088
rect 3677 9100 3709 9128
rect 4122 9108 4156 9386
rect 3677 9080 3682 9100
rect 3703 9080 3709 9100
rect 3677 9073 3709 9080
rect 4100 9103 4156 9108
rect 4100 9083 4107 9103
rect 4127 9083 4156 9103
rect 4100 9076 4156 9083
rect 4100 9075 4135 9076
rect 896 9025 1007 9029
rect 2638 9025 4188 9028
rect 216 9007 4188 9025
rect 216 8987 904 9007
rect 923 8987 981 9007
rect 1000 9002 4188 9007
rect 1000 8987 3399 9002
rect 216 8982 3399 8987
rect 3418 8982 3476 9002
rect 3495 8982 4188 9002
rect 216 8972 4188 8982
rect 216 8969 841 8972
rect 1028 8969 4188 8972
rect 218 8741 325 8969
rect 2638 8968 4188 8969
rect 3391 8965 3502 8968
rect 686 8930 807 8940
rect 686 8928 755 8930
rect 686 8887 699 8928
rect 736 8889 755 8928
rect 792 8889 807 8930
rect 736 8887 807 8889
rect 686 8869 807 8887
rect 692 8767 771 8869
rect 1744 8829 1811 8848
rect 1744 8809 1764 8829
rect 218 8686 326 8741
rect 693 8686 771 8767
rect 1743 8763 1764 8809
rect 1794 8809 1811 8829
rect 1794 8779 1813 8809
rect 1794 8763 1814 8779
rect 1743 8747 1814 8763
rect 1393 8736 1465 8737
rect 1392 8728 1491 8736
rect 1392 8725 1444 8728
rect 1392 8690 1400 8725
rect 1425 8690 1444 8725
rect 1469 8690 1491 8728
rect 218 8257 325 8686
rect 697 8445 769 8686
rect 1392 8678 1491 8690
rect 1393 8659 1461 8678
rect 1394 8656 1427 8659
rect 1629 8656 1661 8657
rect 804 8595 1007 8608
rect 804 8562 828 8595
rect 864 8594 1007 8595
rect 864 8591 975 8594
rect 864 8564 901 8591
rect 930 8567 975 8591
rect 1004 8567 1007 8594
rect 930 8564 1007 8567
rect 864 8562 1007 8564
rect 804 8549 1007 8562
rect 804 8548 905 8549
rect 697 8403 706 8445
rect 755 8403 769 8445
rect 697 8382 769 8403
rect 697 8340 707 8382
rect 756 8340 769 8382
rect 697 8322 769 8340
rect 1182 8486 1214 8493
rect 1182 8466 1189 8486
rect 1210 8466 1214 8486
rect 1182 8401 1214 8466
rect 1394 8457 1425 8656
rect 1626 8651 1661 8656
rect 1626 8631 1633 8651
rect 1653 8631 1661 8651
rect 1626 8623 1661 8631
rect 1394 8427 1400 8457
rect 1421 8427 1425 8457
rect 1394 8419 1425 8427
rect 1552 8401 1592 8402
rect 1182 8399 1594 8401
rect 1182 8373 1562 8399
rect 1588 8373 1594 8399
rect 1182 8365 1594 8373
rect 1182 8337 1214 8365
rect 1627 8345 1661 8623
rect 1743 8436 1813 8747
rect 2440 8738 3782 8743
rect 2440 8736 3739 8738
rect 2437 8710 3739 8736
rect 3767 8710 3782 8738
rect 2437 8702 3782 8710
rect 2437 8677 2476 8702
rect 2437 8660 2478 8677
rect 2437 8653 2476 8660
rect 1852 8591 2055 8604
rect 1852 8558 1876 8591
rect 1912 8590 2055 8591
rect 1912 8587 2023 8590
rect 1912 8560 1949 8587
rect 1978 8563 2023 8587
rect 2052 8563 2055 8590
rect 1978 8560 2055 8563
rect 1912 8558 2055 8560
rect 1852 8545 2055 8558
rect 1852 8544 1953 8545
rect 1182 8317 1187 8337
rect 1208 8317 1214 8337
rect 1182 8310 1214 8317
rect 1605 8340 1661 8345
rect 1605 8320 1612 8340
rect 1632 8320 1661 8340
rect 1738 8430 1813 8436
rect 1738 8397 1746 8430
rect 1799 8397 1813 8430
rect 1738 8372 1813 8397
rect 1738 8339 1751 8372
rect 1804 8339 1813 8372
rect 1738 8330 1813 8339
rect 2230 8482 2262 8489
rect 2230 8462 2237 8482
rect 2258 8462 2262 8482
rect 2230 8397 2262 8462
rect 2442 8453 2473 8653
rect 2677 8652 2709 8653
rect 2674 8647 2709 8652
rect 2674 8627 2681 8647
rect 2701 8627 2709 8647
rect 2674 8619 2709 8627
rect 2442 8423 2448 8453
rect 2469 8423 2473 8453
rect 2442 8415 2473 8423
rect 2600 8397 2640 8398
rect 2230 8395 2642 8397
rect 2230 8369 2610 8395
rect 2636 8369 2642 8395
rect 2230 8361 2642 8369
rect 2230 8333 2262 8361
rect 2675 8341 2709 8619
rect 1738 8325 1796 8330
rect 1605 8313 1661 8320
rect 2230 8313 2235 8333
rect 2256 8313 2262 8333
rect 1605 8312 1640 8313
rect 2230 8306 2262 8313
rect 2653 8336 2709 8341
rect 2653 8316 2660 8336
rect 2680 8316 2709 8336
rect 2653 8309 2709 8316
rect 2653 8308 2688 8309
rect 896 8257 1007 8261
rect 2771 8257 3761 8258
rect 218 8239 3761 8257
rect 218 8219 904 8239
rect 923 8219 981 8239
rect 1000 8235 3761 8239
rect 1000 8219 1952 8235
rect 218 8215 1952 8219
rect 1971 8215 2029 8235
rect 2048 8215 3761 8235
rect 218 8201 3761 8215
rect 218 7578 325 8201
rect 1944 8198 2055 8201
rect 704 8152 768 8156
rect 700 8146 768 8152
rect 700 8113 717 8146
rect 757 8113 768 8146
rect 700 8101 768 8113
rect 1751 8115 1816 8137
rect 700 8099 757 8101
rect 704 7738 755 8099
rect 1751 8076 1768 8115
rect 1813 8076 1816 8115
rect 1392 8031 1427 8033
rect 1392 8022 1496 8031
rect 1392 8021 1443 8022
rect 1392 8001 1395 8021
rect 1420 8002 1443 8021
rect 1475 8002 1496 8022
rect 1420 8001 1496 8002
rect 1392 7994 1496 8001
rect 1392 7982 1427 7994
rect 804 7916 1007 7929
rect 804 7883 828 7916
rect 864 7915 1007 7916
rect 864 7912 975 7915
rect 864 7885 901 7912
rect 930 7888 975 7912
rect 1004 7888 1007 7915
rect 930 7885 1007 7888
rect 864 7883 1007 7885
rect 804 7870 1007 7883
rect 804 7869 905 7870
rect 1182 7807 1214 7814
rect 1182 7787 1189 7807
rect 1210 7787 1214 7807
rect 693 7729 758 7738
rect 693 7692 703 7729
rect 743 7695 758 7729
rect 1182 7722 1214 7787
rect 1394 7778 1425 7982
rect 1629 7977 1661 7978
rect 1626 7972 1661 7977
rect 1626 7952 1633 7972
rect 1653 7952 1661 7972
rect 1626 7944 1661 7952
rect 1394 7748 1400 7778
rect 1421 7748 1425 7778
rect 1394 7740 1425 7748
rect 1552 7722 1592 7723
rect 1182 7720 1594 7722
rect 743 7692 760 7695
rect 693 7673 760 7692
rect 693 7652 707 7673
rect 743 7652 760 7673
rect 693 7645 760 7652
rect 1182 7694 1562 7720
rect 1588 7694 1594 7720
rect 1182 7686 1594 7694
rect 1182 7658 1214 7686
rect 1627 7666 1661 7944
rect 1751 7776 1816 8076
rect 1182 7638 1187 7658
rect 1208 7638 1214 7658
rect 1182 7631 1214 7638
rect 1605 7661 1661 7666
rect 1605 7641 1612 7661
rect 1632 7641 1661 7661
rect 1605 7634 1661 7641
rect 1741 7765 1821 7776
rect 1741 7739 1758 7765
rect 1798 7739 1821 7765
rect 1741 7712 1821 7739
rect 4293 7715 4342 12901
rect 4790 12898 4948 12901
rect 4810 12890 4948 12898
rect 5330 12343 5438 13473
rect 16049 13470 16069 13522
rect 16147 13470 16160 13528
rect 16049 13457 16160 13470
rect 14992 13389 15079 13407
rect 14992 13345 15009 13389
rect 15061 13345 15079 13389
rect 14992 13328 15079 13345
rect 13734 13285 13815 13286
rect 13728 13271 13827 13285
rect 13728 13221 13748 13271
rect 13800 13221 13827 13271
rect 13728 13201 13827 13221
rect 9931 13088 9996 13171
rect 9881 13070 10002 13088
rect 9881 13068 9952 13070
rect 9881 13027 9896 13068
rect 9933 13029 9952 13068
rect 9989 13029 10002 13070
rect 9933 13027 10002 13029
rect 9881 13017 10002 13027
rect 6397 12988 7875 12990
rect 10362 12988 11039 13012
rect 6397 12983 9557 12988
rect 9815 12983 11039 12988
rect 6397 12970 11039 12983
rect 6397 12950 9688 12970
rect 9707 12950 9765 12970
rect 9784 12950 11039 12970
rect 6397 12932 11039 12950
rect 7830 12931 8037 12932
rect 9681 12928 9792 12932
rect 10362 12924 11039 12932
rect 8867 12869 8947 12881
rect 9048 12876 9083 12877
rect 8867 12843 8883 12869
rect 8923 12843 8947 12869
rect 8867 12824 8947 12843
rect 8867 12798 8886 12824
rect 8926 12798 8947 12824
rect 8867 12771 8947 12798
rect 8867 12745 8890 12771
rect 8930 12745 8947 12771
rect 8867 12734 8947 12745
rect 9027 12869 9083 12876
rect 9027 12849 9056 12869
rect 9076 12849 9083 12869
rect 9027 12844 9083 12849
rect 9474 12872 9506 12879
rect 9474 12852 9480 12872
rect 9501 12852 9506 12872
rect 8872 12434 8937 12734
rect 9027 12566 9061 12844
rect 9474 12824 9506 12852
rect 9094 12816 9506 12824
rect 9094 12790 9100 12816
rect 9126 12790 9506 12816
rect 9928 12858 9995 12865
rect 9928 12837 9945 12858
rect 9981 12837 9995 12858
rect 9928 12818 9995 12837
rect 9928 12815 9945 12818
rect 9094 12788 9506 12790
rect 9096 12787 9136 12788
rect 9263 12762 9294 12770
rect 9263 12732 9267 12762
rect 9288 12732 9294 12762
rect 9027 12558 9062 12566
rect 9027 12538 9035 12558
rect 9055 12538 9062 12558
rect 9027 12533 9062 12538
rect 9027 12532 9059 12533
rect 9263 12528 9294 12732
rect 9474 12723 9506 12788
rect 9930 12781 9945 12815
rect 9985 12781 9995 12818
rect 9930 12772 9995 12781
rect 9474 12703 9478 12723
rect 9499 12703 9506 12723
rect 9474 12696 9506 12703
rect 9783 12640 9884 12641
rect 9681 12627 9884 12640
rect 9681 12625 9824 12627
rect 9681 12622 9758 12625
rect 9681 12595 9684 12622
rect 9713 12598 9758 12622
rect 9787 12598 9824 12625
rect 9713 12595 9824 12598
rect 9681 12594 9824 12595
rect 9860 12594 9884 12627
rect 9681 12581 9884 12594
rect 9261 12516 9296 12528
rect 9192 12509 9296 12516
rect 9192 12508 9268 12509
rect 9192 12488 9213 12508
rect 9245 12489 9268 12508
rect 9293 12489 9296 12509
rect 9245 12488 9296 12489
rect 9192 12479 9296 12488
rect 9261 12477 9296 12479
rect 8872 12395 8875 12434
rect 8920 12395 8937 12434
rect 9933 12411 9984 12772
rect 9931 12409 9988 12411
rect 8872 12373 8937 12395
rect 9920 12397 9988 12409
rect 9920 12364 9931 12397
rect 9971 12364 9988 12397
rect 9920 12358 9988 12364
rect 9920 12354 9984 12358
rect 4407 7907 4610 7920
rect 4407 7874 4431 7907
rect 4467 7906 4610 7907
rect 4467 7903 4578 7906
rect 4467 7876 4504 7903
rect 4533 7879 4578 7903
rect 4607 7879 4610 7906
rect 4533 7876 4610 7879
rect 4467 7874 4610 7876
rect 4407 7861 4610 7874
rect 4407 7860 4508 7861
rect 4785 7798 4817 7805
rect 4785 7778 4792 7798
rect 4813 7778 4817 7798
rect 1741 7686 1762 7712
rect 1802 7686 1821 7712
rect 1741 7667 1821 7686
rect 4292 7705 4403 7715
rect 4292 7704 4357 7705
rect 4292 7680 4300 7704
rect 4324 7681 4357 7704
rect 4381 7681 4403 7705
rect 4324 7680 4403 7681
rect 4292 7673 4403 7680
rect 4785 7713 4817 7778
rect 4997 7769 5028 7969
rect 5232 7968 5264 7969
rect 5229 7963 5264 7968
rect 5229 7943 5236 7963
rect 5256 7943 5264 7963
rect 5229 7935 5264 7943
rect 4997 7739 5003 7769
rect 5024 7739 5028 7769
rect 4997 7731 5028 7739
rect 5155 7713 5195 7714
rect 4785 7711 5197 7713
rect 4785 7685 5165 7711
rect 5191 7685 5197 7711
rect 4785 7677 5197 7685
rect 1741 7641 1765 7667
rect 1805 7641 1821 7667
rect 1605 7633 1640 7634
rect 1741 7629 1821 7641
rect 4785 7649 4817 7677
rect 5230 7657 5264 7935
rect 4785 7629 4790 7649
rect 4811 7629 4817 7649
rect 4785 7622 4817 7629
rect 4996 7649 5030 7656
rect 4996 7627 5003 7649
rect 5027 7627 5030 7649
rect 896 7578 1007 7582
rect 2651 7578 2858 7579
rect 216 7573 4291 7578
rect 216 7560 4610 7573
rect 216 7540 904 7560
rect 923 7540 981 7560
rect 1000 7551 4610 7560
rect 1000 7540 4507 7551
rect 216 7531 4507 7540
rect 4526 7531 4584 7551
rect 4603 7531 4610 7551
rect 216 7522 4610 7531
rect 218 7349 325 7522
rect 2813 7520 4610 7522
rect 4499 7514 4610 7520
rect 686 7483 807 7493
rect 686 7481 755 7483
rect 686 7440 699 7481
rect 736 7442 755 7481
rect 792 7442 807 7483
rect 736 7440 807 7442
rect 686 7422 807 7440
rect 4834 7472 4886 7503
rect 4834 7438 4843 7472
rect 4872 7438 4886 7472
rect 209 7322 325 7349
rect 692 7330 757 7422
rect 4834 7412 4886 7438
rect 4996 7421 5030 7627
rect 5208 7652 5264 7657
rect 5208 7632 5215 7652
rect 5235 7632 5264 7652
rect 5208 7625 5264 7632
rect 5208 7624 5243 7625
rect 209 7183 320 7322
rect 690 7284 757 7330
rect 1742 7368 1814 7390
rect 1742 7320 1756 7368
rect 1802 7363 1814 7368
rect 4834 7378 4842 7412
rect 4871 7378 4886 7412
rect 1802 7320 1819 7363
rect 690 7183 755 7284
rect 209 7123 322 7183
rect 690 7145 766 7183
rect 215 6663 322 7123
rect 694 6851 766 7145
rect 1390 7142 1462 7143
rect 1389 7134 1488 7142
rect 1742 7137 1819 7320
rect 3030 7321 3114 7332
rect 3030 7293 3058 7321
rect 3102 7293 3114 7321
rect 2844 7242 2918 7270
rect 2844 7194 2867 7242
rect 2904 7194 2918 7242
rect 3030 7264 3114 7293
rect 3030 7236 3055 7264
rect 3099 7236 3114 7264
rect 3030 7203 3114 7236
rect 2844 7185 2918 7194
rect 2440 7143 2512 7144
rect 1389 7131 1441 7134
rect 1389 7096 1397 7131
rect 1422 7096 1441 7131
rect 1466 7096 1488 7134
rect 1389 7084 1488 7096
rect 1740 7108 1819 7137
rect 2439 7135 2528 7143
rect 2439 7132 2491 7135
rect 1390 7065 1458 7084
rect 1391 7062 1424 7065
rect 1626 7062 1658 7063
rect 801 7001 1004 7014
rect 801 6968 825 7001
rect 861 7000 1004 7001
rect 861 6997 972 7000
rect 861 6970 898 6997
rect 927 6973 972 6997
rect 1001 6973 1004 7000
rect 927 6970 1004 6973
rect 861 6968 1004 6970
rect 801 6955 1004 6968
rect 801 6954 902 6955
rect 694 6809 703 6851
rect 752 6809 766 6851
rect 694 6788 766 6809
rect 694 6746 704 6788
rect 753 6746 766 6788
rect 694 6728 766 6746
rect 1179 6892 1211 6899
rect 1179 6872 1186 6892
rect 1207 6872 1211 6892
rect 1179 6807 1211 6872
rect 1391 6863 1422 7062
rect 1623 7057 1658 7062
rect 1623 7037 1630 7057
rect 1650 7037 1658 7057
rect 1623 7029 1658 7037
rect 1391 6833 1397 6863
rect 1418 6833 1422 6863
rect 1391 6825 1422 6833
rect 1549 6807 1589 6808
rect 1179 6805 1591 6807
rect 1179 6779 1559 6805
rect 1585 6779 1591 6805
rect 1179 6771 1591 6779
rect 1179 6743 1211 6771
rect 1624 6751 1658 7029
rect 1740 6842 1810 7108
rect 2439 7097 2447 7132
rect 2472 7097 2491 7132
rect 2516 7097 2528 7135
rect 2439 7085 2528 7097
rect 2439 7084 2508 7085
rect 2439 7066 2475 7084
rect 1849 6997 2052 7010
rect 1849 6964 1873 6997
rect 1909 6996 2052 6997
rect 1909 6993 2020 6996
rect 1909 6966 1946 6993
rect 1975 6969 2020 6993
rect 2049 6969 2052 6996
rect 1975 6966 2052 6969
rect 1909 6964 2052 6966
rect 1849 6951 2052 6964
rect 1849 6950 1950 6951
rect 1179 6723 1184 6743
rect 1205 6723 1211 6743
rect 1179 6716 1211 6723
rect 1602 6746 1658 6751
rect 1602 6726 1609 6746
rect 1629 6726 1658 6746
rect 1735 6836 1810 6842
rect 1735 6803 1743 6836
rect 1796 6803 1810 6836
rect 1735 6778 1810 6803
rect 1735 6745 1748 6778
rect 1801 6745 1810 6778
rect 1735 6736 1810 6745
rect 2227 6888 2259 6895
rect 2227 6868 2234 6888
rect 2255 6868 2259 6888
rect 2227 6803 2259 6868
rect 2439 6859 2470 7066
rect 2674 7058 2706 7059
rect 2671 7053 2706 7058
rect 2671 7033 2678 7053
rect 2698 7033 2706 7053
rect 2671 7025 2706 7033
rect 2439 6829 2445 6859
rect 2466 6829 2470 6859
rect 2439 6821 2470 6829
rect 2597 6803 2637 6804
rect 2227 6801 2639 6803
rect 2227 6775 2607 6801
rect 2633 6775 2639 6801
rect 2227 6767 2639 6775
rect 2227 6739 2259 6767
rect 2672 6747 2706 7025
rect 2855 6840 2917 7185
rect 3024 7158 3114 7203
rect 3024 6843 3106 7158
rect 2855 6821 2919 6840
rect 2855 6782 2868 6821
rect 2902 6782 2919 6821
rect 2855 6763 2919 6782
rect 3024 6802 3045 6843
rect 3081 6802 3106 6843
rect 3024 6773 3106 6802
rect 1735 6731 1793 6736
rect 1602 6719 1658 6726
rect 2227 6719 2232 6739
rect 2253 6719 2259 6739
rect 1602 6718 1637 6719
rect 2227 6712 2259 6719
rect 2650 6742 2706 6747
rect 2650 6722 2657 6742
rect 2677 6722 2706 6742
rect 2650 6715 2706 6722
rect 2650 6714 2685 6715
rect 893 6663 1004 6667
rect 2676 6663 4246 6664
rect 215 6645 4246 6663
rect 215 6625 901 6645
rect 920 6625 978 6645
rect 997 6641 4246 6645
rect 997 6625 1949 6641
rect 215 6621 1949 6625
rect 1968 6621 2026 6641
rect 2045 6621 4246 6641
rect 215 6607 4246 6621
rect 215 5984 322 6607
rect 1941 6604 2052 6607
rect 701 6558 765 6562
rect 697 6552 765 6558
rect 697 6519 714 6552
rect 754 6519 765 6552
rect 697 6507 765 6519
rect 1748 6521 1813 6543
rect 697 6505 754 6507
rect 701 6144 752 6505
rect 1748 6482 1765 6521
rect 1810 6482 1813 6521
rect 1389 6437 1424 6439
rect 1389 6428 1493 6437
rect 1389 6427 1440 6428
rect 1389 6407 1392 6427
rect 1417 6408 1440 6427
rect 1472 6408 1493 6428
rect 1417 6407 1493 6408
rect 1389 6400 1493 6407
rect 1389 6388 1424 6400
rect 801 6322 1004 6335
rect 801 6289 825 6322
rect 861 6321 1004 6322
rect 861 6318 972 6321
rect 861 6291 898 6318
rect 927 6294 972 6318
rect 1001 6294 1004 6321
rect 927 6291 1004 6294
rect 861 6289 1004 6291
rect 801 6276 1004 6289
rect 801 6275 902 6276
rect 1179 6213 1211 6220
rect 1179 6193 1186 6213
rect 1207 6193 1211 6213
rect 690 6135 755 6144
rect 690 6098 700 6135
rect 740 6101 755 6135
rect 1179 6128 1211 6193
rect 1391 6184 1422 6388
rect 1626 6383 1658 6384
rect 1623 6378 1658 6383
rect 1623 6358 1630 6378
rect 1650 6358 1658 6378
rect 1623 6350 1658 6358
rect 1391 6154 1397 6184
rect 1418 6154 1422 6184
rect 1391 6146 1422 6154
rect 1549 6128 1589 6129
rect 1179 6126 1591 6128
rect 740 6098 757 6101
rect 690 6079 757 6098
rect 690 6058 704 6079
rect 740 6058 757 6079
rect 690 6051 757 6058
rect 1179 6100 1559 6126
rect 1585 6100 1591 6126
rect 1179 6092 1591 6100
rect 1179 6064 1211 6092
rect 1624 6072 1658 6350
rect 1748 6182 1813 6482
rect 3019 6506 3112 6521
rect 3019 6462 3034 6506
rect 3094 6462 3112 6506
rect 1179 6044 1184 6064
rect 1205 6044 1211 6064
rect 1179 6037 1211 6044
rect 1602 6067 1658 6072
rect 1602 6047 1609 6067
rect 1629 6047 1658 6067
rect 1602 6040 1658 6047
rect 1738 6171 1818 6182
rect 1738 6145 1755 6171
rect 1795 6145 1818 6171
rect 1738 6118 1818 6145
rect 1738 6092 1759 6118
rect 1799 6092 1818 6118
rect 1738 6073 1818 6092
rect 1738 6047 1762 6073
rect 1802 6047 1818 6073
rect 1602 6039 1637 6040
rect 1738 6035 1818 6047
rect 3019 6089 3112 6462
rect 3296 6317 3499 6330
rect 3296 6284 3320 6317
rect 3356 6316 3499 6317
rect 3356 6313 3467 6316
rect 3356 6286 3393 6313
rect 3422 6289 3467 6313
rect 3496 6289 3499 6316
rect 3422 6286 3499 6289
rect 3356 6284 3499 6286
rect 3296 6271 3499 6284
rect 3296 6270 3397 6271
rect 3019 6048 3034 6089
rect 3088 6048 3112 6089
rect 3019 6041 3112 6048
rect 3674 6208 3706 6215
rect 3674 6188 3681 6208
rect 3702 6188 3706 6208
rect 3674 6123 3706 6188
rect 3886 6179 3917 6380
rect 4121 6378 4153 6379
rect 4118 6373 4153 6378
rect 4118 6353 4125 6373
rect 4145 6353 4153 6373
rect 4118 6345 4153 6353
rect 3886 6149 3892 6179
rect 3913 6149 3917 6179
rect 3886 6141 3917 6149
rect 4044 6123 4084 6124
rect 3674 6121 4086 6123
rect 3674 6095 4054 6121
rect 4080 6095 4086 6121
rect 3674 6087 4086 6095
rect 3674 6059 3706 6087
rect 4119 6067 4153 6345
rect 3674 6039 3679 6059
rect 3700 6039 3706 6059
rect 3674 6032 3706 6039
rect 4097 6062 4153 6067
rect 4097 6042 4104 6062
rect 4124 6042 4153 6062
rect 4097 6035 4153 6042
rect 4097 6034 4132 6035
rect 893 5984 1004 5988
rect 2635 5984 4279 5987
rect 213 5966 4279 5984
rect 213 5946 901 5966
rect 920 5946 978 5966
rect 997 5961 4279 5966
rect 997 5946 3396 5961
rect 213 5941 3396 5946
rect 3415 5941 3473 5961
rect 3492 5941 4279 5961
rect 213 5931 4279 5941
rect 213 5928 838 5931
rect 1025 5928 4279 5931
rect 215 5700 322 5928
rect 2635 5927 4279 5928
rect 3388 5924 3499 5927
rect 683 5889 804 5899
rect 683 5887 752 5889
rect 683 5846 696 5887
rect 733 5848 752 5887
rect 789 5848 804 5889
rect 733 5846 804 5848
rect 683 5828 804 5846
rect 3888 5869 3974 5873
rect 3888 5851 3903 5869
rect 3955 5851 3974 5869
rect 3888 5842 3974 5851
rect 689 5726 768 5828
rect 1741 5788 1808 5807
rect 1741 5768 1761 5788
rect 215 5645 323 5700
rect 690 5645 768 5726
rect 1740 5722 1761 5768
rect 1791 5768 1808 5788
rect 1791 5738 1810 5768
rect 1791 5722 1811 5738
rect 1740 5706 1811 5722
rect 1390 5695 1462 5696
rect 1389 5687 1488 5695
rect 1389 5684 1441 5687
rect 1389 5649 1397 5684
rect 1422 5649 1441 5684
rect 1466 5649 1488 5687
rect 215 5216 322 5645
rect 694 5404 766 5645
rect 1389 5637 1488 5649
rect 1390 5618 1458 5637
rect 1391 5615 1424 5618
rect 1626 5615 1658 5616
rect 801 5554 1004 5567
rect 801 5521 825 5554
rect 861 5553 1004 5554
rect 861 5550 972 5553
rect 861 5523 898 5550
rect 927 5526 972 5550
rect 1001 5526 1004 5553
rect 927 5523 1004 5526
rect 861 5521 1004 5523
rect 801 5508 1004 5521
rect 801 5507 902 5508
rect 694 5362 703 5404
rect 752 5362 766 5404
rect 694 5341 766 5362
rect 694 5299 704 5341
rect 753 5299 766 5341
rect 694 5281 766 5299
rect 1179 5445 1211 5452
rect 1179 5425 1186 5445
rect 1207 5425 1211 5445
rect 1179 5360 1211 5425
rect 1391 5416 1422 5615
rect 1623 5610 1658 5615
rect 1623 5590 1630 5610
rect 1650 5590 1658 5610
rect 1623 5582 1658 5590
rect 1391 5386 1397 5416
rect 1418 5386 1422 5416
rect 1391 5378 1422 5386
rect 1549 5360 1589 5361
rect 1179 5358 1591 5360
rect 1179 5332 1559 5358
rect 1585 5332 1591 5358
rect 1179 5324 1591 5332
rect 1179 5296 1211 5324
rect 1624 5304 1658 5582
rect 1740 5395 1810 5706
rect 3665 5696 3737 5697
rect 3664 5693 3753 5696
rect 2436 5691 3753 5693
rect 2433 5688 3753 5691
rect 2433 5685 3716 5688
rect 2433 5650 3672 5685
rect 3697 5650 3716 5685
rect 3741 5650 3753 5688
rect 2433 5640 3753 5650
rect 3929 5689 3965 5842
rect 3929 5666 3935 5689
rect 3959 5666 3965 5689
rect 3929 5645 3965 5666
rect 2433 5638 3718 5640
rect 2433 5628 2530 5638
rect 2439 5619 2475 5628
rect 3929 5622 3935 5645
rect 3959 5622 3965 5645
rect 1849 5550 2052 5563
rect 1849 5517 1873 5550
rect 1909 5549 2052 5550
rect 1909 5546 2020 5549
rect 1909 5519 1946 5546
rect 1975 5522 2020 5546
rect 2049 5522 2052 5549
rect 1975 5519 2052 5522
rect 1909 5517 2052 5519
rect 1849 5504 2052 5517
rect 1849 5503 1950 5504
rect 1179 5276 1184 5296
rect 1205 5276 1211 5296
rect 1179 5269 1211 5276
rect 1602 5299 1658 5304
rect 1602 5279 1609 5299
rect 1629 5279 1658 5299
rect 1735 5389 1810 5395
rect 1735 5356 1743 5389
rect 1796 5356 1810 5389
rect 1735 5331 1810 5356
rect 1735 5298 1748 5331
rect 1801 5298 1810 5331
rect 1735 5289 1810 5298
rect 2227 5441 2259 5448
rect 2227 5421 2234 5441
rect 2255 5421 2259 5441
rect 2227 5356 2259 5421
rect 2439 5412 2470 5619
rect 2674 5611 2706 5612
rect 3929 5611 3965 5622
rect 2671 5606 2706 5611
rect 2671 5586 2678 5606
rect 2698 5586 2706 5606
rect 2671 5578 2706 5586
rect 2439 5382 2445 5412
rect 2466 5382 2470 5412
rect 2439 5374 2470 5382
rect 2597 5356 2637 5357
rect 2227 5354 2639 5356
rect 2227 5328 2607 5354
rect 2633 5328 2639 5354
rect 2227 5320 2639 5328
rect 2227 5292 2259 5320
rect 2672 5300 2706 5578
rect 1735 5284 1793 5289
rect 1602 5272 1658 5279
rect 2227 5272 2232 5292
rect 2253 5272 2259 5292
rect 1602 5271 1637 5272
rect 2227 5265 2259 5272
rect 2650 5295 2706 5300
rect 2650 5275 2657 5295
rect 2677 5275 2706 5295
rect 2650 5268 2706 5275
rect 2650 5267 2685 5268
rect 893 5216 1004 5220
rect 2768 5216 3927 5217
rect 215 5198 3927 5216
rect 215 5178 901 5198
rect 920 5178 978 5198
rect 997 5194 3927 5198
rect 997 5178 1949 5194
rect 215 5174 1949 5178
rect 1968 5174 2026 5194
rect 2045 5174 3927 5194
rect 215 5160 3927 5174
rect 215 4537 322 5160
rect 1941 5157 2052 5160
rect 701 5111 765 5115
rect 697 5105 765 5111
rect 697 5072 714 5105
rect 754 5072 765 5105
rect 697 5060 765 5072
rect 1748 5074 1813 5096
rect 697 5058 754 5060
rect 701 4697 752 5058
rect 1748 5035 1765 5074
rect 1810 5035 1813 5074
rect 4834 5072 4886 7378
rect 4995 7355 5030 7421
rect 4995 6039 5029 7355
rect 5333 7208 5438 12343
rect 8633 12309 8744 12312
rect 10363 12309 10470 12924
rect 6397 12295 10470 12309
rect 6397 12275 8640 12295
rect 8659 12275 8717 12295
rect 8736 12291 10470 12295
rect 8736 12275 9688 12291
rect 6397 12271 9688 12275
rect 9707 12271 9765 12291
rect 9784 12271 10470 12291
rect 6397 12253 10470 12271
rect 6397 12252 7917 12253
rect 9681 12249 9792 12253
rect 8000 12201 8035 12202
rect 7979 12194 8035 12201
rect 7979 12174 8008 12194
rect 8028 12174 8035 12194
rect 7979 12169 8035 12174
rect 8426 12197 8458 12204
rect 9048 12197 9083 12198
rect 8426 12177 8432 12197
rect 8453 12177 8458 12197
rect 9027 12190 9083 12197
rect 8892 12180 8950 12185
rect 7979 11891 8013 12169
rect 8426 12149 8458 12177
rect 8046 12141 8458 12149
rect 8046 12115 8052 12141
rect 8078 12115 8458 12141
rect 8046 12113 8458 12115
rect 8048 12112 8088 12113
rect 8215 12087 8246 12095
rect 8215 12057 8219 12087
rect 8240 12057 8246 12087
rect 7979 11883 8014 11891
rect 7979 11863 7987 11883
rect 8007 11863 8014 11883
rect 7979 11858 8014 11863
rect 7979 11857 8011 11858
rect 8215 11857 8246 12057
rect 8426 12048 8458 12113
rect 8426 12028 8430 12048
rect 8451 12028 8458 12048
rect 8426 12021 8458 12028
rect 8875 12171 8950 12180
rect 8875 12138 8884 12171
rect 8937 12138 8950 12171
rect 8875 12113 8950 12138
rect 8875 12080 8889 12113
rect 8942 12080 8950 12113
rect 8875 12074 8950 12080
rect 9027 12170 9056 12190
rect 9076 12170 9083 12190
rect 9027 12165 9083 12170
rect 9474 12193 9506 12200
rect 9474 12173 9480 12193
rect 9501 12173 9506 12193
rect 8735 11965 8836 11966
rect 8633 11952 8836 11965
rect 8633 11950 8776 11952
rect 8633 11947 8710 11950
rect 8633 11920 8636 11947
rect 8665 11923 8710 11947
rect 8739 11923 8776 11950
rect 8665 11920 8776 11923
rect 8633 11919 8776 11920
rect 8812 11919 8836 11952
rect 8633 11906 8836 11919
rect 8212 11850 8251 11857
rect 8210 11833 8251 11850
rect 8212 11808 8251 11833
rect 6906 11800 8251 11808
rect 6906 11772 6921 11800
rect 6949 11774 8251 11800
rect 6949 11772 8248 11774
rect 6906 11767 8248 11772
rect 8875 11763 8945 12074
rect 9027 11887 9061 12165
rect 9474 12145 9506 12173
rect 9094 12137 9506 12145
rect 9094 12111 9100 12137
rect 9126 12111 9506 12137
rect 9094 12109 9506 12111
rect 9096 12108 9136 12109
rect 9263 12083 9294 12091
rect 9263 12053 9267 12083
rect 9288 12053 9294 12083
rect 9027 11879 9062 11887
rect 9027 11859 9035 11879
rect 9055 11859 9062 11879
rect 9027 11854 9062 11859
rect 9263 11854 9294 12053
rect 9474 12044 9506 12109
rect 9474 12024 9478 12044
rect 9499 12024 9506 12044
rect 9474 12017 9506 12024
rect 9919 12170 9991 12188
rect 9919 12128 9932 12170
rect 9981 12128 9991 12170
rect 9919 12107 9991 12128
rect 9919 12065 9933 12107
rect 9982 12065 9991 12107
rect 9783 11961 9884 11962
rect 9681 11948 9884 11961
rect 9681 11946 9824 11948
rect 9681 11943 9758 11946
rect 9681 11916 9684 11943
rect 9713 11919 9758 11943
rect 9787 11919 9824 11946
rect 9713 11916 9824 11919
rect 9681 11915 9824 11916
rect 9860 11915 9884 11948
rect 9681 11902 9884 11915
rect 9027 11853 9059 11854
rect 9261 11851 9294 11854
rect 9227 11832 9295 11851
rect 9197 11820 9296 11832
rect 9919 11824 9991 12065
rect 10363 11824 10470 12253
rect 10925 12665 11032 12924
rect 11404 12853 11476 13154
rect 12100 13144 12172 13145
rect 12099 13136 12198 13144
rect 12099 13133 12151 13136
rect 12099 13098 12107 13133
rect 12132 13098 12151 13133
rect 12176 13098 12198 13136
rect 12099 13086 12198 13098
rect 12100 13067 12168 13086
rect 12101 13064 12134 13067
rect 12336 13064 12368 13065
rect 11511 13003 11714 13016
rect 11511 12970 11535 13003
rect 11571 13002 11714 13003
rect 11571 12999 11682 13002
rect 11571 12972 11608 12999
rect 11637 12975 11682 12999
rect 11711 12975 11714 13002
rect 11637 12972 11714 12975
rect 11571 12970 11714 12972
rect 11511 12957 11714 12970
rect 11511 12956 11612 12957
rect 11404 12811 11413 12853
rect 11462 12811 11476 12853
rect 11404 12790 11476 12811
rect 11404 12748 11414 12790
rect 11463 12748 11476 12790
rect 11404 12730 11476 12748
rect 11889 12894 11921 12901
rect 11889 12874 11896 12894
rect 11917 12874 11921 12894
rect 11889 12809 11921 12874
rect 12101 12865 12132 13064
rect 12333 13059 12368 13064
rect 12333 13039 12340 13059
rect 12360 13039 12368 13059
rect 12333 13031 12368 13039
rect 12101 12835 12107 12865
rect 12128 12835 12132 12865
rect 12101 12827 12132 12835
rect 12259 12809 12299 12810
rect 11889 12807 12301 12809
rect 11889 12781 12269 12807
rect 12295 12781 12301 12807
rect 11889 12773 12301 12781
rect 11889 12745 11921 12773
rect 12334 12753 12368 13031
rect 12450 12844 12520 13144
rect 13149 13137 13238 13144
rect 13149 13134 13201 13137
rect 13149 13099 13157 13134
rect 13182 13099 13201 13134
rect 13226 13099 13238 13137
rect 13149 13087 13238 13099
rect 13149 13086 13218 13087
rect 13149 13068 13185 13086
rect 12559 12999 12762 13012
rect 12559 12966 12583 12999
rect 12619 12998 12762 12999
rect 12619 12995 12730 12998
rect 12619 12968 12656 12995
rect 12685 12971 12730 12995
rect 12759 12971 12762 12998
rect 12685 12968 12762 12971
rect 12619 12966 12762 12968
rect 12559 12953 12762 12966
rect 12559 12952 12660 12953
rect 11889 12725 11894 12745
rect 11915 12725 11921 12745
rect 11889 12718 11921 12725
rect 12312 12748 12368 12753
rect 12312 12728 12319 12748
rect 12339 12728 12368 12748
rect 12445 12838 12520 12844
rect 12445 12805 12453 12838
rect 12506 12805 12520 12838
rect 12445 12780 12520 12805
rect 12445 12747 12458 12780
rect 12511 12747 12520 12780
rect 12445 12738 12520 12747
rect 12937 12890 12969 12897
rect 12937 12870 12944 12890
rect 12965 12870 12969 12890
rect 12937 12805 12969 12870
rect 13149 12861 13180 13068
rect 13384 13060 13416 13061
rect 13381 13055 13416 13060
rect 13381 13035 13388 13055
rect 13408 13035 13416 13055
rect 13381 13027 13416 13035
rect 13149 12831 13155 12861
rect 13176 12831 13180 12861
rect 13149 12823 13180 12831
rect 13307 12805 13347 12806
rect 12937 12803 13349 12805
rect 12937 12777 13317 12803
rect 13343 12777 13349 12803
rect 12937 12769 13349 12777
rect 12937 12741 12969 12769
rect 13382 12749 13416 13027
rect 13565 12842 13627 13144
rect 13734 12845 13816 13201
rect 15001 13041 15050 13328
rect 15001 13009 15170 13041
rect 15001 13003 15116 13009
rect 15001 12994 15056 13003
rect 14991 12906 15056 12994
rect 15094 12912 15116 13003
rect 15154 12912 15170 13009
rect 15094 12906 15170 12912
rect 14991 12895 15170 12906
rect 13565 12823 13629 12842
rect 13565 12784 13578 12823
rect 13612 12784 13629 12823
rect 13565 12765 13629 12784
rect 13734 12804 13755 12845
rect 13791 12804 13816 12845
rect 13734 12775 13816 12804
rect 15001 12890 15170 12895
rect 12445 12733 12503 12738
rect 12312 12721 12368 12728
rect 12937 12721 12942 12741
rect 12963 12721 12969 12741
rect 12312 12720 12347 12721
rect 12937 12714 12969 12721
rect 13360 12744 13416 12749
rect 13360 12724 13367 12744
rect 13387 12724 13416 12744
rect 13360 12717 13416 12724
rect 13360 12716 13395 12717
rect 11603 12665 11714 12669
rect 13386 12665 14499 12666
rect 10925 12647 14499 12665
rect 10925 12627 11611 12647
rect 11630 12627 11688 12647
rect 11707 12643 14499 12647
rect 11707 12627 12659 12643
rect 10925 12623 12659 12627
rect 12678 12623 12736 12643
rect 12755 12623 14499 12643
rect 10925 12609 14499 12623
rect 10925 11986 11032 12609
rect 12651 12606 12762 12609
rect 11411 12560 11475 12564
rect 11407 12554 11475 12560
rect 11407 12521 11424 12554
rect 11464 12521 11475 12554
rect 11407 12509 11475 12521
rect 12458 12523 12523 12545
rect 11407 12507 11464 12509
rect 11411 12146 11462 12507
rect 12458 12484 12475 12523
rect 12520 12484 12523 12523
rect 12099 12439 12134 12441
rect 12099 12430 12203 12439
rect 12099 12429 12150 12430
rect 12099 12409 12102 12429
rect 12127 12410 12150 12429
rect 12182 12410 12203 12430
rect 12127 12409 12203 12410
rect 12099 12402 12203 12409
rect 12099 12390 12134 12402
rect 11511 12324 11714 12337
rect 11511 12291 11535 12324
rect 11571 12323 11714 12324
rect 11571 12320 11682 12323
rect 11571 12293 11608 12320
rect 11637 12296 11682 12320
rect 11711 12296 11714 12323
rect 11637 12293 11714 12296
rect 11571 12291 11714 12293
rect 11511 12278 11714 12291
rect 11511 12277 11612 12278
rect 11889 12215 11921 12222
rect 11889 12195 11896 12215
rect 11917 12195 11921 12215
rect 11400 12137 11465 12146
rect 11400 12100 11410 12137
rect 11450 12103 11465 12137
rect 11889 12130 11921 12195
rect 12101 12186 12132 12390
rect 12336 12385 12368 12386
rect 12333 12380 12368 12385
rect 12333 12360 12340 12380
rect 12360 12360 12368 12380
rect 12333 12352 12368 12360
rect 12101 12156 12107 12186
rect 12128 12156 12132 12186
rect 12101 12148 12132 12156
rect 12259 12130 12299 12131
rect 11889 12128 12301 12130
rect 11450 12100 11467 12103
rect 11400 12081 11467 12100
rect 11400 12060 11414 12081
rect 11450 12060 11467 12081
rect 11400 12053 11467 12060
rect 11889 12102 12269 12128
rect 12295 12102 12301 12128
rect 11889 12094 12301 12102
rect 11889 12066 11921 12094
rect 12334 12074 12368 12352
rect 12458 12184 12523 12484
rect 13729 12508 13822 12523
rect 13729 12464 13744 12508
rect 13804 12464 13822 12508
rect 11889 12046 11894 12066
rect 11915 12046 11921 12066
rect 11889 12039 11921 12046
rect 12312 12069 12368 12074
rect 12312 12049 12319 12069
rect 12339 12049 12368 12069
rect 12312 12042 12368 12049
rect 12448 12173 12528 12184
rect 12448 12147 12465 12173
rect 12505 12147 12528 12173
rect 12448 12120 12528 12147
rect 12448 12094 12469 12120
rect 12509 12094 12528 12120
rect 12448 12075 12528 12094
rect 12448 12049 12472 12075
rect 12512 12049 12528 12075
rect 12312 12041 12347 12042
rect 12448 12037 12528 12049
rect 13729 12091 13822 12464
rect 14006 12319 14209 12332
rect 14006 12286 14030 12319
rect 14066 12318 14209 12319
rect 14066 12315 14177 12318
rect 14066 12288 14103 12315
rect 14132 12291 14177 12315
rect 14206 12291 14209 12318
rect 14132 12288 14209 12291
rect 14066 12286 14209 12288
rect 14006 12273 14209 12286
rect 14006 12272 14107 12273
rect 13729 12050 13744 12091
rect 13798 12050 13822 12091
rect 13729 12043 13822 12050
rect 14384 12210 14416 12217
rect 14384 12190 14391 12210
rect 14412 12190 14416 12210
rect 14384 12125 14416 12190
rect 14596 12181 14627 12382
rect 14831 12380 14863 12381
rect 14828 12375 14863 12380
rect 14828 12355 14835 12375
rect 14855 12355 14863 12375
rect 14828 12347 14863 12355
rect 14596 12151 14602 12181
rect 14623 12151 14627 12181
rect 14596 12143 14627 12151
rect 14754 12125 14794 12126
rect 14384 12123 14796 12125
rect 14384 12097 14764 12123
rect 14790 12097 14796 12123
rect 14384 12089 14796 12097
rect 14384 12061 14416 12089
rect 14829 12069 14863 12347
rect 14384 12041 14389 12061
rect 14410 12041 14416 12061
rect 14384 12034 14416 12041
rect 14807 12064 14863 12069
rect 14807 12044 14814 12064
rect 14834 12044 14863 12064
rect 14807 12037 14863 12044
rect 14807 12036 14842 12037
rect 11603 11986 11714 11990
rect 13345 11986 14894 11989
rect 10923 11968 14894 11986
rect 10923 11948 11611 11968
rect 11630 11948 11688 11968
rect 11707 11963 14894 11968
rect 11707 11948 14106 11963
rect 10923 11943 14106 11948
rect 14125 11943 14183 11963
rect 14202 11943 14894 11963
rect 10923 11933 14894 11943
rect 10923 11930 11548 11933
rect 11735 11930 14894 11933
rect 9197 11782 9219 11820
rect 9244 11785 9263 11820
rect 9288 11785 9296 11820
rect 9244 11782 9296 11785
rect 9197 11774 9296 11782
rect 9223 11773 9295 11774
rect 8874 11747 8945 11763
rect 8874 11731 8894 11747
rect 8875 11701 8894 11731
rect 8877 11681 8894 11701
rect 8924 11701 8945 11747
rect 9917 11743 9995 11824
rect 10362 11769 10470 11824
rect 8924 11681 8944 11701
rect 8877 11662 8944 11681
rect 9917 11641 9996 11743
rect 9881 11623 10002 11641
rect 9881 11621 9952 11623
rect 9881 11580 9896 11621
rect 9933 11582 9952 11621
rect 9989 11582 10002 11623
rect 9933 11580 10002 11582
rect 9881 11570 10002 11580
rect 7186 11542 7297 11545
rect 6397 11541 8050 11542
rect 10363 11541 10470 11769
rect 10925 11702 11032 11930
rect 13345 11929 14894 11930
rect 14098 11926 14209 11929
rect 11393 11891 11514 11901
rect 11393 11889 11462 11891
rect 11393 11848 11406 11889
rect 11443 11850 11462 11889
rect 11499 11850 11514 11891
rect 11443 11848 11514 11850
rect 11393 11830 11514 11848
rect 14598 11871 14684 11875
rect 14598 11853 14613 11871
rect 14665 11853 14684 11871
rect 14598 11844 14684 11853
rect 11399 11728 11478 11830
rect 12451 11790 12518 11809
rect 12451 11770 12471 11790
rect 10925 11647 11033 11702
rect 11400 11647 11478 11728
rect 12450 11724 12471 11770
rect 12501 11770 12518 11790
rect 12501 11740 12520 11770
rect 12501 11724 12521 11740
rect 12450 11708 12521 11724
rect 12100 11697 12172 11698
rect 12099 11689 12198 11697
rect 12099 11686 12151 11689
rect 12099 11651 12107 11686
rect 12132 11651 12151 11686
rect 12176 11651 12198 11689
rect 6397 11538 9660 11541
rect 9847 11538 10472 11541
rect 6397 11528 10472 11538
rect 6397 11508 7193 11528
rect 7212 11508 7270 11528
rect 7289 11523 10472 11528
rect 7289 11508 9688 11523
rect 6397 11503 9688 11508
rect 9707 11503 9765 11523
rect 9784 11503 10472 11523
rect 6397 11485 10472 11503
rect 6397 11482 8050 11485
rect 9681 11481 9792 11485
rect 6553 11434 6588 11435
rect 6532 11427 6588 11434
rect 6532 11407 6561 11427
rect 6581 11407 6588 11427
rect 6532 11402 6588 11407
rect 6979 11430 7011 11437
rect 6979 11410 6985 11430
rect 7006 11410 7011 11430
rect 6532 11124 6566 11402
rect 6979 11382 7011 11410
rect 8867 11422 8947 11434
rect 9048 11429 9083 11430
rect 6599 11374 7011 11382
rect 6599 11348 6605 11374
rect 6631 11348 7011 11374
rect 7397 11388 7834 11401
rect 7397 11365 7410 11388
rect 7436 11381 7834 11388
rect 7436 11365 7790 11381
rect 7397 11358 7790 11365
rect 7816 11358 7834 11381
rect 7397 11352 7834 11358
rect 8867 11396 8883 11422
rect 8923 11396 8947 11422
rect 8867 11377 8947 11396
rect 6599 11346 7011 11348
rect 6601 11345 6641 11346
rect 6768 11320 6799 11328
rect 6768 11290 6772 11320
rect 6793 11290 6799 11320
rect 6532 11116 6567 11124
rect 6532 11096 6540 11116
rect 6560 11096 6567 11116
rect 6532 11091 6567 11096
rect 6532 11090 6564 11091
rect 6768 11083 6799 11290
rect 6979 11281 7011 11346
rect 8867 11351 8886 11377
rect 8926 11351 8947 11377
rect 8867 11324 8947 11351
rect 8867 11298 8890 11324
rect 8930 11298 8947 11324
rect 8867 11287 8947 11298
rect 9027 11422 9083 11429
rect 9027 11402 9056 11422
rect 9076 11402 9083 11422
rect 9027 11397 9083 11402
rect 9474 11425 9506 11432
rect 9474 11405 9480 11425
rect 9501 11405 9506 11425
rect 6979 11261 6983 11281
rect 7004 11261 7011 11281
rect 6979 11254 7011 11261
rect 7288 11198 7389 11199
rect 7186 11185 7389 11198
rect 7186 11183 7329 11185
rect 7186 11180 7263 11183
rect 7186 11153 7189 11180
rect 7218 11156 7263 11180
rect 7292 11156 7329 11183
rect 7218 11153 7329 11156
rect 7186 11152 7329 11153
rect 7365 11152 7389 11185
rect 7186 11139 7389 11152
rect 6766 11077 6799 11083
rect 6762 11073 6799 11077
rect 6762 11063 6800 11073
rect 6762 11050 6772 11063
rect 6763 11026 6772 11050
rect 6789 11026 6800 11063
rect 6763 11005 6800 11026
rect 8872 10987 8937 11287
rect 9027 11119 9061 11397
rect 9474 11377 9506 11405
rect 9094 11369 9506 11377
rect 9094 11343 9100 11369
rect 9126 11343 9506 11369
rect 9928 11411 9995 11418
rect 9928 11390 9945 11411
rect 9981 11390 9995 11411
rect 9928 11371 9995 11390
rect 9928 11368 9945 11371
rect 9094 11341 9506 11343
rect 9096 11340 9136 11341
rect 9263 11315 9294 11323
rect 9263 11285 9267 11315
rect 9288 11285 9294 11315
rect 9027 11111 9062 11119
rect 9027 11091 9035 11111
rect 9055 11091 9062 11111
rect 9027 11086 9062 11091
rect 9027 11085 9059 11086
rect 9263 11081 9294 11285
rect 9474 11276 9506 11341
rect 9930 11334 9945 11368
rect 9985 11334 9995 11371
rect 9930 11325 9995 11334
rect 9474 11256 9478 11276
rect 9499 11256 9506 11276
rect 9474 11249 9506 11256
rect 9783 11193 9884 11194
rect 9681 11180 9884 11193
rect 9681 11178 9824 11180
rect 9681 11175 9758 11178
rect 9681 11148 9684 11175
rect 9713 11151 9758 11175
rect 9787 11151 9824 11178
rect 9713 11148 9824 11151
rect 9681 11147 9824 11148
rect 9860 11147 9884 11180
rect 9681 11134 9884 11147
rect 9261 11069 9296 11081
rect 9192 11062 9296 11069
rect 9192 11061 9268 11062
rect 9192 11041 9213 11061
rect 9245 11042 9268 11061
rect 9293 11042 9296 11062
rect 9245 11041 9296 11042
rect 9192 11032 9296 11041
rect 9261 11030 9296 11032
rect 8872 10948 8875 10987
rect 8920 10948 8937 10987
rect 9933 10964 9984 11325
rect 9931 10962 9988 10964
rect 8872 10926 8937 10948
rect 9920 10950 9988 10962
rect 9920 10917 9931 10950
rect 9971 10917 9988 10950
rect 9920 10911 9988 10917
rect 9920 10907 9984 10911
rect 8633 10862 8744 10865
rect 10363 10862 10470 11485
rect 6020 10848 10470 10862
rect 6020 10828 8640 10848
rect 8659 10828 8717 10848
rect 8736 10844 10470 10848
rect 8736 10828 9688 10844
rect 6020 10824 9688 10828
rect 9707 10824 9765 10844
rect 9784 10824 10470 10844
rect 6020 10810 10470 10824
rect 6439 10806 10470 10810
rect 6439 10805 8009 10806
rect 9681 10802 9792 10806
rect 8000 10754 8035 10755
rect 7979 10747 8035 10754
rect 7979 10727 8008 10747
rect 8028 10727 8035 10747
rect 7979 10722 8035 10727
rect 8426 10750 8458 10757
rect 9048 10750 9083 10751
rect 8426 10730 8432 10750
rect 8453 10730 8458 10750
rect 9027 10743 9083 10750
rect 8892 10733 8950 10738
rect 7979 10444 8013 10722
rect 8426 10702 8458 10730
rect 8046 10694 8458 10702
rect 8046 10668 8052 10694
rect 8078 10668 8458 10694
rect 8046 10666 8458 10668
rect 8048 10665 8088 10666
rect 8215 10640 8246 10648
rect 8215 10610 8219 10640
rect 8240 10610 8246 10640
rect 7979 10436 8014 10444
rect 7979 10416 7987 10436
rect 8007 10416 8014 10436
rect 7979 10411 8014 10416
rect 7979 10410 8011 10411
rect 8215 10403 8246 10610
rect 8426 10601 8458 10666
rect 8426 10581 8430 10601
rect 8451 10581 8458 10601
rect 8426 10574 8458 10581
rect 8875 10724 8950 10733
rect 8875 10691 8884 10724
rect 8937 10691 8950 10724
rect 8875 10666 8950 10691
rect 8875 10633 8889 10666
rect 8942 10633 8950 10666
rect 8875 10627 8950 10633
rect 9027 10723 9056 10743
rect 9076 10723 9083 10743
rect 9027 10718 9083 10723
rect 9474 10746 9506 10753
rect 9474 10726 9480 10746
rect 9501 10726 9506 10746
rect 8735 10518 8836 10519
rect 8633 10505 8836 10518
rect 8633 10503 8776 10505
rect 8633 10500 8710 10503
rect 8633 10473 8636 10500
rect 8665 10476 8710 10500
rect 8739 10476 8776 10503
rect 8665 10473 8776 10476
rect 8633 10472 8776 10473
rect 8812 10472 8836 10505
rect 8633 10459 8836 10472
rect 7713 10390 7877 10393
rect 8210 10390 8246 10403
rect 6912 10372 8251 10390
rect 6912 10334 6922 10372
rect 6947 10357 8251 10372
rect 6947 10334 6957 10357
rect 7713 10350 7877 10357
rect 6912 10326 6957 10334
rect 6926 10325 6957 10326
rect 8875 10311 8945 10627
rect 9027 10440 9061 10718
rect 9474 10698 9506 10726
rect 9094 10690 9506 10698
rect 9094 10664 9100 10690
rect 9126 10664 9506 10690
rect 9094 10662 9506 10664
rect 9096 10661 9136 10662
rect 9263 10636 9294 10644
rect 9263 10606 9267 10636
rect 9288 10606 9294 10636
rect 9027 10432 9062 10440
rect 9027 10412 9035 10432
rect 9055 10412 9062 10432
rect 9027 10407 9062 10412
rect 9263 10407 9294 10606
rect 9474 10597 9506 10662
rect 9474 10577 9478 10597
rect 9499 10577 9506 10597
rect 9474 10570 9506 10577
rect 9919 10723 9991 10741
rect 9919 10681 9932 10723
rect 9981 10681 9991 10723
rect 9919 10660 9991 10681
rect 9919 10618 9933 10660
rect 9982 10618 9991 10660
rect 9783 10514 9884 10515
rect 9681 10501 9884 10514
rect 9681 10499 9824 10501
rect 9681 10496 9758 10499
rect 9681 10469 9684 10496
rect 9713 10472 9758 10496
rect 9787 10472 9824 10499
rect 9713 10469 9824 10472
rect 9681 10468 9824 10469
rect 9860 10468 9884 10501
rect 9681 10455 9884 10468
rect 9027 10406 9059 10407
rect 9261 10404 9294 10407
rect 9227 10385 9295 10404
rect 9197 10373 9296 10385
rect 9197 10335 9219 10373
rect 9244 10338 9263 10373
rect 9288 10338 9296 10373
rect 9244 10335 9296 10338
rect 9197 10327 9296 10335
rect 9223 10326 9295 10327
rect 8875 10292 8954 10311
rect 8878 10272 8954 10292
rect 8871 10248 8954 10272
rect 9919 10307 9991 10618
rect 9919 10264 9995 10307
rect 8871 10182 8883 10248
rect 8937 10182 8954 10248
rect 8871 10162 8954 10182
rect 8871 10125 8888 10162
rect 8932 10148 8954 10162
rect 9920 10213 9995 10264
rect 10363 10213 10470 10806
rect 10925 11218 11032 11647
rect 11404 11406 11476 11647
rect 12099 11639 12198 11651
rect 12100 11620 12168 11639
rect 12101 11617 12134 11620
rect 12336 11617 12368 11618
rect 11511 11556 11714 11569
rect 11511 11523 11535 11556
rect 11571 11555 11714 11556
rect 11571 11552 11682 11555
rect 11571 11525 11608 11552
rect 11637 11528 11682 11552
rect 11711 11528 11714 11555
rect 11637 11525 11714 11528
rect 11571 11523 11714 11525
rect 11511 11510 11714 11523
rect 11511 11509 11612 11510
rect 11404 11364 11413 11406
rect 11462 11364 11476 11406
rect 11404 11343 11476 11364
rect 11404 11301 11414 11343
rect 11463 11301 11476 11343
rect 11404 11283 11476 11301
rect 11889 11447 11921 11454
rect 11889 11427 11896 11447
rect 11917 11427 11921 11447
rect 11889 11362 11921 11427
rect 12101 11418 12132 11617
rect 12333 11612 12368 11617
rect 12333 11592 12340 11612
rect 12360 11592 12368 11612
rect 12333 11584 12368 11592
rect 12101 11388 12107 11418
rect 12128 11388 12132 11418
rect 12101 11380 12132 11388
rect 12259 11362 12299 11363
rect 11889 11360 12301 11362
rect 11889 11334 12269 11360
rect 12295 11334 12301 11360
rect 11889 11326 12301 11334
rect 11889 11298 11921 11326
rect 12334 11306 12368 11584
rect 12450 11397 12520 11708
rect 14375 11698 14447 11699
rect 14374 11695 14463 11698
rect 13146 11693 14463 11695
rect 13143 11690 14463 11693
rect 13143 11687 14426 11690
rect 13143 11652 14382 11687
rect 14407 11652 14426 11687
rect 14451 11652 14463 11690
rect 13143 11642 14463 11652
rect 14639 11691 14675 11844
rect 14639 11668 14645 11691
rect 14669 11668 14675 11691
rect 14639 11647 14675 11668
rect 13143 11640 14428 11642
rect 13143 11630 13240 11640
rect 13149 11621 13185 11630
rect 14639 11624 14645 11647
rect 14669 11624 14675 11647
rect 12559 11552 12762 11565
rect 12559 11519 12583 11552
rect 12619 11551 12762 11552
rect 12619 11548 12730 11551
rect 12619 11521 12656 11548
rect 12685 11524 12730 11548
rect 12759 11524 12762 11551
rect 12685 11521 12762 11524
rect 12619 11519 12762 11521
rect 12559 11506 12762 11519
rect 12559 11505 12660 11506
rect 11889 11278 11894 11298
rect 11915 11278 11921 11298
rect 11889 11271 11921 11278
rect 12312 11301 12368 11306
rect 12312 11281 12319 11301
rect 12339 11281 12368 11301
rect 12445 11391 12520 11397
rect 12445 11358 12453 11391
rect 12506 11358 12520 11391
rect 12445 11333 12520 11358
rect 12445 11300 12458 11333
rect 12511 11300 12520 11333
rect 12445 11291 12520 11300
rect 12937 11443 12969 11450
rect 12937 11423 12944 11443
rect 12965 11423 12969 11443
rect 12937 11358 12969 11423
rect 13149 11414 13180 11621
rect 13384 11613 13416 11614
rect 14639 11613 14675 11624
rect 13381 11608 13416 11613
rect 13381 11588 13388 11608
rect 13408 11588 13416 11608
rect 13381 11580 13416 11588
rect 13149 11384 13155 11414
rect 13176 11384 13180 11414
rect 13149 11376 13180 11384
rect 13307 11358 13347 11359
rect 12937 11356 13349 11358
rect 12937 11330 13317 11356
rect 13343 11330 13349 11356
rect 12937 11322 13349 11330
rect 12937 11294 12969 11322
rect 13382 11302 13416 11580
rect 12445 11286 12503 11291
rect 12312 11274 12368 11281
rect 12937 11274 12942 11294
rect 12963 11274 12969 11294
rect 12312 11273 12347 11274
rect 12937 11267 12969 11274
rect 13360 11297 13416 11302
rect 13360 11277 13367 11297
rect 13387 11277 13416 11297
rect 13360 11270 13416 11277
rect 13360 11269 13395 11270
rect 11603 11218 11714 11222
rect 13478 11218 14719 11219
rect 10925 11200 14719 11218
rect 10925 11180 11611 11200
rect 11630 11180 11688 11200
rect 11707 11196 14719 11200
rect 11707 11180 12659 11196
rect 10925 11176 12659 11180
rect 12678 11176 12736 11196
rect 12755 11176 14719 11196
rect 10925 11162 14719 11176
rect 10925 10539 11032 11162
rect 12651 11159 12762 11162
rect 11411 11113 11475 11117
rect 11407 11107 11475 11113
rect 11407 11074 11424 11107
rect 11464 11074 11475 11107
rect 11407 11062 11475 11074
rect 12458 11076 12523 11098
rect 11407 11060 11464 11062
rect 11411 10699 11462 11060
rect 12458 11037 12475 11076
rect 12520 11037 12523 11076
rect 12099 10992 12134 10994
rect 12099 10983 12203 10992
rect 12099 10982 12150 10983
rect 12099 10962 12102 10982
rect 12127 10963 12150 10982
rect 12182 10963 12203 10983
rect 12127 10962 12203 10963
rect 12099 10955 12203 10962
rect 12099 10943 12134 10955
rect 11511 10877 11714 10890
rect 11511 10844 11535 10877
rect 11571 10876 11714 10877
rect 11571 10873 11682 10876
rect 11571 10846 11608 10873
rect 11637 10849 11682 10873
rect 11711 10849 11714 10876
rect 11637 10846 11714 10849
rect 11571 10844 11714 10846
rect 11511 10831 11714 10844
rect 11511 10830 11612 10831
rect 11889 10768 11921 10775
rect 11889 10748 11896 10768
rect 11917 10748 11921 10768
rect 11400 10690 11465 10699
rect 11400 10653 11410 10690
rect 11450 10656 11465 10690
rect 11889 10683 11921 10748
rect 12101 10739 12132 10943
rect 12336 10938 12368 10939
rect 12333 10933 12368 10938
rect 12333 10913 12340 10933
rect 12360 10913 12368 10933
rect 12333 10905 12368 10913
rect 12101 10709 12107 10739
rect 12128 10709 12132 10739
rect 12101 10701 12132 10709
rect 12259 10683 12299 10684
rect 11889 10681 12301 10683
rect 11450 10653 11467 10656
rect 11400 10634 11467 10653
rect 11400 10613 11414 10634
rect 11450 10613 11467 10634
rect 11400 10606 11467 10613
rect 11889 10655 12269 10681
rect 12295 10655 12301 10681
rect 11889 10647 12301 10655
rect 11889 10619 11921 10647
rect 12334 10627 12368 10905
rect 12458 10737 12523 11037
rect 14637 11031 14742 11040
rect 14637 11026 14691 11031
rect 14637 11005 14650 11026
rect 14670 11010 14691 11026
rect 14711 11010 14742 11031
rect 14670 11005 14742 11010
rect 14637 10974 14742 11005
rect 14640 10957 14675 10974
rect 14639 10939 14675 10957
rect 14049 10874 14252 10887
rect 14049 10841 14073 10874
rect 14109 10873 14252 10874
rect 14109 10870 14220 10873
rect 14109 10843 14146 10870
rect 14175 10846 14220 10870
rect 14249 10846 14252 10873
rect 14175 10843 14252 10846
rect 14109 10841 14252 10843
rect 14049 10828 14252 10841
rect 14049 10827 14150 10828
rect 14427 10765 14459 10772
rect 14427 10745 14434 10765
rect 14455 10745 14459 10765
rect 11889 10599 11894 10619
rect 11915 10599 11921 10619
rect 11889 10592 11921 10599
rect 12312 10622 12368 10627
rect 12312 10602 12319 10622
rect 12339 10602 12368 10622
rect 12312 10595 12368 10602
rect 12448 10726 12528 10737
rect 12448 10700 12465 10726
rect 12505 10700 12528 10726
rect 12448 10673 12528 10700
rect 12448 10647 12469 10673
rect 12509 10647 12528 10673
rect 12448 10628 12528 10647
rect 12448 10602 12472 10628
rect 12512 10602 12528 10628
rect 12312 10594 12347 10595
rect 12448 10590 12528 10602
rect 14427 10680 14459 10745
rect 14639 10736 14670 10939
rect 14874 10935 14906 10936
rect 14871 10930 14906 10935
rect 14871 10910 14878 10930
rect 14898 10910 14906 10930
rect 14871 10902 14906 10910
rect 14639 10706 14645 10736
rect 14666 10706 14670 10736
rect 14639 10698 14670 10706
rect 14797 10680 14837 10681
rect 14427 10678 14839 10680
rect 14427 10652 14807 10678
rect 14833 10652 14839 10678
rect 14427 10644 14839 10652
rect 14427 10616 14459 10644
rect 14872 10624 14906 10902
rect 14427 10596 14432 10616
rect 14453 10596 14459 10616
rect 14427 10589 14459 10596
rect 14850 10619 14906 10624
rect 14850 10599 14857 10619
rect 14877 10599 14906 10619
rect 14850 10592 14906 10599
rect 14850 10591 14885 10592
rect 11603 10539 11714 10543
rect 13358 10539 13565 10540
rect 14141 10539 14252 10540
rect 10923 10521 14943 10539
rect 10923 10501 11611 10521
rect 11630 10501 11688 10521
rect 11707 10518 14943 10521
rect 11707 10501 14149 10518
rect 10923 10498 14149 10501
rect 14168 10498 14226 10518
rect 14245 10498 14943 10518
rect 10923 10483 14943 10498
rect 10925 10295 11032 10483
rect 13520 10481 14943 10483
rect 11393 10444 11514 10454
rect 11393 10442 11462 10444
rect 11393 10401 11406 10442
rect 11443 10403 11462 10442
rect 11499 10403 11514 10444
rect 11443 10401 11514 10403
rect 11393 10383 11514 10401
rect 10925 10291 11033 10295
rect 11399 10291 11476 10383
rect 12449 10379 12525 10395
rect 12449 10356 12464 10379
rect 8932 10125 8947 10148
rect 8871 10109 8947 10125
rect 9920 10121 9997 10213
rect 10363 10209 10471 10213
rect 9882 10103 10003 10121
rect 9882 10101 9953 10103
rect 9882 10060 9897 10101
rect 9934 10062 9953 10101
rect 9990 10062 10003 10103
rect 9934 10060 10003 10062
rect 9882 10050 10003 10060
rect 6407 10021 7876 10023
rect 10364 10021 10471 10209
rect 6407 10006 10473 10021
rect 6407 9986 7151 10006
rect 7170 9986 7228 10006
rect 7247 10003 10473 10006
rect 7247 9986 9689 10003
rect 6407 9983 9689 9986
rect 9708 9983 9766 10003
rect 9785 9983 10473 10003
rect 6407 9965 10473 9983
rect 7144 9964 7255 9965
rect 7831 9964 8038 9965
rect 9682 9961 9793 9965
rect 6511 9912 6546 9913
rect 6490 9905 6546 9912
rect 6490 9885 6519 9905
rect 6539 9885 6546 9905
rect 6490 9880 6546 9885
rect 6937 9908 6969 9915
rect 6937 9888 6943 9908
rect 6964 9888 6969 9908
rect 6490 9602 6524 9880
rect 6937 9860 6969 9888
rect 6557 9852 6969 9860
rect 6557 9826 6563 9852
rect 6589 9826 6969 9852
rect 6557 9824 6969 9826
rect 6559 9823 6599 9824
rect 6726 9798 6757 9806
rect 6726 9768 6730 9798
rect 6751 9768 6757 9798
rect 6490 9594 6525 9602
rect 6490 9574 6498 9594
rect 6518 9574 6525 9594
rect 6490 9569 6525 9574
rect 6726 9572 6757 9768
rect 6937 9759 6969 9824
rect 8868 9902 8948 9914
rect 9049 9909 9084 9910
rect 8868 9876 8884 9902
rect 8924 9876 8948 9902
rect 8868 9857 8948 9876
rect 8868 9831 8887 9857
rect 8927 9831 8948 9857
rect 8868 9804 8948 9831
rect 8868 9778 8891 9804
rect 8931 9778 8948 9804
rect 8868 9767 8948 9778
rect 9028 9902 9084 9909
rect 9028 9882 9057 9902
rect 9077 9882 9084 9902
rect 9028 9877 9084 9882
rect 9475 9905 9507 9912
rect 9475 9885 9481 9905
rect 9502 9885 9507 9905
rect 6937 9739 6941 9759
rect 6962 9739 6969 9759
rect 6937 9732 6969 9739
rect 7246 9676 7347 9677
rect 7144 9663 7347 9676
rect 7144 9661 7287 9663
rect 7144 9658 7221 9661
rect 7144 9631 7147 9658
rect 7176 9634 7221 9658
rect 7250 9634 7287 9661
rect 7176 9631 7287 9634
rect 7144 9630 7287 9631
rect 7323 9630 7347 9663
rect 7144 9617 7347 9630
rect 6490 9568 6522 9569
rect 6726 9483 6760 9572
rect 6347 9479 6760 9483
rect 5333 7154 5350 7208
rect 5413 7154 5438 7208
rect 5333 7133 5438 7154
rect 5800 9434 6760 9479
rect 8873 9467 8938 9767
rect 9028 9599 9062 9877
rect 9475 9857 9507 9885
rect 9095 9849 9507 9857
rect 9095 9823 9101 9849
rect 9127 9823 9507 9849
rect 9929 9891 9996 9898
rect 9929 9870 9946 9891
rect 9982 9870 9996 9891
rect 9929 9851 9996 9870
rect 9929 9848 9946 9851
rect 9095 9821 9507 9823
rect 9097 9820 9137 9821
rect 9264 9795 9295 9803
rect 9264 9765 9268 9795
rect 9289 9765 9295 9795
rect 9028 9591 9063 9599
rect 9028 9571 9036 9591
rect 9056 9571 9063 9591
rect 9028 9566 9063 9571
rect 9028 9565 9060 9566
rect 9264 9561 9295 9765
rect 9475 9756 9507 9821
rect 9931 9814 9946 9848
rect 9986 9814 9996 9851
rect 9931 9805 9996 9814
rect 9475 9736 9479 9756
rect 9500 9736 9507 9756
rect 9475 9729 9507 9736
rect 9784 9673 9885 9674
rect 9682 9660 9885 9673
rect 9682 9658 9825 9660
rect 9682 9655 9759 9658
rect 9682 9628 9685 9655
rect 9714 9631 9759 9655
rect 9788 9631 9825 9658
rect 9714 9628 9825 9631
rect 9682 9627 9825 9628
rect 9861 9627 9885 9660
rect 9682 9614 9885 9627
rect 9262 9549 9297 9561
rect 9193 9542 9297 9549
rect 9193 9541 9269 9542
rect 9193 9521 9214 9541
rect 9246 9522 9269 9541
rect 9294 9522 9297 9542
rect 9246 9521 9297 9522
rect 9193 9512 9297 9521
rect 9262 9510 9297 9512
rect 5800 9430 6397 9434
rect 5800 7124 5852 9430
rect 8873 9428 8876 9467
rect 8921 9428 8938 9467
rect 9934 9444 9985 9805
rect 9932 9442 9989 9444
rect 8873 9406 8938 9428
rect 9921 9430 9989 9442
rect 9921 9397 9932 9430
rect 9972 9397 9989 9430
rect 9921 9391 9989 9397
rect 9921 9387 9985 9391
rect 8634 9342 8745 9345
rect 10364 9342 10471 9965
rect 6759 9328 10471 9342
rect 6759 9308 8641 9328
rect 8660 9308 8718 9328
rect 8737 9324 10471 9328
rect 8737 9308 9689 9324
rect 6759 9304 9689 9308
rect 9708 9304 9766 9324
rect 9785 9304 10471 9324
rect 6759 9286 10471 9304
rect 6759 9285 7918 9286
rect 9682 9282 9793 9286
rect 8001 9234 8036 9235
rect 7980 9227 8036 9234
rect 7980 9207 8009 9227
rect 8029 9207 8036 9227
rect 7980 9202 8036 9207
rect 8427 9230 8459 9237
rect 9049 9230 9084 9231
rect 8427 9210 8433 9230
rect 8454 9210 8459 9230
rect 9028 9223 9084 9230
rect 8893 9213 8951 9218
rect 7980 8924 8014 9202
rect 8427 9182 8459 9210
rect 8047 9174 8459 9182
rect 8047 9148 8053 9174
rect 8079 9148 8459 9174
rect 8047 9146 8459 9148
rect 8049 9145 8089 9146
rect 8216 9120 8247 9128
rect 8216 9090 8220 9120
rect 8241 9090 8247 9120
rect 7980 8916 8015 8924
rect 7980 8896 7988 8916
rect 8008 8896 8015 8916
rect 7980 8891 8015 8896
rect 6721 8880 6757 8891
rect 7980 8890 8012 8891
rect 8216 8883 8247 9090
rect 8427 9081 8459 9146
rect 8427 9061 8431 9081
rect 8452 9061 8459 9081
rect 8427 9054 8459 9061
rect 8876 9204 8951 9213
rect 8876 9171 8885 9204
rect 8938 9171 8951 9204
rect 8876 9146 8951 9171
rect 8876 9113 8890 9146
rect 8943 9113 8951 9146
rect 8876 9107 8951 9113
rect 9028 9203 9057 9223
rect 9077 9203 9084 9223
rect 9028 9198 9084 9203
rect 9475 9226 9507 9233
rect 9475 9206 9481 9226
rect 9502 9206 9507 9226
rect 8736 8998 8837 8999
rect 8634 8985 8837 8998
rect 8634 8983 8777 8985
rect 8634 8980 8711 8983
rect 8634 8953 8637 8980
rect 8666 8956 8711 8980
rect 8740 8956 8777 8983
rect 8666 8953 8777 8956
rect 8634 8952 8777 8953
rect 8813 8952 8837 8985
rect 8634 8939 8837 8952
rect 6721 8857 6727 8880
rect 6751 8857 6757 8880
rect 8211 8874 8247 8883
rect 8156 8864 8253 8874
rect 6968 8862 8253 8864
rect 6721 8836 6757 8857
rect 6721 8813 6727 8836
rect 6751 8813 6757 8836
rect 6721 8660 6757 8813
rect 6933 8852 8253 8862
rect 6933 8814 6945 8852
rect 6970 8817 6989 8852
rect 7014 8817 8253 8852
rect 6970 8814 8253 8817
rect 6933 8811 8253 8814
rect 6933 8809 8250 8811
rect 6933 8806 7022 8809
rect 6949 8805 7021 8806
rect 8876 8796 8946 9107
rect 9028 8920 9062 9198
rect 9475 9178 9507 9206
rect 9095 9170 9507 9178
rect 9095 9144 9101 9170
rect 9127 9144 9507 9170
rect 9095 9142 9507 9144
rect 9097 9141 9137 9142
rect 9264 9116 9295 9124
rect 9264 9086 9268 9116
rect 9289 9086 9295 9116
rect 9028 8912 9063 8920
rect 9028 8892 9036 8912
rect 9056 8892 9063 8912
rect 9028 8887 9063 8892
rect 9264 8887 9295 9086
rect 9475 9077 9507 9142
rect 9475 9057 9479 9077
rect 9500 9057 9507 9077
rect 9475 9050 9507 9057
rect 9920 9203 9992 9221
rect 9920 9161 9933 9203
rect 9982 9161 9992 9203
rect 9920 9140 9992 9161
rect 9920 9098 9934 9140
rect 9983 9098 9992 9140
rect 9784 8994 9885 8995
rect 9682 8981 9885 8994
rect 9682 8979 9825 8981
rect 9682 8976 9759 8979
rect 9682 8949 9685 8976
rect 9714 8952 9759 8976
rect 9788 8952 9825 8979
rect 9714 8949 9825 8952
rect 9682 8948 9825 8949
rect 9861 8948 9885 8981
rect 9682 8935 9885 8948
rect 9028 8886 9060 8887
rect 9262 8884 9295 8887
rect 9228 8865 9296 8884
rect 9198 8853 9297 8865
rect 9920 8857 9992 9098
rect 10364 8857 10471 9286
rect 10926 9698 11033 10291
rect 11401 10240 11476 10291
rect 12442 10342 12464 10356
rect 12508 10342 12525 10379
rect 12442 10322 12525 10342
rect 12442 10256 12459 10322
rect 12513 10256 12525 10322
rect 11401 10197 11477 10240
rect 11405 9886 11477 10197
rect 12442 10232 12525 10256
rect 12442 10212 12518 10232
rect 12442 10193 12521 10212
rect 12101 10177 12173 10178
rect 12100 10169 12199 10177
rect 12100 10166 12152 10169
rect 12100 10131 12108 10166
rect 12133 10131 12152 10166
rect 12177 10131 12199 10169
rect 12100 10119 12199 10131
rect 12101 10100 12169 10119
rect 12102 10097 12135 10100
rect 12337 10097 12369 10098
rect 11512 10036 11715 10049
rect 11512 10003 11536 10036
rect 11572 10035 11715 10036
rect 11572 10032 11683 10035
rect 11572 10005 11609 10032
rect 11638 10008 11683 10032
rect 11712 10008 11715 10035
rect 11638 10005 11715 10008
rect 11572 10003 11715 10005
rect 11512 9990 11715 10003
rect 11512 9989 11613 9990
rect 11405 9844 11414 9886
rect 11463 9844 11477 9886
rect 11405 9823 11477 9844
rect 11405 9781 11415 9823
rect 11464 9781 11477 9823
rect 11405 9763 11477 9781
rect 11890 9927 11922 9934
rect 11890 9907 11897 9927
rect 11918 9907 11922 9927
rect 11890 9842 11922 9907
rect 12102 9898 12133 10097
rect 12334 10092 12369 10097
rect 12334 10072 12341 10092
rect 12361 10072 12369 10092
rect 12334 10064 12369 10072
rect 12102 9868 12108 9898
rect 12129 9868 12133 9898
rect 12102 9860 12133 9868
rect 12260 9842 12300 9843
rect 11890 9840 12302 9842
rect 11890 9814 12270 9840
rect 12296 9814 12302 9840
rect 11890 9806 12302 9814
rect 11890 9778 11922 9806
rect 12335 9786 12369 10064
rect 12451 9877 12521 10193
rect 14439 10178 14470 10179
rect 14439 10170 14484 10178
rect 13519 10147 13683 10154
rect 14439 10147 14449 10170
rect 13145 10132 14449 10147
rect 14474 10132 14484 10170
rect 13145 10114 14484 10132
rect 13150 10101 13186 10114
rect 13519 10111 13683 10114
rect 12560 10032 12763 10045
rect 12560 9999 12584 10032
rect 12620 10031 12763 10032
rect 12620 10028 12731 10031
rect 12620 10001 12657 10028
rect 12686 10004 12731 10028
rect 12760 10004 12763 10031
rect 12686 10001 12763 10004
rect 12620 9999 12763 10001
rect 12560 9986 12763 9999
rect 12560 9985 12661 9986
rect 11890 9758 11895 9778
rect 11916 9758 11922 9778
rect 11890 9751 11922 9758
rect 12313 9781 12369 9786
rect 12313 9761 12320 9781
rect 12340 9761 12369 9781
rect 12446 9871 12521 9877
rect 12446 9838 12454 9871
rect 12507 9838 12521 9871
rect 12446 9813 12521 9838
rect 12446 9780 12459 9813
rect 12512 9780 12521 9813
rect 12446 9771 12521 9780
rect 12938 9923 12970 9930
rect 12938 9903 12945 9923
rect 12966 9903 12970 9923
rect 12938 9838 12970 9903
rect 13150 9894 13181 10101
rect 13385 10093 13417 10094
rect 13382 10088 13417 10093
rect 13382 10068 13389 10088
rect 13409 10068 13417 10088
rect 13382 10060 13417 10068
rect 13150 9864 13156 9894
rect 13177 9864 13181 9894
rect 13150 9856 13181 9864
rect 13308 9838 13348 9839
rect 12938 9836 13350 9838
rect 12938 9810 13318 9836
rect 13344 9810 13350 9836
rect 12938 9802 13350 9810
rect 12938 9774 12970 9802
rect 13383 9782 13417 10060
rect 12446 9766 12504 9771
rect 12313 9754 12369 9761
rect 12938 9754 12943 9774
rect 12964 9754 12970 9774
rect 12313 9753 12348 9754
rect 12938 9747 12970 9754
rect 13361 9777 13417 9782
rect 13361 9757 13368 9777
rect 13388 9757 13417 9777
rect 13361 9750 13417 9757
rect 13361 9749 13396 9750
rect 11604 9698 11715 9702
rect 13387 9698 14687 9699
rect 10926 9680 14687 9698
rect 10926 9660 11612 9680
rect 11631 9660 11689 9680
rect 11708 9676 14687 9680
rect 11708 9660 12660 9676
rect 10926 9656 12660 9660
rect 12679 9656 12737 9676
rect 12756 9656 14687 9676
rect 10926 9642 14687 9656
rect 10926 9019 11033 9642
rect 12652 9639 12763 9642
rect 11412 9593 11476 9597
rect 11408 9587 11476 9593
rect 11408 9554 11425 9587
rect 11465 9554 11476 9587
rect 11408 9542 11476 9554
rect 12459 9556 12524 9578
rect 11408 9540 11465 9542
rect 11412 9179 11463 9540
rect 12459 9517 12476 9556
rect 12521 9517 12524 9556
rect 12100 9472 12135 9474
rect 12100 9463 12204 9472
rect 12100 9462 12151 9463
rect 12100 9442 12103 9462
rect 12128 9443 12151 9462
rect 12183 9443 12204 9463
rect 12128 9442 12204 9443
rect 12100 9435 12204 9442
rect 12100 9423 12135 9435
rect 11512 9357 11715 9370
rect 11512 9324 11536 9357
rect 11572 9356 11715 9357
rect 11572 9353 11683 9356
rect 11572 9326 11609 9353
rect 11638 9329 11683 9353
rect 11712 9329 11715 9356
rect 11638 9326 11715 9329
rect 11572 9324 11715 9326
rect 11512 9311 11715 9324
rect 11512 9310 11613 9311
rect 11890 9248 11922 9255
rect 11890 9228 11897 9248
rect 11918 9228 11922 9248
rect 11401 9170 11466 9179
rect 11401 9133 11411 9170
rect 11451 9136 11466 9170
rect 11890 9163 11922 9228
rect 12102 9219 12133 9423
rect 12337 9418 12369 9419
rect 12334 9413 12369 9418
rect 12334 9393 12341 9413
rect 12361 9393 12369 9413
rect 12334 9385 12369 9393
rect 12102 9189 12108 9219
rect 12129 9189 12133 9219
rect 12102 9181 12133 9189
rect 12260 9163 12300 9164
rect 11890 9161 12302 9163
rect 11451 9133 11468 9136
rect 11401 9114 11468 9133
rect 11401 9093 11415 9114
rect 11451 9093 11468 9114
rect 11401 9086 11468 9093
rect 11890 9135 12270 9161
rect 12296 9135 12302 9161
rect 11890 9127 12302 9135
rect 11890 9099 11922 9127
rect 12335 9107 12369 9385
rect 12459 9217 12524 9517
rect 14596 9478 14633 9499
rect 14596 9441 14607 9478
rect 14624 9454 14633 9478
rect 14624 9441 14634 9454
rect 14596 9431 14634 9441
rect 14597 9427 14634 9431
rect 14597 9421 14630 9427
rect 14007 9352 14210 9365
rect 14007 9319 14031 9352
rect 14067 9351 14210 9352
rect 14067 9348 14178 9351
rect 14067 9321 14104 9348
rect 14133 9324 14178 9348
rect 14207 9324 14210 9351
rect 14133 9321 14210 9324
rect 14067 9319 14210 9321
rect 14007 9306 14210 9319
rect 14007 9305 14108 9306
rect 14385 9243 14417 9250
rect 14385 9223 14392 9243
rect 14413 9223 14417 9243
rect 11890 9079 11895 9099
rect 11916 9079 11922 9099
rect 11890 9072 11922 9079
rect 12313 9102 12369 9107
rect 12313 9082 12320 9102
rect 12340 9082 12369 9102
rect 12313 9075 12369 9082
rect 12449 9206 12529 9217
rect 12449 9180 12466 9206
rect 12506 9180 12529 9206
rect 12449 9153 12529 9180
rect 12449 9127 12470 9153
rect 12510 9127 12529 9153
rect 14385 9158 14417 9223
rect 14597 9214 14628 9421
rect 14832 9413 14864 9414
rect 14829 9408 14864 9413
rect 14829 9388 14836 9408
rect 14856 9388 14864 9408
rect 14829 9380 14864 9388
rect 14597 9184 14603 9214
rect 14624 9184 14628 9214
rect 14597 9176 14628 9184
rect 14755 9158 14795 9159
rect 14385 9156 14797 9158
rect 12449 9108 12529 9127
rect 12449 9082 12473 9108
rect 12513 9082 12529 9108
rect 13562 9146 13999 9152
rect 13562 9123 13580 9146
rect 13606 9139 13999 9146
rect 13606 9123 13960 9139
rect 13562 9116 13960 9123
rect 13986 9116 13999 9139
rect 13562 9103 13999 9116
rect 14385 9130 14765 9156
rect 14791 9130 14797 9156
rect 14385 9122 14797 9130
rect 12313 9074 12348 9075
rect 12449 9070 12529 9082
rect 14385 9094 14417 9122
rect 14830 9102 14864 9380
rect 14385 9074 14390 9094
rect 14411 9074 14417 9094
rect 14385 9067 14417 9074
rect 14808 9097 14864 9102
rect 14808 9077 14815 9097
rect 14835 9077 14864 9097
rect 14808 9070 14864 9077
rect 14808 9069 14843 9070
rect 11604 9019 11715 9023
rect 13346 9019 14896 9022
rect 10924 9001 14896 9019
rect 10924 8981 11612 9001
rect 11631 8981 11689 9001
rect 11708 8996 14896 9001
rect 11708 8981 14107 8996
rect 10924 8976 14107 8981
rect 14126 8976 14184 8996
rect 14203 8976 14896 8996
rect 10924 8966 14896 8976
rect 10924 8963 11549 8966
rect 11736 8963 14896 8966
rect 9198 8815 9220 8853
rect 9245 8818 9264 8853
rect 9289 8818 9297 8853
rect 9245 8815 9297 8818
rect 9198 8807 9297 8815
rect 9224 8806 9296 8807
rect 8875 8780 8946 8796
rect 8875 8764 8895 8780
rect 8876 8734 8895 8764
rect 8878 8714 8895 8734
rect 8925 8734 8946 8780
rect 9918 8776 9996 8857
rect 10363 8802 10471 8857
rect 8925 8714 8945 8734
rect 8878 8695 8945 8714
rect 9918 8674 9997 8776
rect 6712 8651 6798 8660
rect 6712 8633 6731 8651
rect 6783 8633 6798 8651
rect 6712 8629 6798 8633
rect 9882 8656 10003 8674
rect 9882 8654 9953 8656
rect 9882 8613 9897 8654
rect 9934 8615 9953 8654
rect 9990 8615 10003 8656
rect 9934 8613 10003 8615
rect 9882 8603 10003 8613
rect 7187 8575 7298 8578
rect 6407 8574 8051 8575
rect 10364 8574 10471 8802
rect 10926 8735 11033 8963
rect 13346 8962 14896 8963
rect 14099 8959 14210 8962
rect 11394 8924 11515 8934
rect 11394 8922 11463 8924
rect 11394 8881 11407 8922
rect 11444 8883 11463 8922
rect 11500 8883 11515 8924
rect 11444 8881 11515 8883
rect 11394 8863 11515 8881
rect 11400 8761 11479 8863
rect 12452 8823 12519 8842
rect 12452 8803 12472 8823
rect 10926 8680 11034 8735
rect 11401 8680 11479 8761
rect 12451 8757 12472 8803
rect 12502 8803 12519 8823
rect 12502 8773 12521 8803
rect 12502 8757 12522 8773
rect 12451 8741 12522 8757
rect 12101 8730 12173 8731
rect 12100 8722 12199 8730
rect 12100 8719 12152 8722
rect 12100 8684 12108 8719
rect 12133 8684 12152 8719
rect 12177 8684 12199 8722
rect 6407 8571 9661 8574
rect 9848 8571 10473 8574
rect 6407 8561 10473 8571
rect 6407 8541 7194 8561
rect 7213 8541 7271 8561
rect 7290 8556 10473 8561
rect 7290 8541 9689 8556
rect 6407 8536 9689 8541
rect 9708 8536 9766 8556
rect 9785 8536 10473 8556
rect 6407 8518 10473 8536
rect 6407 8515 8051 8518
rect 9682 8514 9793 8518
rect 6554 8467 6589 8468
rect 6533 8460 6589 8467
rect 6533 8440 6562 8460
rect 6582 8440 6589 8460
rect 6533 8435 6589 8440
rect 6980 8463 7012 8470
rect 6980 8443 6986 8463
rect 7007 8443 7012 8463
rect 6533 8157 6567 8435
rect 6980 8415 7012 8443
rect 6600 8407 7012 8415
rect 6600 8381 6606 8407
rect 6632 8381 7012 8407
rect 6600 8379 7012 8381
rect 6602 8378 6642 8379
rect 6769 8353 6800 8361
rect 6769 8323 6773 8353
rect 6794 8323 6800 8353
rect 6533 8149 6568 8157
rect 6533 8129 6541 8149
rect 6561 8129 6568 8149
rect 6533 8124 6568 8129
rect 6533 8123 6565 8124
rect 6769 8122 6800 8323
rect 6980 8314 7012 8379
rect 6980 8294 6984 8314
rect 7005 8294 7012 8314
rect 6980 8287 7012 8294
rect 7574 8454 7667 8461
rect 7574 8413 7598 8454
rect 7652 8413 7667 8454
rect 7289 8231 7390 8232
rect 7187 8218 7390 8231
rect 7187 8216 7330 8218
rect 7187 8213 7264 8216
rect 7187 8186 7190 8213
rect 7219 8189 7264 8213
rect 7293 8189 7330 8216
rect 7219 8186 7330 8189
rect 7187 8185 7330 8186
rect 7366 8185 7390 8218
rect 7187 8172 7390 8185
rect 7574 8040 7667 8413
rect 8868 8455 8948 8467
rect 9049 8462 9084 8463
rect 8868 8429 8884 8455
rect 8924 8429 8948 8455
rect 8868 8410 8948 8429
rect 8868 8384 8887 8410
rect 8927 8384 8948 8410
rect 8868 8357 8948 8384
rect 8868 8331 8891 8357
rect 8931 8331 8948 8357
rect 8868 8320 8948 8331
rect 9028 8455 9084 8462
rect 9028 8435 9057 8455
rect 9077 8435 9084 8455
rect 9028 8430 9084 8435
rect 9475 8458 9507 8465
rect 9475 8438 9481 8458
rect 9502 8438 9507 8458
rect 7574 7996 7592 8040
rect 7652 7996 7667 8040
rect 7574 7981 7667 7996
rect 8873 8020 8938 8320
rect 9028 8152 9062 8430
rect 9475 8410 9507 8438
rect 9095 8402 9507 8410
rect 9095 8376 9101 8402
rect 9127 8376 9507 8402
rect 9929 8444 9996 8451
rect 9929 8423 9946 8444
rect 9982 8423 9996 8444
rect 9929 8404 9996 8423
rect 9929 8401 9946 8404
rect 9095 8374 9507 8376
rect 9097 8373 9137 8374
rect 9264 8348 9295 8356
rect 9264 8318 9268 8348
rect 9289 8318 9295 8348
rect 9028 8144 9063 8152
rect 9028 8124 9036 8144
rect 9056 8124 9063 8144
rect 9028 8119 9063 8124
rect 9028 8118 9060 8119
rect 9264 8114 9295 8318
rect 9475 8309 9507 8374
rect 9931 8367 9946 8401
rect 9986 8367 9996 8404
rect 9931 8358 9996 8367
rect 9475 8289 9479 8309
rect 9500 8289 9507 8309
rect 9475 8282 9507 8289
rect 9784 8226 9885 8227
rect 9682 8213 9885 8226
rect 9682 8211 9825 8213
rect 9682 8208 9759 8211
rect 9682 8181 9685 8208
rect 9714 8184 9759 8208
rect 9788 8184 9825 8211
rect 9714 8181 9825 8184
rect 9682 8180 9825 8181
rect 9861 8180 9885 8213
rect 9682 8167 9885 8180
rect 9262 8102 9297 8114
rect 9193 8095 9297 8102
rect 9193 8094 9269 8095
rect 9193 8074 9214 8094
rect 9246 8075 9269 8094
rect 9294 8075 9297 8095
rect 9246 8074 9297 8075
rect 9193 8065 9297 8074
rect 9262 8063 9297 8065
rect 8873 7981 8876 8020
rect 8921 7981 8938 8020
rect 9934 7997 9985 8358
rect 9932 7995 9989 7997
rect 8873 7959 8938 7981
rect 9921 7983 9989 7995
rect 9921 7950 9932 7983
rect 9972 7950 9989 7983
rect 9921 7944 9989 7950
rect 9921 7940 9985 7944
rect 8634 7895 8745 7898
rect 10364 7895 10471 8518
rect 6440 7881 10471 7895
rect 6440 7861 8641 7881
rect 8660 7861 8718 7881
rect 8737 7877 10471 7881
rect 8737 7861 9689 7877
rect 6440 7857 9689 7861
rect 9708 7857 9766 7877
rect 9785 7857 10471 7877
rect 6440 7839 10471 7857
rect 6440 7838 8010 7839
rect 9682 7835 9793 7839
rect 8001 7787 8036 7788
rect 7980 7780 8036 7787
rect 7980 7760 8009 7780
rect 8029 7760 8036 7780
rect 7980 7755 8036 7760
rect 8427 7783 8459 7790
rect 9049 7783 9084 7784
rect 8427 7763 8433 7783
rect 8454 7763 8459 7783
rect 9028 7776 9084 7783
rect 8893 7766 8951 7771
rect 7580 7700 7662 7729
rect 7580 7659 7605 7700
rect 7641 7659 7662 7700
rect 7767 7720 7831 7739
rect 7767 7681 7784 7720
rect 7818 7681 7831 7720
rect 7767 7662 7831 7681
rect 7580 7344 7662 7659
rect 7572 7299 7662 7344
rect 7769 7317 7831 7662
rect 7980 7477 8014 7755
rect 8427 7735 8459 7763
rect 8047 7727 8459 7735
rect 8047 7701 8053 7727
rect 8079 7701 8459 7727
rect 8047 7699 8459 7701
rect 8049 7698 8089 7699
rect 8216 7673 8247 7681
rect 8216 7643 8220 7673
rect 8241 7643 8247 7673
rect 7980 7469 8015 7477
rect 7980 7449 7988 7469
rect 8008 7449 8015 7469
rect 7980 7444 8015 7449
rect 7980 7443 8012 7444
rect 8216 7436 8247 7643
rect 8427 7634 8459 7699
rect 8427 7614 8431 7634
rect 8452 7614 8459 7634
rect 8427 7607 8459 7614
rect 8876 7757 8951 7766
rect 8876 7724 8885 7757
rect 8938 7724 8951 7757
rect 8876 7699 8951 7724
rect 8876 7666 8890 7699
rect 8943 7666 8951 7699
rect 8876 7660 8951 7666
rect 9028 7756 9057 7776
rect 9077 7756 9084 7776
rect 9028 7751 9084 7756
rect 9475 7779 9507 7786
rect 9475 7759 9481 7779
rect 9502 7759 9507 7779
rect 8736 7551 8837 7552
rect 8634 7538 8837 7551
rect 8634 7536 8777 7538
rect 8634 7533 8711 7536
rect 8634 7506 8637 7533
rect 8666 7509 8711 7533
rect 8740 7509 8777 7536
rect 8666 7506 8777 7509
rect 8634 7505 8777 7506
rect 8813 7505 8837 7538
rect 8634 7492 8837 7505
rect 8211 7418 8247 7436
rect 8178 7417 8247 7418
rect 8158 7405 8247 7417
rect 8158 7367 8170 7405
rect 8195 7370 8214 7405
rect 8239 7370 8247 7405
rect 8876 7394 8946 7660
rect 9028 7473 9062 7751
rect 9475 7731 9507 7759
rect 9095 7723 9507 7731
rect 9095 7697 9101 7723
rect 9127 7697 9507 7723
rect 9095 7695 9507 7697
rect 9097 7694 9137 7695
rect 9264 7669 9295 7677
rect 9264 7639 9268 7669
rect 9289 7639 9295 7669
rect 9028 7465 9063 7473
rect 9028 7445 9036 7465
rect 9056 7445 9063 7465
rect 9028 7440 9063 7445
rect 9264 7440 9295 7639
rect 9475 7630 9507 7695
rect 9475 7610 9479 7630
rect 9500 7610 9507 7630
rect 9475 7603 9507 7610
rect 9920 7756 9992 7774
rect 9920 7714 9933 7756
rect 9982 7714 9992 7756
rect 9920 7693 9992 7714
rect 9920 7651 9934 7693
rect 9983 7651 9992 7693
rect 9784 7547 9885 7548
rect 9682 7534 9885 7547
rect 9682 7532 9825 7534
rect 9682 7529 9759 7532
rect 9682 7502 9685 7529
rect 9714 7505 9759 7529
rect 9788 7505 9825 7532
rect 9714 7502 9825 7505
rect 9682 7501 9825 7502
rect 9861 7501 9885 7534
rect 9682 7488 9885 7501
rect 9028 7439 9060 7440
rect 9262 7437 9295 7440
rect 9228 7418 9296 7437
rect 8195 7367 8247 7370
rect 8158 7359 8247 7367
rect 8867 7365 8946 7394
rect 9198 7406 9297 7418
rect 9198 7368 9220 7406
rect 9245 7371 9264 7406
rect 9289 7371 9297 7406
rect 9245 7368 9297 7371
rect 8174 7358 8246 7359
rect 7768 7308 7842 7317
rect 7572 7266 7656 7299
rect 7572 7238 7587 7266
rect 7631 7238 7656 7266
rect 7572 7209 7656 7238
rect 7768 7260 7782 7308
rect 7819 7260 7842 7308
rect 7768 7232 7842 7260
rect 7572 7181 7584 7209
rect 7628 7181 7656 7209
rect 7572 7170 7656 7181
rect 8867 7182 8944 7365
rect 9198 7360 9297 7368
rect 9224 7359 9296 7360
rect 9920 7357 9992 7651
rect 10364 7379 10471 7839
rect 10926 8251 11033 8680
rect 11405 8439 11477 8680
rect 12100 8672 12199 8684
rect 12101 8653 12169 8672
rect 12102 8650 12135 8653
rect 12337 8650 12369 8651
rect 11512 8589 11715 8602
rect 11512 8556 11536 8589
rect 11572 8588 11715 8589
rect 11572 8585 11683 8588
rect 11572 8558 11609 8585
rect 11638 8561 11683 8585
rect 11712 8561 11715 8588
rect 11638 8558 11715 8561
rect 11572 8556 11715 8558
rect 11512 8543 11715 8556
rect 11512 8542 11613 8543
rect 11405 8397 11414 8439
rect 11463 8397 11477 8439
rect 11405 8376 11477 8397
rect 11405 8334 11415 8376
rect 11464 8334 11477 8376
rect 11405 8316 11477 8334
rect 11890 8480 11922 8487
rect 11890 8460 11897 8480
rect 11918 8460 11922 8480
rect 11890 8395 11922 8460
rect 12102 8451 12133 8650
rect 12334 8645 12369 8650
rect 12334 8625 12341 8645
rect 12361 8625 12369 8645
rect 12334 8617 12369 8625
rect 12102 8421 12108 8451
rect 12129 8421 12133 8451
rect 12102 8413 12133 8421
rect 12260 8395 12300 8396
rect 11890 8393 12302 8395
rect 11890 8367 12270 8393
rect 12296 8367 12302 8393
rect 11890 8359 12302 8367
rect 11890 8331 11922 8359
rect 12335 8339 12369 8617
rect 12451 8430 12521 8741
rect 13148 8732 14490 8737
rect 13148 8730 14447 8732
rect 13145 8704 14447 8730
rect 14475 8704 14490 8732
rect 13145 8696 14490 8704
rect 13145 8671 13184 8696
rect 13145 8654 13186 8671
rect 13145 8647 13184 8654
rect 12560 8585 12763 8598
rect 12560 8552 12584 8585
rect 12620 8584 12763 8585
rect 12620 8581 12731 8584
rect 12620 8554 12657 8581
rect 12686 8557 12731 8581
rect 12760 8557 12763 8584
rect 12686 8554 12763 8557
rect 12620 8552 12763 8554
rect 12560 8539 12763 8552
rect 12560 8538 12661 8539
rect 11890 8311 11895 8331
rect 11916 8311 11922 8331
rect 11890 8304 11922 8311
rect 12313 8334 12369 8339
rect 12313 8314 12320 8334
rect 12340 8314 12369 8334
rect 12446 8424 12521 8430
rect 12446 8391 12454 8424
rect 12507 8391 12521 8424
rect 12446 8366 12521 8391
rect 12446 8333 12459 8366
rect 12512 8333 12521 8366
rect 12446 8324 12521 8333
rect 12938 8476 12970 8483
rect 12938 8456 12945 8476
rect 12966 8456 12970 8476
rect 12938 8391 12970 8456
rect 13150 8447 13181 8647
rect 13385 8646 13417 8647
rect 13382 8641 13417 8646
rect 13382 8621 13389 8641
rect 13409 8621 13417 8641
rect 13382 8613 13417 8621
rect 13150 8417 13156 8447
rect 13177 8417 13181 8447
rect 13150 8409 13181 8417
rect 13308 8391 13348 8392
rect 12938 8389 13350 8391
rect 12938 8363 13318 8389
rect 13344 8363 13350 8389
rect 12938 8355 13350 8363
rect 12938 8327 12970 8355
rect 13383 8335 13417 8613
rect 12446 8319 12504 8324
rect 12313 8307 12369 8314
rect 12938 8307 12943 8327
rect 12964 8307 12970 8327
rect 12313 8306 12348 8307
rect 12938 8300 12970 8307
rect 13361 8330 13417 8335
rect 13361 8310 13368 8330
rect 13388 8310 13417 8330
rect 13361 8303 13417 8310
rect 13361 8302 13396 8303
rect 11604 8251 11715 8255
rect 13479 8251 14469 8252
rect 10926 8233 14469 8251
rect 10926 8213 11612 8233
rect 11631 8213 11689 8233
rect 11708 8229 14469 8233
rect 11708 8213 12660 8229
rect 10926 8209 12660 8213
rect 12679 8209 12737 8229
rect 12756 8209 14469 8229
rect 10926 8195 14469 8209
rect 10926 7572 11033 8195
rect 12652 8192 12763 8195
rect 11412 8146 11476 8150
rect 11408 8140 11476 8146
rect 11408 8107 11425 8140
rect 11465 8107 11476 8140
rect 11408 8095 11476 8107
rect 12459 8109 12524 8131
rect 11408 8093 11465 8095
rect 11412 7732 11463 8093
rect 12459 8070 12476 8109
rect 12521 8070 12524 8109
rect 12100 8025 12135 8027
rect 12100 8016 12204 8025
rect 12100 8015 12151 8016
rect 12100 7995 12103 8015
rect 12128 7996 12151 8015
rect 12183 7996 12204 8016
rect 12128 7995 12204 7996
rect 12100 7988 12204 7995
rect 12100 7976 12135 7988
rect 11512 7910 11715 7923
rect 11512 7877 11536 7910
rect 11572 7909 11715 7910
rect 11572 7906 11683 7909
rect 11572 7879 11609 7906
rect 11638 7882 11683 7906
rect 11712 7882 11715 7909
rect 11638 7879 11715 7882
rect 11572 7877 11715 7879
rect 11512 7864 11715 7877
rect 11512 7863 11613 7864
rect 11890 7801 11922 7808
rect 11890 7781 11897 7801
rect 11918 7781 11922 7801
rect 11401 7723 11466 7732
rect 11401 7686 11411 7723
rect 11451 7689 11466 7723
rect 11890 7716 11922 7781
rect 12102 7772 12133 7976
rect 12337 7971 12369 7972
rect 12334 7966 12369 7971
rect 12334 7946 12341 7966
rect 12361 7946 12369 7966
rect 12334 7938 12369 7946
rect 12102 7742 12108 7772
rect 12129 7742 12133 7772
rect 12102 7734 12133 7742
rect 12260 7716 12300 7717
rect 11890 7714 12302 7716
rect 11451 7686 11468 7689
rect 11401 7667 11468 7686
rect 11401 7646 11415 7667
rect 11451 7646 11468 7667
rect 11401 7639 11468 7646
rect 11890 7688 12270 7714
rect 12296 7688 12302 7714
rect 11890 7680 12302 7688
rect 11890 7652 11922 7680
rect 12335 7660 12369 7938
rect 12459 7770 12524 8070
rect 11890 7632 11895 7652
rect 11916 7632 11922 7652
rect 11890 7625 11922 7632
rect 12313 7655 12369 7660
rect 12313 7635 12320 7655
rect 12340 7635 12369 7655
rect 12313 7628 12369 7635
rect 12449 7759 12529 7770
rect 12449 7733 12466 7759
rect 12506 7733 12529 7759
rect 12449 7706 12529 7733
rect 15001 7709 15050 12890
rect 16049 12302 16136 13457
rect 20639 13082 20704 13220
rect 20589 13064 20710 13082
rect 20589 13062 20660 13064
rect 20589 13021 20604 13062
rect 20641 13023 20660 13062
rect 20697 13023 20710 13064
rect 20641 13021 20710 13023
rect 20589 13011 20710 13021
rect 17105 12982 18583 12984
rect 21071 12982 21178 13182
rect 17105 12964 21180 12982
rect 17105 12944 20396 12964
rect 20415 12944 20473 12964
rect 20492 12944 21180 12964
rect 17105 12926 21180 12944
rect 18538 12925 18745 12926
rect 20389 12922 20500 12926
rect 19575 12863 19655 12875
rect 19756 12870 19791 12871
rect 19575 12837 19591 12863
rect 19631 12837 19655 12863
rect 19575 12818 19655 12837
rect 19575 12792 19594 12818
rect 19634 12792 19655 12818
rect 19575 12765 19655 12792
rect 19575 12739 19598 12765
rect 19638 12739 19655 12765
rect 19575 12728 19655 12739
rect 19735 12863 19791 12870
rect 19735 12843 19764 12863
rect 19784 12843 19791 12863
rect 19735 12838 19791 12843
rect 20182 12866 20214 12873
rect 20182 12846 20188 12866
rect 20209 12846 20214 12866
rect 19580 12428 19645 12728
rect 19735 12560 19769 12838
rect 20182 12818 20214 12846
rect 19802 12810 20214 12818
rect 19802 12784 19808 12810
rect 19834 12784 20214 12810
rect 20636 12852 20703 12859
rect 20636 12831 20653 12852
rect 20689 12831 20703 12852
rect 20636 12812 20703 12831
rect 20636 12809 20653 12812
rect 19802 12782 20214 12784
rect 19804 12781 19844 12782
rect 19971 12756 20002 12764
rect 19971 12726 19975 12756
rect 19996 12726 20002 12756
rect 19735 12552 19770 12560
rect 19735 12532 19743 12552
rect 19763 12532 19770 12552
rect 19735 12527 19770 12532
rect 19735 12526 19767 12527
rect 19971 12522 20002 12726
rect 20182 12717 20214 12782
rect 20638 12775 20653 12809
rect 20693 12775 20703 12812
rect 20638 12766 20703 12775
rect 20182 12697 20186 12717
rect 20207 12697 20214 12717
rect 20182 12690 20214 12697
rect 20491 12634 20592 12635
rect 20389 12621 20592 12634
rect 20389 12619 20532 12621
rect 20389 12616 20466 12619
rect 20389 12589 20392 12616
rect 20421 12592 20466 12616
rect 20495 12592 20532 12619
rect 20421 12589 20532 12592
rect 20389 12588 20532 12589
rect 20568 12588 20592 12621
rect 20389 12575 20592 12588
rect 19969 12510 20004 12522
rect 19900 12503 20004 12510
rect 19900 12502 19976 12503
rect 19900 12482 19921 12502
rect 19953 12483 19976 12502
rect 20001 12483 20004 12503
rect 19953 12482 20004 12483
rect 19900 12473 20004 12482
rect 19969 12471 20004 12473
rect 19580 12389 19583 12428
rect 19628 12389 19645 12428
rect 20641 12405 20692 12766
rect 20639 12403 20696 12405
rect 19580 12367 19645 12389
rect 20628 12391 20696 12403
rect 20628 12358 20639 12391
rect 20679 12358 20696 12391
rect 20628 12352 20696 12358
rect 20628 12348 20692 12352
rect 19341 12303 19452 12306
rect 21071 12303 21178 12926
rect 15115 7901 15318 7914
rect 15115 7868 15139 7901
rect 15175 7900 15318 7901
rect 15175 7897 15286 7900
rect 15175 7870 15212 7897
rect 15241 7873 15286 7897
rect 15315 7873 15318 7900
rect 15241 7870 15318 7873
rect 15175 7868 15318 7870
rect 15115 7855 15318 7868
rect 15115 7854 15216 7855
rect 15493 7792 15525 7799
rect 15493 7772 15500 7792
rect 15521 7772 15525 7792
rect 12449 7680 12470 7706
rect 12510 7680 12529 7706
rect 12449 7661 12529 7680
rect 15000 7699 15111 7709
rect 15000 7698 15065 7699
rect 15000 7674 15008 7698
rect 15032 7675 15065 7698
rect 15089 7675 15111 7699
rect 15032 7674 15111 7675
rect 15000 7667 15111 7674
rect 15493 7707 15525 7772
rect 15705 7763 15736 7963
rect 15940 7962 15972 7963
rect 15937 7957 15972 7962
rect 15937 7937 15944 7957
rect 15964 7937 15972 7957
rect 15937 7929 15972 7937
rect 15705 7733 15711 7763
rect 15732 7733 15736 7763
rect 15705 7725 15736 7733
rect 15863 7707 15903 7708
rect 15493 7705 15905 7707
rect 15493 7679 15873 7705
rect 15899 7679 15905 7705
rect 15493 7671 15905 7679
rect 12449 7635 12473 7661
rect 12513 7635 12529 7661
rect 12313 7627 12348 7628
rect 12449 7623 12529 7635
rect 15493 7643 15525 7671
rect 15938 7651 15972 7929
rect 15493 7623 15498 7643
rect 15519 7623 15525 7643
rect 15493 7616 15525 7623
rect 15704 7643 15738 7650
rect 15704 7621 15711 7643
rect 15735 7621 15738 7643
rect 11604 7572 11715 7576
rect 13359 7572 13566 7573
rect 10924 7567 14999 7572
rect 10924 7554 15318 7567
rect 10924 7534 11612 7554
rect 11631 7534 11689 7554
rect 11708 7545 15318 7554
rect 11708 7534 15215 7545
rect 10924 7525 15215 7534
rect 15234 7525 15292 7545
rect 15311 7525 15318 7545
rect 10924 7516 15318 7525
rect 9920 7319 9996 7357
rect 10364 7319 10477 7379
rect 10926 7343 11033 7516
rect 13521 7514 15318 7516
rect 15207 7508 15318 7514
rect 11394 7477 11515 7487
rect 11394 7475 11463 7477
rect 11394 7434 11407 7475
rect 11444 7436 11463 7475
rect 11500 7436 11515 7477
rect 11444 7434 11515 7436
rect 11394 7416 11515 7434
rect 15542 7466 15594 7497
rect 15542 7432 15551 7466
rect 15580 7432 15594 7466
rect 9931 7218 9996 7319
rect 8867 7139 8884 7182
rect 5800 7090 5815 7124
rect 5844 7090 5852 7124
rect 8872 7134 8884 7139
rect 8930 7134 8944 7182
rect 8872 7112 8944 7134
rect 9929 7172 9996 7218
rect 10366 7180 10477 7319
rect 5800 7064 5852 7090
rect 9929 7080 9994 7172
rect 10361 7153 10477 7180
rect 10917 7316 11033 7343
rect 11400 7324 11465 7416
rect 15542 7406 15594 7432
rect 15704 7415 15738 7621
rect 15916 7646 15972 7651
rect 15916 7626 15923 7646
rect 15943 7626 15972 7646
rect 15916 7619 15972 7626
rect 15916 7618 15951 7619
rect 10917 7177 11028 7316
rect 11398 7278 11465 7324
rect 12450 7362 12522 7384
rect 12450 7314 12464 7362
rect 12510 7357 12522 7362
rect 15542 7372 15550 7406
rect 15579 7372 15594 7406
rect 12510 7314 12527 7357
rect 11398 7177 11463 7278
rect 5800 7030 5814 7064
rect 5843 7030 5852 7064
rect 5800 6999 5852 7030
rect 9879 7062 10000 7080
rect 9879 7060 9950 7062
rect 9879 7019 9894 7060
rect 9931 7021 9950 7060
rect 9987 7021 10000 7062
rect 9931 7019 10000 7021
rect 9879 7009 10000 7019
rect 6076 6982 6187 6988
rect 6076 6980 7873 6982
rect 10361 6980 10468 7153
rect 10917 7117 11030 7177
rect 11398 7139 11474 7177
rect 6076 6971 10470 6980
rect 6076 6951 6083 6971
rect 6102 6951 6160 6971
rect 6179 6962 10470 6971
rect 6179 6951 9686 6962
rect 6076 6942 9686 6951
rect 9705 6942 9763 6962
rect 9782 6942 10470 6962
rect 6076 6929 10470 6942
rect 6395 6924 10470 6929
rect 7828 6923 8035 6924
rect 9679 6920 9790 6924
rect 5443 6877 5478 6878
rect 5422 6870 5478 6877
rect 5422 6850 5451 6870
rect 5471 6850 5478 6870
rect 5422 6845 5478 6850
rect 5869 6873 5901 6880
rect 5869 6853 5875 6873
rect 5896 6853 5901 6873
rect 5422 6567 5456 6845
rect 5869 6825 5901 6853
rect 8865 6861 8945 6873
rect 9046 6868 9081 6869
rect 8865 6835 8881 6861
rect 8921 6835 8945 6861
rect 5489 6817 5901 6825
rect 5489 6791 5495 6817
rect 5521 6791 5901 6817
rect 5489 6789 5901 6791
rect 5491 6788 5531 6789
rect 5658 6763 5689 6771
rect 5658 6733 5662 6763
rect 5683 6733 5689 6763
rect 5422 6559 5457 6567
rect 5422 6539 5430 6559
rect 5450 6539 5457 6559
rect 5658 6548 5689 6733
rect 5869 6724 5901 6789
rect 6283 6822 6394 6829
rect 6283 6821 6362 6822
rect 6283 6797 6305 6821
rect 6329 6798 6362 6821
rect 6386 6798 6394 6822
rect 6329 6797 6394 6798
rect 6283 6787 6394 6797
rect 8865 6816 8945 6835
rect 8865 6790 8884 6816
rect 8924 6790 8945 6816
rect 6344 6770 6393 6787
rect 8865 6763 8945 6790
rect 8865 6737 8888 6763
rect 8928 6737 8945 6763
rect 8865 6726 8945 6737
rect 9025 6861 9081 6868
rect 9025 6841 9054 6861
rect 9074 6841 9081 6861
rect 9025 6836 9081 6841
rect 9472 6864 9504 6871
rect 9472 6844 9478 6864
rect 9499 6844 9504 6864
rect 5869 6704 5873 6724
rect 5894 6704 5901 6724
rect 5869 6697 5901 6704
rect 6178 6641 6279 6642
rect 6076 6628 6279 6641
rect 6076 6626 6219 6628
rect 6076 6623 6153 6626
rect 6076 6596 6079 6623
rect 6108 6599 6153 6623
rect 6182 6599 6219 6626
rect 6108 6596 6219 6599
rect 6076 6595 6219 6596
rect 6255 6595 6279 6628
rect 6076 6582 6279 6595
rect 5422 6534 5457 6539
rect 5422 6533 5454 6534
rect 5656 6471 5690 6548
rect 4289 5068 4886 5072
rect 1389 4990 1424 4992
rect 1389 4981 1493 4990
rect 1389 4980 1440 4981
rect 1389 4960 1392 4980
rect 1417 4961 1440 4980
rect 1472 4961 1493 4981
rect 1417 4960 1493 4961
rect 1389 4953 1493 4960
rect 1389 4941 1424 4953
rect 801 4875 1004 4888
rect 801 4842 825 4875
rect 861 4874 1004 4875
rect 861 4871 972 4874
rect 861 4844 898 4871
rect 927 4847 972 4871
rect 1001 4847 1004 4874
rect 927 4844 1004 4847
rect 861 4842 1004 4844
rect 801 4829 1004 4842
rect 801 4828 902 4829
rect 1179 4766 1211 4773
rect 1179 4746 1186 4766
rect 1207 4746 1211 4766
rect 690 4688 755 4697
rect 690 4651 700 4688
rect 740 4654 755 4688
rect 1179 4681 1211 4746
rect 1391 4737 1422 4941
rect 1626 4936 1658 4937
rect 1623 4931 1658 4936
rect 1623 4911 1630 4931
rect 1650 4911 1658 4931
rect 1623 4903 1658 4911
rect 1391 4707 1397 4737
rect 1418 4707 1422 4737
rect 1391 4699 1422 4707
rect 1549 4681 1589 4682
rect 1179 4679 1591 4681
rect 740 4651 757 4654
rect 690 4632 757 4651
rect 690 4611 704 4632
rect 740 4611 757 4632
rect 690 4604 757 4611
rect 1179 4653 1559 4679
rect 1585 4653 1591 4679
rect 1179 4645 1591 4653
rect 1179 4617 1211 4645
rect 1624 4625 1658 4903
rect 1748 4735 1813 5035
rect 3926 5023 4886 5068
rect 4993 5411 5029 6039
rect 3926 5019 4339 5023
rect 3926 4930 3960 5019
rect 4164 4933 4196 4934
rect 3339 4872 3542 4885
rect 3339 4839 3363 4872
rect 3399 4871 3542 4872
rect 3399 4868 3510 4871
rect 3399 4841 3436 4868
rect 3465 4844 3510 4868
rect 3539 4844 3542 4871
rect 3465 4841 3542 4844
rect 3399 4839 3542 4841
rect 3339 4826 3542 4839
rect 3339 4825 3440 4826
rect 3717 4763 3749 4770
rect 3717 4743 3724 4763
rect 3745 4743 3749 4763
rect 1179 4597 1184 4617
rect 1205 4597 1211 4617
rect 1179 4590 1211 4597
rect 1602 4620 1658 4625
rect 1602 4600 1609 4620
rect 1629 4600 1658 4620
rect 1602 4593 1658 4600
rect 1738 4724 1818 4735
rect 1738 4698 1755 4724
rect 1795 4698 1818 4724
rect 1738 4671 1818 4698
rect 1738 4645 1759 4671
rect 1799 4645 1818 4671
rect 1738 4626 1818 4645
rect 1738 4600 1762 4626
rect 1802 4600 1818 4626
rect 1602 4592 1637 4593
rect 1738 4588 1818 4600
rect 3717 4678 3749 4743
rect 3929 4734 3960 4930
rect 4161 4928 4196 4933
rect 4161 4908 4168 4928
rect 4188 4908 4196 4928
rect 4161 4900 4196 4908
rect 3929 4704 3935 4734
rect 3956 4704 3960 4734
rect 3929 4696 3960 4704
rect 4087 4678 4127 4679
rect 3717 4676 4129 4678
rect 3717 4650 4097 4676
rect 4123 4650 4129 4676
rect 3717 4642 4129 4650
rect 3717 4614 3749 4642
rect 4162 4622 4196 4900
rect 3717 4594 3722 4614
rect 3743 4594 3749 4614
rect 3717 4587 3749 4594
rect 4140 4617 4196 4622
rect 4140 4597 4147 4617
rect 4167 4597 4196 4617
rect 4140 4590 4196 4597
rect 4140 4589 4175 4590
rect 893 4537 1004 4541
rect 2648 4537 2855 4538
rect 3431 4537 3542 4538
rect 213 4519 4279 4537
rect 213 4499 901 4519
rect 920 4499 978 4519
rect 997 4516 4279 4519
rect 997 4499 3439 4516
rect 213 4496 3439 4499
rect 3458 4496 3516 4516
rect 3535 4496 4279 4516
rect 213 4481 4279 4496
rect 215 4293 322 4481
rect 2810 4479 4279 4481
rect 683 4442 804 4452
rect 683 4440 752 4442
rect 683 4399 696 4440
rect 733 4401 752 4440
rect 789 4401 804 4442
rect 733 4399 804 4401
rect 683 4381 804 4399
rect 215 4289 323 4293
rect 689 4289 766 4381
rect 1739 4377 1815 4393
rect 1739 4354 1754 4377
rect 216 3696 323 4289
rect 691 4238 766 4289
rect 1732 4340 1754 4354
rect 1798 4340 1815 4377
rect 1732 4320 1815 4340
rect 1732 4254 1749 4320
rect 1803 4254 1815 4320
rect 691 4195 767 4238
rect 695 3884 767 4195
rect 1732 4230 1815 4254
rect 1732 4210 1808 4230
rect 1732 4191 1811 4210
rect 1391 4175 1463 4176
rect 1390 4167 1489 4175
rect 1390 4164 1442 4167
rect 1390 4129 1398 4164
rect 1423 4129 1442 4164
rect 1467 4129 1489 4167
rect 1390 4117 1489 4129
rect 1391 4098 1459 4117
rect 1392 4095 1425 4098
rect 1627 4095 1659 4096
rect 802 4034 1005 4047
rect 802 4001 826 4034
rect 862 4033 1005 4034
rect 862 4030 973 4033
rect 862 4003 899 4030
rect 928 4006 973 4030
rect 1002 4006 1005 4033
rect 928 4003 1005 4006
rect 862 4001 1005 4003
rect 802 3988 1005 4001
rect 802 3987 903 3988
rect 695 3842 704 3884
rect 753 3842 767 3884
rect 695 3821 767 3842
rect 695 3779 705 3821
rect 754 3779 767 3821
rect 695 3761 767 3779
rect 1180 3925 1212 3932
rect 1180 3905 1187 3925
rect 1208 3905 1212 3925
rect 1180 3840 1212 3905
rect 1392 3896 1423 4095
rect 1624 4090 1659 4095
rect 1624 4070 1631 4090
rect 1651 4070 1659 4090
rect 1624 4062 1659 4070
rect 1392 3866 1398 3896
rect 1419 3866 1423 3896
rect 1392 3858 1423 3866
rect 1550 3840 1590 3841
rect 1180 3838 1592 3840
rect 1180 3812 1560 3838
rect 1586 3812 1592 3838
rect 1180 3804 1592 3812
rect 1180 3776 1212 3804
rect 1625 3784 1659 4062
rect 1741 3875 1811 4191
rect 3729 4176 3760 4177
rect 3729 4168 3774 4176
rect 2809 4145 2973 4152
rect 3729 4145 3739 4168
rect 2435 4130 3739 4145
rect 3764 4130 3774 4168
rect 4993 4171 5027 5411
rect 4993 4167 5223 4171
rect 4993 4141 5192 4167
rect 5217 4141 5223 4167
rect 4993 4133 5223 4141
rect 2435 4112 3774 4130
rect 2440 4099 2476 4112
rect 2809 4109 2973 4112
rect 1850 4030 2053 4043
rect 1850 3997 1874 4030
rect 1910 4029 2053 4030
rect 1910 4026 2021 4029
rect 1910 3999 1947 4026
rect 1976 4002 2021 4026
rect 2050 4002 2053 4029
rect 1976 3999 2053 4002
rect 1910 3997 2053 3999
rect 1850 3984 2053 3997
rect 1850 3983 1951 3984
rect 1180 3756 1185 3776
rect 1206 3756 1212 3776
rect 1180 3749 1212 3756
rect 1603 3779 1659 3784
rect 1603 3759 1610 3779
rect 1630 3759 1659 3779
rect 1736 3869 1811 3875
rect 1736 3836 1744 3869
rect 1797 3836 1811 3869
rect 1736 3811 1811 3836
rect 1736 3778 1749 3811
rect 1802 3778 1811 3811
rect 1736 3769 1811 3778
rect 2228 3921 2260 3928
rect 2228 3901 2235 3921
rect 2256 3901 2260 3921
rect 2228 3836 2260 3901
rect 2440 3892 2471 4099
rect 2675 4091 2707 4092
rect 2672 4086 2707 4091
rect 2672 4066 2679 4086
rect 2699 4066 2707 4086
rect 2672 4058 2707 4066
rect 2440 3862 2446 3892
rect 2467 3862 2471 3892
rect 2440 3854 2471 3862
rect 2598 3836 2638 3837
rect 2228 3834 2640 3836
rect 2228 3808 2608 3834
rect 2634 3808 2640 3834
rect 2228 3800 2640 3808
rect 2228 3772 2260 3800
rect 2673 3780 2707 4058
rect 4752 4036 4955 4049
rect 4752 4003 4776 4036
rect 4812 4035 4955 4036
rect 4812 4032 4923 4035
rect 4812 4005 4849 4032
rect 4878 4008 4923 4032
rect 4952 4008 4955 4035
rect 4878 4005 4955 4008
rect 4812 4003 4955 4005
rect 4752 3990 4955 4003
rect 4752 3989 4853 3990
rect 1736 3764 1794 3769
rect 1603 3752 1659 3759
rect 2228 3752 2233 3772
rect 2254 3752 2260 3772
rect 1603 3751 1638 3752
rect 2228 3745 2260 3752
rect 2651 3775 2707 3780
rect 2651 3755 2658 3775
rect 2678 3755 2707 3775
rect 2651 3748 2707 3755
rect 5130 3927 5162 3934
rect 5130 3907 5137 3927
rect 5158 3907 5162 3927
rect 5130 3842 5162 3907
rect 5342 3898 5373 4098
rect 5577 4097 5609 4098
rect 5574 4092 5609 4097
rect 5574 4072 5581 4092
rect 5601 4072 5609 4092
rect 5574 4064 5609 4072
rect 5342 3868 5348 3898
rect 5369 3868 5373 3898
rect 5342 3860 5373 3868
rect 5500 3842 5540 3843
rect 5130 3840 5542 3842
rect 5130 3814 5510 3840
rect 5536 3814 5542 3840
rect 5130 3806 5542 3814
rect 5130 3778 5162 3806
rect 5130 3758 5135 3778
rect 5156 3758 5162 3778
rect 5130 3751 5162 3758
rect 5332 3780 5380 3787
rect 5575 3786 5609 4064
rect 5332 3760 5339 3780
rect 5372 3760 5380 3780
rect 2651 3747 2686 3748
rect 894 3696 1005 3700
rect 2677 3696 4247 3697
rect 216 3692 4247 3696
rect 4572 3692 4990 3705
rect 216 3680 4990 3692
rect 216 3678 4852 3680
rect 216 3658 902 3678
rect 921 3658 979 3678
rect 998 3674 4852 3678
rect 998 3658 1950 3674
rect 216 3654 1950 3658
rect 1969 3654 2027 3674
rect 2046 3660 4852 3674
rect 4871 3660 4929 3680
rect 4948 3660 4990 3680
rect 2046 3654 4990 3660
rect 216 3640 4990 3654
rect 216 3017 323 3640
rect 1942 3637 2053 3640
rect 4572 3634 4990 3640
rect 702 3591 766 3595
rect 698 3585 766 3591
rect 698 3552 715 3585
rect 755 3552 766 3585
rect 698 3540 766 3552
rect 1749 3554 1814 3576
rect 698 3538 755 3540
rect 702 3177 753 3538
rect 1749 3515 1766 3554
rect 1811 3515 1814 3554
rect 1390 3470 1425 3472
rect 1390 3461 1494 3470
rect 1390 3460 1441 3461
rect 1390 3440 1393 3460
rect 1418 3441 1441 3460
rect 1473 3441 1494 3461
rect 1418 3440 1494 3441
rect 1390 3433 1494 3440
rect 1390 3421 1425 3433
rect 802 3355 1005 3368
rect 802 3322 826 3355
rect 862 3354 1005 3355
rect 862 3351 973 3354
rect 862 3324 899 3351
rect 928 3327 973 3351
rect 1002 3327 1005 3354
rect 928 3324 1005 3327
rect 862 3322 1005 3324
rect 802 3309 1005 3322
rect 802 3308 903 3309
rect 1180 3246 1212 3253
rect 1180 3226 1187 3246
rect 1208 3226 1212 3246
rect 691 3168 756 3177
rect 691 3131 701 3168
rect 741 3134 756 3168
rect 1180 3161 1212 3226
rect 1392 3217 1423 3421
rect 1627 3416 1659 3417
rect 1624 3411 1659 3416
rect 1624 3391 1631 3411
rect 1651 3391 1659 3411
rect 1624 3383 1659 3391
rect 1392 3187 1398 3217
rect 1419 3187 1423 3217
rect 1392 3179 1423 3187
rect 1550 3161 1590 3162
rect 1180 3159 1592 3161
rect 741 3131 758 3134
rect 691 3112 758 3131
rect 691 3091 705 3112
rect 741 3091 758 3112
rect 691 3084 758 3091
rect 1180 3133 1560 3159
rect 1586 3133 1592 3159
rect 1180 3125 1592 3133
rect 1180 3097 1212 3125
rect 1625 3105 1659 3383
rect 1749 3215 1814 3515
rect 3886 3476 3923 3497
rect 3886 3439 3897 3476
rect 3914 3452 3923 3476
rect 3914 3439 3924 3452
rect 3886 3429 3924 3439
rect 3887 3425 3924 3429
rect 3887 3419 3920 3425
rect 3297 3350 3500 3363
rect 3297 3317 3321 3350
rect 3357 3349 3500 3350
rect 3357 3346 3468 3349
rect 3357 3319 3394 3346
rect 3423 3322 3468 3346
rect 3497 3322 3500 3349
rect 3423 3319 3500 3322
rect 3357 3317 3500 3319
rect 3297 3304 3500 3317
rect 3297 3303 3398 3304
rect 3675 3241 3707 3248
rect 3675 3221 3682 3241
rect 3703 3221 3707 3241
rect 1180 3077 1185 3097
rect 1206 3077 1212 3097
rect 1180 3070 1212 3077
rect 1603 3100 1659 3105
rect 1603 3080 1610 3100
rect 1630 3080 1659 3100
rect 1603 3073 1659 3080
rect 1739 3204 1819 3215
rect 1739 3178 1756 3204
rect 1796 3178 1819 3204
rect 1739 3151 1819 3178
rect 1739 3125 1760 3151
rect 1800 3125 1819 3151
rect 1739 3106 1819 3125
rect 1739 3080 1763 3106
rect 1803 3080 1819 3106
rect 2813 3150 2918 3171
rect 3675 3156 3707 3221
rect 3887 3212 3918 3419
rect 4122 3411 4154 3412
rect 4119 3406 4154 3411
rect 4119 3386 4126 3406
rect 4146 3386 4154 3406
rect 4119 3378 4154 3386
rect 3887 3182 3893 3212
rect 3914 3182 3918 3212
rect 3887 3174 3918 3182
rect 4045 3156 4085 3157
rect 3675 3154 4087 3156
rect 2813 3144 3289 3150
rect 2813 3142 2870 3144
rect 2813 3111 2825 3142
rect 2850 3121 2870 3142
rect 2896 3137 3289 3144
rect 2896 3121 3250 3137
rect 2850 3114 3250 3121
rect 3276 3114 3289 3137
rect 2850 3111 3289 3114
rect 2813 3101 3289 3111
rect 3675 3128 4055 3154
rect 4081 3128 4087 3154
rect 3675 3120 4087 3128
rect 2813 3099 2918 3101
rect 1603 3072 1638 3073
rect 1739 3068 1819 3080
rect 3675 3092 3707 3120
rect 4120 3100 4154 3378
rect 3675 3072 3680 3092
rect 3701 3072 3707 3092
rect 3675 3065 3707 3072
rect 4098 3095 4154 3100
rect 4098 3075 4105 3095
rect 4125 3075 4154 3095
rect 4098 3068 4154 3075
rect 4098 3067 4133 3068
rect 894 3017 1005 3021
rect 2636 3017 4289 3020
rect 214 2999 4289 3017
rect 214 2979 902 2999
rect 921 2979 979 2999
rect 998 2994 4289 2999
rect 998 2979 3397 2994
rect 214 2974 3397 2979
rect 3416 2974 3474 2994
rect 3493 2974 4289 2994
rect 214 2964 4289 2974
rect 214 2961 839 2964
rect 1026 2961 4289 2964
rect 216 2733 323 2961
rect 2636 2960 4289 2961
rect 3389 2957 3500 2960
rect 684 2922 805 2932
rect 684 2920 753 2922
rect 684 2879 697 2920
rect 734 2881 753 2920
rect 790 2881 805 2922
rect 734 2879 805 2881
rect 684 2861 805 2879
rect 690 2759 769 2861
rect 1742 2821 1809 2840
rect 1742 2801 1762 2821
rect 216 2678 324 2733
rect 691 2678 769 2759
rect 1741 2755 1762 2801
rect 1792 2801 1809 2821
rect 1792 2771 1811 2801
rect 1792 2755 1812 2771
rect 1741 2739 1812 2755
rect 1391 2728 1463 2729
rect 1390 2720 1489 2728
rect 1390 2717 1442 2720
rect 1390 2682 1398 2717
rect 1423 2682 1442 2717
rect 1467 2682 1489 2720
rect 216 2249 323 2678
rect 695 2437 767 2678
rect 1390 2670 1489 2682
rect 1391 2651 1459 2670
rect 1392 2648 1425 2651
rect 1627 2648 1659 2649
rect 802 2587 1005 2600
rect 802 2554 826 2587
rect 862 2586 1005 2587
rect 862 2583 973 2586
rect 862 2556 899 2583
rect 928 2559 973 2583
rect 1002 2559 1005 2586
rect 928 2556 1005 2559
rect 862 2554 1005 2556
rect 802 2541 1005 2554
rect 802 2540 903 2541
rect 695 2395 704 2437
rect 753 2395 767 2437
rect 695 2374 767 2395
rect 695 2332 705 2374
rect 754 2332 767 2374
rect 695 2314 767 2332
rect 1180 2478 1212 2485
rect 1180 2458 1187 2478
rect 1208 2458 1212 2478
rect 1180 2393 1212 2458
rect 1392 2449 1423 2648
rect 1624 2643 1659 2648
rect 1624 2623 1631 2643
rect 1651 2623 1659 2643
rect 1624 2615 1659 2623
rect 1392 2419 1398 2449
rect 1419 2419 1423 2449
rect 1392 2411 1423 2419
rect 1550 2393 1590 2394
rect 1180 2391 1592 2393
rect 1180 2365 1560 2391
rect 1586 2365 1592 2391
rect 1180 2357 1592 2365
rect 1180 2329 1212 2357
rect 1625 2337 1659 2615
rect 1741 2428 1811 2739
rect 2438 2730 3780 2735
rect 2438 2728 3737 2730
rect 2435 2702 3737 2728
rect 3765 2702 3780 2730
rect 2435 2694 3780 2702
rect 2435 2669 2474 2694
rect 2435 2652 2476 2669
rect 2435 2645 2474 2652
rect 1850 2583 2053 2596
rect 1850 2550 1874 2583
rect 1910 2582 2053 2583
rect 1910 2579 2021 2582
rect 1910 2552 1947 2579
rect 1976 2555 2021 2579
rect 2050 2555 2053 2582
rect 1976 2552 2053 2555
rect 1910 2550 2053 2552
rect 1850 2537 2053 2550
rect 1850 2536 1951 2537
rect 1180 2309 1185 2329
rect 1206 2309 1212 2329
rect 1180 2302 1212 2309
rect 1603 2332 1659 2337
rect 1603 2312 1610 2332
rect 1630 2312 1659 2332
rect 1736 2422 1811 2428
rect 1736 2389 1744 2422
rect 1797 2389 1811 2422
rect 1736 2364 1811 2389
rect 1736 2331 1749 2364
rect 1802 2331 1811 2364
rect 1736 2322 1811 2331
rect 2228 2474 2260 2481
rect 2228 2454 2235 2474
rect 2256 2454 2260 2474
rect 2228 2389 2260 2454
rect 2440 2445 2471 2645
rect 2675 2644 2707 2645
rect 2672 2639 2707 2644
rect 2672 2619 2679 2639
rect 2699 2619 2707 2639
rect 2672 2611 2707 2619
rect 2440 2415 2446 2445
rect 2467 2415 2471 2445
rect 2440 2407 2471 2415
rect 2598 2389 2638 2390
rect 2228 2387 2640 2389
rect 2228 2361 2608 2387
rect 2634 2361 2640 2387
rect 2228 2353 2640 2361
rect 2228 2325 2260 2353
rect 2673 2333 2707 2611
rect 1736 2317 1794 2322
rect 1603 2305 1659 2312
rect 2228 2305 2233 2325
rect 2254 2305 2260 2325
rect 1603 2304 1638 2305
rect 2228 2298 2260 2305
rect 2651 2328 2707 2333
rect 2651 2308 2658 2328
rect 2678 2308 2707 2328
rect 2651 2301 2707 2308
rect 2651 2300 2686 2301
rect 894 2249 1005 2253
rect 2769 2249 4289 2250
rect 216 2231 4289 2249
rect 216 2211 902 2231
rect 921 2211 979 2231
rect 998 2227 4289 2231
rect 998 2211 1950 2227
rect 216 2207 1950 2211
rect 1969 2207 2027 2227
rect 2046 2207 4289 2227
rect 216 2193 4289 2207
rect 216 1570 323 2193
rect 1942 2190 2053 2193
rect 702 2144 766 2148
rect 698 2138 766 2144
rect 698 2105 715 2138
rect 755 2105 766 2138
rect 698 2093 766 2105
rect 1749 2107 1814 2129
rect 698 2091 755 2093
rect 702 1730 753 2091
rect 1749 2068 1766 2107
rect 1811 2068 1814 2107
rect 1390 2023 1425 2025
rect 1390 2014 1494 2023
rect 1390 2013 1441 2014
rect 1390 1993 1393 2013
rect 1418 1994 1441 2013
rect 1473 1994 1494 2014
rect 1418 1993 1494 1994
rect 1390 1986 1494 1993
rect 1390 1974 1425 1986
rect 802 1908 1005 1921
rect 802 1875 826 1908
rect 862 1907 1005 1908
rect 862 1904 973 1907
rect 862 1877 899 1904
rect 928 1880 973 1904
rect 1002 1880 1005 1907
rect 928 1877 1005 1880
rect 862 1875 1005 1877
rect 802 1862 1005 1875
rect 802 1861 903 1862
rect 1180 1799 1212 1806
rect 1180 1779 1187 1799
rect 1208 1779 1212 1799
rect 691 1721 756 1730
rect 691 1684 701 1721
rect 741 1687 756 1721
rect 1180 1714 1212 1779
rect 1392 1770 1423 1974
rect 1627 1969 1659 1970
rect 1624 1964 1659 1969
rect 1624 1944 1631 1964
rect 1651 1944 1659 1964
rect 1624 1936 1659 1944
rect 1392 1740 1398 1770
rect 1419 1740 1423 1770
rect 1392 1732 1423 1740
rect 1550 1714 1590 1715
rect 1180 1712 1592 1714
rect 741 1684 758 1687
rect 691 1665 758 1684
rect 691 1644 705 1665
rect 741 1644 758 1665
rect 691 1637 758 1644
rect 1180 1686 1560 1712
rect 1586 1686 1592 1712
rect 1180 1678 1592 1686
rect 1180 1650 1212 1678
rect 1625 1658 1659 1936
rect 1749 1805 1814 2068
rect 1749 1801 1810 1805
rect 1180 1630 1185 1650
rect 1206 1630 1212 1650
rect 1180 1623 1212 1630
rect 1603 1653 1659 1658
rect 1603 1633 1610 1653
rect 1630 1633 1659 1653
rect 1603 1626 1659 1633
rect 1603 1625 1638 1626
rect 894 1570 1005 1574
rect 214 1552 1533 1570
rect 214 1532 902 1552
rect 921 1532 979 1552
rect 998 1532 1533 1552
rect 214 1514 1533 1532
rect 216 1394 323 1514
rect 684 1475 805 1485
rect 684 1473 753 1475
rect 684 1432 697 1473
rect 734 1434 753 1473
rect 790 1434 805 1475
rect 734 1432 805 1434
rect 684 1414 805 1432
rect 15 1321 149 1350
rect 15 1209 53 1321
rect 132 1209 149 1321
rect 216 1314 324 1394
rect 15 256 149 1209
rect 217 502 324 1314
rect 690 1342 755 1414
rect 690 1276 758 1342
rect 691 730 758 1276
rect 1745 914 1810 1801
rect 2788 1531 2925 1535
rect 2775 1527 2932 1531
rect 2775 1420 2812 1527
rect 2912 1420 2932 1527
rect 2775 1378 2932 1420
rect 2788 1130 2925 1378
rect 2778 1088 2944 1130
rect 2778 1013 2807 1088
rect 2924 1013 2944 1088
rect 2778 997 2944 1013
rect 1734 893 1871 914
rect 1734 818 1759 893
rect 1829 818 1871 893
rect 1734 787 1871 818
rect 677 681 852 730
rect 677 602 710 681
rect 810 602 852 681
rect 677 597 852 602
rect 217 460 365 502
rect 217 452 257 460
rect 219 373 257 452
rect 327 373 365 460
rect 219 335 365 373
rect 11 220 150 256
rect 11 125 25 220
rect 115 125 150 220
rect 11 107 150 125
rect 5332 30 5380 3760
rect 5553 3781 5609 3786
rect 5553 3761 5560 3781
rect 5580 3761 5609 3781
rect 5553 3754 5609 3761
rect 5553 3753 5588 3754
rect 5657 3663 5685 6471
rect 8870 6426 8935 6726
rect 9025 6558 9059 6836
rect 9472 6816 9504 6844
rect 9092 6808 9504 6816
rect 9092 6782 9098 6808
rect 9124 6782 9504 6808
rect 9926 6850 9993 6857
rect 9926 6829 9943 6850
rect 9979 6829 9993 6850
rect 9926 6810 9993 6829
rect 9926 6807 9943 6810
rect 9092 6780 9504 6782
rect 9094 6779 9134 6780
rect 9261 6754 9292 6762
rect 9261 6724 9265 6754
rect 9286 6724 9292 6754
rect 9025 6550 9060 6558
rect 9025 6530 9033 6550
rect 9053 6530 9060 6550
rect 9025 6525 9060 6530
rect 9025 6524 9057 6525
rect 9261 6520 9292 6724
rect 9472 6715 9504 6780
rect 9928 6773 9943 6807
rect 9983 6773 9993 6810
rect 9928 6764 9993 6773
rect 9472 6695 9476 6715
rect 9497 6695 9504 6715
rect 9472 6688 9504 6695
rect 9781 6632 9882 6633
rect 9679 6619 9882 6632
rect 9679 6617 9822 6619
rect 9679 6614 9756 6617
rect 9679 6587 9682 6614
rect 9711 6590 9756 6614
rect 9785 6590 9822 6617
rect 9711 6587 9822 6590
rect 9679 6586 9822 6587
rect 9858 6586 9882 6619
rect 9679 6573 9882 6586
rect 9259 6508 9294 6520
rect 9190 6501 9294 6508
rect 9190 6500 9266 6501
rect 9190 6480 9211 6500
rect 9243 6481 9266 6500
rect 9291 6481 9294 6501
rect 9243 6480 9294 6481
rect 9190 6471 9294 6480
rect 9259 6469 9294 6471
rect 8870 6387 8873 6426
rect 8918 6387 8935 6426
rect 9931 6403 9982 6764
rect 9929 6401 9986 6403
rect 8870 6365 8935 6387
rect 9918 6389 9986 6401
rect 9918 6356 9929 6389
rect 9969 6356 9986 6389
rect 9918 6350 9986 6356
rect 9918 6346 9982 6350
rect 8631 6301 8742 6304
rect 10361 6301 10468 6924
rect 6925 6287 10468 6301
rect 6925 6267 8638 6287
rect 8657 6267 8715 6287
rect 8734 6283 10468 6287
rect 8734 6267 9686 6283
rect 6925 6263 9686 6267
rect 9705 6263 9763 6283
rect 9782 6263 10468 6283
rect 6925 6245 10468 6263
rect 6925 6244 7915 6245
rect 9679 6241 9790 6245
rect 7998 6193 8033 6194
rect 7977 6186 8033 6193
rect 7977 6166 8006 6186
rect 8026 6166 8033 6186
rect 7977 6161 8033 6166
rect 8424 6189 8456 6196
rect 9046 6189 9081 6190
rect 8424 6169 8430 6189
rect 8451 6169 8456 6189
rect 9025 6182 9081 6189
rect 8890 6172 8948 6177
rect 7977 5883 8011 6161
rect 8424 6141 8456 6169
rect 8044 6133 8456 6141
rect 8044 6107 8050 6133
rect 8076 6107 8456 6133
rect 8044 6105 8456 6107
rect 8046 6104 8086 6105
rect 8213 6079 8244 6087
rect 8213 6049 8217 6079
rect 8238 6049 8244 6079
rect 7977 5875 8012 5883
rect 7977 5855 7985 5875
rect 8005 5855 8012 5875
rect 7977 5850 8012 5855
rect 7977 5849 8009 5850
rect 8213 5849 8244 6049
rect 8424 6040 8456 6105
rect 8424 6020 8428 6040
rect 8449 6020 8456 6040
rect 8424 6013 8456 6020
rect 8873 6163 8948 6172
rect 8873 6130 8882 6163
rect 8935 6130 8948 6163
rect 8873 6105 8948 6130
rect 8873 6072 8887 6105
rect 8940 6072 8948 6105
rect 8873 6066 8948 6072
rect 9025 6162 9054 6182
rect 9074 6162 9081 6182
rect 9025 6157 9081 6162
rect 9472 6185 9504 6192
rect 9472 6165 9478 6185
rect 9499 6165 9504 6185
rect 8733 5957 8834 5958
rect 8631 5944 8834 5957
rect 8631 5942 8774 5944
rect 8631 5939 8708 5942
rect 8631 5912 8634 5939
rect 8663 5915 8708 5939
rect 8737 5915 8774 5942
rect 8663 5912 8774 5915
rect 8631 5911 8774 5912
rect 8810 5911 8834 5944
rect 8631 5898 8834 5911
rect 8210 5842 8249 5849
rect 8208 5825 8249 5842
rect 8210 5800 8249 5825
rect 6904 5792 8249 5800
rect 6904 5764 6919 5792
rect 6947 5766 8249 5792
rect 6947 5764 8246 5766
rect 6904 5759 8246 5764
rect 8873 5755 8943 6066
rect 9025 5879 9059 6157
rect 9472 6137 9504 6165
rect 9092 6129 9504 6137
rect 9092 6103 9098 6129
rect 9124 6103 9504 6129
rect 9092 6101 9504 6103
rect 9094 6100 9134 6101
rect 9261 6075 9292 6083
rect 9261 6045 9265 6075
rect 9286 6045 9292 6075
rect 9025 5871 9060 5879
rect 9025 5851 9033 5871
rect 9053 5851 9060 5871
rect 9025 5846 9060 5851
rect 9261 5846 9292 6045
rect 9472 6036 9504 6101
rect 9472 6016 9476 6036
rect 9497 6016 9504 6036
rect 9472 6009 9504 6016
rect 9917 6162 9989 6180
rect 9917 6120 9930 6162
rect 9979 6120 9989 6162
rect 9917 6099 9989 6120
rect 9917 6057 9931 6099
rect 9980 6057 9989 6099
rect 9781 5953 9882 5954
rect 9679 5940 9882 5953
rect 9679 5938 9822 5940
rect 9679 5935 9756 5938
rect 9679 5908 9682 5935
rect 9711 5911 9756 5935
rect 9785 5911 9822 5938
rect 9711 5908 9822 5911
rect 9679 5907 9822 5908
rect 9858 5907 9882 5940
rect 9679 5894 9882 5907
rect 9025 5845 9057 5846
rect 9259 5843 9292 5846
rect 9225 5824 9293 5843
rect 9195 5812 9294 5824
rect 9917 5816 9989 6057
rect 10361 5816 10468 6245
rect 10923 6657 11030 7117
rect 11402 6845 11474 7139
rect 12098 7136 12170 7137
rect 12097 7128 12196 7136
rect 12450 7131 12527 7314
rect 13738 7315 13822 7326
rect 13738 7287 13766 7315
rect 13810 7287 13822 7315
rect 13552 7236 13626 7264
rect 13552 7188 13575 7236
rect 13612 7188 13626 7236
rect 13738 7258 13822 7287
rect 13738 7230 13763 7258
rect 13807 7230 13822 7258
rect 13738 7197 13822 7230
rect 13552 7179 13626 7188
rect 13148 7137 13220 7138
rect 12097 7125 12149 7128
rect 12097 7090 12105 7125
rect 12130 7090 12149 7125
rect 12174 7090 12196 7128
rect 12097 7078 12196 7090
rect 12448 7102 12527 7131
rect 13147 7129 13236 7137
rect 13147 7126 13199 7129
rect 12098 7059 12166 7078
rect 12099 7056 12132 7059
rect 12334 7056 12366 7057
rect 11509 6995 11712 7008
rect 11509 6962 11533 6995
rect 11569 6994 11712 6995
rect 11569 6991 11680 6994
rect 11569 6964 11606 6991
rect 11635 6967 11680 6991
rect 11709 6967 11712 6994
rect 11635 6964 11712 6967
rect 11569 6962 11712 6964
rect 11509 6949 11712 6962
rect 11509 6948 11610 6949
rect 11402 6803 11411 6845
rect 11460 6803 11474 6845
rect 11402 6782 11474 6803
rect 11402 6740 11412 6782
rect 11461 6740 11474 6782
rect 11402 6722 11474 6740
rect 11887 6886 11919 6893
rect 11887 6866 11894 6886
rect 11915 6866 11919 6886
rect 11887 6801 11919 6866
rect 12099 6857 12130 7056
rect 12331 7051 12366 7056
rect 12331 7031 12338 7051
rect 12358 7031 12366 7051
rect 12331 7023 12366 7031
rect 12099 6827 12105 6857
rect 12126 6827 12130 6857
rect 12099 6819 12130 6827
rect 12257 6801 12297 6802
rect 11887 6799 12299 6801
rect 11887 6773 12267 6799
rect 12293 6773 12299 6799
rect 11887 6765 12299 6773
rect 11887 6737 11919 6765
rect 12332 6745 12366 7023
rect 12448 6836 12518 7102
rect 13147 7091 13155 7126
rect 13180 7091 13199 7126
rect 13224 7091 13236 7129
rect 13147 7079 13236 7091
rect 13147 7078 13216 7079
rect 13147 7060 13183 7078
rect 12557 6991 12760 7004
rect 12557 6958 12581 6991
rect 12617 6990 12760 6991
rect 12617 6987 12728 6990
rect 12617 6960 12654 6987
rect 12683 6963 12728 6987
rect 12757 6963 12760 6990
rect 12683 6960 12760 6963
rect 12617 6958 12760 6960
rect 12557 6945 12760 6958
rect 12557 6944 12658 6945
rect 11887 6717 11892 6737
rect 11913 6717 11919 6737
rect 11887 6710 11919 6717
rect 12310 6740 12366 6745
rect 12310 6720 12317 6740
rect 12337 6720 12366 6740
rect 12443 6830 12518 6836
rect 12443 6797 12451 6830
rect 12504 6797 12518 6830
rect 12443 6772 12518 6797
rect 12443 6739 12456 6772
rect 12509 6739 12518 6772
rect 12443 6730 12518 6739
rect 12935 6882 12967 6889
rect 12935 6862 12942 6882
rect 12963 6862 12967 6882
rect 12935 6797 12967 6862
rect 13147 6853 13178 7060
rect 13382 7052 13414 7053
rect 13379 7047 13414 7052
rect 13379 7027 13386 7047
rect 13406 7027 13414 7047
rect 13379 7019 13414 7027
rect 13147 6823 13153 6853
rect 13174 6823 13178 6853
rect 13147 6815 13178 6823
rect 13305 6797 13345 6798
rect 12935 6795 13347 6797
rect 12935 6769 13315 6795
rect 13341 6769 13347 6795
rect 12935 6761 13347 6769
rect 12935 6733 12967 6761
rect 13380 6741 13414 7019
rect 13563 6834 13625 7179
rect 13732 7152 13822 7197
rect 13732 6837 13814 7152
rect 13563 6815 13627 6834
rect 13563 6776 13576 6815
rect 13610 6776 13627 6815
rect 13563 6757 13627 6776
rect 13732 6796 13753 6837
rect 13789 6796 13814 6837
rect 13732 6767 13814 6796
rect 12443 6725 12501 6730
rect 12310 6713 12366 6720
rect 12935 6713 12940 6733
rect 12961 6713 12967 6733
rect 12310 6712 12345 6713
rect 12935 6706 12967 6713
rect 13358 6736 13414 6741
rect 13358 6716 13365 6736
rect 13385 6716 13414 6736
rect 13358 6709 13414 6716
rect 13358 6708 13393 6709
rect 11601 6657 11712 6661
rect 13384 6657 14954 6658
rect 10923 6639 14954 6657
rect 10923 6619 11609 6639
rect 11628 6619 11686 6639
rect 11705 6635 14954 6639
rect 11705 6619 12657 6635
rect 10923 6615 12657 6619
rect 12676 6615 12734 6635
rect 12753 6615 14954 6635
rect 10923 6601 14954 6615
rect 10923 5978 11030 6601
rect 12649 6598 12760 6601
rect 11409 6552 11473 6556
rect 11405 6546 11473 6552
rect 11405 6513 11422 6546
rect 11462 6513 11473 6546
rect 11405 6501 11473 6513
rect 12456 6515 12521 6537
rect 11405 6499 11462 6501
rect 11409 6138 11460 6499
rect 12456 6476 12473 6515
rect 12518 6476 12521 6515
rect 12097 6431 12132 6433
rect 12097 6422 12201 6431
rect 12097 6421 12148 6422
rect 12097 6401 12100 6421
rect 12125 6402 12148 6421
rect 12180 6402 12201 6422
rect 12125 6401 12201 6402
rect 12097 6394 12201 6401
rect 12097 6382 12132 6394
rect 11509 6316 11712 6329
rect 11509 6283 11533 6316
rect 11569 6315 11712 6316
rect 11569 6312 11680 6315
rect 11569 6285 11606 6312
rect 11635 6288 11680 6312
rect 11709 6288 11712 6315
rect 11635 6285 11712 6288
rect 11569 6283 11712 6285
rect 11509 6270 11712 6283
rect 11509 6269 11610 6270
rect 11887 6207 11919 6214
rect 11887 6187 11894 6207
rect 11915 6187 11919 6207
rect 11398 6129 11463 6138
rect 11398 6092 11408 6129
rect 11448 6095 11463 6129
rect 11887 6122 11919 6187
rect 12099 6178 12130 6382
rect 12334 6377 12366 6378
rect 12331 6372 12366 6377
rect 12331 6352 12338 6372
rect 12358 6352 12366 6372
rect 12331 6344 12366 6352
rect 12099 6148 12105 6178
rect 12126 6148 12130 6178
rect 12099 6140 12130 6148
rect 12257 6122 12297 6123
rect 11887 6120 12299 6122
rect 11448 6092 11465 6095
rect 11398 6073 11465 6092
rect 11398 6052 11412 6073
rect 11448 6052 11465 6073
rect 11398 6045 11465 6052
rect 11887 6094 12267 6120
rect 12293 6094 12299 6120
rect 11887 6086 12299 6094
rect 11887 6058 11919 6086
rect 12332 6066 12366 6344
rect 12456 6176 12521 6476
rect 13727 6500 13820 6515
rect 13727 6456 13742 6500
rect 13802 6456 13820 6500
rect 11887 6038 11892 6058
rect 11913 6038 11919 6058
rect 11887 6031 11919 6038
rect 12310 6061 12366 6066
rect 12310 6041 12317 6061
rect 12337 6041 12366 6061
rect 12310 6034 12366 6041
rect 12446 6165 12526 6176
rect 12446 6139 12463 6165
rect 12503 6139 12526 6165
rect 12446 6112 12526 6139
rect 12446 6086 12467 6112
rect 12507 6086 12526 6112
rect 12446 6067 12526 6086
rect 12446 6041 12470 6067
rect 12510 6041 12526 6067
rect 12310 6033 12345 6034
rect 12446 6029 12526 6041
rect 13727 6083 13820 6456
rect 14004 6311 14207 6324
rect 14004 6278 14028 6311
rect 14064 6310 14207 6311
rect 14064 6307 14175 6310
rect 14064 6280 14101 6307
rect 14130 6283 14175 6307
rect 14204 6283 14207 6310
rect 14130 6280 14207 6283
rect 14064 6278 14207 6280
rect 14004 6265 14207 6278
rect 14004 6264 14105 6265
rect 13727 6042 13742 6083
rect 13796 6042 13820 6083
rect 13727 6035 13820 6042
rect 14382 6202 14414 6209
rect 14382 6182 14389 6202
rect 14410 6182 14414 6202
rect 14382 6117 14414 6182
rect 14594 6173 14625 6374
rect 14829 6372 14861 6373
rect 14826 6367 14861 6372
rect 14826 6347 14833 6367
rect 14853 6347 14861 6367
rect 14826 6339 14861 6347
rect 14594 6143 14600 6173
rect 14621 6143 14625 6173
rect 14594 6135 14625 6143
rect 14752 6117 14792 6118
rect 14382 6115 14794 6117
rect 14382 6089 14762 6115
rect 14788 6089 14794 6115
rect 14382 6081 14794 6089
rect 14382 6053 14414 6081
rect 14827 6061 14861 6339
rect 14382 6033 14387 6053
rect 14408 6033 14414 6053
rect 14382 6026 14414 6033
rect 14805 6056 14861 6061
rect 14805 6036 14812 6056
rect 14832 6036 14861 6056
rect 14805 6029 14861 6036
rect 14805 6028 14840 6029
rect 11601 5978 11712 5982
rect 13343 5978 14987 5981
rect 10921 5960 14987 5978
rect 10921 5940 11609 5960
rect 11628 5940 11686 5960
rect 11705 5955 14987 5960
rect 11705 5940 14104 5955
rect 10921 5935 14104 5940
rect 14123 5935 14181 5955
rect 14200 5935 14987 5955
rect 10921 5925 14987 5935
rect 10921 5922 11546 5925
rect 11733 5922 14987 5925
rect 9195 5774 9217 5812
rect 9242 5777 9261 5812
rect 9286 5777 9294 5812
rect 9242 5774 9294 5777
rect 9195 5766 9294 5774
rect 9221 5765 9293 5766
rect 8872 5739 8943 5755
rect 8872 5723 8892 5739
rect 8873 5693 8892 5723
rect 8875 5673 8892 5693
rect 8922 5693 8943 5739
rect 9915 5735 9993 5816
rect 10360 5761 10468 5816
rect 8922 5673 8942 5693
rect 8875 5654 8942 5673
rect 9915 5633 9994 5735
rect 9879 5615 10000 5633
rect 9879 5613 9950 5615
rect 9879 5572 9894 5613
rect 9931 5574 9950 5613
rect 9987 5574 10000 5615
rect 9931 5572 10000 5574
rect 9879 5562 10000 5572
rect 7184 5534 7295 5537
rect 6498 5533 8048 5534
rect 10361 5533 10468 5761
rect 10923 5694 11030 5922
rect 13343 5921 14987 5922
rect 14096 5918 14207 5921
rect 11391 5883 11512 5893
rect 11391 5881 11460 5883
rect 11391 5840 11404 5881
rect 11441 5842 11460 5881
rect 11497 5842 11512 5883
rect 11441 5840 11512 5842
rect 11391 5822 11512 5840
rect 14596 5863 14682 5867
rect 14596 5845 14611 5863
rect 14663 5845 14682 5863
rect 14596 5836 14682 5845
rect 11397 5720 11476 5822
rect 12449 5782 12516 5801
rect 12449 5762 12469 5782
rect 10923 5639 11031 5694
rect 11398 5639 11476 5720
rect 12448 5716 12469 5762
rect 12499 5762 12516 5782
rect 12499 5732 12518 5762
rect 12499 5716 12519 5732
rect 12448 5700 12519 5716
rect 12098 5689 12170 5690
rect 12097 5681 12196 5689
rect 12097 5678 12149 5681
rect 12097 5643 12105 5678
rect 12130 5643 12149 5678
rect 12174 5643 12196 5681
rect 6498 5530 9658 5533
rect 9845 5530 10470 5533
rect 6498 5520 10470 5530
rect 6498 5500 7191 5520
rect 7210 5500 7268 5520
rect 7287 5515 10470 5520
rect 7287 5500 9686 5515
rect 6498 5495 9686 5500
rect 9705 5495 9763 5515
rect 9782 5495 10470 5515
rect 6498 5477 10470 5495
rect 6498 5474 8048 5477
rect 9679 5473 9790 5477
rect 6551 5426 6586 5427
rect 6530 5419 6586 5426
rect 6530 5399 6559 5419
rect 6579 5399 6586 5419
rect 6530 5394 6586 5399
rect 6977 5422 7009 5429
rect 6977 5402 6983 5422
rect 7004 5402 7009 5422
rect 6530 5116 6564 5394
rect 6977 5374 7009 5402
rect 8865 5414 8945 5426
rect 9046 5421 9081 5422
rect 6597 5366 7009 5374
rect 6597 5340 6603 5366
rect 6629 5340 7009 5366
rect 7395 5380 7832 5393
rect 7395 5357 7408 5380
rect 7434 5373 7832 5380
rect 7434 5357 7788 5373
rect 7395 5350 7788 5357
rect 7814 5350 7832 5373
rect 7395 5344 7832 5350
rect 8865 5388 8881 5414
rect 8921 5388 8945 5414
rect 8865 5369 8945 5388
rect 6597 5338 7009 5340
rect 6599 5337 6639 5338
rect 6766 5312 6797 5320
rect 6766 5282 6770 5312
rect 6791 5282 6797 5312
rect 6530 5108 6565 5116
rect 6530 5088 6538 5108
rect 6558 5088 6565 5108
rect 6530 5083 6565 5088
rect 6530 5082 6562 5083
rect 6766 5075 6797 5282
rect 6977 5273 7009 5338
rect 8865 5343 8884 5369
rect 8924 5343 8945 5369
rect 8865 5316 8945 5343
rect 8865 5290 8888 5316
rect 8928 5290 8945 5316
rect 8865 5279 8945 5290
rect 9025 5414 9081 5421
rect 9025 5394 9054 5414
rect 9074 5394 9081 5414
rect 9025 5389 9081 5394
rect 9472 5417 9504 5424
rect 9472 5397 9478 5417
rect 9499 5397 9504 5417
rect 6977 5253 6981 5273
rect 7002 5253 7009 5273
rect 6977 5246 7009 5253
rect 7286 5190 7387 5191
rect 7184 5177 7387 5190
rect 7184 5175 7327 5177
rect 7184 5172 7261 5175
rect 7184 5145 7187 5172
rect 7216 5148 7261 5172
rect 7290 5148 7327 5175
rect 7216 5145 7327 5148
rect 7184 5144 7327 5145
rect 7363 5144 7387 5177
rect 7184 5131 7387 5144
rect 6764 5069 6797 5075
rect 6760 5065 6797 5069
rect 6760 5055 6798 5065
rect 6760 5042 6770 5055
rect 6761 5018 6770 5042
rect 6787 5018 6798 5055
rect 6761 4997 6798 5018
rect 8870 4979 8935 5279
rect 9025 5111 9059 5389
rect 9472 5369 9504 5397
rect 9092 5361 9504 5369
rect 9092 5335 9098 5361
rect 9124 5335 9504 5361
rect 9926 5403 9993 5410
rect 9926 5382 9943 5403
rect 9979 5382 9993 5403
rect 9926 5363 9993 5382
rect 9926 5360 9943 5363
rect 9092 5333 9504 5335
rect 9094 5332 9134 5333
rect 9261 5307 9292 5315
rect 9261 5277 9265 5307
rect 9286 5277 9292 5307
rect 9025 5103 9060 5111
rect 9025 5083 9033 5103
rect 9053 5083 9060 5103
rect 9025 5078 9060 5083
rect 9025 5077 9057 5078
rect 9261 5073 9292 5277
rect 9472 5268 9504 5333
rect 9928 5326 9943 5360
rect 9983 5326 9993 5363
rect 9928 5317 9993 5326
rect 9472 5248 9476 5268
rect 9497 5248 9504 5268
rect 9472 5241 9504 5248
rect 9781 5185 9882 5186
rect 9679 5172 9882 5185
rect 9679 5170 9822 5172
rect 9679 5167 9756 5170
rect 9679 5140 9682 5167
rect 9711 5143 9756 5167
rect 9785 5143 9822 5170
rect 9711 5140 9822 5143
rect 9679 5139 9822 5140
rect 9858 5139 9882 5172
rect 9679 5126 9882 5139
rect 9259 5061 9294 5073
rect 9190 5054 9294 5061
rect 9190 5053 9266 5054
rect 9190 5033 9211 5053
rect 9243 5034 9266 5053
rect 9291 5034 9294 5054
rect 9243 5033 9294 5034
rect 9190 5024 9294 5033
rect 9259 5022 9294 5024
rect 8870 4940 8873 4979
rect 8918 4940 8935 4979
rect 9931 4956 9982 5317
rect 9929 4954 9986 4956
rect 8870 4918 8935 4940
rect 9918 4942 9986 4954
rect 9918 4909 9929 4942
rect 9969 4909 9986 4942
rect 9918 4903 9986 4909
rect 9918 4899 9982 4903
rect 8631 4854 8742 4857
rect 10361 4854 10468 5477
rect 6707 4840 10468 4854
rect 6707 4820 8638 4840
rect 8657 4820 8715 4840
rect 8734 4836 10468 4840
rect 8734 4820 9686 4836
rect 6707 4816 9686 4820
rect 9705 4816 9763 4836
rect 9782 4816 10468 4836
rect 6707 4798 10468 4816
rect 6707 4797 8007 4798
rect 9679 4794 9790 4798
rect 7998 4746 8033 4747
rect 7977 4739 8033 4746
rect 7977 4719 8006 4739
rect 8026 4719 8033 4739
rect 7977 4714 8033 4719
rect 8424 4742 8456 4749
rect 9046 4742 9081 4743
rect 8424 4722 8430 4742
rect 8451 4722 8456 4742
rect 9025 4735 9081 4742
rect 8890 4725 8948 4730
rect 7977 4436 8011 4714
rect 8424 4694 8456 4722
rect 8044 4686 8456 4694
rect 8044 4660 8050 4686
rect 8076 4660 8456 4686
rect 8044 4658 8456 4660
rect 8046 4657 8086 4658
rect 8213 4632 8244 4640
rect 8213 4602 8217 4632
rect 8238 4602 8244 4632
rect 7977 4428 8012 4436
rect 7977 4408 7985 4428
rect 8005 4408 8012 4428
rect 7977 4403 8012 4408
rect 7977 4402 8009 4403
rect 8213 4395 8244 4602
rect 8424 4593 8456 4658
rect 8424 4573 8428 4593
rect 8449 4573 8456 4593
rect 8424 4566 8456 4573
rect 8873 4716 8948 4725
rect 8873 4683 8882 4716
rect 8935 4683 8948 4716
rect 8873 4658 8948 4683
rect 8873 4625 8887 4658
rect 8940 4625 8948 4658
rect 8873 4619 8948 4625
rect 9025 4715 9054 4735
rect 9074 4715 9081 4735
rect 9025 4710 9081 4715
rect 9472 4738 9504 4745
rect 9472 4718 9478 4738
rect 9499 4718 9504 4738
rect 8733 4510 8834 4511
rect 8631 4497 8834 4510
rect 8631 4495 8774 4497
rect 8631 4492 8708 4495
rect 8631 4465 8634 4492
rect 8663 4468 8708 4492
rect 8737 4468 8774 4495
rect 8663 4465 8774 4468
rect 8631 4464 8774 4465
rect 8810 4464 8834 4497
rect 8631 4451 8834 4464
rect 7711 4382 7875 4385
rect 8208 4382 8244 4395
rect 6910 4364 8249 4382
rect 6910 4326 6920 4364
rect 6945 4349 8249 4364
rect 6945 4326 6955 4349
rect 7711 4342 7875 4349
rect 6910 4318 6955 4326
rect 6924 4317 6955 4318
rect 8873 4303 8943 4619
rect 9025 4432 9059 4710
rect 9472 4690 9504 4718
rect 9092 4682 9504 4690
rect 9092 4656 9098 4682
rect 9124 4656 9504 4682
rect 9092 4654 9504 4656
rect 9094 4653 9134 4654
rect 9261 4628 9292 4636
rect 9261 4598 9265 4628
rect 9286 4598 9292 4628
rect 9025 4424 9060 4432
rect 9025 4404 9033 4424
rect 9053 4404 9060 4424
rect 9025 4399 9060 4404
rect 9261 4399 9292 4598
rect 9472 4589 9504 4654
rect 9472 4569 9476 4589
rect 9497 4569 9504 4589
rect 9472 4562 9504 4569
rect 9917 4715 9989 4733
rect 9917 4673 9930 4715
rect 9979 4673 9989 4715
rect 9917 4652 9989 4673
rect 9917 4610 9931 4652
rect 9980 4610 9989 4652
rect 9781 4506 9882 4507
rect 9679 4493 9882 4506
rect 9679 4491 9822 4493
rect 9679 4488 9756 4491
rect 9679 4461 9682 4488
rect 9711 4464 9756 4488
rect 9785 4464 9822 4491
rect 9711 4461 9822 4464
rect 9679 4460 9822 4461
rect 9858 4460 9882 4493
rect 9679 4447 9882 4460
rect 9025 4398 9057 4399
rect 9259 4396 9292 4399
rect 9225 4377 9293 4396
rect 9195 4365 9294 4377
rect 9195 4327 9217 4365
rect 9242 4330 9261 4365
rect 9286 4330 9294 4365
rect 9242 4327 9294 4330
rect 9195 4319 9294 4327
rect 9221 4318 9293 4319
rect 8873 4284 8952 4303
rect 8876 4264 8952 4284
rect 8869 4240 8952 4264
rect 9917 4299 9989 4610
rect 9917 4256 9993 4299
rect 8869 4174 8881 4240
rect 8935 4174 8952 4240
rect 8869 4154 8952 4174
rect 8869 4117 8886 4154
rect 8930 4140 8952 4154
rect 9918 4205 9993 4256
rect 10361 4205 10468 4798
rect 10923 5210 11030 5639
rect 11402 5398 11474 5639
rect 12097 5631 12196 5643
rect 12098 5612 12166 5631
rect 12099 5609 12132 5612
rect 12334 5609 12366 5610
rect 11509 5548 11712 5561
rect 11509 5515 11533 5548
rect 11569 5547 11712 5548
rect 11569 5544 11680 5547
rect 11569 5517 11606 5544
rect 11635 5520 11680 5544
rect 11709 5520 11712 5547
rect 11635 5517 11712 5520
rect 11569 5515 11712 5517
rect 11509 5502 11712 5515
rect 11509 5501 11610 5502
rect 11402 5356 11411 5398
rect 11460 5356 11474 5398
rect 11402 5335 11474 5356
rect 11402 5293 11412 5335
rect 11461 5293 11474 5335
rect 11402 5275 11474 5293
rect 11887 5439 11919 5446
rect 11887 5419 11894 5439
rect 11915 5419 11919 5439
rect 11887 5354 11919 5419
rect 12099 5410 12130 5609
rect 12331 5604 12366 5609
rect 12331 5584 12338 5604
rect 12358 5584 12366 5604
rect 12331 5576 12366 5584
rect 12099 5380 12105 5410
rect 12126 5380 12130 5410
rect 12099 5372 12130 5380
rect 12257 5354 12297 5355
rect 11887 5352 12299 5354
rect 11887 5326 12267 5352
rect 12293 5326 12299 5352
rect 11887 5318 12299 5326
rect 11887 5290 11919 5318
rect 12332 5298 12366 5576
rect 12448 5389 12518 5700
rect 14373 5690 14445 5691
rect 14372 5687 14461 5690
rect 13144 5685 14461 5687
rect 13141 5682 14461 5685
rect 13141 5679 14424 5682
rect 13141 5644 14380 5679
rect 14405 5644 14424 5679
rect 14449 5644 14461 5682
rect 13141 5634 14461 5644
rect 14637 5683 14673 5836
rect 14637 5660 14643 5683
rect 14667 5660 14673 5683
rect 14637 5639 14673 5660
rect 13141 5632 14426 5634
rect 13141 5622 13238 5632
rect 13147 5613 13183 5622
rect 14637 5616 14643 5639
rect 14667 5616 14673 5639
rect 12557 5544 12760 5557
rect 12557 5511 12581 5544
rect 12617 5543 12760 5544
rect 12617 5540 12728 5543
rect 12617 5513 12654 5540
rect 12683 5516 12728 5540
rect 12757 5516 12760 5543
rect 12683 5513 12760 5516
rect 12617 5511 12760 5513
rect 12557 5498 12760 5511
rect 12557 5497 12658 5498
rect 11887 5270 11892 5290
rect 11913 5270 11919 5290
rect 11887 5263 11919 5270
rect 12310 5293 12366 5298
rect 12310 5273 12317 5293
rect 12337 5273 12366 5293
rect 12443 5383 12518 5389
rect 12443 5350 12451 5383
rect 12504 5350 12518 5383
rect 12443 5325 12518 5350
rect 12443 5292 12456 5325
rect 12509 5292 12518 5325
rect 12443 5283 12518 5292
rect 12935 5435 12967 5442
rect 12935 5415 12942 5435
rect 12963 5415 12967 5435
rect 12935 5350 12967 5415
rect 13147 5406 13178 5613
rect 13382 5605 13414 5606
rect 14637 5605 14673 5616
rect 13379 5600 13414 5605
rect 13379 5580 13386 5600
rect 13406 5580 13414 5600
rect 13379 5572 13414 5580
rect 13147 5376 13153 5406
rect 13174 5376 13178 5406
rect 13147 5368 13178 5376
rect 13305 5350 13345 5351
rect 12935 5348 13347 5350
rect 12935 5322 13315 5348
rect 13341 5322 13347 5348
rect 12935 5314 13347 5322
rect 12935 5286 12967 5314
rect 13380 5294 13414 5572
rect 12443 5278 12501 5283
rect 12310 5266 12366 5273
rect 12935 5266 12940 5286
rect 12961 5266 12967 5286
rect 12310 5265 12345 5266
rect 12935 5259 12967 5266
rect 13358 5289 13414 5294
rect 13358 5269 13365 5289
rect 13385 5269 13414 5289
rect 13358 5262 13414 5269
rect 13358 5261 13393 5262
rect 11601 5210 11712 5214
rect 13476 5210 14635 5211
rect 10923 5192 14635 5210
rect 10923 5172 11609 5192
rect 11628 5172 11686 5192
rect 11705 5188 14635 5192
rect 11705 5172 12657 5188
rect 10923 5168 12657 5172
rect 12676 5168 12734 5188
rect 12753 5168 14635 5188
rect 10923 5154 14635 5168
rect 10923 4531 11030 5154
rect 12649 5151 12760 5154
rect 11409 5105 11473 5109
rect 11405 5099 11473 5105
rect 11405 5066 11422 5099
rect 11462 5066 11473 5099
rect 11405 5054 11473 5066
rect 12456 5068 12521 5090
rect 11405 5052 11462 5054
rect 11409 4691 11460 5052
rect 12456 5029 12473 5068
rect 12518 5029 12521 5068
rect 15542 5066 15594 7372
rect 15703 7349 15738 7415
rect 15703 6033 15737 7349
rect 16041 7202 16146 12302
rect 17105 12289 21178 12303
rect 17105 12269 19348 12289
rect 19367 12269 19425 12289
rect 19444 12285 21178 12289
rect 19444 12269 20396 12285
rect 17105 12265 20396 12269
rect 20415 12265 20473 12285
rect 20492 12265 21178 12285
rect 17105 12247 21178 12265
rect 17105 12246 18625 12247
rect 20389 12243 20500 12247
rect 18708 12195 18743 12196
rect 18687 12188 18743 12195
rect 18687 12168 18716 12188
rect 18736 12168 18743 12188
rect 18687 12163 18743 12168
rect 19134 12191 19166 12198
rect 19756 12191 19791 12192
rect 19134 12171 19140 12191
rect 19161 12171 19166 12191
rect 19735 12184 19791 12191
rect 19600 12174 19658 12179
rect 18687 11885 18721 12163
rect 19134 12143 19166 12171
rect 18754 12135 19166 12143
rect 18754 12109 18760 12135
rect 18786 12109 19166 12135
rect 18754 12107 19166 12109
rect 18756 12106 18796 12107
rect 18923 12081 18954 12089
rect 18923 12051 18927 12081
rect 18948 12051 18954 12081
rect 18687 11877 18722 11885
rect 18687 11857 18695 11877
rect 18715 11857 18722 11877
rect 18687 11852 18722 11857
rect 18687 11851 18719 11852
rect 18923 11851 18954 12051
rect 19134 12042 19166 12107
rect 19134 12022 19138 12042
rect 19159 12022 19166 12042
rect 19134 12015 19166 12022
rect 19583 12165 19658 12174
rect 19583 12132 19592 12165
rect 19645 12132 19658 12165
rect 19583 12107 19658 12132
rect 19583 12074 19597 12107
rect 19650 12074 19658 12107
rect 19583 12068 19658 12074
rect 19735 12164 19764 12184
rect 19784 12164 19791 12184
rect 19735 12159 19791 12164
rect 20182 12187 20214 12194
rect 20182 12167 20188 12187
rect 20209 12167 20214 12187
rect 19443 11959 19544 11960
rect 19341 11946 19544 11959
rect 19341 11944 19484 11946
rect 19341 11941 19418 11944
rect 19341 11914 19344 11941
rect 19373 11917 19418 11941
rect 19447 11917 19484 11944
rect 19373 11914 19484 11917
rect 19341 11913 19484 11914
rect 19520 11913 19544 11946
rect 19341 11900 19544 11913
rect 18920 11844 18959 11851
rect 18918 11827 18959 11844
rect 18920 11802 18959 11827
rect 17614 11794 18959 11802
rect 17614 11766 17629 11794
rect 17657 11768 18959 11794
rect 17657 11766 18956 11768
rect 17614 11761 18956 11766
rect 19583 11757 19653 12068
rect 19735 11881 19769 12159
rect 20182 12139 20214 12167
rect 19802 12131 20214 12139
rect 19802 12105 19808 12131
rect 19834 12105 20214 12131
rect 19802 12103 20214 12105
rect 19804 12102 19844 12103
rect 19971 12077 20002 12085
rect 19971 12047 19975 12077
rect 19996 12047 20002 12077
rect 19735 11873 19770 11881
rect 19735 11853 19743 11873
rect 19763 11853 19770 11873
rect 19735 11848 19770 11853
rect 19971 11848 20002 12047
rect 20182 12038 20214 12103
rect 20182 12018 20186 12038
rect 20207 12018 20214 12038
rect 20182 12011 20214 12018
rect 20627 12164 20699 12182
rect 20627 12122 20640 12164
rect 20689 12122 20699 12164
rect 20627 12101 20699 12122
rect 20627 12059 20641 12101
rect 20690 12059 20699 12101
rect 20491 11955 20592 11956
rect 20389 11942 20592 11955
rect 20389 11940 20532 11942
rect 20389 11937 20466 11940
rect 20389 11910 20392 11937
rect 20421 11913 20466 11937
rect 20495 11913 20532 11940
rect 20421 11910 20532 11913
rect 20389 11909 20532 11910
rect 20568 11909 20592 11942
rect 20389 11896 20592 11909
rect 19735 11847 19767 11848
rect 19969 11845 20002 11848
rect 19935 11826 20003 11845
rect 19905 11814 20004 11826
rect 20627 11818 20699 12059
rect 21071 11818 21178 12247
rect 19905 11776 19927 11814
rect 19952 11779 19971 11814
rect 19996 11779 20004 11814
rect 19952 11776 20004 11779
rect 19905 11768 20004 11776
rect 19931 11767 20003 11768
rect 19582 11741 19653 11757
rect 19582 11725 19602 11741
rect 19583 11695 19602 11725
rect 19585 11675 19602 11695
rect 19632 11695 19653 11741
rect 20625 11737 20703 11818
rect 21070 11763 21178 11818
rect 19632 11675 19652 11695
rect 19585 11656 19652 11675
rect 20625 11635 20704 11737
rect 20589 11617 20710 11635
rect 20589 11615 20660 11617
rect 20589 11574 20604 11615
rect 20641 11576 20660 11615
rect 20697 11576 20710 11617
rect 20641 11574 20710 11576
rect 20589 11564 20710 11574
rect 17894 11536 18005 11539
rect 17105 11535 18758 11536
rect 21071 11535 21178 11763
rect 17105 11532 20368 11535
rect 20555 11532 21180 11535
rect 17105 11522 21180 11532
rect 17105 11502 17901 11522
rect 17920 11502 17978 11522
rect 17997 11517 21180 11522
rect 17997 11502 20396 11517
rect 17105 11497 20396 11502
rect 20415 11497 20473 11517
rect 20492 11497 21180 11517
rect 17105 11479 21180 11497
rect 17105 11476 18758 11479
rect 20389 11475 20500 11479
rect 17261 11428 17296 11429
rect 17240 11421 17296 11428
rect 17240 11401 17269 11421
rect 17289 11401 17296 11421
rect 17240 11396 17296 11401
rect 17687 11424 17719 11431
rect 17687 11404 17693 11424
rect 17714 11404 17719 11424
rect 17240 11118 17274 11396
rect 17687 11376 17719 11404
rect 19575 11416 19655 11428
rect 19756 11423 19791 11424
rect 17307 11368 17719 11376
rect 17307 11342 17313 11368
rect 17339 11342 17719 11368
rect 18105 11382 18542 11395
rect 18105 11359 18118 11382
rect 18144 11375 18542 11382
rect 18144 11359 18498 11375
rect 18105 11352 18498 11359
rect 18524 11352 18542 11375
rect 18105 11346 18542 11352
rect 19575 11390 19591 11416
rect 19631 11390 19655 11416
rect 19575 11371 19655 11390
rect 17307 11340 17719 11342
rect 17309 11339 17349 11340
rect 17476 11314 17507 11322
rect 17476 11284 17480 11314
rect 17501 11284 17507 11314
rect 17240 11110 17275 11118
rect 17240 11090 17248 11110
rect 17268 11090 17275 11110
rect 17240 11085 17275 11090
rect 17240 11084 17272 11085
rect 17476 11077 17507 11284
rect 17687 11275 17719 11340
rect 19575 11345 19594 11371
rect 19634 11345 19655 11371
rect 19575 11318 19655 11345
rect 19575 11292 19598 11318
rect 19638 11292 19655 11318
rect 19575 11281 19655 11292
rect 19735 11416 19791 11423
rect 19735 11396 19764 11416
rect 19784 11396 19791 11416
rect 19735 11391 19791 11396
rect 20182 11419 20214 11426
rect 20182 11399 20188 11419
rect 20209 11399 20214 11419
rect 17687 11255 17691 11275
rect 17712 11255 17719 11275
rect 17687 11248 17719 11255
rect 17996 11192 18097 11193
rect 17894 11179 18097 11192
rect 17894 11177 18037 11179
rect 17894 11174 17971 11177
rect 17894 11147 17897 11174
rect 17926 11150 17971 11174
rect 18000 11150 18037 11177
rect 17926 11147 18037 11150
rect 17894 11146 18037 11147
rect 18073 11146 18097 11179
rect 17894 11133 18097 11146
rect 17474 11071 17507 11077
rect 17470 11067 17507 11071
rect 17470 11057 17508 11067
rect 17470 11044 17480 11057
rect 17471 11020 17480 11044
rect 17497 11020 17508 11057
rect 17471 10999 17508 11020
rect 19580 10981 19645 11281
rect 19735 11113 19769 11391
rect 20182 11371 20214 11399
rect 19802 11363 20214 11371
rect 19802 11337 19808 11363
rect 19834 11337 20214 11363
rect 20636 11405 20703 11412
rect 20636 11384 20653 11405
rect 20689 11384 20703 11405
rect 20636 11365 20703 11384
rect 20636 11362 20653 11365
rect 19802 11335 20214 11337
rect 19804 11334 19844 11335
rect 19971 11309 20002 11317
rect 19971 11279 19975 11309
rect 19996 11279 20002 11309
rect 19735 11105 19770 11113
rect 19735 11085 19743 11105
rect 19763 11085 19770 11105
rect 19735 11080 19770 11085
rect 19735 11079 19767 11080
rect 19971 11075 20002 11279
rect 20182 11270 20214 11335
rect 20638 11328 20653 11362
rect 20693 11328 20703 11365
rect 20638 11319 20703 11328
rect 20182 11250 20186 11270
rect 20207 11250 20214 11270
rect 20182 11243 20214 11250
rect 20491 11187 20592 11188
rect 20389 11174 20592 11187
rect 20389 11172 20532 11174
rect 20389 11169 20466 11172
rect 20389 11142 20392 11169
rect 20421 11145 20466 11169
rect 20495 11145 20532 11172
rect 20421 11142 20532 11145
rect 20389 11141 20532 11142
rect 20568 11141 20592 11174
rect 20389 11128 20592 11141
rect 19969 11063 20004 11075
rect 19900 11056 20004 11063
rect 19900 11055 19976 11056
rect 19900 11035 19921 11055
rect 19953 11036 19976 11055
rect 20001 11036 20004 11056
rect 19953 11035 20004 11036
rect 19900 11026 20004 11035
rect 19969 11024 20004 11026
rect 19580 10942 19583 10981
rect 19628 10942 19645 10981
rect 20641 10958 20692 11319
rect 20639 10956 20696 10958
rect 19580 10920 19645 10942
rect 20628 10944 20696 10956
rect 20628 10911 20639 10944
rect 20679 10911 20696 10944
rect 20628 10905 20696 10911
rect 20628 10901 20692 10905
rect 19341 10856 19452 10859
rect 21071 10856 21178 11479
rect 16728 10842 21178 10856
rect 16728 10822 19348 10842
rect 19367 10822 19425 10842
rect 19444 10838 21178 10842
rect 19444 10822 20396 10838
rect 16728 10818 20396 10822
rect 20415 10818 20473 10838
rect 20492 10818 21178 10838
rect 16728 10804 21178 10818
rect 17147 10800 21178 10804
rect 17147 10799 18717 10800
rect 20389 10796 20500 10800
rect 18708 10748 18743 10749
rect 18687 10741 18743 10748
rect 18687 10721 18716 10741
rect 18736 10721 18743 10741
rect 18687 10716 18743 10721
rect 19134 10744 19166 10751
rect 19756 10744 19791 10745
rect 19134 10724 19140 10744
rect 19161 10724 19166 10744
rect 19735 10737 19791 10744
rect 19600 10727 19658 10732
rect 18687 10438 18721 10716
rect 19134 10696 19166 10724
rect 18754 10688 19166 10696
rect 18754 10662 18760 10688
rect 18786 10662 19166 10688
rect 18754 10660 19166 10662
rect 18756 10659 18796 10660
rect 18923 10634 18954 10642
rect 18923 10604 18927 10634
rect 18948 10604 18954 10634
rect 18687 10430 18722 10438
rect 18687 10410 18695 10430
rect 18715 10410 18722 10430
rect 18687 10405 18722 10410
rect 18687 10404 18719 10405
rect 18923 10397 18954 10604
rect 19134 10595 19166 10660
rect 19134 10575 19138 10595
rect 19159 10575 19166 10595
rect 19134 10568 19166 10575
rect 19583 10718 19658 10727
rect 19583 10685 19592 10718
rect 19645 10685 19658 10718
rect 19583 10660 19658 10685
rect 19583 10627 19597 10660
rect 19650 10627 19658 10660
rect 19583 10621 19658 10627
rect 19735 10717 19764 10737
rect 19784 10717 19791 10737
rect 19735 10712 19791 10717
rect 20182 10740 20214 10747
rect 20182 10720 20188 10740
rect 20209 10720 20214 10740
rect 19443 10512 19544 10513
rect 19341 10499 19544 10512
rect 19341 10497 19484 10499
rect 19341 10494 19418 10497
rect 19341 10467 19344 10494
rect 19373 10470 19418 10494
rect 19447 10470 19484 10497
rect 19373 10467 19484 10470
rect 19341 10466 19484 10467
rect 19520 10466 19544 10499
rect 19341 10453 19544 10466
rect 18421 10384 18585 10387
rect 18918 10384 18954 10397
rect 17620 10366 18959 10384
rect 17620 10328 17630 10366
rect 17655 10351 18959 10366
rect 17655 10328 17665 10351
rect 18421 10344 18585 10351
rect 17620 10320 17665 10328
rect 17634 10319 17665 10320
rect 19583 10305 19653 10621
rect 19735 10434 19769 10712
rect 20182 10692 20214 10720
rect 19802 10684 20214 10692
rect 19802 10658 19808 10684
rect 19834 10658 20214 10684
rect 19802 10656 20214 10658
rect 19804 10655 19844 10656
rect 19971 10630 20002 10638
rect 19971 10600 19975 10630
rect 19996 10600 20002 10630
rect 19735 10426 19770 10434
rect 19735 10406 19743 10426
rect 19763 10406 19770 10426
rect 19735 10401 19770 10406
rect 19971 10401 20002 10600
rect 20182 10591 20214 10656
rect 20182 10571 20186 10591
rect 20207 10571 20214 10591
rect 20182 10564 20214 10571
rect 20627 10717 20699 10735
rect 20627 10675 20640 10717
rect 20689 10675 20699 10717
rect 20627 10654 20699 10675
rect 20627 10612 20641 10654
rect 20690 10612 20699 10654
rect 20491 10508 20592 10509
rect 20389 10495 20592 10508
rect 20389 10493 20532 10495
rect 20389 10490 20466 10493
rect 20389 10463 20392 10490
rect 20421 10466 20466 10490
rect 20495 10466 20532 10493
rect 20421 10463 20532 10466
rect 20389 10462 20532 10463
rect 20568 10462 20592 10495
rect 20389 10449 20592 10462
rect 19735 10400 19767 10401
rect 19969 10398 20002 10401
rect 19935 10379 20003 10398
rect 19905 10367 20004 10379
rect 19905 10329 19927 10367
rect 19952 10332 19971 10367
rect 19996 10332 20004 10367
rect 19952 10329 20004 10332
rect 19905 10321 20004 10329
rect 19931 10320 20003 10321
rect 19583 10286 19662 10305
rect 19586 10266 19662 10286
rect 19579 10242 19662 10266
rect 20627 10301 20699 10612
rect 20627 10258 20703 10301
rect 19579 10176 19591 10242
rect 19645 10176 19662 10242
rect 19579 10156 19662 10176
rect 19579 10119 19596 10156
rect 19640 10142 19662 10156
rect 20628 10207 20703 10258
rect 21071 10207 21178 10800
rect 19640 10119 19655 10142
rect 19579 10103 19655 10119
rect 20628 10115 20705 10207
rect 21071 10203 21179 10207
rect 20590 10097 20711 10115
rect 20590 10095 20661 10097
rect 20590 10054 20605 10095
rect 20642 10056 20661 10095
rect 20698 10056 20711 10097
rect 20642 10054 20711 10056
rect 20590 10044 20711 10054
rect 17115 10015 18584 10017
rect 21072 10015 21179 10203
rect 17115 10000 21181 10015
rect 17115 9980 17859 10000
rect 17878 9980 17936 10000
rect 17955 9997 21181 10000
rect 17955 9980 20397 9997
rect 17115 9977 20397 9980
rect 20416 9977 20474 9997
rect 20493 9977 21181 9997
rect 17115 9959 21181 9977
rect 17852 9958 17963 9959
rect 18539 9958 18746 9959
rect 20390 9955 20501 9959
rect 17219 9906 17254 9907
rect 17198 9899 17254 9906
rect 17198 9879 17227 9899
rect 17247 9879 17254 9899
rect 17198 9874 17254 9879
rect 17645 9902 17677 9909
rect 17645 9882 17651 9902
rect 17672 9882 17677 9902
rect 17198 9596 17232 9874
rect 17645 9854 17677 9882
rect 17265 9846 17677 9854
rect 17265 9820 17271 9846
rect 17297 9820 17677 9846
rect 17265 9818 17677 9820
rect 17267 9817 17307 9818
rect 17434 9792 17465 9800
rect 17434 9762 17438 9792
rect 17459 9762 17465 9792
rect 17198 9588 17233 9596
rect 17198 9568 17206 9588
rect 17226 9568 17233 9588
rect 17198 9563 17233 9568
rect 17434 9566 17465 9762
rect 17645 9753 17677 9818
rect 19576 9896 19656 9908
rect 19757 9903 19792 9904
rect 19576 9870 19592 9896
rect 19632 9870 19656 9896
rect 19576 9851 19656 9870
rect 19576 9825 19595 9851
rect 19635 9825 19656 9851
rect 19576 9798 19656 9825
rect 19576 9772 19599 9798
rect 19639 9772 19656 9798
rect 19576 9761 19656 9772
rect 19736 9896 19792 9903
rect 19736 9876 19765 9896
rect 19785 9876 19792 9896
rect 19736 9871 19792 9876
rect 20183 9899 20215 9906
rect 20183 9879 20189 9899
rect 20210 9879 20215 9899
rect 17645 9733 17649 9753
rect 17670 9733 17677 9753
rect 17645 9726 17677 9733
rect 17954 9670 18055 9671
rect 17852 9657 18055 9670
rect 17852 9655 17995 9657
rect 17852 9652 17929 9655
rect 17852 9625 17855 9652
rect 17884 9628 17929 9652
rect 17958 9628 17995 9655
rect 17884 9625 17995 9628
rect 17852 9624 17995 9625
rect 18031 9624 18055 9657
rect 17852 9611 18055 9624
rect 17198 9562 17230 9563
rect 17434 9477 17468 9566
rect 17055 9473 17468 9477
rect 16041 7148 16058 7202
rect 16121 7148 16146 7202
rect 16041 7127 16146 7148
rect 16508 9428 17468 9473
rect 19581 9461 19646 9761
rect 19736 9593 19770 9871
rect 20183 9851 20215 9879
rect 19803 9843 20215 9851
rect 19803 9817 19809 9843
rect 19835 9817 20215 9843
rect 20637 9885 20704 9892
rect 20637 9864 20654 9885
rect 20690 9864 20704 9885
rect 20637 9845 20704 9864
rect 20637 9842 20654 9845
rect 19803 9815 20215 9817
rect 19805 9814 19845 9815
rect 19972 9789 20003 9797
rect 19972 9759 19976 9789
rect 19997 9759 20003 9789
rect 19736 9585 19771 9593
rect 19736 9565 19744 9585
rect 19764 9565 19771 9585
rect 19736 9560 19771 9565
rect 19736 9559 19768 9560
rect 19972 9555 20003 9759
rect 20183 9750 20215 9815
rect 20639 9808 20654 9842
rect 20694 9808 20704 9845
rect 20639 9799 20704 9808
rect 20183 9730 20187 9750
rect 20208 9730 20215 9750
rect 20183 9723 20215 9730
rect 20492 9667 20593 9668
rect 20390 9654 20593 9667
rect 20390 9652 20533 9654
rect 20390 9649 20467 9652
rect 20390 9622 20393 9649
rect 20422 9625 20467 9649
rect 20496 9625 20533 9652
rect 20422 9622 20533 9625
rect 20390 9621 20533 9622
rect 20569 9621 20593 9654
rect 20390 9608 20593 9621
rect 19970 9543 20005 9555
rect 19901 9536 20005 9543
rect 19901 9535 19977 9536
rect 19901 9515 19922 9535
rect 19954 9516 19977 9535
rect 20002 9516 20005 9536
rect 19954 9515 20005 9516
rect 19901 9506 20005 9515
rect 19970 9504 20005 9506
rect 16508 9424 17105 9428
rect 16508 7118 16560 9424
rect 19581 9422 19584 9461
rect 19629 9422 19646 9461
rect 20642 9438 20693 9799
rect 20640 9436 20697 9438
rect 19581 9400 19646 9422
rect 20629 9424 20697 9436
rect 20629 9391 20640 9424
rect 20680 9391 20697 9424
rect 20629 9385 20697 9391
rect 20629 9381 20693 9385
rect 19342 9336 19453 9339
rect 21072 9336 21179 9959
rect 17467 9322 21179 9336
rect 17467 9302 19349 9322
rect 19368 9302 19426 9322
rect 19445 9318 21179 9322
rect 19445 9302 20397 9318
rect 17467 9298 20397 9302
rect 20416 9298 20474 9318
rect 20493 9298 21179 9318
rect 17467 9280 21179 9298
rect 17467 9279 18626 9280
rect 20390 9276 20501 9280
rect 18709 9228 18744 9229
rect 18688 9221 18744 9228
rect 18688 9201 18717 9221
rect 18737 9201 18744 9221
rect 18688 9196 18744 9201
rect 19135 9224 19167 9231
rect 19757 9224 19792 9225
rect 19135 9204 19141 9224
rect 19162 9204 19167 9224
rect 19736 9217 19792 9224
rect 19601 9207 19659 9212
rect 18688 8918 18722 9196
rect 19135 9176 19167 9204
rect 18755 9168 19167 9176
rect 18755 9142 18761 9168
rect 18787 9142 19167 9168
rect 18755 9140 19167 9142
rect 18757 9139 18797 9140
rect 18924 9114 18955 9122
rect 18924 9084 18928 9114
rect 18949 9084 18955 9114
rect 18688 8910 18723 8918
rect 18688 8890 18696 8910
rect 18716 8890 18723 8910
rect 18688 8885 18723 8890
rect 17429 8874 17465 8885
rect 18688 8884 18720 8885
rect 18924 8877 18955 9084
rect 19135 9075 19167 9140
rect 19135 9055 19139 9075
rect 19160 9055 19167 9075
rect 19135 9048 19167 9055
rect 19584 9198 19659 9207
rect 19584 9165 19593 9198
rect 19646 9165 19659 9198
rect 19584 9140 19659 9165
rect 19584 9107 19598 9140
rect 19651 9107 19659 9140
rect 19584 9101 19659 9107
rect 19736 9197 19765 9217
rect 19785 9197 19792 9217
rect 19736 9192 19792 9197
rect 20183 9220 20215 9227
rect 20183 9200 20189 9220
rect 20210 9200 20215 9220
rect 19444 8992 19545 8993
rect 19342 8979 19545 8992
rect 19342 8977 19485 8979
rect 19342 8974 19419 8977
rect 19342 8947 19345 8974
rect 19374 8950 19419 8974
rect 19448 8950 19485 8977
rect 19374 8947 19485 8950
rect 19342 8946 19485 8947
rect 19521 8946 19545 8979
rect 19342 8933 19545 8946
rect 17429 8851 17435 8874
rect 17459 8851 17465 8874
rect 18919 8868 18955 8877
rect 18864 8858 18961 8868
rect 17676 8856 18961 8858
rect 17429 8830 17465 8851
rect 17429 8807 17435 8830
rect 17459 8807 17465 8830
rect 17429 8654 17465 8807
rect 17641 8846 18961 8856
rect 17641 8808 17653 8846
rect 17678 8811 17697 8846
rect 17722 8811 18961 8846
rect 17678 8808 18961 8811
rect 17641 8805 18961 8808
rect 17641 8803 18958 8805
rect 17641 8800 17730 8803
rect 17657 8799 17729 8800
rect 19584 8790 19654 9101
rect 19736 8914 19770 9192
rect 20183 9172 20215 9200
rect 19803 9164 20215 9172
rect 19803 9138 19809 9164
rect 19835 9138 20215 9164
rect 19803 9136 20215 9138
rect 19805 9135 19845 9136
rect 19972 9110 20003 9118
rect 19972 9080 19976 9110
rect 19997 9080 20003 9110
rect 19736 8906 19771 8914
rect 19736 8886 19744 8906
rect 19764 8886 19771 8906
rect 19736 8881 19771 8886
rect 19972 8881 20003 9080
rect 20183 9071 20215 9136
rect 20183 9051 20187 9071
rect 20208 9051 20215 9071
rect 20183 9044 20215 9051
rect 20628 9197 20700 9215
rect 20628 9155 20641 9197
rect 20690 9155 20700 9197
rect 20628 9134 20700 9155
rect 20628 9092 20642 9134
rect 20691 9092 20700 9134
rect 20492 8988 20593 8989
rect 20390 8975 20593 8988
rect 20390 8973 20533 8975
rect 20390 8970 20467 8973
rect 20390 8943 20393 8970
rect 20422 8946 20467 8970
rect 20496 8946 20533 8973
rect 20422 8943 20533 8946
rect 20390 8942 20533 8943
rect 20569 8942 20593 8975
rect 20390 8929 20593 8942
rect 19736 8880 19768 8881
rect 19970 8878 20003 8881
rect 19936 8859 20004 8878
rect 19906 8847 20005 8859
rect 20628 8851 20700 9092
rect 21072 8851 21179 9280
rect 19906 8809 19928 8847
rect 19953 8812 19972 8847
rect 19997 8812 20005 8847
rect 19953 8809 20005 8812
rect 19906 8801 20005 8809
rect 19932 8800 20004 8801
rect 19583 8774 19654 8790
rect 19583 8758 19603 8774
rect 19584 8728 19603 8758
rect 19586 8708 19603 8728
rect 19633 8728 19654 8774
rect 20626 8770 20704 8851
rect 21071 8796 21179 8851
rect 19633 8708 19653 8728
rect 19586 8689 19653 8708
rect 20626 8668 20705 8770
rect 17420 8645 17506 8654
rect 17420 8627 17439 8645
rect 17491 8627 17506 8645
rect 17420 8623 17506 8627
rect 20590 8650 20711 8668
rect 20590 8648 20661 8650
rect 20590 8607 20605 8648
rect 20642 8609 20661 8648
rect 20698 8609 20711 8650
rect 20642 8607 20711 8609
rect 20590 8597 20711 8607
rect 17895 8569 18006 8572
rect 17115 8568 18759 8569
rect 21072 8568 21179 8796
rect 17115 8565 20369 8568
rect 20556 8565 21181 8568
rect 17115 8555 21181 8565
rect 17115 8535 17902 8555
rect 17921 8535 17979 8555
rect 17998 8550 21181 8555
rect 17998 8535 20397 8550
rect 17115 8530 20397 8535
rect 20416 8530 20474 8550
rect 20493 8530 21181 8550
rect 17115 8512 21181 8530
rect 17115 8509 18759 8512
rect 20390 8508 20501 8512
rect 17262 8461 17297 8462
rect 17241 8454 17297 8461
rect 17241 8434 17270 8454
rect 17290 8434 17297 8454
rect 17241 8429 17297 8434
rect 17688 8457 17720 8464
rect 17688 8437 17694 8457
rect 17715 8437 17720 8457
rect 17241 8151 17275 8429
rect 17688 8409 17720 8437
rect 17308 8401 17720 8409
rect 17308 8375 17314 8401
rect 17340 8375 17720 8401
rect 17308 8373 17720 8375
rect 17310 8372 17350 8373
rect 17477 8347 17508 8355
rect 17477 8317 17481 8347
rect 17502 8317 17508 8347
rect 17241 8143 17276 8151
rect 17241 8123 17249 8143
rect 17269 8123 17276 8143
rect 17241 8118 17276 8123
rect 17241 8117 17273 8118
rect 17477 8116 17508 8317
rect 17688 8308 17720 8373
rect 17688 8288 17692 8308
rect 17713 8288 17720 8308
rect 17688 8281 17720 8288
rect 18282 8448 18375 8455
rect 18282 8407 18306 8448
rect 18360 8407 18375 8448
rect 17997 8225 18098 8226
rect 17895 8212 18098 8225
rect 17895 8210 18038 8212
rect 17895 8207 17972 8210
rect 17895 8180 17898 8207
rect 17927 8183 17972 8207
rect 18001 8183 18038 8210
rect 17927 8180 18038 8183
rect 17895 8179 18038 8180
rect 18074 8179 18098 8212
rect 17895 8166 18098 8179
rect 18282 8034 18375 8407
rect 19576 8449 19656 8461
rect 19757 8456 19792 8457
rect 19576 8423 19592 8449
rect 19632 8423 19656 8449
rect 19576 8404 19656 8423
rect 19576 8378 19595 8404
rect 19635 8378 19656 8404
rect 19576 8351 19656 8378
rect 19576 8325 19599 8351
rect 19639 8325 19656 8351
rect 19576 8314 19656 8325
rect 19736 8449 19792 8456
rect 19736 8429 19765 8449
rect 19785 8429 19792 8449
rect 19736 8424 19792 8429
rect 20183 8452 20215 8459
rect 20183 8432 20189 8452
rect 20210 8432 20215 8452
rect 18282 7990 18300 8034
rect 18360 7990 18375 8034
rect 18282 7975 18375 7990
rect 19581 8014 19646 8314
rect 19736 8146 19770 8424
rect 20183 8404 20215 8432
rect 19803 8396 20215 8404
rect 19803 8370 19809 8396
rect 19835 8370 20215 8396
rect 20637 8438 20704 8445
rect 20637 8417 20654 8438
rect 20690 8417 20704 8438
rect 20637 8398 20704 8417
rect 20637 8395 20654 8398
rect 19803 8368 20215 8370
rect 19805 8367 19845 8368
rect 19972 8342 20003 8350
rect 19972 8312 19976 8342
rect 19997 8312 20003 8342
rect 19736 8138 19771 8146
rect 19736 8118 19744 8138
rect 19764 8118 19771 8138
rect 19736 8113 19771 8118
rect 19736 8112 19768 8113
rect 19972 8108 20003 8312
rect 20183 8303 20215 8368
rect 20639 8361 20654 8395
rect 20694 8361 20704 8398
rect 20639 8352 20704 8361
rect 20183 8283 20187 8303
rect 20208 8283 20215 8303
rect 20183 8276 20215 8283
rect 20492 8220 20593 8221
rect 20390 8207 20593 8220
rect 20390 8205 20533 8207
rect 20390 8202 20467 8205
rect 20390 8175 20393 8202
rect 20422 8178 20467 8202
rect 20496 8178 20533 8205
rect 20422 8175 20533 8178
rect 20390 8174 20533 8175
rect 20569 8174 20593 8207
rect 20390 8161 20593 8174
rect 19970 8096 20005 8108
rect 19901 8089 20005 8096
rect 19901 8088 19977 8089
rect 19901 8068 19922 8088
rect 19954 8069 19977 8088
rect 20002 8069 20005 8089
rect 19954 8068 20005 8069
rect 19901 8059 20005 8068
rect 19970 8057 20005 8059
rect 19581 7975 19584 8014
rect 19629 7975 19646 8014
rect 20642 7991 20693 8352
rect 20640 7989 20697 7991
rect 19581 7953 19646 7975
rect 20629 7977 20697 7989
rect 20629 7944 20640 7977
rect 20680 7944 20697 7977
rect 20629 7938 20697 7944
rect 20629 7934 20693 7938
rect 19342 7889 19453 7892
rect 21072 7889 21179 8512
rect 17148 7875 21179 7889
rect 17148 7855 19349 7875
rect 19368 7855 19426 7875
rect 19445 7871 21179 7875
rect 19445 7855 20397 7871
rect 17148 7851 20397 7855
rect 20416 7851 20474 7871
rect 20493 7851 21179 7871
rect 17148 7833 21179 7851
rect 17148 7832 18718 7833
rect 20390 7829 20501 7833
rect 18709 7781 18744 7782
rect 18688 7774 18744 7781
rect 18688 7754 18717 7774
rect 18737 7754 18744 7774
rect 18688 7749 18744 7754
rect 19135 7777 19167 7784
rect 19757 7777 19792 7778
rect 19135 7757 19141 7777
rect 19162 7757 19167 7777
rect 19736 7770 19792 7777
rect 19601 7760 19659 7765
rect 18288 7694 18370 7723
rect 18288 7653 18313 7694
rect 18349 7653 18370 7694
rect 18475 7714 18539 7733
rect 18475 7675 18492 7714
rect 18526 7675 18539 7714
rect 18475 7656 18539 7675
rect 18288 7338 18370 7653
rect 18280 7293 18370 7338
rect 18477 7311 18539 7656
rect 18688 7471 18722 7749
rect 19135 7729 19167 7757
rect 18755 7721 19167 7729
rect 18755 7695 18761 7721
rect 18787 7695 19167 7721
rect 18755 7693 19167 7695
rect 18757 7692 18797 7693
rect 18924 7667 18955 7675
rect 18924 7637 18928 7667
rect 18949 7637 18955 7667
rect 18688 7463 18723 7471
rect 18688 7443 18696 7463
rect 18716 7443 18723 7463
rect 18688 7438 18723 7443
rect 18688 7437 18720 7438
rect 18924 7430 18955 7637
rect 19135 7628 19167 7693
rect 19135 7608 19139 7628
rect 19160 7608 19167 7628
rect 19135 7601 19167 7608
rect 19584 7751 19659 7760
rect 19584 7718 19593 7751
rect 19646 7718 19659 7751
rect 19584 7693 19659 7718
rect 19584 7660 19598 7693
rect 19651 7660 19659 7693
rect 19584 7654 19659 7660
rect 19736 7750 19765 7770
rect 19785 7750 19792 7770
rect 19736 7745 19792 7750
rect 20183 7773 20215 7780
rect 20183 7753 20189 7773
rect 20210 7753 20215 7773
rect 19444 7545 19545 7546
rect 19342 7532 19545 7545
rect 19342 7530 19485 7532
rect 19342 7527 19419 7530
rect 19342 7500 19345 7527
rect 19374 7503 19419 7527
rect 19448 7503 19485 7530
rect 19374 7500 19485 7503
rect 19342 7499 19485 7500
rect 19521 7499 19545 7532
rect 19342 7486 19545 7499
rect 18919 7412 18955 7430
rect 18886 7411 18955 7412
rect 18866 7399 18955 7411
rect 18866 7361 18878 7399
rect 18903 7364 18922 7399
rect 18947 7364 18955 7399
rect 19584 7388 19654 7654
rect 19736 7467 19770 7745
rect 20183 7725 20215 7753
rect 19803 7717 20215 7725
rect 19803 7691 19809 7717
rect 19835 7691 20215 7717
rect 19803 7689 20215 7691
rect 19805 7688 19845 7689
rect 19972 7663 20003 7671
rect 19972 7633 19976 7663
rect 19997 7633 20003 7663
rect 19736 7459 19771 7467
rect 19736 7439 19744 7459
rect 19764 7439 19771 7459
rect 19736 7434 19771 7439
rect 19972 7434 20003 7633
rect 20183 7624 20215 7689
rect 20183 7604 20187 7624
rect 20208 7604 20215 7624
rect 20183 7597 20215 7604
rect 20628 7750 20700 7768
rect 20628 7708 20641 7750
rect 20690 7708 20700 7750
rect 20628 7687 20700 7708
rect 20628 7645 20642 7687
rect 20691 7645 20700 7687
rect 20492 7541 20593 7542
rect 20390 7528 20593 7541
rect 20390 7526 20533 7528
rect 20390 7523 20467 7526
rect 20390 7496 20393 7523
rect 20422 7499 20467 7523
rect 20496 7499 20533 7526
rect 20422 7496 20533 7499
rect 20390 7495 20533 7496
rect 20569 7495 20593 7528
rect 20390 7482 20593 7495
rect 19736 7433 19768 7434
rect 19970 7431 20003 7434
rect 19936 7412 20004 7431
rect 18903 7361 18955 7364
rect 18866 7353 18955 7361
rect 19575 7359 19654 7388
rect 19906 7400 20005 7412
rect 19906 7362 19928 7400
rect 19953 7365 19972 7400
rect 19997 7365 20005 7400
rect 19953 7362 20005 7365
rect 18882 7352 18954 7353
rect 18476 7302 18550 7311
rect 18280 7260 18364 7293
rect 18280 7232 18295 7260
rect 18339 7232 18364 7260
rect 18280 7203 18364 7232
rect 18476 7254 18490 7302
rect 18527 7254 18550 7302
rect 18476 7226 18550 7254
rect 18280 7175 18292 7203
rect 18336 7175 18364 7203
rect 18280 7164 18364 7175
rect 19575 7176 19652 7359
rect 19906 7354 20005 7362
rect 19932 7353 20004 7354
rect 20628 7351 20700 7645
rect 21072 7373 21179 7833
rect 20628 7313 20704 7351
rect 21072 7313 21185 7373
rect 20639 7212 20704 7313
rect 19575 7133 19592 7176
rect 16508 7084 16523 7118
rect 16552 7084 16560 7118
rect 19580 7128 19592 7133
rect 19638 7128 19652 7176
rect 19580 7106 19652 7128
rect 20637 7166 20704 7212
rect 21074 7174 21185 7313
rect 16508 7058 16560 7084
rect 20637 7074 20702 7166
rect 21069 7147 21185 7174
rect 16508 7024 16522 7058
rect 16551 7024 16560 7058
rect 16508 6993 16560 7024
rect 20587 7056 20708 7074
rect 20587 7054 20658 7056
rect 20587 7013 20602 7054
rect 20639 7015 20658 7054
rect 20695 7015 20708 7056
rect 20639 7013 20708 7015
rect 20587 7003 20708 7013
rect 16784 6976 16895 6982
rect 16784 6974 18581 6976
rect 21069 6974 21176 7147
rect 16784 6965 21178 6974
rect 16784 6945 16791 6965
rect 16810 6945 16868 6965
rect 16887 6956 21178 6965
rect 16887 6945 20394 6956
rect 16784 6936 20394 6945
rect 20413 6936 20471 6956
rect 20490 6936 21178 6956
rect 16784 6923 21178 6936
rect 17103 6918 21178 6923
rect 18536 6917 18743 6918
rect 20387 6914 20498 6918
rect 16151 6871 16186 6872
rect 16130 6864 16186 6871
rect 16130 6844 16159 6864
rect 16179 6844 16186 6864
rect 16130 6839 16186 6844
rect 16577 6867 16609 6874
rect 16577 6847 16583 6867
rect 16604 6847 16609 6867
rect 16130 6561 16164 6839
rect 16577 6819 16609 6847
rect 19573 6855 19653 6867
rect 19754 6862 19789 6863
rect 19573 6829 19589 6855
rect 19629 6829 19653 6855
rect 16197 6811 16609 6819
rect 16197 6785 16203 6811
rect 16229 6785 16609 6811
rect 16197 6783 16609 6785
rect 16199 6782 16239 6783
rect 16366 6757 16397 6765
rect 16366 6727 16370 6757
rect 16391 6727 16397 6757
rect 16130 6553 16165 6561
rect 16130 6533 16138 6553
rect 16158 6533 16165 6553
rect 16366 6542 16397 6727
rect 16577 6718 16609 6783
rect 16991 6816 17102 6823
rect 16991 6815 17070 6816
rect 16991 6791 17013 6815
rect 17037 6792 17070 6815
rect 17094 6792 17102 6816
rect 17037 6791 17102 6792
rect 16991 6781 17102 6791
rect 19573 6810 19653 6829
rect 19573 6784 19592 6810
rect 19632 6784 19653 6810
rect 17052 6764 17101 6781
rect 19573 6757 19653 6784
rect 19573 6731 19596 6757
rect 19636 6731 19653 6757
rect 19573 6720 19653 6731
rect 19733 6855 19789 6862
rect 19733 6835 19762 6855
rect 19782 6835 19789 6855
rect 19733 6830 19789 6835
rect 20180 6858 20212 6865
rect 20180 6838 20186 6858
rect 20207 6838 20212 6858
rect 16577 6698 16581 6718
rect 16602 6698 16609 6718
rect 16577 6691 16609 6698
rect 16886 6635 16987 6636
rect 16784 6622 16987 6635
rect 16784 6620 16927 6622
rect 16784 6617 16861 6620
rect 16784 6590 16787 6617
rect 16816 6593 16861 6617
rect 16890 6593 16927 6620
rect 16816 6590 16927 6593
rect 16784 6589 16927 6590
rect 16963 6589 16987 6622
rect 16784 6576 16987 6589
rect 16130 6528 16165 6533
rect 16130 6527 16162 6528
rect 16364 6465 16398 6542
rect 14997 5062 15594 5066
rect 12097 4984 12132 4986
rect 12097 4975 12201 4984
rect 12097 4974 12148 4975
rect 12097 4954 12100 4974
rect 12125 4955 12148 4974
rect 12180 4955 12201 4975
rect 12125 4954 12201 4955
rect 12097 4947 12201 4954
rect 12097 4935 12132 4947
rect 11509 4869 11712 4882
rect 11509 4836 11533 4869
rect 11569 4868 11712 4869
rect 11569 4865 11680 4868
rect 11569 4838 11606 4865
rect 11635 4841 11680 4865
rect 11709 4841 11712 4868
rect 11635 4838 11712 4841
rect 11569 4836 11712 4838
rect 11509 4823 11712 4836
rect 11509 4822 11610 4823
rect 11887 4760 11919 4767
rect 11887 4740 11894 4760
rect 11915 4740 11919 4760
rect 11398 4682 11463 4691
rect 11398 4645 11408 4682
rect 11448 4648 11463 4682
rect 11887 4675 11919 4740
rect 12099 4731 12130 4935
rect 12334 4930 12366 4931
rect 12331 4925 12366 4930
rect 12331 4905 12338 4925
rect 12358 4905 12366 4925
rect 12331 4897 12366 4905
rect 12099 4701 12105 4731
rect 12126 4701 12130 4731
rect 12099 4693 12130 4701
rect 12257 4675 12297 4676
rect 11887 4673 12299 4675
rect 11448 4645 11465 4648
rect 11398 4626 11465 4645
rect 11398 4605 11412 4626
rect 11448 4605 11465 4626
rect 11398 4598 11465 4605
rect 11887 4647 12267 4673
rect 12293 4647 12299 4673
rect 11887 4639 12299 4647
rect 11887 4611 11919 4639
rect 12332 4619 12366 4897
rect 12456 4729 12521 5029
rect 14634 5017 15594 5062
rect 15701 5405 15737 6033
rect 14634 5013 15047 5017
rect 14634 4924 14668 5013
rect 14872 4927 14904 4928
rect 14047 4866 14250 4879
rect 14047 4833 14071 4866
rect 14107 4865 14250 4866
rect 14107 4862 14218 4865
rect 14107 4835 14144 4862
rect 14173 4838 14218 4862
rect 14247 4838 14250 4865
rect 14173 4835 14250 4838
rect 14107 4833 14250 4835
rect 14047 4820 14250 4833
rect 14047 4819 14148 4820
rect 14425 4757 14457 4764
rect 14425 4737 14432 4757
rect 14453 4737 14457 4757
rect 11887 4591 11892 4611
rect 11913 4591 11919 4611
rect 11887 4584 11919 4591
rect 12310 4614 12366 4619
rect 12310 4594 12317 4614
rect 12337 4594 12366 4614
rect 12310 4587 12366 4594
rect 12446 4718 12526 4729
rect 12446 4692 12463 4718
rect 12503 4692 12526 4718
rect 12446 4665 12526 4692
rect 12446 4639 12467 4665
rect 12507 4639 12526 4665
rect 12446 4620 12526 4639
rect 12446 4594 12470 4620
rect 12510 4594 12526 4620
rect 12310 4586 12345 4587
rect 12446 4582 12526 4594
rect 14425 4672 14457 4737
rect 14637 4728 14668 4924
rect 14869 4922 14904 4927
rect 14869 4902 14876 4922
rect 14896 4902 14904 4922
rect 14869 4894 14904 4902
rect 14637 4698 14643 4728
rect 14664 4698 14668 4728
rect 14637 4690 14668 4698
rect 14795 4672 14835 4673
rect 14425 4670 14837 4672
rect 14425 4644 14805 4670
rect 14831 4644 14837 4670
rect 14425 4636 14837 4644
rect 14425 4608 14457 4636
rect 14870 4616 14904 4894
rect 14425 4588 14430 4608
rect 14451 4588 14457 4608
rect 14425 4581 14457 4588
rect 14848 4611 14904 4616
rect 14848 4591 14855 4611
rect 14875 4591 14904 4611
rect 14848 4584 14904 4591
rect 14848 4583 14883 4584
rect 11601 4531 11712 4535
rect 13356 4531 13563 4532
rect 14139 4531 14250 4532
rect 10921 4513 14987 4531
rect 10921 4493 11609 4513
rect 11628 4493 11686 4513
rect 11705 4510 14987 4513
rect 11705 4493 14147 4510
rect 10921 4490 14147 4493
rect 14166 4490 14224 4510
rect 14243 4490 14987 4510
rect 10921 4475 14987 4490
rect 10923 4287 11030 4475
rect 13518 4473 14987 4475
rect 11391 4436 11512 4446
rect 11391 4434 11460 4436
rect 11391 4393 11404 4434
rect 11441 4395 11460 4434
rect 11497 4395 11512 4436
rect 11441 4393 11512 4395
rect 11391 4375 11512 4393
rect 10923 4283 11031 4287
rect 11397 4283 11474 4375
rect 12447 4371 12523 4387
rect 12447 4348 12462 4371
rect 8930 4117 8945 4140
rect 8869 4101 8945 4117
rect 9918 4113 9995 4205
rect 10361 4201 10469 4205
rect 9880 4095 10001 4113
rect 9880 4093 9951 4095
rect 9880 4052 9895 4093
rect 9932 4054 9951 4093
rect 9988 4054 10001 4095
rect 9932 4052 10001 4054
rect 9880 4042 10001 4052
rect 6451 4013 7874 4015
rect 10362 4013 10469 4201
rect 6451 3998 10471 4013
rect 6451 3978 7149 3998
rect 7168 3978 7226 3998
rect 7245 3995 10471 3998
rect 7245 3978 9687 3995
rect 6451 3975 9687 3978
rect 9706 3975 9764 3995
rect 9783 3975 10471 3995
rect 6451 3957 10471 3975
rect 7142 3956 7253 3957
rect 7829 3956 8036 3957
rect 9680 3953 9791 3957
rect 6509 3904 6544 3905
rect 6488 3897 6544 3904
rect 6488 3877 6517 3897
rect 6537 3877 6544 3897
rect 6488 3872 6544 3877
rect 6935 3900 6967 3907
rect 6935 3880 6941 3900
rect 6962 3880 6967 3900
rect 5657 3648 5683 3663
rect 5654 3641 5690 3648
rect 5654 3603 5660 3641
rect 5683 3603 5690 3641
rect 5654 3597 5690 3603
rect 6488 3594 6522 3872
rect 6935 3852 6967 3880
rect 6555 3844 6967 3852
rect 6555 3818 6561 3844
rect 6587 3818 6967 3844
rect 6555 3816 6967 3818
rect 6557 3815 6597 3816
rect 6724 3790 6755 3798
rect 6724 3760 6728 3790
rect 6749 3760 6755 3790
rect 6488 3586 6523 3594
rect 6488 3566 6496 3586
rect 6516 3566 6523 3586
rect 6488 3561 6523 3566
rect 6488 3560 6520 3561
rect 6724 3557 6755 3760
rect 6935 3751 6967 3816
rect 8866 3894 8946 3906
rect 9047 3901 9082 3902
rect 8866 3868 8882 3894
rect 8922 3868 8946 3894
rect 8866 3849 8946 3868
rect 8866 3823 8885 3849
rect 8925 3823 8946 3849
rect 8866 3796 8946 3823
rect 8866 3770 8889 3796
rect 8929 3770 8946 3796
rect 8866 3759 8946 3770
rect 9026 3894 9082 3901
rect 9026 3874 9055 3894
rect 9075 3874 9082 3894
rect 9026 3869 9082 3874
rect 9473 3897 9505 3904
rect 9473 3877 9479 3897
rect 9500 3877 9505 3897
rect 6935 3731 6939 3751
rect 6960 3731 6967 3751
rect 6935 3724 6967 3731
rect 7244 3668 7345 3669
rect 7142 3655 7345 3668
rect 7142 3653 7285 3655
rect 7142 3650 7219 3653
rect 7142 3623 7145 3650
rect 7174 3626 7219 3650
rect 7248 3626 7285 3653
rect 7174 3623 7285 3626
rect 7142 3622 7285 3623
rect 7321 3622 7345 3655
rect 7142 3609 7345 3622
rect 6719 3539 6755 3557
rect 6719 3522 6754 3539
rect 6652 3491 6757 3522
rect 6652 3486 6724 3491
rect 6652 3465 6683 3486
rect 6703 3470 6724 3486
rect 6744 3470 6757 3491
rect 6703 3465 6757 3470
rect 6652 3456 6757 3465
rect 8871 3459 8936 3759
rect 9026 3591 9060 3869
rect 9473 3849 9505 3877
rect 9093 3841 9505 3849
rect 9093 3815 9099 3841
rect 9125 3815 9505 3841
rect 9927 3883 9994 3890
rect 9927 3862 9944 3883
rect 9980 3862 9994 3883
rect 9927 3843 9994 3862
rect 9927 3840 9944 3843
rect 9093 3813 9505 3815
rect 9095 3812 9135 3813
rect 9262 3787 9293 3795
rect 9262 3757 9266 3787
rect 9287 3757 9293 3787
rect 9026 3583 9061 3591
rect 9026 3563 9034 3583
rect 9054 3563 9061 3583
rect 9026 3558 9061 3563
rect 9026 3557 9058 3558
rect 9262 3553 9293 3757
rect 9473 3748 9505 3813
rect 9929 3806 9944 3840
rect 9984 3806 9994 3843
rect 9929 3797 9994 3806
rect 9473 3728 9477 3748
rect 9498 3728 9505 3748
rect 9473 3721 9505 3728
rect 9782 3665 9883 3666
rect 9680 3652 9883 3665
rect 9680 3650 9823 3652
rect 9680 3647 9757 3650
rect 9680 3620 9683 3647
rect 9712 3623 9757 3647
rect 9786 3623 9823 3650
rect 9712 3620 9823 3623
rect 9680 3619 9823 3620
rect 9859 3619 9883 3652
rect 9680 3606 9883 3619
rect 9260 3541 9295 3553
rect 9191 3534 9295 3541
rect 9191 3533 9267 3534
rect 9191 3513 9212 3533
rect 9244 3514 9267 3533
rect 9292 3514 9295 3534
rect 9244 3513 9295 3514
rect 9191 3504 9295 3513
rect 9260 3502 9295 3504
rect 8871 3420 8874 3459
rect 8919 3420 8936 3459
rect 9932 3436 9983 3797
rect 9930 3434 9987 3436
rect 8871 3398 8936 3420
rect 9919 3422 9987 3434
rect 9919 3389 9930 3422
rect 9970 3389 9987 3422
rect 9919 3383 9987 3389
rect 9919 3379 9983 3383
rect 8632 3334 8743 3337
rect 10362 3334 10469 3957
rect 6675 3320 10469 3334
rect 6675 3300 8639 3320
rect 8658 3300 8716 3320
rect 8735 3316 10469 3320
rect 8735 3300 9687 3316
rect 6675 3296 9687 3300
rect 9706 3296 9764 3316
rect 9783 3296 10469 3316
rect 6675 3278 10469 3296
rect 6675 3277 7916 3278
rect 9680 3274 9791 3278
rect 7999 3226 8034 3227
rect 7978 3219 8034 3226
rect 7978 3199 8007 3219
rect 8027 3199 8034 3219
rect 7978 3194 8034 3199
rect 8425 3222 8457 3229
rect 9047 3222 9082 3223
rect 8425 3202 8431 3222
rect 8452 3202 8457 3222
rect 9026 3215 9082 3222
rect 8891 3205 8949 3210
rect 7978 2916 8012 3194
rect 8425 3174 8457 3202
rect 8045 3166 8457 3174
rect 8045 3140 8051 3166
rect 8077 3140 8457 3166
rect 8045 3138 8457 3140
rect 8047 3137 8087 3138
rect 8214 3112 8245 3120
rect 8214 3082 8218 3112
rect 8239 3082 8245 3112
rect 7978 2908 8013 2916
rect 7978 2888 7986 2908
rect 8006 2888 8013 2908
rect 7978 2883 8013 2888
rect 6719 2872 6755 2883
rect 7978 2882 8010 2883
rect 8214 2875 8245 3082
rect 8425 3073 8457 3138
rect 8425 3053 8429 3073
rect 8450 3053 8457 3073
rect 8425 3046 8457 3053
rect 8874 3196 8949 3205
rect 8874 3163 8883 3196
rect 8936 3163 8949 3196
rect 8874 3138 8949 3163
rect 8874 3105 8888 3138
rect 8941 3105 8949 3138
rect 8874 3099 8949 3105
rect 9026 3195 9055 3215
rect 9075 3195 9082 3215
rect 9026 3190 9082 3195
rect 9473 3218 9505 3225
rect 9473 3198 9479 3218
rect 9500 3198 9505 3218
rect 8734 2990 8835 2991
rect 8632 2977 8835 2990
rect 8632 2975 8775 2977
rect 8632 2972 8709 2975
rect 8632 2945 8635 2972
rect 8664 2948 8709 2972
rect 8738 2948 8775 2975
rect 8664 2945 8775 2948
rect 8632 2944 8775 2945
rect 8811 2944 8835 2977
rect 8632 2931 8835 2944
rect 6719 2849 6725 2872
rect 6749 2849 6755 2872
rect 8209 2866 8245 2875
rect 8154 2856 8251 2866
rect 6966 2854 8251 2856
rect 6719 2828 6755 2849
rect 6719 2805 6725 2828
rect 6749 2805 6755 2828
rect 6719 2652 6755 2805
rect 6931 2844 8251 2854
rect 6931 2806 6943 2844
rect 6968 2809 6987 2844
rect 7012 2809 8251 2844
rect 6968 2806 8251 2809
rect 6931 2803 8251 2806
rect 6931 2801 8248 2803
rect 6931 2798 7020 2801
rect 6947 2797 7019 2798
rect 8874 2788 8944 3099
rect 9026 2912 9060 3190
rect 9473 3170 9505 3198
rect 9093 3162 9505 3170
rect 9093 3136 9099 3162
rect 9125 3136 9505 3162
rect 9093 3134 9505 3136
rect 9095 3133 9135 3134
rect 9262 3108 9293 3116
rect 9262 3078 9266 3108
rect 9287 3078 9293 3108
rect 9026 2904 9061 2912
rect 9026 2884 9034 2904
rect 9054 2884 9061 2904
rect 9026 2879 9061 2884
rect 9262 2879 9293 3078
rect 9473 3069 9505 3134
rect 9473 3049 9477 3069
rect 9498 3049 9505 3069
rect 9473 3042 9505 3049
rect 9918 3195 9990 3213
rect 9918 3153 9931 3195
rect 9980 3153 9990 3195
rect 9918 3132 9990 3153
rect 9918 3090 9932 3132
rect 9981 3090 9990 3132
rect 9782 2986 9883 2987
rect 9680 2973 9883 2986
rect 9680 2971 9823 2973
rect 9680 2968 9757 2971
rect 9680 2941 9683 2968
rect 9712 2944 9757 2968
rect 9786 2944 9823 2971
rect 9712 2941 9823 2944
rect 9680 2940 9823 2941
rect 9859 2940 9883 2973
rect 9680 2927 9883 2940
rect 9026 2878 9058 2879
rect 9260 2876 9293 2879
rect 9226 2857 9294 2876
rect 9196 2845 9295 2857
rect 9918 2849 9990 3090
rect 10362 2849 10469 3278
rect 10924 3690 11031 4283
rect 11399 4232 11474 4283
rect 12440 4334 12462 4348
rect 12506 4334 12523 4371
rect 12440 4314 12523 4334
rect 12440 4248 12457 4314
rect 12511 4248 12523 4314
rect 11399 4189 11475 4232
rect 11403 3878 11475 4189
rect 12440 4224 12523 4248
rect 12440 4204 12516 4224
rect 12440 4185 12519 4204
rect 12099 4169 12171 4170
rect 12098 4161 12197 4169
rect 12098 4158 12150 4161
rect 12098 4123 12106 4158
rect 12131 4123 12150 4158
rect 12175 4123 12197 4161
rect 12098 4111 12197 4123
rect 12099 4092 12167 4111
rect 12100 4089 12133 4092
rect 12335 4089 12367 4090
rect 11510 4028 11713 4041
rect 11510 3995 11534 4028
rect 11570 4027 11713 4028
rect 11570 4024 11681 4027
rect 11570 3997 11607 4024
rect 11636 4000 11681 4024
rect 11710 4000 11713 4027
rect 11636 3997 11713 4000
rect 11570 3995 11713 3997
rect 11510 3982 11713 3995
rect 11510 3981 11611 3982
rect 11403 3836 11412 3878
rect 11461 3836 11475 3878
rect 11403 3815 11475 3836
rect 11403 3773 11413 3815
rect 11462 3773 11475 3815
rect 11403 3755 11475 3773
rect 11888 3919 11920 3926
rect 11888 3899 11895 3919
rect 11916 3899 11920 3919
rect 11888 3834 11920 3899
rect 12100 3890 12131 4089
rect 12332 4084 12367 4089
rect 12332 4064 12339 4084
rect 12359 4064 12367 4084
rect 12332 4056 12367 4064
rect 12100 3860 12106 3890
rect 12127 3860 12131 3890
rect 12100 3852 12131 3860
rect 12258 3834 12298 3835
rect 11888 3832 12300 3834
rect 11888 3806 12268 3832
rect 12294 3806 12300 3832
rect 11888 3798 12300 3806
rect 11888 3770 11920 3798
rect 12333 3778 12367 4056
rect 12449 3869 12519 4185
rect 14437 4170 14468 4171
rect 14437 4162 14482 4170
rect 13517 4139 13681 4146
rect 14437 4139 14447 4162
rect 13143 4124 14447 4139
rect 14472 4124 14482 4162
rect 15701 4165 15735 5405
rect 15701 4161 15931 4165
rect 15701 4135 15900 4161
rect 15925 4135 15931 4161
rect 15701 4127 15931 4135
rect 13143 4106 14482 4124
rect 13148 4093 13184 4106
rect 13517 4103 13681 4106
rect 12558 4024 12761 4037
rect 12558 3991 12582 4024
rect 12618 4023 12761 4024
rect 12618 4020 12729 4023
rect 12618 3993 12655 4020
rect 12684 3996 12729 4020
rect 12758 3996 12761 4023
rect 12684 3993 12761 3996
rect 12618 3991 12761 3993
rect 12558 3978 12761 3991
rect 12558 3977 12659 3978
rect 11888 3750 11893 3770
rect 11914 3750 11920 3770
rect 11888 3743 11920 3750
rect 12311 3773 12367 3778
rect 12311 3753 12318 3773
rect 12338 3753 12367 3773
rect 12444 3863 12519 3869
rect 12444 3830 12452 3863
rect 12505 3830 12519 3863
rect 12444 3805 12519 3830
rect 12444 3772 12457 3805
rect 12510 3772 12519 3805
rect 12444 3763 12519 3772
rect 12936 3915 12968 3922
rect 12936 3895 12943 3915
rect 12964 3895 12968 3915
rect 12936 3830 12968 3895
rect 13148 3886 13179 4093
rect 16285 4091 16317 4092
rect 13383 4085 13415 4086
rect 13380 4080 13415 4085
rect 13380 4060 13387 4080
rect 13407 4060 13415 4080
rect 13380 4052 13415 4060
rect 13148 3856 13154 3886
rect 13175 3856 13179 3886
rect 13148 3848 13179 3856
rect 13306 3830 13346 3831
rect 12936 3828 13348 3830
rect 12936 3802 13316 3828
rect 13342 3802 13348 3828
rect 12936 3794 13348 3802
rect 12936 3766 12968 3794
rect 13381 3774 13415 4052
rect 15460 4030 15663 4043
rect 15460 3997 15484 4030
rect 15520 4029 15663 4030
rect 15520 4026 15631 4029
rect 15520 3999 15557 4026
rect 15586 4002 15631 4026
rect 15660 4002 15663 4029
rect 15586 3999 15663 4002
rect 15520 3997 15663 3999
rect 15460 3984 15663 3997
rect 15460 3983 15561 3984
rect 12444 3758 12502 3763
rect 12311 3746 12367 3753
rect 12936 3746 12941 3766
rect 12962 3746 12968 3766
rect 12311 3745 12346 3746
rect 12936 3739 12968 3746
rect 13359 3769 13415 3774
rect 13359 3749 13366 3769
rect 13386 3749 13415 3769
rect 13359 3742 13415 3749
rect 15838 3921 15870 3928
rect 15838 3901 15845 3921
rect 15866 3901 15870 3921
rect 15838 3836 15870 3901
rect 16050 3892 16081 4089
rect 16282 4086 16317 4091
rect 16282 4066 16289 4086
rect 16309 4066 16317 4086
rect 16282 4058 16317 4066
rect 16050 3862 16056 3892
rect 16077 3862 16081 3892
rect 16050 3854 16081 3862
rect 16208 3836 16248 3837
rect 15838 3834 16250 3836
rect 15838 3808 16218 3834
rect 16244 3808 16250 3834
rect 15838 3800 16250 3808
rect 15838 3772 15870 3800
rect 15838 3752 15843 3772
rect 15864 3752 15870 3772
rect 15838 3745 15870 3752
rect 16040 3774 16088 3781
rect 16283 3780 16317 4058
rect 16040 3754 16047 3774
rect 16080 3754 16088 3774
rect 13359 3741 13394 3742
rect 11602 3690 11713 3694
rect 13385 3690 14955 3691
rect 10924 3686 14955 3690
rect 15280 3686 15698 3699
rect 10924 3674 15698 3686
rect 10924 3672 15560 3674
rect 10924 3652 11610 3672
rect 11629 3652 11687 3672
rect 11706 3668 15560 3672
rect 11706 3652 12658 3668
rect 10924 3648 12658 3652
rect 12677 3648 12735 3668
rect 12754 3654 15560 3668
rect 15579 3654 15637 3674
rect 15656 3654 15698 3674
rect 12754 3648 15698 3654
rect 10924 3634 15698 3648
rect 10924 3011 11031 3634
rect 12650 3631 12761 3634
rect 15280 3628 15698 3634
rect 11410 3585 11474 3589
rect 11406 3579 11474 3585
rect 11406 3546 11423 3579
rect 11463 3546 11474 3579
rect 11406 3534 11474 3546
rect 12457 3548 12522 3570
rect 11406 3532 11463 3534
rect 11410 3171 11461 3532
rect 12457 3509 12474 3548
rect 12519 3509 12522 3548
rect 12098 3464 12133 3466
rect 12098 3455 12202 3464
rect 12098 3454 12149 3455
rect 12098 3434 12101 3454
rect 12126 3435 12149 3454
rect 12181 3435 12202 3455
rect 12126 3434 12202 3435
rect 12098 3427 12202 3434
rect 12098 3415 12133 3427
rect 11510 3349 11713 3362
rect 11510 3316 11534 3349
rect 11570 3348 11713 3349
rect 11570 3345 11681 3348
rect 11570 3318 11607 3345
rect 11636 3321 11681 3345
rect 11710 3321 11713 3348
rect 11636 3318 11713 3321
rect 11570 3316 11713 3318
rect 11510 3303 11713 3316
rect 11510 3302 11611 3303
rect 11888 3240 11920 3247
rect 11888 3220 11895 3240
rect 11916 3220 11920 3240
rect 11399 3162 11464 3171
rect 11399 3125 11409 3162
rect 11449 3128 11464 3162
rect 11888 3155 11920 3220
rect 12100 3211 12131 3415
rect 12335 3410 12367 3411
rect 12332 3405 12367 3410
rect 12332 3385 12339 3405
rect 12359 3385 12367 3405
rect 12332 3377 12367 3385
rect 12100 3181 12106 3211
rect 12127 3181 12131 3211
rect 12100 3173 12131 3181
rect 12258 3155 12298 3156
rect 11888 3153 12300 3155
rect 11449 3125 11466 3128
rect 11399 3106 11466 3125
rect 11399 3085 11413 3106
rect 11449 3085 11466 3106
rect 11399 3078 11466 3085
rect 11888 3127 12268 3153
rect 12294 3127 12300 3153
rect 11888 3119 12300 3127
rect 11888 3091 11920 3119
rect 12333 3099 12367 3377
rect 12457 3209 12522 3509
rect 14594 3470 14631 3491
rect 14594 3433 14605 3470
rect 14622 3446 14631 3470
rect 14622 3433 14632 3446
rect 14594 3423 14632 3433
rect 14595 3419 14632 3423
rect 14595 3413 14628 3419
rect 14005 3344 14208 3357
rect 14005 3311 14029 3344
rect 14065 3343 14208 3344
rect 14065 3340 14176 3343
rect 14065 3313 14102 3340
rect 14131 3316 14176 3340
rect 14205 3316 14208 3343
rect 14131 3313 14208 3316
rect 14065 3311 14208 3313
rect 14005 3298 14208 3311
rect 14005 3297 14106 3298
rect 14383 3235 14415 3242
rect 14383 3215 14390 3235
rect 14411 3215 14415 3235
rect 11888 3071 11893 3091
rect 11914 3071 11920 3091
rect 11888 3064 11920 3071
rect 12311 3094 12367 3099
rect 12311 3074 12318 3094
rect 12338 3074 12367 3094
rect 12311 3067 12367 3074
rect 12447 3198 12527 3209
rect 12447 3172 12464 3198
rect 12504 3172 12527 3198
rect 12447 3145 12527 3172
rect 12447 3119 12468 3145
rect 12508 3119 12527 3145
rect 12447 3100 12527 3119
rect 12447 3074 12471 3100
rect 12511 3074 12527 3100
rect 13521 3144 13626 3165
rect 14383 3150 14415 3215
rect 14595 3206 14626 3413
rect 14830 3405 14862 3406
rect 14827 3400 14862 3405
rect 14827 3380 14834 3400
rect 14854 3380 14862 3400
rect 14827 3372 14862 3380
rect 14595 3176 14601 3206
rect 14622 3176 14626 3206
rect 14595 3168 14626 3176
rect 14753 3150 14793 3151
rect 14383 3148 14795 3150
rect 13521 3138 13997 3144
rect 13521 3136 13578 3138
rect 13521 3105 13533 3136
rect 13558 3115 13578 3136
rect 13604 3131 13997 3138
rect 13604 3115 13958 3131
rect 13558 3108 13958 3115
rect 13984 3108 13997 3131
rect 13558 3105 13997 3108
rect 13521 3095 13997 3105
rect 14383 3122 14763 3148
rect 14789 3122 14795 3148
rect 14383 3114 14795 3122
rect 13521 3093 13626 3095
rect 12311 3066 12346 3067
rect 12447 3062 12527 3074
rect 14383 3086 14415 3114
rect 14828 3094 14862 3372
rect 14383 3066 14388 3086
rect 14409 3066 14415 3086
rect 14383 3059 14415 3066
rect 14806 3089 14862 3094
rect 14806 3069 14813 3089
rect 14833 3069 14862 3089
rect 14806 3062 14862 3069
rect 14806 3061 14841 3062
rect 11602 3011 11713 3015
rect 13344 3011 14997 3014
rect 10922 2993 14997 3011
rect 10922 2973 11610 2993
rect 11629 2973 11687 2993
rect 11706 2988 14997 2993
rect 11706 2973 14105 2988
rect 10922 2968 14105 2973
rect 14124 2968 14182 2988
rect 14201 2968 14997 2988
rect 10922 2958 14997 2968
rect 10922 2955 11547 2958
rect 11734 2955 14997 2958
rect 9196 2807 9218 2845
rect 9243 2810 9262 2845
rect 9287 2810 9295 2845
rect 9243 2807 9295 2810
rect 9196 2799 9295 2807
rect 9222 2798 9294 2799
rect 8873 2772 8944 2788
rect 8873 2756 8893 2772
rect 8874 2726 8893 2756
rect 8876 2706 8893 2726
rect 8923 2726 8944 2772
rect 9916 2768 9994 2849
rect 10361 2794 10469 2849
rect 8923 2706 8943 2726
rect 8876 2687 8943 2706
rect 9916 2666 9995 2768
rect 6710 2643 6796 2652
rect 6710 2625 6729 2643
rect 6781 2625 6796 2643
rect 6710 2621 6796 2625
rect 9880 2648 10001 2666
rect 9880 2646 9951 2648
rect 9880 2605 9895 2646
rect 9932 2607 9951 2646
rect 9988 2607 10001 2648
rect 9932 2605 10001 2607
rect 9880 2595 10001 2605
rect 7185 2567 7296 2570
rect 6500 2566 8049 2567
rect 10362 2566 10469 2794
rect 10924 2727 11031 2955
rect 13344 2954 14997 2955
rect 14097 2951 14208 2954
rect 11392 2916 11513 2926
rect 11392 2914 11461 2916
rect 11392 2873 11405 2914
rect 11442 2875 11461 2914
rect 11498 2875 11513 2916
rect 11442 2873 11513 2875
rect 11392 2855 11513 2873
rect 11398 2753 11477 2855
rect 12450 2815 12517 2834
rect 12450 2795 12470 2815
rect 10924 2672 11032 2727
rect 11399 2672 11477 2753
rect 12449 2749 12470 2795
rect 12500 2795 12517 2815
rect 12500 2765 12519 2795
rect 12500 2749 12520 2765
rect 12449 2733 12520 2749
rect 12099 2722 12171 2723
rect 12098 2714 12197 2722
rect 12098 2711 12150 2714
rect 12098 2676 12106 2711
rect 12131 2676 12150 2711
rect 12175 2676 12197 2714
rect 6500 2563 9659 2566
rect 9846 2563 10471 2566
rect 6500 2553 10471 2563
rect 6500 2533 7192 2553
rect 7211 2533 7269 2553
rect 7288 2548 10471 2553
rect 7288 2533 9687 2548
rect 6500 2528 9687 2533
rect 9706 2528 9764 2548
rect 9783 2528 10471 2548
rect 6500 2510 10471 2528
rect 6500 2507 8049 2510
rect 9680 2506 9791 2510
rect 6552 2459 6587 2460
rect 6531 2452 6587 2459
rect 6531 2432 6560 2452
rect 6580 2432 6587 2452
rect 6531 2427 6587 2432
rect 6978 2455 7010 2462
rect 6978 2435 6984 2455
rect 7005 2435 7010 2455
rect 6531 2149 6565 2427
rect 6978 2407 7010 2435
rect 6598 2399 7010 2407
rect 6598 2373 6604 2399
rect 6630 2373 7010 2399
rect 6598 2371 7010 2373
rect 6600 2370 6640 2371
rect 6767 2345 6798 2353
rect 6767 2315 6771 2345
rect 6792 2315 6798 2345
rect 6531 2141 6566 2149
rect 6531 2121 6539 2141
rect 6559 2121 6566 2141
rect 6531 2116 6566 2121
rect 6531 2115 6563 2116
rect 6767 2114 6798 2315
rect 6978 2306 7010 2371
rect 6978 2286 6982 2306
rect 7003 2286 7010 2306
rect 6978 2279 7010 2286
rect 7572 2446 7665 2453
rect 7572 2405 7596 2446
rect 7650 2405 7665 2446
rect 7287 2223 7388 2224
rect 7185 2210 7388 2223
rect 7185 2208 7328 2210
rect 7185 2205 7262 2208
rect 7185 2178 7188 2205
rect 7217 2181 7262 2205
rect 7291 2181 7328 2208
rect 7217 2178 7328 2181
rect 7185 2177 7328 2178
rect 7364 2177 7388 2210
rect 7185 2164 7388 2177
rect 7572 2032 7665 2405
rect 8866 2447 8946 2459
rect 9047 2454 9082 2455
rect 8866 2421 8882 2447
rect 8922 2421 8946 2447
rect 8866 2402 8946 2421
rect 8866 2376 8885 2402
rect 8925 2376 8946 2402
rect 8866 2349 8946 2376
rect 8866 2323 8889 2349
rect 8929 2323 8946 2349
rect 8866 2312 8946 2323
rect 9026 2447 9082 2454
rect 9026 2427 9055 2447
rect 9075 2427 9082 2447
rect 9026 2422 9082 2427
rect 9473 2450 9505 2457
rect 9473 2430 9479 2450
rect 9500 2430 9505 2450
rect 7572 1988 7590 2032
rect 7650 1988 7665 2032
rect 7572 1973 7665 1988
rect 8871 2012 8936 2312
rect 9026 2144 9060 2422
rect 9473 2402 9505 2430
rect 9093 2394 9505 2402
rect 9093 2368 9099 2394
rect 9125 2368 9505 2394
rect 9927 2436 9994 2443
rect 9927 2415 9944 2436
rect 9980 2415 9994 2436
rect 9927 2396 9994 2415
rect 9927 2393 9944 2396
rect 9093 2366 9505 2368
rect 9095 2365 9135 2366
rect 9262 2340 9293 2348
rect 9262 2310 9266 2340
rect 9287 2310 9293 2340
rect 9026 2136 9061 2144
rect 9026 2116 9034 2136
rect 9054 2116 9061 2136
rect 9026 2111 9061 2116
rect 9026 2110 9058 2111
rect 9262 2106 9293 2310
rect 9473 2301 9505 2366
rect 9929 2359 9944 2393
rect 9984 2359 9994 2396
rect 9929 2350 9994 2359
rect 9473 2281 9477 2301
rect 9498 2281 9505 2301
rect 9473 2274 9505 2281
rect 9782 2218 9883 2219
rect 9680 2205 9883 2218
rect 9680 2203 9823 2205
rect 9680 2200 9757 2203
rect 9680 2173 9683 2200
rect 9712 2176 9757 2200
rect 9786 2176 9823 2203
rect 9712 2173 9823 2176
rect 9680 2172 9823 2173
rect 9859 2172 9883 2205
rect 9680 2159 9883 2172
rect 9260 2094 9295 2106
rect 9191 2087 9295 2094
rect 9191 2086 9267 2087
rect 9191 2066 9212 2086
rect 9244 2067 9267 2086
rect 9292 2067 9295 2087
rect 9244 2066 9295 2067
rect 9191 2057 9295 2066
rect 9260 2055 9295 2057
rect 8871 1973 8874 2012
rect 8919 1973 8936 2012
rect 9932 1989 9983 2350
rect 9930 1987 9987 1989
rect 8871 1951 8936 1973
rect 9919 1975 9987 1987
rect 9919 1942 9930 1975
rect 9970 1942 9987 1975
rect 9919 1936 9987 1942
rect 9919 1932 9983 1936
rect 8632 1887 8743 1890
rect 10362 1887 10469 2510
rect 6895 1873 10469 1887
rect 6895 1853 8639 1873
rect 8658 1853 8716 1873
rect 8735 1869 10469 1873
rect 8735 1853 9687 1869
rect 6895 1849 9687 1853
rect 9706 1849 9764 1869
rect 9783 1849 10469 1869
rect 6895 1831 10469 1849
rect 6895 1830 8008 1831
rect 9680 1827 9791 1831
rect 7999 1779 8034 1780
rect 7978 1772 8034 1779
rect 7978 1752 8007 1772
rect 8027 1752 8034 1772
rect 7978 1747 8034 1752
rect 8425 1775 8457 1782
rect 9047 1775 9082 1776
rect 8425 1755 8431 1775
rect 8452 1755 8457 1775
rect 9026 1768 9082 1775
rect 8891 1758 8949 1763
rect 5814 1712 7667 1745
rect 5814 1647 5879 1712
rect 6010 1692 7667 1712
rect 6010 1651 7603 1692
rect 7639 1651 7667 1692
rect 7765 1712 7829 1731
rect 7765 1673 7782 1712
rect 7816 1673 7829 1712
rect 7765 1654 7829 1673
rect 6010 1647 7667 1651
rect 5814 1622 7667 1647
rect 7578 1619 7660 1622
rect 7767 1142 7829 1654
rect 7978 1469 8012 1747
rect 8425 1727 8457 1755
rect 8045 1719 8457 1727
rect 8045 1693 8051 1719
rect 8077 1693 8457 1719
rect 8045 1691 8457 1693
rect 8047 1690 8087 1691
rect 8214 1665 8245 1673
rect 8214 1635 8218 1665
rect 8239 1635 8245 1665
rect 7978 1461 8013 1469
rect 7978 1441 7986 1461
rect 8006 1441 8013 1461
rect 7978 1436 8013 1441
rect 7978 1435 8010 1436
rect 8214 1428 8245 1635
rect 8425 1626 8457 1691
rect 8425 1606 8429 1626
rect 8450 1606 8457 1626
rect 8425 1599 8457 1606
rect 8874 1749 8949 1758
rect 8874 1716 8883 1749
rect 8936 1716 8949 1749
rect 8874 1691 8949 1716
rect 8874 1658 8888 1691
rect 8941 1658 8949 1691
rect 8874 1652 8949 1658
rect 9026 1748 9055 1768
rect 9075 1748 9082 1768
rect 9026 1743 9082 1748
rect 9473 1771 9505 1778
rect 9473 1751 9479 1771
rect 9500 1751 9505 1771
rect 8734 1543 8835 1544
rect 8632 1530 8835 1543
rect 8632 1528 8775 1530
rect 8632 1525 8709 1528
rect 8632 1498 8635 1525
rect 8664 1501 8709 1525
rect 8738 1501 8775 1528
rect 8664 1498 8775 1501
rect 8632 1497 8775 1498
rect 8811 1497 8835 1530
rect 8632 1484 8835 1497
rect 8209 1410 8245 1428
rect 8176 1409 8245 1410
rect 8156 1397 8245 1409
rect 8156 1359 8168 1397
rect 8193 1362 8212 1397
rect 8237 1362 8245 1397
rect 8193 1359 8245 1362
rect 8156 1351 8245 1359
rect 8172 1350 8244 1351
rect 7725 1084 7841 1142
rect 8874 1131 8944 1652
rect 9026 1465 9060 1743
rect 9473 1723 9505 1751
rect 9093 1715 9505 1723
rect 9093 1689 9099 1715
rect 9125 1689 9505 1715
rect 9093 1687 9505 1689
rect 9095 1686 9135 1687
rect 9262 1661 9293 1669
rect 9262 1631 9266 1661
rect 9287 1631 9293 1661
rect 9026 1457 9061 1465
rect 9026 1437 9034 1457
rect 9054 1437 9061 1457
rect 9026 1432 9061 1437
rect 9262 1432 9293 1631
rect 9473 1622 9505 1687
rect 9473 1602 9477 1622
rect 9498 1602 9505 1622
rect 9473 1595 9505 1602
rect 9918 1748 9990 1766
rect 9918 1706 9931 1748
rect 9980 1706 9990 1748
rect 9918 1685 9990 1706
rect 9918 1643 9932 1685
rect 9981 1643 9990 1685
rect 9782 1539 9883 1540
rect 9680 1526 9883 1539
rect 9680 1524 9823 1526
rect 9680 1521 9757 1524
rect 9680 1494 9683 1521
rect 9712 1497 9757 1521
rect 9786 1497 9823 1524
rect 9712 1494 9823 1497
rect 9680 1493 9823 1494
rect 9859 1493 9883 1526
rect 9680 1480 9883 1493
rect 9026 1431 9058 1432
rect 9260 1429 9293 1432
rect 9226 1410 9294 1429
rect 9196 1398 9295 1410
rect 9196 1360 9218 1398
rect 9243 1363 9262 1398
rect 9287 1363 9295 1398
rect 9243 1360 9295 1363
rect 9196 1352 9295 1360
rect 9222 1351 9294 1352
rect 7725 1013 7737 1084
rect 7816 1013 7841 1084
rect 7725 993 7841 1013
rect 8855 930 8957 1131
rect 9918 1123 9990 1643
rect 10362 1219 10469 1831
rect 10924 2243 11031 2672
rect 11403 2431 11475 2672
rect 12098 2664 12197 2676
rect 12099 2645 12167 2664
rect 12100 2642 12133 2645
rect 12335 2642 12367 2643
rect 11510 2581 11713 2594
rect 11510 2548 11534 2581
rect 11570 2580 11713 2581
rect 11570 2577 11681 2580
rect 11570 2550 11607 2577
rect 11636 2553 11681 2577
rect 11710 2553 11713 2580
rect 11636 2550 11713 2553
rect 11570 2548 11713 2550
rect 11510 2535 11713 2548
rect 11510 2534 11611 2535
rect 11403 2389 11412 2431
rect 11461 2389 11475 2431
rect 11403 2368 11475 2389
rect 11403 2326 11413 2368
rect 11462 2326 11475 2368
rect 11403 2308 11475 2326
rect 11888 2472 11920 2479
rect 11888 2452 11895 2472
rect 11916 2452 11920 2472
rect 11888 2387 11920 2452
rect 12100 2443 12131 2642
rect 12332 2637 12367 2642
rect 12332 2617 12339 2637
rect 12359 2617 12367 2637
rect 12332 2609 12367 2617
rect 12100 2413 12106 2443
rect 12127 2413 12131 2443
rect 12100 2405 12131 2413
rect 12258 2387 12298 2388
rect 11888 2385 12300 2387
rect 11888 2359 12268 2385
rect 12294 2359 12300 2385
rect 11888 2351 12300 2359
rect 11888 2323 11920 2351
rect 12333 2331 12367 2609
rect 12449 2422 12519 2733
rect 13146 2724 14488 2729
rect 13146 2722 14445 2724
rect 13143 2696 14445 2722
rect 14473 2696 14488 2724
rect 13143 2688 14488 2696
rect 13143 2663 13182 2688
rect 13143 2646 13184 2663
rect 13143 2639 13182 2646
rect 12558 2577 12761 2590
rect 12558 2544 12582 2577
rect 12618 2576 12761 2577
rect 12618 2573 12729 2576
rect 12618 2546 12655 2573
rect 12684 2549 12729 2573
rect 12758 2549 12761 2576
rect 12684 2546 12761 2549
rect 12618 2544 12761 2546
rect 12558 2531 12761 2544
rect 12558 2530 12659 2531
rect 11888 2303 11893 2323
rect 11914 2303 11920 2323
rect 11888 2296 11920 2303
rect 12311 2326 12367 2331
rect 12311 2306 12318 2326
rect 12338 2306 12367 2326
rect 12444 2416 12519 2422
rect 12444 2383 12452 2416
rect 12505 2383 12519 2416
rect 12444 2358 12519 2383
rect 12444 2325 12457 2358
rect 12510 2325 12519 2358
rect 12444 2316 12519 2325
rect 12936 2468 12968 2475
rect 12936 2448 12943 2468
rect 12964 2448 12968 2468
rect 12936 2383 12968 2448
rect 13148 2439 13179 2639
rect 13383 2638 13415 2639
rect 13380 2633 13415 2638
rect 13380 2613 13387 2633
rect 13407 2613 13415 2633
rect 13380 2605 13415 2613
rect 13148 2409 13154 2439
rect 13175 2409 13179 2439
rect 13148 2401 13179 2409
rect 13306 2383 13346 2384
rect 12936 2381 13348 2383
rect 12936 2355 13316 2381
rect 13342 2355 13348 2381
rect 12936 2347 13348 2355
rect 12936 2319 12968 2347
rect 13381 2327 13415 2605
rect 12444 2311 12502 2316
rect 12311 2299 12367 2306
rect 12936 2299 12941 2319
rect 12962 2299 12968 2319
rect 12311 2298 12346 2299
rect 12936 2292 12968 2299
rect 13359 2322 13415 2327
rect 13359 2302 13366 2322
rect 13386 2302 13415 2322
rect 13359 2295 13415 2302
rect 13359 2294 13394 2295
rect 11602 2243 11713 2247
rect 13477 2243 14997 2244
rect 10924 2225 14997 2243
rect 10924 2205 11610 2225
rect 11629 2205 11687 2225
rect 11706 2221 14997 2225
rect 11706 2205 12658 2221
rect 10924 2201 12658 2205
rect 12677 2201 12735 2221
rect 12754 2201 14997 2221
rect 10924 2187 14997 2201
rect 10924 1564 11031 2187
rect 12650 2184 12761 2187
rect 11410 2138 11474 2142
rect 11406 2132 11474 2138
rect 11406 2099 11423 2132
rect 11463 2099 11474 2132
rect 11406 2087 11474 2099
rect 12457 2101 12522 2123
rect 11406 2085 11463 2087
rect 11410 1724 11461 2085
rect 12457 2062 12474 2101
rect 12519 2062 12522 2101
rect 12098 2017 12133 2019
rect 12098 2008 12202 2017
rect 12098 2007 12149 2008
rect 12098 1987 12101 2007
rect 12126 1988 12149 2007
rect 12181 1988 12202 2008
rect 12126 1987 12202 1988
rect 12098 1980 12202 1987
rect 12098 1968 12133 1980
rect 11510 1902 11713 1915
rect 11510 1869 11534 1902
rect 11570 1901 11713 1902
rect 11570 1898 11681 1901
rect 11570 1871 11607 1898
rect 11636 1874 11681 1898
rect 11710 1874 11713 1901
rect 11636 1871 11713 1874
rect 11570 1869 11713 1871
rect 11510 1856 11713 1869
rect 11510 1855 11611 1856
rect 11888 1793 11920 1800
rect 11888 1773 11895 1793
rect 11916 1773 11920 1793
rect 11399 1715 11464 1724
rect 11399 1678 11409 1715
rect 11449 1681 11464 1715
rect 11888 1708 11920 1773
rect 12100 1764 12131 1968
rect 12335 1963 12367 1964
rect 12332 1958 12367 1963
rect 12332 1938 12339 1958
rect 12359 1938 12367 1958
rect 12332 1930 12367 1938
rect 12100 1734 12106 1764
rect 12127 1734 12131 1764
rect 12100 1726 12131 1734
rect 12258 1708 12298 1709
rect 11888 1706 12300 1708
rect 11449 1678 11466 1681
rect 11399 1659 11466 1678
rect 11399 1638 11413 1659
rect 11449 1638 11466 1659
rect 11399 1631 11466 1638
rect 11888 1680 12268 1706
rect 12294 1680 12300 1706
rect 11888 1672 12300 1680
rect 11888 1644 11920 1672
rect 12333 1652 12367 1930
rect 12457 1799 12522 2062
rect 12457 1795 12518 1799
rect 11888 1624 11893 1644
rect 11914 1624 11920 1644
rect 11888 1617 11920 1624
rect 12311 1647 12367 1652
rect 12311 1627 12318 1647
rect 12338 1627 12367 1647
rect 12311 1620 12367 1627
rect 12311 1619 12346 1620
rect 11602 1564 11713 1568
rect 10922 1546 12241 1564
rect 10922 1526 11610 1546
rect 11629 1526 11687 1546
rect 11706 1526 12241 1546
rect 10922 1508 12241 1526
rect 10924 1388 11031 1508
rect 11392 1469 11513 1479
rect 11392 1467 11461 1469
rect 11392 1426 11405 1467
rect 11442 1428 11461 1467
rect 11498 1428 11513 1469
rect 11442 1426 11513 1428
rect 11392 1408 11513 1426
rect 10361 1183 10469 1219
rect 10516 1342 10670 1367
rect 10516 1230 10529 1342
rect 10650 1230 10670 1342
rect 8819 893 8985 930
rect 8819 814 8856 893
rect 8940 814 8985 893
rect 8819 776 8985 814
rect 9896 722 9993 1123
rect 10354 1047 10474 1183
rect 10361 1041 10469 1047
rect 9826 693 10001 722
rect 9826 614 9872 693
rect 9972 614 10001 693
rect 9826 589 10001 614
rect 10361 498 10465 1041
rect 10204 468 10475 498
rect 10204 381 10238 468
rect 10308 460 10475 468
rect 10308 381 10371 460
rect 10204 373 10371 381
rect 10441 373 10475 460
rect 10204 327 10475 373
rect 5328 12 10237 30
rect 5328 -34 10139 12
rect 10215 -34 10237 12
rect 5328 -45 10237 -34
rect 10089 -430 10218 -423
rect 10089 -434 10113 -430
rect -74 -489 10113 -434
rect 10144 -489 10175 -430
rect 10206 -489 10218 -430
rect -74 -498 10218 -489
rect 10089 -502 10218 -498
rect 10309 -606 10381 327
rect 10516 256 10670 1230
rect 10514 240 10670 256
rect 10723 1315 10857 1344
rect 10723 1203 10761 1315
rect 10840 1203 10857 1315
rect 10924 1308 11032 1388
rect 10723 250 10857 1203
rect 10925 496 11032 1308
rect 11398 1336 11463 1408
rect 11398 1270 11466 1336
rect 11399 724 11466 1270
rect 12453 908 12518 1795
rect 13496 1525 13633 1529
rect 13483 1521 13640 1525
rect 13483 1414 13520 1521
rect 13620 1414 13640 1521
rect 13483 1372 13640 1414
rect 13496 1124 13633 1372
rect 13486 1082 13652 1124
rect 13486 1007 13515 1082
rect 13632 1007 13652 1082
rect 13486 991 13652 1007
rect 12442 887 12579 908
rect 12442 812 12467 887
rect 12537 812 12579 887
rect 12442 781 12579 812
rect 11385 675 11560 724
rect 11385 596 11418 675
rect 11518 596 11560 675
rect 11385 591 11560 596
rect 10925 454 11073 496
rect 10925 446 10965 454
rect 10927 367 10965 446
rect 11035 367 11073 454
rect 10927 329 11073 367
rect 10514 215 10666 240
rect 10514 120 10544 215
rect 10634 120 10666 215
rect 10514 107 10666 120
rect 10719 214 10858 250
rect 10719 119 10733 214
rect 10823 119 10858 214
rect 10719 101 10858 119
rect 16040 34 16088 3754
rect 16261 3775 16317 3780
rect 16261 3755 16268 3775
rect 16288 3755 16317 3775
rect 16261 3748 16317 3755
rect 16261 3747 16296 3748
rect 16365 3657 16393 6465
rect 19578 6420 19643 6720
rect 19733 6552 19767 6830
rect 20180 6810 20212 6838
rect 19800 6802 20212 6810
rect 19800 6776 19806 6802
rect 19832 6776 20212 6802
rect 20634 6844 20701 6851
rect 20634 6823 20651 6844
rect 20687 6823 20701 6844
rect 20634 6804 20701 6823
rect 20634 6801 20651 6804
rect 19800 6774 20212 6776
rect 19802 6773 19842 6774
rect 19969 6748 20000 6756
rect 19969 6718 19973 6748
rect 19994 6718 20000 6748
rect 19733 6544 19768 6552
rect 19733 6524 19741 6544
rect 19761 6524 19768 6544
rect 19733 6519 19768 6524
rect 19733 6518 19765 6519
rect 19969 6514 20000 6718
rect 20180 6709 20212 6774
rect 20636 6767 20651 6801
rect 20691 6767 20701 6804
rect 20636 6758 20701 6767
rect 20180 6689 20184 6709
rect 20205 6689 20212 6709
rect 20180 6682 20212 6689
rect 20489 6626 20590 6627
rect 20387 6613 20590 6626
rect 20387 6611 20530 6613
rect 20387 6608 20464 6611
rect 20387 6581 20390 6608
rect 20419 6584 20464 6608
rect 20493 6584 20530 6611
rect 20419 6581 20530 6584
rect 20387 6580 20530 6581
rect 20566 6580 20590 6613
rect 20387 6567 20590 6580
rect 19967 6502 20002 6514
rect 19898 6495 20002 6502
rect 19898 6494 19974 6495
rect 19898 6474 19919 6494
rect 19951 6475 19974 6494
rect 19999 6475 20002 6495
rect 19951 6474 20002 6475
rect 19898 6465 20002 6474
rect 19967 6463 20002 6465
rect 19578 6381 19581 6420
rect 19626 6381 19643 6420
rect 20639 6397 20690 6758
rect 20637 6395 20694 6397
rect 19578 6359 19643 6381
rect 20626 6383 20694 6395
rect 20626 6350 20637 6383
rect 20677 6350 20694 6383
rect 20626 6344 20694 6350
rect 20626 6340 20690 6344
rect 19339 6295 19450 6298
rect 21069 6295 21176 6918
rect 17633 6281 21176 6295
rect 17633 6261 19346 6281
rect 19365 6261 19423 6281
rect 19442 6277 21176 6281
rect 19442 6261 20394 6277
rect 17633 6257 20394 6261
rect 20413 6257 20471 6277
rect 20490 6257 21176 6277
rect 17633 6239 21176 6257
rect 17633 6238 18623 6239
rect 20387 6235 20498 6239
rect 18706 6187 18741 6188
rect 18685 6180 18741 6187
rect 18685 6160 18714 6180
rect 18734 6160 18741 6180
rect 18685 6155 18741 6160
rect 19132 6183 19164 6190
rect 19754 6183 19789 6184
rect 19132 6163 19138 6183
rect 19159 6163 19164 6183
rect 19733 6176 19789 6183
rect 19598 6166 19656 6171
rect 18685 5877 18719 6155
rect 19132 6135 19164 6163
rect 18752 6127 19164 6135
rect 18752 6101 18758 6127
rect 18784 6101 19164 6127
rect 18752 6099 19164 6101
rect 18754 6098 18794 6099
rect 18921 6073 18952 6081
rect 18921 6043 18925 6073
rect 18946 6043 18952 6073
rect 18685 5869 18720 5877
rect 18685 5849 18693 5869
rect 18713 5849 18720 5869
rect 18685 5844 18720 5849
rect 18685 5843 18717 5844
rect 18921 5843 18952 6043
rect 19132 6034 19164 6099
rect 19132 6014 19136 6034
rect 19157 6014 19164 6034
rect 19132 6007 19164 6014
rect 19581 6157 19656 6166
rect 19581 6124 19590 6157
rect 19643 6124 19656 6157
rect 19581 6099 19656 6124
rect 19581 6066 19595 6099
rect 19648 6066 19656 6099
rect 19581 6060 19656 6066
rect 19733 6156 19762 6176
rect 19782 6156 19789 6176
rect 19733 6151 19789 6156
rect 20180 6179 20212 6186
rect 20180 6159 20186 6179
rect 20207 6159 20212 6179
rect 19441 5951 19542 5952
rect 19339 5938 19542 5951
rect 19339 5936 19482 5938
rect 19339 5933 19416 5936
rect 19339 5906 19342 5933
rect 19371 5909 19416 5933
rect 19445 5909 19482 5936
rect 19371 5906 19482 5909
rect 19339 5905 19482 5906
rect 19518 5905 19542 5938
rect 19339 5892 19542 5905
rect 18918 5836 18957 5843
rect 18916 5819 18957 5836
rect 18918 5794 18957 5819
rect 17612 5786 18957 5794
rect 17612 5758 17627 5786
rect 17655 5760 18957 5786
rect 17655 5758 18954 5760
rect 17612 5753 18954 5758
rect 19581 5749 19651 6060
rect 19733 5873 19767 6151
rect 20180 6131 20212 6159
rect 19800 6123 20212 6131
rect 19800 6097 19806 6123
rect 19832 6097 20212 6123
rect 19800 6095 20212 6097
rect 19802 6094 19842 6095
rect 19969 6069 20000 6077
rect 19969 6039 19973 6069
rect 19994 6039 20000 6069
rect 19733 5865 19768 5873
rect 19733 5845 19741 5865
rect 19761 5845 19768 5865
rect 19733 5840 19768 5845
rect 19969 5840 20000 6039
rect 20180 6030 20212 6095
rect 20180 6010 20184 6030
rect 20205 6010 20212 6030
rect 20180 6003 20212 6010
rect 20625 6156 20697 6174
rect 20625 6114 20638 6156
rect 20687 6114 20697 6156
rect 20625 6093 20697 6114
rect 20625 6051 20639 6093
rect 20688 6051 20697 6093
rect 20489 5947 20590 5948
rect 20387 5934 20590 5947
rect 20387 5932 20530 5934
rect 20387 5929 20464 5932
rect 20387 5902 20390 5929
rect 20419 5905 20464 5929
rect 20493 5905 20530 5932
rect 20419 5902 20530 5905
rect 20387 5901 20530 5902
rect 20566 5901 20590 5934
rect 20387 5888 20590 5901
rect 19733 5839 19765 5840
rect 19967 5837 20000 5840
rect 19933 5818 20001 5837
rect 19903 5806 20002 5818
rect 20625 5810 20697 6051
rect 21069 5810 21176 6239
rect 19903 5768 19925 5806
rect 19950 5771 19969 5806
rect 19994 5771 20002 5806
rect 19950 5768 20002 5771
rect 19903 5760 20002 5768
rect 19929 5759 20001 5760
rect 19580 5733 19651 5749
rect 19580 5717 19600 5733
rect 19581 5687 19600 5717
rect 19583 5667 19600 5687
rect 19630 5687 19651 5733
rect 20623 5729 20701 5810
rect 21068 5755 21176 5810
rect 19630 5667 19650 5687
rect 19583 5648 19650 5667
rect 20623 5627 20702 5729
rect 20587 5609 20708 5627
rect 20587 5607 20658 5609
rect 20587 5566 20602 5607
rect 20639 5568 20658 5607
rect 20695 5568 20708 5609
rect 20639 5566 20708 5568
rect 20587 5556 20708 5566
rect 17892 5528 18003 5531
rect 17206 5527 18756 5528
rect 21069 5527 21176 5755
rect 17206 5524 20366 5527
rect 20553 5524 21178 5527
rect 17206 5514 21178 5524
rect 17206 5494 17899 5514
rect 17918 5494 17976 5514
rect 17995 5509 21178 5514
rect 17995 5494 20394 5509
rect 17206 5489 20394 5494
rect 20413 5489 20471 5509
rect 20490 5489 21178 5509
rect 17206 5471 21178 5489
rect 17206 5468 18756 5471
rect 20387 5467 20498 5471
rect 17259 5420 17294 5421
rect 17238 5413 17294 5420
rect 17238 5393 17267 5413
rect 17287 5393 17294 5413
rect 17238 5388 17294 5393
rect 17685 5416 17717 5423
rect 17685 5396 17691 5416
rect 17712 5396 17717 5416
rect 17238 5110 17272 5388
rect 17685 5368 17717 5396
rect 19573 5408 19653 5420
rect 19754 5415 19789 5416
rect 17305 5360 17717 5368
rect 17305 5334 17311 5360
rect 17337 5334 17717 5360
rect 18103 5374 18540 5387
rect 18103 5351 18116 5374
rect 18142 5367 18540 5374
rect 18142 5351 18496 5367
rect 18103 5344 18496 5351
rect 18522 5344 18540 5367
rect 18103 5338 18540 5344
rect 19573 5382 19589 5408
rect 19629 5382 19653 5408
rect 19573 5363 19653 5382
rect 17305 5332 17717 5334
rect 17307 5331 17347 5332
rect 17474 5306 17505 5314
rect 17474 5276 17478 5306
rect 17499 5276 17505 5306
rect 17238 5102 17273 5110
rect 17238 5082 17246 5102
rect 17266 5082 17273 5102
rect 17238 5077 17273 5082
rect 17238 5076 17270 5077
rect 17474 5069 17505 5276
rect 17685 5267 17717 5332
rect 19573 5337 19592 5363
rect 19632 5337 19653 5363
rect 19573 5310 19653 5337
rect 19573 5284 19596 5310
rect 19636 5284 19653 5310
rect 19573 5273 19653 5284
rect 19733 5408 19789 5415
rect 19733 5388 19762 5408
rect 19782 5388 19789 5408
rect 19733 5383 19789 5388
rect 20180 5411 20212 5418
rect 20180 5391 20186 5411
rect 20207 5391 20212 5411
rect 17685 5247 17689 5267
rect 17710 5247 17717 5267
rect 17685 5240 17717 5247
rect 17994 5184 18095 5185
rect 17892 5171 18095 5184
rect 17892 5169 18035 5171
rect 17892 5166 17969 5169
rect 17892 5139 17895 5166
rect 17924 5142 17969 5166
rect 17998 5142 18035 5169
rect 17924 5139 18035 5142
rect 17892 5138 18035 5139
rect 18071 5138 18095 5171
rect 17892 5125 18095 5138
rect 17472 5063 17505 5069
rect 17468 5059 17505 5063
rect 17468 5049 17506 5059
rect 17468 5036 17478 5049
rect 17469 5012 17478 5036
rect 17495 5012 17506 5049
rect 17469 4991 17506 5012
rect 19578 4973 19643 5273
rect 19733 5105 19767 5383
rect 20180 5363 20212 5391
rect 19800 5355 20212 5363
rect 19800 5329 19806 5355
rect 19832 5329 20212 5355
rect 20634 5397 20701 5404
rect 20634 5376 20651 5397
rect 20687 5376 20701 5397
rect 20634 5357 20701 5376
rect 20634 5354 20651 5357
rect 19800 5327 20212 5329
rect 19802 5326 19842 5327
rect 19969 5301 20000 5309
rect 19969 5271 19973 5301
rect 19994 5271 20000 5301
rect 19733 5097 19768 5105
rect 19733 5077 19741 5097
rect 19761 5077 19768 5097
rect 19733 5072 19768 5077
rect 19733 5071 19765 5072
rect 19969 5067 20000 5271
rect 20180 5262 20212 5327
rect 20636 5320 20651 5354
rect 20691 5320 20701 5357
rect 20636 5311 20701 5320
rect 20180 5242 20184 5262
rect 20205 5242 20212 5262
rect 20180 5235 20212 5242
rect 20489 5179 20590 5180
rect 20387 5166 20590 5179
rect 20387 5164 20530 5166
rect 20387 5161 20464 5164
rect 20387 5134 20390 5161
rect 20419 5137 20464 5161
rect 20493 5137 20530 5164
rect 20419 5134 20530 5137
rect 20387 5133 20530 5134
rect 20566 5133 20590 5166
rect 20387 5120 20590 5133
rect 19967 5055 20002 5067
rect 19898 5048 20002 5055
rect 19898 5047 19974 5048
rect 19898 5027 19919 5047
rect 19951 5028 19974 5047
rect 19999 5028 20002 5048
rect 19951 5027 20002 5028
rect 19898 5018 20002 5027
rect 19967 5016 20002 5018
rect 19578 4934 19581 4973
rect 19626 4934 19643 4973
rect 20639 4950 20690 5311
rect 20637 4948 20694 4950
rect 19578 4912 19643 4934
rect 20626 4936 20694 4948
rect 20626 4903 20637 4936
rect 20677 4903 20694 4936
rect 20626 4897 20694 4903
rect 20626 4893 20690 4897
rect 19339 4848 19450 4851
rect 21069 4848 21176 5471
rect 17415 4834 21176 4848
rect 17415 4814 19346 4834
rect 19365 4814 19423 4834
rect 19442 4830 21176 4834
rect 19442 4814 20394 4830
rect 17415 4810 20394 4814
rect 20413 4810 20471 4830
rect 20490 4810 21176 4830
rect 17415 4792 21176 4810
rect 17415 4791 18715 4792
rect 20387 4788 20498 4792
rect 18706 4740 18741 4741
rect 18685 4733 18741 4740
rect 18685 4713 18714 4733
rect 18734 4713 18741 4733
rect 18685 4708 18741 4713
rect 19132 4736 19164 4743
rect 19754 4736 19789 4737
rect 19132 4716 19138 4736
rect 19159 4716 19164 4736
rect 19733 4729 19789 4736
rect 19598 4719 19656 4724
rect 18685 4430 18719 4708
rect 19132 4688 19164 4716
rect 18752 4680 19164 4688
rect 18752 4654 18758 4680
rect 18784 4654 19164 4680
rect 18752 4652 19164 4654
rect 18754 4651 18794 4652
rect 18921 4626 18952 4634
rect 18921 4596 18925 4626
rect 18946 4596 18952 4626
rect 18685 4422 18720 4430
rect 18685 4402 18693 4422
rect 18713 4402 18720 4422
rect 18685 4397 18720 4402
rect 18685 4396 18717 4397
rect 18921 4389 18952 4596
rect 19132 4587 19164 4652
rect 19132 4567 19136 4587
rect 19157 4567 19164 4587
rect 19132 4560 19164 4567
rect 19581 4710 19656 4719
rect 19581 4677 19590 4710
rect 19643 4677 19656 4710
rect 19581 4652 19656 4677
rect 19581 4619 19595 4652
rect 19648 4619 19656 4652
rect 19581 4613 19656 4619
rect 19733 4709 19762 4729
rect 19782 4709 19789 4729
rect 19733 4704 19789 4709
rect 20180 4732 20212 4739
rect 20180 4712 20186 4732
rect 20207 4712 20212 4732
rect 19441 4504 19542 4505
rect 19339 4491 19542 4504
rect 19339 4489 19482 4491
rect 19339 4486 19416 4489
rect 19339 4459 19342 4486
rect 19371 4462 19416 4486
rect 19445 4462 19482 4489
rect 19371 4459 19482 4462
rect 19339 4458 19482 4459
rect 19518 4458 19542 4491
rect 19339 4445 19542 4458
rect 18419 4376 18583 4379
rect 18916 4376 18952 4389
rect 17618 4358 18957 4376
rect 17618 4320 17628 4358
rect 17653 4343 18957 4358
rect 17653 4320 17663 4343
rect 18419 4336 18583 4343
rect 17618 4312 17663 4320
rect 17632 4311 17663 4312
rect 19581 4297 19651 4613
rect 19733 4426 19767 4704
rect 20180 4684 20212 4712
rect 19800 4676 20212 4684
rect 19800 4650 19806 4676
rect 19832 4650 20212 4676
rect 19800 4648 20212 4650
rect 19802 4647 19842 4648
rect 19969 4622 20000 4630
rect 19969 4592 19973 4622
rect 19994 4592 20000 4622
rect 19733 4418 19768 4426
rect 19733 4398 19741 4418
rect 19761 4398 19768 4418
rect 19733 4393 19768 4398
rect 19969 4393 20000 4592
rect 20180 4583 20212 4648
rect 20180 4563 20184 4583
rect 20205 4563 20212 4583
rect 20180 4556 20212 4563
rect 20625 4709 20697 4727
rect 20625 4667 20638 4709
rect 20687 4667 20697 4709
rect 20625 4646 20697 4667
rect 20625 4604 20639 4646
rect 20688 4604 20697 4646
rect 20489 4500 20590 4501
rect 20387 4487 20590 4500
rect 20387 4485 20530 4487
rect 20387 4482 20464 4485
rect 20387 4455 20390 4482
rect 20419 4458 20464 4482
rect 20493 4458 20530 4485
rect 20419 4455 20530 4458
rect 20387 4454 20530 4455
rect 20566 4454 20590 4487
rect 20387 4441 20590 4454
rect 19733 4392 19765 4393
rect 19967 4390 20000 4393
rect 19933 4371 20001 4390
rect 19903 4359 20002 4371
rect 19903 4321 19925 4359
rect 19950 4324 19969 4359
rect 19994 4324 20002 4359
rect 19950 4321 20002 4324
rect 19903 4313 20002 4321
rect 19929 4312 20001 4313
rect 19581 4278 19660 4297
rect 19584 4258 19660 4278
rect 19577 4234 19660 4258
rect 20625 4293 20697 4604
rect 20625 4250 20701 4293
rect 19577 4168 19589 4234
rect 19643 4168 19660 4234
rect 19577 4148 19660 4168
rect 19577 4111 19594 4148
rect 19638 4134 19660 4148
rect 20626 4199 20701 4250
rect 21069 4199 21176 4792
rect 19638 4111 19653 4134
rect 19577 4095 19653 4111
rect 20626 4107 20703 4199
rect 21069 4195 21177 4199
rect 20588 4089 20709 4107
rect 20588 4087 20659 4089
rect 20588 4046 20603 4087
rect 20640 4048 20659 4087
rect 20696 4048 20709 4089
rect 20640 4046 20709 4048
rect 20588 4036 20709 4046
rect 17159 4007 18582 4009
rect 21070 4007 21177 4195
rect 17159 3992 21179 4007
rect 17159 3972 17857 3992
rect 17876 3972 17934 3992
rect 17953 3989 21179 3992
rect 17953 3972 20395 3989
rect 17159 3969 20395 3972
rect 20414 3969 20472 3989
rect 20491 3969 21179 3989
rect 17159 3951 21179 3969
rect 17850 3950 17961 3951
rect 18537 3950 18744 3951
rect 20388 3947 20499 3951
rect 17217 3898 17252 3899
rect 17196 3891 17252 3898
rect 17196 3871 17225 3891
rect 17245 3871 17252 3891
rect 17196 3866 17252 3871
rect 17643 3894 17675 3901
rect 17643 3874 17649 3894
rect 17670 3874 17675 3894
rect 16365 3642 16391 3657
rect 16362 3635 16398 3642
rect 16362 3597 16368 3635
rect 16391 3597 16398 3635
rect 16362 3591 16398 3597
rect 17196 3588 17230 3866
rect 17643 3846 17675 3874
rect 17263 3838 17675 3846
rect 17263 3812 17269 3838
rect 17295 3812 17675 3838
rect 17263 3810 17675 3812
rect 17265 3809 17305 3810
rect 17432 3784 17463 3792
rect 17432 3754 17436 3784
rect 17457 3754 17463 3784
rect 17196 3580 17231 3588
rect 17196 3560 17204 3580
rect 17224 3560 17231 3580
rect 17196 3555 17231 3560
rect 17196 3554 17228 3555
rect 17432 3551 17463 3754
rect 17643 3745 17675 3810
rect 19574 3888 19654 3900
rect 19755 3895 19790 3896
rect 19574 3862 19590 3888
rect 19630 3862 19654 3888
rect 19574 3843 19654 3862
rect 19574 3817 19593 3843
rect 19633 3817 19654 3843
rect 19574 3790 19654 3817
rect 19574 3764 19597 3790
rect 19637 3764 19654 3790
rect 19574 3753 19654 3764
rect 19734 3888 19790 3895
rect 19734 3868 19763 3888
rect 19783 3868 19790 3888
rect 19734 3863 19790 3868
rect 20181 3891 20213 3898
rect 20181 3871 20187 3891
rect 20208 3871 20213 3891
rect 17643 3725 17647 3745
rect 17668 3725 17675 3745
rect 17643 3718 17675 3725
rect 17952 3662 18053 3663
rect 17850 3649 18053 3662
rect 17850 3647 17993 3649
rect 17850 3644 17927 3647
rect 17850 3617 17853 3644
rect 17882 3620 17927 3644
rect 17956 3620 17993 3647
rect 17882 3617 17993 3620
rect 17850 3616 17993 3617
rect 18029 3616 18053 3649
rect 17850 3603 18053 3616
rect 17427 3533 17463 3551
rect 17427 3516 17462 3533
rect 17360 3485 17465 3516
rect 17360 3480 17432 3485
rect 17360 3459 17391 3480
rect 17411 3464 17432 3480
rect 17452 3464 17465 3485
rect 17411 3459 17465 3464
rect 17360 3450 17465 3459
rect 19579 3453 19644 3753
rect 19734 3585 19768 3863
rect 20181 3843 20213 3871
rect 19801 3835 20213 3843
rect 19801 3809 19807 3835
rect 19833 3809 20213 3835
rect 20635 3877 20702 3884
rect 20635 3856 20652 3877
rect 20688 3856 20702 3877
rect 20635 3837 20702 3856
rect 20635 3834 20652 3837
rect 19801 3807 20213 3809
rect 19803 3806 19843 3807
rect 19970 3781 20001 3789
rect 19970 3751 19974 3781
rect 19995 3751 20001 3781
rect 19734 3577 19769 3585
rect 19734 3557 19742 3577
rect 19762 3557 19769 3577
rect 19734 3552 19769 3557
rect 19734 3551 19766 3552
rect 19970 3547 20001 3751
rect 20181 3742 20213 3807
rect 20637 3800 20652 3834
rect 20692 3800 20702 3837
rect 20637 3791 20702 3800
rect 20181 3722 20185 3742
rect 20206 3722 20213 3742
rect 20181 3715 20213 3722
rect 20490 3659 20591 3660
rect 20388 3646 20591 3659
rect 20388 3644 20531 3646
rect 20388 3641 20465 3644
rect 20388 3614 20391 3641
rect 20420 3617 20465 3641
rect 20494 3617 20531 3644
rect 20420 3614 20531 3617
rect 20388 3613 20531 3614
rect 20567 3613 20591 3646
rect 20388 3600 20591 3613
rect 19968 3535 20003 3547
rect 19899 3528 20003 3535
rect 19899 3527 19975 3528
rect 19899 3507 19920 3527
rect 19952 3508 19975 3527
rect 20000 3508 20003 3528
rect 19952 3507 20003 3508
rect 19899 3498 20003 3507
rect 19968 3496 20003 3498
rect 19579 3414 19582 3453
rect 19627 3414 19644 3453
rect 20640 3430 20691 3791
rect 20638 3428 20695 3430
rect 19579 3392 19644 3414
rect 20627 3416 20695 3428
rect 20627 3383 20638 3416
rect 20678 3383 20695 3416
rect 20627 3377 20695 3383
rect 20627 3373 20691 3377
rect 19340 3328 19451 3331
rect 21070 3328 21177 3951
rect 17383 3314 21177 3328
rect 17383 3294 19347 3314
rect 19366 3294 19424 3314
rect 19443 3310 21177 3314
rect 19443 3294 20395 3310
rect 17383 3290 20395 3294
rect 20414 3290 20472 3310
rect 20491 3290 21177 3310
rect 17383 3272 21177 3290
rect 17383 3271 18624 3272
rect 20388 3268 20499 3272
rect 18707 3220 18742 3221
rect 18686 3213 18742 3220
rect 18686 3193 18715 3213
rect 18735 3193 18742 3213
rect 18686 3188 18742 3193
rect 19133 3216 19165 3223
rect 19755 3216 19790 3217
rect 19133 3196 19139 3216
rect 19160 3196 19165 3216
rect 19734 3209 19790 3216
rect 19599 3199 19657 3204
rect 18686 2910 18720 3188
rect 19133 3168 19165 3196
rect 18753 3160 19165 3168
rect 18753 3134 18759 3160
rect 18785 3134 19165 3160
rect 18753 3132 19165 3134
rect 18755 3131 18795 3132
rect 18922 3106 18953 3114
rect 18922 3076 18926 3106
rect 18947 3076 18953 3106
rect 18686 2902 18721 2910
rect 18686 2882 18694 2902
rect 18714 2882 18721 2902
rect 18686 2877 18721 2882
rect 17427 2866 17463 2877
rect 18686 2876 18718 2877
rect 18922 2869 18953 3076
rect 19133 3067 19165 3132
rect 19133 3047 19137 3067
rect 19158 3047 19165 3067
rect 19133 3040 19165 3047
rect 19582 3190 19657 3199
rect 19582 3157 19591 3190
rect 19644 3157 19657 3190
rect 19582 3132 19657 3157
rect 19582 3099 19596 3132
rect 19649 3099 19657 3132
rect 19582 3093 19657 3099
rect 19734 3189 19763 3209
rect 19783 3189 19790 3209
rect 19734 3184 19790 3189
rect 20181 3212 20213 3219
rect 20181 3192 20187 3212
rect 20208 3192 20213 3212
rect 19442 2984 19543 2985
rect 19340 2971 19543 2984
rect 19340 2969 19483 2971
rect 19340 2966 19417 2969
rect 19340 2939 19343 2966
rect 19372 2942 19417 2966
rect 19446 2942 19483 2969
rect 19372 2939 19483 2942
rect 19340 2938 19483 2939
rect 19519 2938 19543 2971
rect 19340 2925 19543 2938
rect 17427 2843 17433 2866
rect 17457 2843 17463 2866
rect 18917 2860 18953 2869
rect 18862 2850 18959 2860
rect 17674 2848 18959 2850
rect 17427 2822 17463 2843
rect 17427 2799 17433 2822
rect 17457 2799 17463 2822
rect 17427 2646 17463 2799
rect 17639 2838 18959 2848
rect 17639 2800 17651 2838
rect 17676 2803 17695 2838
rect 17720 2803 18959 2838
rect 17676 2800 18959 2803
rect 17639 2797 18959 2800
rect 17639 2795 18956 2797
rect 17639 2792 17728 2795
rect 17655 2791 17727 2792
rect 19582 2782 19652 3093
rect 19734 2906 19768 3184
rect 20181 3164 20213 3192
rect 19801 3156 20213 3164
rect 19801 3130 19807 3156
rect 19833 3130 20213 3156
rect 19801 3128 20213 3130
rect 19803 3127 19843 3128
rect 19970 3102 20001 3110
rect 19970 3072 19974 3102
rect 19995 3072 20001 3102
rect 19734 2898 19769 2906
rect 19734 2878 19742 2898
rect 19762 2878 19769 2898
rect 19734 2873 19769 2878
rect 19970 2873 20001 3072
rect 20181 3063 20213 3128
rect 20181 3043 20185 3063
rect 20206 3043 20213 3063
rect 20181 3036 20213 3043
rect 20626 3189 20698 3207
rect 20626 3147 20639 3189
rect 20688 3147 20698 3189
rect 20626 3126 20698 3147
rect 20626 3084 20640 3126
rect 20689 3084 20698 3126
rect 20490 2980 20591 2981
rect 20388 2967 20591 2980
rect 20388 2965 20531 2967
rect 20388 2962 20465 2965
rect 20388 2935 20391 2962
rect 20420 2938 20465 2962
rect 20494 2938 20531 2965
rect 20420 2935 20531 2938
rect 20388 2934 20531 2935
rect 20567 2934 20591 2967
rect 20388 2921 20591 2934
rect 19734 2872 19766 2873
rect 19968 2870 20001 2873
rect 19934 2851 20002 2870
rect 19904 2839 20003 2851
rect 20626 2843 20698 3084
rect 21070 2843 21177 3272
rect 19904 2801 19926 2839
rect 19951 2804 19970 2839
rect 19995 2804 20003 2839
rect 19951 2801 20003 2804
rect 19904 2793 20003 2801
rect 19930 2792 20002 2793
rect 19581 2766 19652 2782
rect 19581 2750 19601 2766
rect 19582 2720 19601 2750
rect 19584 2700 19601 2720
rect 19631 2720 19652 2766
rect 20624 2762 20702 2843
rect 21069 2788 21177 2843
rect 19631 2700 19651 2720
rect 19584 2681 19651 2700
rect 20624 2660 20703 2762
rect 17418 2637 17504 2646
rect 17418 2619 17437 2637
rect 17489 2619 17504 2637
rect 17418 2615 17504 2619
rect 20588 2642 20709 2660
rect 20588 2640 20659 2642
rect 20588 2599 20603 2640
rect 20640 2601 20659 2640
rect 20696 2601 20709 2642
rect 20640 2599 20709 2601
rect 20588 2589 20709 2599
rect 17893 2561 18004 2564
rect 17208 2560 18757 2561
rect 21070 2560 21177 2788
rect 17208 2557 20367 2560
rect 20554 2557 21179 2560
rect 17208 2547 21179 2557
rect 17208 2527 17900 2547
rect 17919 2527 17977 2547
rect 17996 2542 21179 2547
rect 17996 2527 20395 2542
rect 17208 2522 20395 2527
rect 20414 2522 20472 2542
rect 20491 2522 21179 2542
rect 17208 2504 21179 2522
rect 17208 2501 18757 2504
rect 20388 2500 20499 2504
rect 17260 2453 17295 2454
rect 17239 2446 17295 2453
rect 17239 2426 17268 2446
rect 17288 2426 17295 2446
rect 17239 2421 17295 2426
rect 17686 2449 17718 2456
rect 17686 2429 17692 2449
rect 17713 2429 17718 2449
rect 17239 2143 17273 2421
rect 17686 2401 17718 2429
rect 17306 2393 17718 2401
rect 17306 2367 17312 2393
rect 17338 2367 17718 2393
rect 17306 2365 17718 2367
rect 17308 2364 17348 2365
rect 17475 2339 17506 2347
rect 17475 2309 17479 2339
rect 17500 2309 17506 2339
rect 17239 2135 17274 2143
rect 17239 2115 17247 2135
rect 17267 2115 17274 2135
rect 17239 2110 17274 2115
rect 17239 2109 17271 2110
rect 17475 2108 17506 2309
rect 17686 2300 17718 2365
rect 17686 2280 17690 2300
rect 17711 2280 17718 2300
rect 17686 2273 17718 2280
rect 18280 2440 18373 2447
rect 18280 2399 18304 2440
rect 18358 2399 18373 2440
rect 17995 2217 18096 2218
rect 17893 2204 18096 2217
rect 17893 2202 18036 2204
rect 17893 2199 17970 2202
rect 17893 2172 17896 2199
rect 17925 2175 17970 2199
rect 17999 2175 18036 2202
rect 17925 2172 18036 2175
rect 17893 2171 18036 2172
rect 18072 2171 18096 2204
rect 17893 2158 18096 2171
rect 18280 2026 18373 2399
rect 19574 2441 19654 2453
rect 19755 2448 19790 2449
rect 19574 2415 19590 2441
rect 19630 2415 19654 2441
rect 19574 2396 19654 2415
rect 19574 2370 19593 2396
rect 19633 2370 19654 2396
rect 19574 2343 19654 2370
rect 19574 2317 19597 2343
rect 19637 2317 19654 2343
rect 19574 2306 19654 2317
rect 19734 2441 19790 2448
rect 19734 2421 19763 2441
rect 19783 2421 19790 2441
rect 19734 2416 19790 2421
rect 20181 2444 20213 2451
rect 20181 2424 20187 2444
rect 20208 2424 20213 2444
rect 18280 1982 18298 2026
rect 18358 1982 18373 2026
rect 18280 1967 18373 1982
rect 19579 2006 19644 2306
rect 19734 2138 19768 2416
rect 20181 2396 20213 2424
rect 19801 2388 20213 2396
rect 19801 2362 19807 2388
rect 19833 2362 20213 2388
rect 20635 2430 20702 2437
rect 20635 2409 20652 2430
rect 20688 2409 20702 2430
rect 20635 2390 20702 2409
rect 20635 2387 20652 2390
rect 19801 2360 20213 2362
rect 19803 2359 19843 2360
rect 19970 2334 20001 2342
rect 19970 2304 19974 2334
rect 19995 2304 20001 2334
rect 19734 2130 19769 2138
rect 19734 2110 19742 2130
rect 19762 2110 19769 2130
rect 19734 2105 19769 2110
rect 19734 2104 19766 2105
rect 19970 2100 20001 2304
rect 20181 2295 20213 2360
rect 20637 2353 20652 2387
rect 20692 2353 20702 2390
rect 20637 2344 20702 2353
rect 20181 2275 20185 2295
rect 20206 2275 20213 2295
rect 20181 2268 20213 2275
rect 20490 2212 20591 2213
rect 20388 2199 20591 2212
rect 20388 2197 20531 2199
rect 20388 2194 20465 2197
rect 20388 2167 20391 2194
rect 20420 2170 20465 2194
rect 20494 2170 20531 2197
rect 20420 2167 20531 2170
rect 20388 2166 20531 2167
rect 20567 2166 20591 2199
rect 20388 2153 20591 2166
rect 19968 2088 20003 2100
rect 19899 2081 20003 2088
rect 19899 2080 19975 2081
rect 19899 2060 19920 2080
rect 19952 2061 19975 2080
rect 20000 2061 20003 2081
rect 19952 2060 20003 2061
rect 19899 2051 20003 2060
rect 19968 2049 20003 2051
rect 19579 1967 19582 2006
rect 19627 1967 19644 2006
rect 20640 1983 20691 2344
rect 20638 1981 20695 1983
rect 19579 1945 19644 1967
rect 20627 1969 20695 1981
rect 20627 1936 20638 1969
rect 20678 1936 20695 1969
rect 20627 1930 20695 1936
rect 20627 1926 20691 1930
rect 19340 1881 19451 1884
rect 21070 1881 21177 2504
rect 17603 1867 21177 1881
rect 17603 1847 19347 1867
rect 19366 1847 19424 1867
rect 19443 1863 21177 1867
rect 19443 1847 20395 1863
rect 17603 1843 20395 1847
rect 20414 1843 20472 1863
rect 20491 1843 21177 1863
rect 17603 1825 21177 1843
rect 17603 1824 18716 1825
rect 20388 1821 20499 1825
rect 18707 1773 18742 1774
rect 18686 1766 18742 1773
rect 18686 1746 18715 1766
rect 18735 1746 18742 1766
rect 18686 1741 18742 1746
rect 19133 1769 19165 1776
rect 19755 1769 19790 1770
rect 19133 1749 19139 1769
rect 19160 1749 19165 1769
rect 19734 1762 19790 1769
rect 19599 1752 19657 1757
rect 16522 1706 18375 1739
rect 16522 1641 16587 1706
rect 16718 1686 18375 1706
rect 16718 1645 18311 1686
rect 18347 1645 18375 1686
rect 18473 1706 18537 1725
rect 18473 1667 18490 1706
rect 18524 1667 18537 1706
rect 18473 1648 18537 1667
rect 16718 1641 18375 1645
rect 16522 1616 18375 1641
rect 18286 1613 18368 1616
rect 18475 1136 18537 1648
rect 18686 1463 18720 1741
rect 19133 1721 19165 1749
rect 18753 1713 19165 1721
rect 18753 1687 18759 1713
rect 18785 1687 19165 1713
rect 18753 1685 19165 1687
rect 18755 1684 18795 1685
rect 18922 1659 18953 1667
rect 18922 1629 18926 1659
rect 18947 1629 18953 1659
rect 18686 1455 18721 1463
rect 18686 1435 18694 1455
rect 18714 1435 18721 1455
rect 18686 1430 18721 1435
rect 18686 1429 18718 1430
rect 18922 1422 18953 1629
rect 19133 1620 19165 1685
rect 19133 1600 19137 1620
rect 19158 1600 19165 1620
rect 19133 1593 19165 1600
rect 19582 1743 19657 1752
rect 19582 1710 19591 1743
rect 19644 1710 19657 1743
rect 19582 1685 19657 1710
rect 19582 1652 19596 1685
rect 19649 1652 19657 1685
rect 19582 1646 19657 1652
rect 19734 1742 19763 1762
rect 19783 1742 19790 1762
rect 19734 1737 19790 1742
rect 20181 1765 20213 1772
rect 20181 1745 20187 1765
rect 20208 1745 20213 1765
rect 19442 1537 19543 1538
rect 19340 1524 19543 1537
rect 19340 1522 19483 1524
rect 19340 1519 19417 1522
rect 19340 1492 19343 1519
rect 19372 1495 19417 1519
rect 19446 1495 19483 1522
rect 19372 1492 19483 1495
rect 19340 1491 19483 1492
rect 19519 1491 19543 1524
rect 19340 1478 19543 1491
rect 18917 1404 18953 1422
rect 18884 1403 18953 1404
rect 18864 1391 18953 1403
rect 18864 1353 18876 1391
rect 18901 1356 18920 1391
rect 18945 1356 18953 1391
rect 18901 1353 18953 1356
rect 18864 1345 18953 1353
rect 18880 1344 18952 1345
rect 18433 1078 18549 1136
rect 19582 1125 19652 1646
rect 19734 1459 19768 1737
rect 20181 1717 20213 1745
rect 19801 1709 20213 1717
rect 19801 1683 19807 1709
rect 19833 1683 20213 1709
rect 19801 1681 20213 1683
rect 19803 1680 19843 1681
rect 19970 1655 20001 1663
rect 19970 1625 19974 1655
rect 19995 1625 20001 1655
rect 19734 1451 19769 1459
rect 19734 1431 19742 1451
rect 19762 1431 19769 1451
rect 19734 1426 19769 1431
rect 19970 1426 20001 1625
rect 20181 1616 20213 1681
rect 20181 1596 20185 1616
rect 20206 1596 20213 1616
rect 20181 1589 20213 1596
rect 20626 1742 20698 1760
rect 20626 1700 20639 1742
rect 20688 1700 20698 1742
rect 20626 1679 20698 1700
rect 20626 1637 20640 1679
rect 20689 1637 20698 1679
rect 20490 1533 20591 1534
rect 20388 1520 20591 1533
rect 20388 1518 20531 1520
rect 20388 1515 20465 1518
rect 20388 1488 20391 1515
rect 20420 1491 20465 1515
rect 20494 1491 20531 1518
rect 20420 1488 20531 1491
rect 20388 1487 20531 1488
rect 20567 1487 20591 1520
rect 20388 1474 20591 1487
rect 19734 1425 19766 1426
rect 19968 1423 20001 1426
rect 19934 1404 20002 1423
rect 19904 1392 20003 1404
rect 19904 1354 19926 1392
rect 19951 1357 19970 1392
rect 19995 1357 20003 1392
rect 19951 1354 20003 1357
rect 19904 1346 20003 1354
rect 19930 1345 20002 1346
rect 18433 1007 18445 1078
rect 18524 1007 18549 1078
rect 18433 987 18549 1007
rect 19563 924 19665 1125
rect 20626 1117 20698 1637
rect 21070 1213 21177 1825
rect 21069 1177 21177 1213
rect 21224 1336 21378 1361
rect 21224 1224 21237 1336
rect 21358 1224 21378 1336
rect 19527 887 19693 924
rect 19527 808 19564 887
rect 19648 808 19693 887
rect 19527 770 19693 808
rect 20604 716 20701 1117
rect 21062 1041 21182 1177
rect 21069 1035 21177 1041
rect 20534 687 20709 716
rect 20534 608 20580 687
rect 20680 608 20709 687
rect 20534 583 20709 608
rect 21069 492 21173 1035
rect 20912 462 21183 492
rect 20912 375 20946 462
rect 21016 454 21183 462
rect 21016 375 21079 454
rect 20912 367 21079 375
rect 21149 367 21183 454
rect 20912 321 21183 367
rect 21224 250 21378 1224
rect 21222 234 21378 250
rect 21222 209 21374 234
rect 21222 114 21252 209
rect 21342 114 21374 209
rect 21222 101 21374 114
rect 16040 -6 16092 34
rect 16042 -53 16092 -6
rect 11586 -64 16092 -53
rect 11586 -112 11601 -64
rect 11642 -112 16092 -64
rect 11586 -117 16092 -112
rect 11586 -132 11651 -117
rect 16042 -123 16092 -117
rect 10513 -251 10716 -238
rect 10513 -284 10537 -251
rect 10573 -252 10716 -251
rect 10573 -255 10684 -252
rect 10573 -282 10610 -255
rect 10639 -279 10684 -255
rect 10713 -279 10716 -252
rect 10639 -282 10716 -279
rect 10573 -284 10716 -282
rect 10513 -297 10716 -284
rect 10513 -298 10614 -297
rect 10891 -360 10923 -353
rect 10891 -380 10898 -360
rect 10919 -380 10923 -360
rect 10891 -445 10923 -380
rect 11103 -389 11134 -163
rect 11338 -190 11370 -189
rect 11335 -195 11370 -190
rect 11335 -215 11342 -195
rect 11362 -215 11370 -195
rect 11335 -223 11370 -215
rect 11103 -419 11109 -389
rect 11130 -419 11134 -389
rect 11103 -427 11134 -419
rect 11261 -445 11301 -444
rect 10891 -447 11303 -445
rect 10891 -473 11271 -447
rect 11297 -473 11303 -447
rect 10891 -481 11303 -473
rect 10891 -509 10923 -481
rect 11336 -501 11370 -223
rect 10891 -529 10896 -509
rect 10917 -529 10923 -509
rect 10891 -536 10923 -529
rect 11102 -508 11135 -501
rect 11102 -531 11110 -508
rect 11130 -531 11135 -508
rect 10605 -606 10716 -585
rect 10309 -607 10716 -606
rect 10309 -627 10613 -607
rect 10632 -627 10690 -607
rect 10709 -627 10716 -607
rect 10309 -644 10716 -627
rect 10309 -678 10710 -644
rect 11102 -763 11135 -531
rect 11314 -506 11370 -501
rect 11314 -526 11321 -506
rect 11341 -526 11370 -506
rect 11314 -533 11370 -526
rect 11314 -534 11349 -533
<< via1 >>
rect 827 12976 863 13009
rect 1875 12972 1911 13005
rect 5350 13473 5428 13531
rect 4287 13351 4353 13406
rect 3025 13222 3095 13295
rect 827 12297 863 12330
rect 3322 12292 3358 12325
rect 827 11529 863 11562
rect 1875 11525 1911 11558
rect 827 10850 863 10883
rect 3365 10847 3401 10880
rect 828 10009 864 10042
rect 1876 10005 1912 10038
rect 828 9330 864 9363
rect 3323 9325 3359 9358
rect 828 8562 864 8595
rect 1876 8558 1912 8591
rect 828 7883 864 7916
rect 16069 13470 16147 13528
rect 15009 13345 15061 13389
rect 13748 13221 13800 13271
rect 9824 12594 9860 12627
rect 4431 7874 4467 7907
rect 825 6968 861 7001
rect 1873 6964 1909 6997
rect 825 6289 861 6322
rect 3320 6284 3356 6317
rect 825 5521 861 5554
rect 1873 5517 1909 5550
rect 8776 11919 8812 11952
rect 9824 11915 9860 11948
rect 11535 12970 11571 13003
rect 12583 12966 12619 12999
rect 11535 12291 11571 12324
rect 14030 12286 14066 12319
rect 7329 11152 7365 11185
rect 9824 11147 9860 11180
rect 8776 10472 8812 10505
rect 9824 10468 9860 10501
rect 11535 11523 11571 11556
rect 12583 11519 12619 11552
rect 11535 10844 11571 10877
rect 14073 10841 14109 10874
rect 7287 9630 7323 9663
rect 9825 9627 9861 9660
rect 8777 8952 8813 8985
rect 9825 8948 9861 8981
rect 11536 10003 11572 10036
rect 12584 9999 12620 10032
rect 11536 9324 11572 9357
rect 14031 9319 14067 9352
rect 7330 8185 7366 8218
rect 9825 8180 9861 8213
rect 8777 7505 8813 7538
rect 9825 7501 9861 7534
rect 11536 8556 11572 8589
rect 12584 8552 12620 8585
rect 11536 7877 11572 7910
rect 20532 12588 20568 12621
rect 15139 7868 15175 7901
rect 6219 6595 6255 6628
rect 825 4842 861 4875
rect 3363 4839 3399 4872
rect 826 4001 862 4034
rect 1874 3997 1910 4030
rect 4776 4003 4812 4036
rect 826 3322 862 3355
rect 3321 3317 3357 3350
rect 826 2554 862 2587
rect 1874 2550 1910 2583
rect 826 1875 862 1908
rect 53 1209 132 1321
rect 2807 1013 2924 1088
rect 1759 818 1829 893
rect 710 602 810 681
rect 257 373 327 460
rect 25 125 115 220
rect 9822 6586 9858 6619
rect 8774 5911 8810 5944
rect 9822 5907 9858 5940
rect 11533 6962 11569 6995
rect 12581 6958 12617 6991
rect 11533 6283 11569 6316
rect 14028 6278 14064 6311
rect 7327 5144 7363 5177
rect 9822 5139 9858 5172
rect 8774 4464 8810 4497
rect 9822 4460 9858 4493
rect 11533 5515 11569 5548
rect 12581 5511 12617 5544
rect 19484 11913 19520 11946
rect 20532 11909 20568 11942
rect 18037 11146 18073 11179
rect 20532 11141 20568 11174
rect 19484 10466 19520 10499
rect 20532 10462 20568 10495
rect 17995 9624 18031 9657
rect 20533 9621 20569 9654
rect 19485 8946 19521 8979
rect 20533 8942 20569 8975
rect 18038 8179 18074 8212
rect 20533 8174 20569 8207
rect 19485 7499 19521 7532
rect 20533 7495 20569 7528
rect 16927 6589 16963 6622
rect 11533 4836 11569 4869
rect 14071 4833 14107 4866
rect 7285 3622 7321 3655
rect 9823 3619 9859 3652
rect 8775 2944 8811 2977
rect 9823 2940 9859 2973
rect 11534 3995 11570 4028
rect 12582 3991 12618 4024
rect 15484 3997 15520 4030
rect 11534 3316 11570 3349
rect 14029 3311 14065 3344
rect 7328 2177 7364 2210
rect 9823 2172 9859 2205
rect 8775 1497 8811 1530
rect 9823 1493 9859 1526
rect 7737 1013 7816 1084
rect 11534 2548 11570 2581
rect 12582 2544 12618 2577
rect 11534 1869 11570 1902
rect 10529 1230 10650 1342
rect 8856 814 8940 893
rect 9872 614 9972 693
rect 10238 381 10308 468
rect 10371 373 10441 460
rect 10761 1203 10840 1315
rect 13515 1007 13632 1082
rect 12467 812 12537 887
rect 11418 596 11518 675
rect 10965 367 11035 454
rect 10544 120 10634 215
rect 10733 119 10823 214
rect 20530 6580 20566 6613
rect 19482 5905 19518 5938
rect 20530 5901 20566 5934
rect 18035 5138 18071 5171
rect 20530 5133 20566 5166
rect 19482 4458 19518 4491
rect 20530 4454 20566 4487
rect 17993 3616 18029 3649
rect 20531 3613 20567 3646
rect 19483 2938 19519 2971
rect 20531 2934 20567 2967
rect 18036 2171 18072 2204
rect 20531 2166 20567 2199
rect 19483 1491 19519 1524
rect 20531 1487 20567 1520
rect 18445 1007 18524 1078
rect 21237 1224 21358 1336
rect 19564 808 19648 887
rect 20580 608 20680 687
rect 20946 375 21016 462
rect 21079 367 21149 454
rect 21252 114 21342 209
rect 10537 -284 10573 -251
<< metal2 >>
rect 16052 13545 16160 13548
rect 5319 13531 16160 13545
rect 5319 13473 5350 13531
rect 5428 13528 16160 13531
rect 5428 13473 16069 13528
rect 5319 13470 16069 13473
rect 16147 13470 16160 13528
rect 5319 13458 16160 13470
rect 46 13024 153 13458
rect 16052 13457 16160 13458
rect 4271 13406 4370 13417
rect 4271 13351 4287 13406
rect 4353 13393 4370 13406
rect 14992 13393 15079 13407
rect 4353 13389 15079 13393
rect 4353 13351 15009 13389
rect 4271 13345 15009 13351
rect 15061 13345 15079 13389
rect 4271 13337 15079 13345
rect 4288 13336 15079 13337
rect 14992 13328 15079 13336
rect 3011 13295 3132 13316
rect 3011 13222 3025 13295
rect 3095 13279 3132 13295
rect 13728 13279 13827 13285
rect 3095 13271 13827 13279
rect 3095 13222 13748 13271
rect 3011 13221 13748 13222
rect 13800 13221 13827 13271
rect 3011 13209 13827 13221
rect 3011 13206 3132 13209
rect 13728 13201 13827 13209
rect 46 13009 3791 13024
rect 46 12976 827 13009
rect 863 13005 3791 13009
rect 863 12976 1875 13005
rect 46 12972 1875 12976
rect 1911 12972 3791 13005
rect 46 12955 3791 12972
rect 46 12349 153 12955
rect 2653 12953 3791 12955
rect 10518 13018 10862 13021
rect 10518 13003 14499 13018
rect 10518 12970 11535 13003
rect 11571 12999 14499 13003
rect 11571 12970 12583 12999
rect 10518 12966 12583 12970
rect 12619 12966 14499 12999
rect 10518 12949 14499 12966
rect 10518 12940 10862 12949
rect 13361 12947 14499 12949
rect 6397 12644 7902 12645
rect 10534 12644 10641 12940
rect 6397 12627 10641 12644
rect 6397 12594 9824 12627
rect 9860 12594 10641 12627
rect 6397 12575 10641 12594
rect 6397 12573 7902 12575
rect 46 12330 4186 12349
rect 46 12297 827 12330
rect 863 12325 4186 12330
rect 863 12297 3322 12325
rect 46 12292 3322 12297
rect 3358 12292 4186 12325
rect 46 12280 4186 12292
rect 46 11577 153 12280
rect 2574 12279 4186 12280
rect 10534 11969 10641 12575
rect 6397 11952 10641 11969
rect 6397 11919 8776 11952
rect 8812 11948 10641 11952
rect 8812 11919 9824 11948
rect 6397 11915 9824 11919
rect 9860 11915 10641 11948
rect 6397 11900 10641 11915
rect 6397 11897 7936 11900
rect 2803 11580 3046 11585
rect 2751 11577 4011 11580
rect 46 11562 4011 11577
rect 46 11529 827 11562
rect 863 11558 4011 11562
rect 863 11529 1875 11558
rect 46 11525 1875 11529
rect 1911 11525 4011 11558
rect 46 11508 4011 11525
rect 46 10902 153 11508
rect 2803 11499 3046 11508
rect 6398 11197 8113 11198
rect 10534 11197 10641 11900
rect 6398 11185 10641 11197
rect 6398 11152 7329 11185
rect 7365 11180 10641 11185
rect 7365 11152 9824 11180
rect 6398 11147 9824 11152
rect 9860 11147 10641 11180
rect 6398 11128 10641 11147
rect 2785 10902 4235 10904
rect 46 10883 4235 10902
rect 46 10850 827 10883
rect 863 10880 4235 10883
rect 863 10850 3365 10880
rect 46 10847 3365 10850
rect 3401 10847 4235 10880
rect 46 10833 4235 10847
rect 46 10298 153 10833
rect 2785 10832 4235 10833
rect 6020 10522 8034 10524
rect 10534 10522 10641 11128
rect 6020 10505 10641 10522
rect 6020 10472 8776 10505
rect 8812 10501 10641 10505
rect 8812 10472 9824 10501
rect 6020 10468 9824 10472
rect 9860 10468 10641 10501
rect 6020 10453 10641 10468
rect 7705 10451 7893 10453
rect 46 10297 154 10298
rect 47 10274 154 10297
rect 45 10230 154 10274
rect 47 10057 154 10230
rect 10534 10280 10641 10453
rect 10754 12343 10861 12940
rect 17105 12638 18610 12639
rect 21242 12638 21349 13184
rect 17105 12621 21349 12638
rect 17105 12588 20532 12621
rect 20568 12588 21349 12621
rect 17105 12569 21349 12588
rect 17105 12567 18610 12569
rect 10754 12324 14894 12343
rect 10754 12291 11535 12324
rect 11571 12319 14894 12324
rect 11571 12291 14030 12319
rect 10754 12286 14030 12291
rect 14066 12286 14894 12319
rect 10754 12274 14894 12286
rect 10754 11571 10861 12274
rect 13282 12273 14894 12274
rect 21242 11963 21349 12569
rect 17105 11946 21349 11963
rect 17105 11913 19484 11946
rect 19520 11942 21349 11946
rect 19520 11913 20532 11942
rect 17105 11909 20532 11913
rect 20568 11909 21349 11942
rect 17105 11894 21349 11909
rect 17105 11891 18644 11894
rect 13511 11574 13754 11579
rect 13459 11571 14719 11574
rect 10754 11556 14719 11571
rect 10754 11523 11535 11556
rect 11571 11552 14719 11556
rect 11571 11523 12583 11552
rect 10754 11519 12583 11523
rect 12619 11519 14719 11552
rect 10754 11502 14719 11519
rect 10754 10896 10861 11502
rect 13511 11493 13754 11502
rect 17106 11191 18821 11192
rect 21242 11191 21349 11894
rect 17106 11179 21349 11191
rect 17106 11146 18037 11179
rect 18073 11174 21349 11179
rect 18073 11146 20532 11174
rect 17106 11141 20532 11146
rect 20568 11141 21349 11174
rect 17106 11122 21349 11141
rect 13493 10896 14943 10898
rect 10754 10877 14943 10896
rect 10754 10844 11535 10877
rect 11571 10874 14943 10877
rect 11571 10844 14073 10874
rect 10754 10841 14073 10844
rect 14109 10841 14943 10874
rect 10754 10827 14943 10841
rect 10754 10292 10861 10827
rect 13493 10826 14943 10827
rect 16728 10516 18742 10518
rect 21242 10516 21349 11122
rect 16728 10499 21349 10516
rect 16728 10466 19484 10499
rect 19520 10495 21349 10499
rect 19520 10466 20532 10495
rect 16728 10462 20532 10466
rect 20568 10462 21349 10495
rect 16728 10447 21349 10462
rect 18413 10445 18601 10447
rect 10754 10291 10862 10292
rect 10534 10236 10643 10280
rect 10755 10268 10862 10291
rect 10534 10213 10641 10236
rect 10753 10224 10862 10268
rect 10534 10212 10642 10213
rect 2795 10057 2983 10059
rect 47 10042 3979 10057
rect 47 10009 828 10042
rect 864 10038 3979 10042
rect 864 10009 1876 10038
rect 47 10005 1876 10009
rect 1912 10005 3979 10038
rect 47 9988 3979 10005
rect 47 9382 154 9988
rect 2654 9986 3979 9988
rect 6407 9677 7903 9678
rect 10535 9677 10642 10212
rect 6407 9663 10642 9677
rect 6407 9630 7287 9663
rect 7323 9660 10642 9663
rect 7323 9630 9825 9660
rect 6407 9627 9825 9630
rect 9861 9627 10642 9660
rect 6407 9608 10642 9627
rect 6407 9606 7903 9608
rect 47 9363 4188 9382
rect 47 9330 828 9363
rect 864 9358 4188 9363
rect 864 9330 3323 9358
rect 47 9325 3323 9330
rect 3359 9325 4188 9358
rect 47 9313 4188 9325
rect 47 8610 154 9313
rect 2575 9312 4188 9313
rect 7642 9002 7885 9011
rect 10535 9002 10642 9608
rect 6407 8985 10642 9002
rect 6407 8952 8777 8985
rect 8813 8981 10642 8985
rect 8813 8952 9825 8981
rect 6407 8948 9825 8952
rect 9861 8948 10642 8981
rect 6407 8933 10642 8948
rect 6407 8930 7937 8933
rect 7642 8925 7885 8930
rect 2752 8610 3761 8613
rect 47 8595 3761 8610
rect 47 8562 828 8595
rect 864 8591 3761 8595
rect 864 8562 1876 8591
rect 47 8558 1876 8562
rect 1912 8558 3761 8591
rect 47 8541 3761 8558
rect 47 7935 154 8541
rect 6407 8230 8114 8231
rect 10535 8230 10642 8933
rect 6407 8218 10642 8230
rect 6407 8185 7330 8218
rect 7366 8213 10642 8218
rect 7366 8185 9825 8213
rect 6407 8180 9825 8185
rect 9861 8180 10642 8213
rect 6407 8161 10642 8180
rect 2786 7936 4291 7937
rect 2786 7935 4491 7936
rect 47 7920 4491 7935
rect 47 7916 4494 7920
rect 47 7883 828 7916
rect 864 7907 4494 7916
rect 864 7883 4431 7907
rect 47 7874 4431 7883
rect 4467 7874 4494 7907
rect 47 7866 4494 7874
rect 47 7349 154 7866
rect 2786 7865 4494 7866
rect 4256 7862 4494 7865
rect 6463 7555 8035 7557
rect 10535 7555 10642 8161
rect 6463 7538 10642 7555
rect 6463 7505 8777 7538
rect 8813 7534 10642 7538
rect 8813 7505 9825 7534
rect 6463 7501 9825 7505
rect 9861 7501 10642 7534
rect 6463 7486 10642 7501
rect 40 7157 156 7349
rect 10535 7345 10642 7486
rect 10755 10051 10862 10224
rect 21242 10274 21349 10447
rect 21242 10230 21351 10274
rect 21242 10207 21349 10230
rect 21242 10206 21350 10207
rect 13503 10051 13691 10053
rect 10755 10036 14687 10051
rect 10755 10003 11536 10036
rect 11572 10032 14687 10036
rect 11572 10003 12584 10032
rect 10755 9999 12584 10003
rect 12620 9999 14687 10032
rect 10755 9982 14687 9999
rect 10755 9376 10862 9982
rect 13362 9980 14687 9982
rect 17115 9671 18611 9672
rect 21243 9671 21350 10206
rect 17115 9657 21350 9671
rect 17115 9624 17995 9657
rect 18031 9654 21350 9657
rect 18031 9624 20533 9654
rect 17115 9621 20533 9624
rect 20569 9621 21350 9654
rect 17115 9602 21350 9621
rect 17115 9600 18611 9602
rect 10755 9357 14896 9376
rect 10755 9324 11536 9357
rect 11572 9352 14896 9357
rect 11572 9324 14031 9352
rect 10755 9319 14031 9324
rect 14067 9319 14896 9352
rect 10755 9307 14896 9319
rect 10755 8604 10862 9307
rect 13283 9306 14896 9307
rect 18350 8996 18593 9005
rect 21243 8996 21350 9602
rect 17115 8979 21350 8996
rect 17115 8946 19485 8979
rect 19521 8975 21350 8979
rect 19521 8946 20533 8975
rect 17115 8942 20533 8946
rect 20569 8942 21350 8975
rect 17115 8927 21350 8942
rect 17115 8924 18645 8927
rect 18350 8919 18593 8924
rect 13460 8604 14469 8607
rect 10755 8589 14469 8604
rect 10755 8556 11536 8589
rect 11572 8585 14469 8589
rect 11572 8556 12584 8585
rect 10755 8552 12584 8556
rect 12620 8552 14469 8585
rect 10755 8535 14469 8552
rect 10755 7929 10862 8535
rect 17115 8224 18822 8225
rect 21243 8224 21350 8927
rect 17115 8212 21350 8224
rect 17115 8179 18038 8212
rect 18074 8207 21350 8212
rect 18074 8179 20533 8207
rect 17115 8174 20533 8179
rect 20569 8174 21350 8207
rect 17115 8155 21350 8174
rect 13494 7930 14999 7931
rect 13494 7929 15199 7930
rect 10755 7914 15199 7929
rect 10755 7910 15202 7914
rect 10755 7877 11536 7910
rect 11572 7901 15202 7910
rect 11572 7877 15139 7901
rect 10755 7868 15139 7877
rect 15175 7868 15202 7901
rect 10755 7860 15202 7868
rect 44 7016 151 7157
rect 10530 7153 10646 7345
rect 10755 7343 10862 7860
rect 13494 7859 15202 7860
rect 14964 7856 15202 7859
rect 17171 7549 18743 7551
rect 21243 7549 21350 8155
rect 17171 7532 21350 7549
rect 17171 7499 19485 7532
rect 19521 7528 21350 7532
rect 19521 7499 20533 7528
rect 17171 7495 20533 7499
rect 20569 7495 21350 7528
rect 17171 7480 21350 7495
rect 44 7001 4223 7016
rect 44 6968 825 7001
rect 861 6997 4223 7001
rect 861 6968 1873 6997
rect 44 6964 1873 6968
rect 1909 6964 4223 6997
rect 44 6947 4223 6964
rect 44 6341 151 6947
rect 2651 6945 4223 6947
rect 6192 6637 6326 6640
rect 6413 6637 6430 6640
rect 6192 6636 7900 6637
rect 10532 6636 10639 7153
rect 10748 7151 10864 7343
rect 21243 7339 21350 7480
rect 6192 6628 10639 6636
rect 6192 6595 6219 6628
rect 6255 6619 10639 6628
rect 6255 6595 9822 6619
rect 6192 6586 9822 6595
rect 9858 6586 10639 6619
rect 6192 6582 10639 6586
rect 6195 6567 10639 6582
rect 6195 6566 7900 6567
rect 6311 6565 7900 6566
rect 6311 6550 6433 6565
rect 44 6322 4279 6341
rect 44 6289 825 6322
rect 861 6317 4279 6322
rect 861 6289 3320 6317
rect 44 6284 3320 6289
rect 3356 6284 4279 6317
rect 44 6272 4279 6284
rect 44 5569 151 6272
rect 2572 6271 4279 6272
rect 10532 5961 10639 6567
rect 6925 5944 10639 5961
rect 6925 5911 8774 5944
rect 8810 5940 10639 5944
rect 8810 5911 9822 5940
rect 6925 5907 9822 5911
rect 9858 5907 10639 5940
rect 6925 5892 10639 5907
rect 6925 5889 7934 5892
rect 2801 5572 3044 5577
rect 2749 5569 4279 5572
rect 44 5554 4279 5569
rect 44 5521 825 5554
rect 861 5550 4279 5554
rect 861 5521 1873 5550
rect 44 5517 1873 5521
rect 1909 5517 4279 5550
rect 44 5500 4279 5517
rect 44 4894 151 5500
rect 2801 5491 3044 5500
rect 6498 5189 8111 5190
rect 10532 5189 10639 5892
rect 6498 5177 10639 5189
rect 6498 5144 7327 5177
rect 7363 5172 10639 5177
rect 7363 5144 9822 5172
rect 6498 5139 9822 5144
rect 9858 5139 10639 5172
rect 6498 5120 10639 5139
rect 2783 4894 4279 4896
rect 44 4875 4279 4894
rect 44 4842 825 4875
rect 861 4872 4279 4875
rect 861 4842 3363 4872
rect 44 4839 3363 4842
rect 3399 4839 4279 4872
rect 44 4825 4279 4839
rect 44 4290 151 4825
rect 2783 4824 4279 4825
rect 6707 4514 8032 4516
rect 10532 4514 10639 5120
rect 6707 4497 10639 4514
rect 6707 4464 8774 4497
rect 8810 4493 10639 4497
rect 8810 4464 9822 4493
rect 6707 4460 9822 4464
rect 9858 4460 10639 4493
rect 6707 4445 10639 4460
rect 7703 4443 7891 4445
rect 44 4289 152 4290
rect 45 4266 152 4289
rect 43 4222 152 4266
rect 45 4049 152 4222
rect 10532 4272 10639 4445
rect 10752 7010 10859 7151
rect 21238 7147 21354 7339
rect 10752 6995 14931 7010
rect 10752 6962 11533 6995
rect 11569 6991 14931 6995
rect 11569 6962 12581 6991
rect 10752 6958 12581 6962
rect 12617 6958 14931 6991
rect 10752 6941 14931 6958
rect 10752 6335 10859 6941
rect 13359 6939 14931 6941
rect 16900 6631 17034 6634
rect 17121 6631 17138 6634
rect 16900 6630 18608 6631
rect 21240 6630 21347 7147
rect 16900 6622 21347 6630
rect 16900 6589 16927 6622
rect 16963 6613 21347 6622
rect 16963 6589 20530 6613
rect 16900 6580 20530 6589
rect 20566 6580 21347 6613
rect 16900 6576 21347 6580
rect 16903 6561 21347 6576
rect 16903 6560 18608 6561
rect 17019 6559 18608 6560
rect 17019 6544 17141 6559
rect 10752 6316 14987 6335
rect 10752 6283 11533 6316
rect 11569 6311 14987 6316
rect 11569 6283 14028 6311
rect 10752 6278 14028 6283
rect 14064 6278 14987 6311
rect 10752 6266 14987 6278
rect 10752 5563 10859 6266
rect 13280 6265 14987 6266
rect 21240 5955 21347 6561
rect 17633 5938 21347 5955
rect 17633 5905 19482 5938
rect 19518 5934 21347 5938
rect 19518 5905 20530 5934
rect 17633 5901 20530 5905
rect 20566 5901 21347 5934
rect 17633 5886 21347 5901
rect 17633 5883 18642 5886
rect 13509 5566 13752 5571
rect 13457 5563 14987 5566
rect 10752 5548 14987 5563
rect 10752 5515 11533 5548
rect 11569 5544 14987 5548
rect 11569 5515 12581 5544
rect 10752 5511 12581 5515
rect 12617 5511 14987 5544
rect 10752 5494 14987 5511
rect 10752 4888 10859 5494
rect 13509 5485 13752 5494
rect 17206 5183 18819 5184
rect 21240 5183 21347 5886
rect 17206 5171 21347 5183
rect 17206 5138 18035 5171
rect 18071 5166 21347 5171
rect 18071 5138 20530 5166
rect 17206 5133 20530 5138
rect 20566 5133 21347 5166
rect 17206 5114 21347 5133
rect 13491 4888 14987 4890
rect 10752 4869 14987 4888
rect 10752 4836 11533 4869
rect 11569 4866 14987 4869
rect 11569 4836 14071 4866
rect 10752 4833 14071 4836
rect 14107 4833 14987 4866
rect 10752 4819 14987 4833
rect 10752 4284 10859 4819
rect 13491 4818 14987 4819
rect 17415 4508 18740 4510
rect 21240 4508 21347 5114
rect 17415 4491 21347 4508
rect 17415 4458 19482 4491
rect 19518 4487 21347 4491
rect 19518 4458 20530 4487
rect 17415 4454 20530 4458
rect 20566 4454 21347 4487
rect 17415 4439 21347 4454
rect 18411 4437 18599 4439
rect 10752 4283 10860 4284
rect 10532 4228 10641 4272
rect 10753 4260 10860 4283
rect 10532 4205 10639 4228
rect 10751 4216 10860 4260
rect 10532 4204 10640 4205
rect 2793 4049 2981 4051
rect 4572 4049 4990 4056
rect 45 4036 4990 4049
rect 45 4034 4776 4036
rect 45 4001 826 4034
rect 862 4030 4776 4034
rect 862 4001 1874 4030
rect 45 3997 1874 4001
rect 1910 4003 4776 4030
rect 4812 4003 4990 4036
rect 1910 3997 4990 4003
rect 45 3985 4990 3997
rect 45 3980 4666 3985
rect 45 3374 152 3980
rect 2652 3978 4666 3980
rect 6451 3669 7901 3670
rect 10533 3669 10640 4204
rect 6451 3655 10640 3669
rect 6451 3622 7285 3655
rect 7321 3652 10640 3655
rect 7321 3622 9823 3652
rect 6451 3619 9823 3622
rect 9859 3619 10640 3652
rect 6451 3600 10640 3619
rect 6451 3598 7901 3600
rect 45 3355 4288 3374
rect 45 3322 826 3355
rect 862 3350 4288 3355
rect 862 3322 3321 3350
rect 45 3317 3321 3322
rect 3357 3317 4288 3350
rect 45 3305 4288 3317
rect 45 2602 152 3305
rect 2573 3304 4288 3305
rect 7640 2994 7883 3003
rect 10533 2994 10640 3600
rect 6675 2977 10640 2994
rect 6675 2944 8775 2977
rect 8811 2973 10640 2977
rect 8811 2944 9823 2973
rect 6675 2940 9823 2944
rect 9859 2940 10640 2973
rect 6675 2925 10640 2940
rect 6675 2922 7935 2925
rect 7640 2917 7883 2922
rect 2750 2602 4289 2605
rect 45 2587 4289 2602
rect 45 2554 826 2587
rect 862 2583 4289 2587
rect 862 2554 1874 2583
rect 45 2550 1874 2554
rect 1910 2550 4289 2583
rect 45 2533 4289 2550
rect 45 1927 152 2533
rect 6500 2222 8112 2223
rect 10533 2222 10640 2925
rect 6500 2210 10640 2222
rect 6500 2177 7328 2210
rect 7364 2205 10640 2210
rect 7364 2177 9823 2205
rect 6500 2172 9823 2177
rect 9859 2172 10640 2205
rect 6500 2153 10640 2172
rect 2784 1927 4289 1929
rect 45 1908 4289 1927
rect 45 1875 826 1908
rect 862 1875 4289 1908
rect 45 1858 4289 1875
rect 45 1359 152 1858
rect 2784 1857 4289 1858
rect 7675 1547 8033 1549
rect 10533 1547 10640 2153
rect 7675 1530 10640 1547
rect 7675 1497 8775 1530
rect 8811 1526 10640 1530
rect 8811 1497 9823 1526
rect 7675 1493 9823 1497
rect 9859 1496 10640 1526
rect 10753 4043 10860 4216
rect 21240 4266 21347 4439
rect 21240 4222 21349 4266
rect 21240 4199 21347 4222
rect 21240 4198 21348 4199
rect 13501 4043 13689 4045
rect 15280 4043 15698 4050
rect 10753 4030 15698 4043
rect 10753 4028 15484 4030
rect 10753 3995 11534 4028
rect 11570 4024 15484 4028
rect 11570 3995 12582 4024
rect 10753 3991 12582 3995
rect 12618 3997 15484 4024
rect 15520 3997 15698 4030
rect 12618 3991 15698 3997
rect 10753 3979 15698 3991
rect 10753 3974 15374 3979
rect 10753 3368 10860 3974
rect 13360 3972 15374 3974
rect 17159 3663 18609 3664
rect 21241 3663 21348 4198
rect 17159 3649 21348 3663
rect 17159 3616 17993 3649
rect 18029 3646 21348 3649
rect 18029 3616 20531 3646
rect 17159 3613 20531 3616
rect 20567 3613 21348 3646
rect 17159 3594 21348 3613
rect 17159 3592 18609 3594
rect 10753 3349 14996 3368
rect 10753 3316 11534 3349
rect 11570 3344 14996 3349
rect 11570 3316 14029 3344
rect 10753 3311 14029 3316
rect 14065 3311 14996 3344
rect 10753 3299 14996 3311
rect 10753 2596 10860 3299
rect 13281 3298 14996 3299
rect 18348 2988 18591 2997
rect 21241 2988 21348 3594
rect 17383 2971 21348 2988
rect 17383 2938 19483 2971
rect 19519 2967 21348 2971
rect 19519 2938 20531 2967
rect 17383 2934 20531 2938
rect 20567 2934 21348 2967
rect 17383 2919 21348 2934
rect 17383 2916 18643 2919
rect 18348 2911 18591 2916
rect 13458 2596 14997 2599
rect 10753 2581 14997 2596
rect 10753 2548 11534 2581
rect 11570 2577 14997 2581
rect 11570 2548 12582 2577
rect 10753 2544 12582 2548
rect 12618 2544 14997 2577
rect 10753 2527 14997 2544
rect 10753 1921 10860 2527
rect 17208 2216 18820 2217
rect 21241 2216 21348 2919
rect 17208 2204 21348 2216
rect 17208 2171 18036 2204
rect 18072 2199 21348 2204
rect 18072 2171 20531 2199
rect 17208 2166 20531 2171
rect 20567 2166 21348 2199
rect 17208 2147 21348 2166
rect 13492 1921 14997 1923
rect 10753 1902 14997 1921
rect 10753 1869 11534 1902
rect 11570 1869 14997 1902
rect 10753 1852 14997 1869
rect 9859 1493 10679 1496
rect 7675 1478 10679 1493
rect 20 1321 153 1359
rect 20 1209 53 1321
rect 132 1290 153 1321
rect 10508 1342 10679 1478
rect 10753 1353 10860 1852
rect 13492 1851 14997 1852
rect 18383 1541 18741 1543
rect 21241 1541 21348 2147
rect 18383 1524 21348 1541
rect 18383 1491 19483 1524
rect 19519 1520 21348 1524
rect 19519 1491 20531 1520
rect 18383 1487 20531 1491
rect 20567 1490 21348 1520
rect 20567 1487 21387 1490
rect 18383 1472 21387 1487
rect 132 1246 165 1290
rect 132 1209 153 1246
rect 20 1192 153 1209
rect 10508 1230 10529 1342
rect 10650 1230 10679 1342
rect 10508 1180 10679 1230
rect 10728 1315 10861 1353
rect 10728 1203 10761 1315
rect 10840 1284 10861 1315
rect 21216 1336 21387 1472
rect 10840 1240 10873 1284
rect 10840 1203 10861 1240
rect 10728 1186 10861 1203
rect 21216 1224 21237 1336
rect 21358 1224 21387 1336
rect 21216 1174 21387 1224
rect 2778 1088 7841 1097
rect 2778 1013 2807 1088
rect 2924 1084 7841 1088
rect 2924 1013 7737 1084
rect 7816 1076 7841 1084
rect 13486 1082 18549 1091
rect 13486 1076 13515 1082
rect 7816 1013 13515 1076
rect 2778 1007 13515 1013
rect 13632 1078 18549 1082
rect 13632 1007 18445 1078
rect 18524 1007 18549 1078
rect 2778 1006 18549 1007
rect 2778 997 7841 1006
rect 13486 991 18549 1006
rect 1734 894 8965 920
rect 12442 894 19673 914
rect 1734 893 19673 894
rect 1734 818 1759 893
rect 1829 818 8856 893
rect 1734 814 8856 818
rect 8940 887 19673 893
rect 8940 814 12467 887
rect 1734 812 12467 814
rect 12537 812 19564 887
rect 1734 808 19564 812
rect 19648 808 19673 887
rect 1734 787 8965 808
rect 12442 781 19673 808
rect 685 700 9992 710
rect 11393 700 20700 704
rect 685 693 20700 700
rect 685 681 9872 693
rect 685 602 710 681
rect 810 614 9872 681
rect 9972 687 20700 693
rect 9972 675 20580 687
rect 9972 614 11418 675
rect 810 602 11418 614
rect 685 598 11418 602
rect 685 593 9992 598
rect 11393 596 11418 598
rect 11518 608 20580 675
rect 20680 608 20700 687
rect 11518 596 20700 608
rect 11393 587 20700 596
rect 219 491 10479 493
rect 219 487 11308 491
rect 219 468 21187 487
rect 219 460 10238 468
rect 219 373 257 460
rect 327 381 10238 460
rect 10308 462 21187 468
rect 10308 460 20946 462
rect 10308 381 10371 460
rect 327 373 10371 381
rect 10441 454 20946 460
rect 10441 373 10965 454
rect 219 367 10965 373
rect 11035 375 20946 454
rect 21016 454 21187 462
rect 21016 375 21079 454
rect 11035 367 21079 375
rect 21149 367 21187 454
rect 219 335 21187 367
rect 219 331 10479 335
rect 10927 325 21187 335
rect 0 244 10673 249
rect 0 243 11189 244
rect 0 220 21381 243
rect 0 125 25 220
rect 115 215 21381 220
rect 115 125 10544 215
rect 0 120 10544 125
rect 10634 214 21381 215
rect 10634 120 10733 214
rect 0 119 10733 120
rect 10823 209 21381 214
rect 10823 119 21252 209
rect 0 114 21252 119
rect 21342 114 21381 209
rect 0 95 21381 114
rect 10233 89 21381 95
rect 10233 88 11189 89
rect 10512 -251 10621 88
rect 10512 -284 10537 -251
rect 10573 -284 10621 -251
rect 10512 -297 10621 -284
<< labels >>
rlabel metal1 1750 13395 1803 13417 1 d1
rlabel metal1 704 13413 766 13440 1 d0
rlabel metal2 49 13398 145 13431 1 vdd
rlabel metal1 225 13398 321 13431 1 gnd
rlabel locali 489 13409 533 13431 1 vref
rlabel metal1 4298 13736 4333 13750 1 d4
rlabel metal1 3036 13691 3088 13710 1 d3
rlabel metal1 2860 13708 2910 13721 1 d2
rlabel metal1 5347 13711 5417 13755 1 d5
rlabel metal1 -56 -497 -25 -438 1 d6
rlabel metal1 11105 -755 11134 -737 1 vout
<< end >>
