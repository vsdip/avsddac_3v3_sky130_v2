magic
tech sky130A
timestamp 1616160868
<< nwell >>
rect 278 7913 1089 8063
rect 4103 7937 4914 8087
rect 5559 7892 6370 8042
rect 9384 7916 10195 8066
rect 1290 7732 2101 7882
rect 3090 7703 3901 7853
rect 6571 7711 7382 7861
rect 8371 7682 9182 7832
rect 277 7498 1088 7648
rect 4102 7522 4913 7672
rect 5558 7477 6369 7627
rect 9383 7501 10194 7651
rect 1345 7171 2156 7321
rect 3040 7283 3851 7433
rect 6626 7150 7437 7300
rect 8321 7262 9132 7412
rect 283 6932 1094 7082
rect 4108 6956 4919 7106
rect 5564 6911 6375 7061
rect 9389 6935 10200 7085
rect 1295 6751 2106 6901
rect 3095 6722 3906 6872
rect 6576 6730 7387 6880
rect 8376 6701 9187 6851
rect 282 6517 1093 6667
rect 4107 6541 4918 6691
rect 5563 6496 6374 6646
rect 9388 6520 10199 6670
rect 1510 6239 2321 6389
rect 2887 6255 3698 6405
rect 6791 6218 7602 6368
rect 8168 6234 8979 6384
rect 290 5953 1101 6103
rect 4115 5977 4926 6127
rect 5571 5932 6382 6082
rect 9396 5956 10207 6106
rect 1302 5772 2113 5922
rect 3102 5743 3913 5893
rect 6583 5751 7394 5901
rect 8383 5722 9194 5872
rect 289 5538 1100 5688
rect 4114 5562 4925 5712
rect 5570 5517 6381 5667
rect 9395 5541 10206 5691
rect 1357 5211 2168 5361
rect 3052 5323 3863 5473
rect 6638 5190 7449 5340
rect 8333 5302 9144 5452
rect 295 4972 1106 5122
rect 4120 4996 4931 5146
rect 5576 4951 6387 5101
rect 9401 4975 10212 5125
rect 1307 4791 2118 4941
rect 3107 4762 3918 4912
rect 6588 4770 7399 4920
rect 8388 4741 9199 4891
rect 294 4557 1105 4707
rect 4119 4581 4930 4731
rect 5575 4536 6386 4686
rect 9400 4560 10211 4710
rect 1605 4247 2416 4397
rect 2812 4330 3623 4480
rect 6886 4226 7697 4376
rect 8093 4309 8904 4459
rect 298 3996 1109 4146
rect 4123 4020 4934 4170
rect 5579 3975 6390 4125
rect 9404 3999 10215 4149
rect 1310 3815 2121 3965
rect 3110 3786 3921 3936
rect 6591 3794 7402 3944
rect 8391 3765 9202 3915
rect 297 3581 1108 3731
rect 4122 3605 4933 3755
rect 5578 3560 6389 3710
rect 9403 3584 10214 3734
rect 1365 3254 2176 3404
rect 3060 3366 3871 3516
rect 6646 3233 7457 3383
rect 8341 3345 9152 3495
rect 303 3015 1114 3165
rect 4128 3039 4939 3189
rect 5584 2994 6395 3144
rect 9409 3018 10220 3168
rect 1315 2834 2126 2984
rect 3115 2805 3926 2955
rect 6596 2813 7407 2963
rect 8396 2784 9207 2934
rect 302 2600 1113 2750
rect 4127 2624 4938 2774
rect 5583 2579 6394 2729
rect 9408 2603 10219 2753
rect 1530 2322 2341 2472
rect 2907 2338 3718 2488
rect 6811 2301 7622 2451
rect 8188 2317 8999 2467
rect 310 2036 1121 2186
rect 4135 2060 4946 2210
rect 5591 2015 6402 2165
rect 9416 2039 10227 2189
rect 1322 1855 2133 2005
rect 3122 1826 3933 1976
rect 6603 1834 7414 1984
rect 8403 1805 9214 1955
rect 309 1621 1120 1771
rect 4134 1645 4945 1795
rect 5590 1600 6401 1750
rect 9415 1624 10226 1774
rect 1377 1294 2188 1444
rect 3072 1406 3883 1556
rect 6658 1273 7469 1423
rect 8353 1385 9164 1535
rect 315 1055 1126 1205
rect 4140 1079 4951 1229
rect 5596 1034 6407 1184
rect 9421 1058 10232 1208
rect 1327 874 2138 1024
rect 3127 845 3938 995
rect 6608 853 7419 1003
rect 8408 824 9219 974
rect 314 640 1125 790
rect 4139 664 4950 814
rect 5595 619 6406 769
rect 9420 643 10231 793
rect 1717 159 2528 309
rect 4807 71 5618 221
rect 6998 138 7809 288
<< nmos >>
rect 4171 8146 4221 8188
rect 4379 8146 4429 8188
rect 4587 8146 4637 8188
rect 4800 8146 4850 8188
rect 9452 8125 9502 8167
rect 9660 8125 9710 8167
rect 9868 8125 9918 8167
rect 10081 8125 10131 8167
rect 3158 7912 3208 7954
rect 3366 7912 3416 7954
rect 3574 7912 3624 7954
rect 3787 7912 3837 7954
rect 342 7812 392 7854
rect 555 7812 605 7854
rect 763 7812 813 7854
rect 971 7812 1021 7854
rect 8439 7891 8489 7933
rect 8647 7891 8697 7933
rect 8855 7891 8905 7933
rect 9068 7891 9118 7933
rect 5623 7791 5673 7833
rect 5836 7791 5886 7833
rect 6044 7791 6094 7833
rect 6252 7791 6302 7833
rect 4170 7731 4220 7773
rect 4378 7731 4428 7773
rect 4586 7731 4636 7773
rect 4799 7731 4849 7773
rect 1354 7631 1404 7673
rect 1567 7631 1617 7673
rect 1775 7631 1825 7673
rect 1983 7631 2033 7673
rect 9451 7710 9501 7752
rect 9659 7710 9709 7752
rect 9867 7710 9917 7752
rect 10080 7710 10130 7752
rect 6635 7610 6685 7652
rect 6848 7610 6898 7652
rect 7056 7610 7106 7652
rect 7264 7610 7314 7652
rect 3108 7492 3158 7534
rect 3316 7492 3366 7534
rect 3524 7492 3574 7534
rect 3737 7492 3787 7534
rect 341 7397 391 7439
rect 554 7397 604 7439
rect 762 7397 812 7439
rect 970 7397 1020 7439
rect 8389 7471 8439 7513
rect 8597 7471 8647 7513
rect 8805 7471 8855 7513
rect 9018 7471 9068 7513
rect 5622 7376 5672 7418
rect 5835 7376 5885 7418
rect 6043 7376 6093 7418
rect 6251 7376 6301 7418
rect 4176 7165 4226 7207
rect 4384 7165 4434 7207
rect 4592 7165 4642 7207
rect 4805 7165 4855 7207
rect 1409 7070 1459 7112
rect 1622 7070 1672 7112
rect 1830 7070 1880 7112
rect 2038 7070 2088 7112
rect 9457 7144 9507 7186
rect 9665 7144 9715 7186
rect 9873 7144 9923 7186
rect 10086 7144 10136 7186
rect 6690 7049 6740 7091
rect 6903 7049 6953 7091
rect 7111 7049 7161 7091
rect 7319 7049 7369 7091
rect 3163 6931 3213 6973
rect 3371 6931 3421 6973
rect 3579 6931 3629 6973
rect 3792 6931 3842 6973
rect 347 6831 397 6873
rect 560 6831 610 6873
rect 768 6831 818 6873
rect 976 6831 1026 6873
rect 8444 6910 8494 6952
rect 8652 6910 8702 6952
rect 8860 6910 8910 6952
rect 9073 6910 9123 6952
rect 5628 6810 5678 6852
rect 5841 6810 5891 6852
rect 6049 6810 6099 6852
rect 6257 6810 6307 6852
rect 4175 6750 4225 6792
rect 4383 6750 4433 6792
rect 4591 6750 4641 6792
rect 4804 6750 4854 6792
rect 1359 6650 1409 6692
rect 1572 6650 1622 6692
rect 1780 6650 1830 6692
rect 1988 6650 2038 6692
rect 9456 6729 9506 6771
rect 9664 6729 9714 6771
rect 9872 6729 9922 6771
rect 10085 6729 10135 6771
rect 6640 6629 6690 6671
rect 6853 6629 6903 6671
rect 7061 6629 7111 6671
rect 7269 6629 7319 6671
rect 2955 6464 3005 6506
rect 3163 6464 3213 6506
rect 3371 6464 3421 6506
rect 3584 6464 3634 6506
rect 346 6416 396 6458
rect 559 6416 609 6458
rect 767 6416 817 6458
rect 975 6416 1025 6458
rect 8236 6443 8286 6485
rect 8444 6443 8494 6485
rect 8652 6443 8702 6485
rect 8865 6443 8915 6485
rect 5627 6395 5677 6437
rect 5840 6395 5890 6437
rect 6048 6395 6098 6437
rect 6256 6395 6306 6437
rect 4183 6186 4233 6228
rect 4391 6186 4441 6228
rect 4599 6186 4649 6228
rect 4812 6186 4862 6228
rect 1574 6138 1624 6180
rect 1787 6138 1837 6180
rect 1995 6138 2045 6180
rect 2203 6138 2253 6180
rect 9464 6165 9514 6207
rect 9672 6165 9722 6207
rect 9880 6165 9930 6207
rect 10093 6165 10143 6207
rect 6855 6117 6905 6159
rect 7068 6117 7118 6159
rect 7276 6117 7326 6159
rect 7484 6117 7534 6159
rect 3170 5952 3220 5994
rect 3378 5952 3428 5994
rect 3586 5952 3636 5994
rect 3799 5952 3849 5994
rect 354 5852 404 5894
rect 567 5852 617 5894
rect 775 5852 825 5894
rect 983 5852 1033 5894
rect 8451 5931 8501 5973
rect 8659 5931 8709 5973
rect 8867 5931 8917 5973
rect 9080 5931 9130 5973
rect 5635 5831 5685 5873
rect 5848 5831 5898 5873
rect 6056 5831 6106 5873
rect 6264 5831 6314 5873
rect 4182 5771 4232 5813
rect 4390 5771 4440 5813
rect 4598 5771 4648 5813
rect 4811 5771 4861 5813
rect 1366 5671 1416 5713
rect 1579 5671 1629 5713
rect 1787 5671 1837 5713
rect 1995 5671 2045 5713
rect 9463 5750 9513 5792
rect 9671 5750 9721 5792
rect 9879 5750 9929 5792
rect 10092 5750 10142 5792
rect 6647 5650 6697 5692
rect 6860 5650 6910 5692
rect 7068 5650 7118 5692
rect 7276 5650 7326 5692
rect 3120 5532 3170 5574
rect 3328 5532 3378 5574
rect 3536 5532 3586 5574
rect 3749 5532 3799 5574
rect 353 5437 403 5479
rect 566 5437 616 5479
rect 774 5437 824 5479
rect 982 5437 1032 5479
rect 8401 5511 8451 5553
rect 8609 5511 8659 5553
rect 8817 5511 8867 5553
rect 9030 5511 9080 5553
rect 5634 5416 5684 5458
rect 5847 5416 5897 5458
rect 6055 5416 6105 5458
rect 6263 5416 6313 5458
rect 4188 5205 4238 5247
rect 4396 5205 4446 5247
rect 4604 5205 4654 5247
rect 4817 5205 4867 5247
rect 1421 5110 1471 5152
rect 1634 5110 1684 5152
rect 1842 5110 1892 5152
rect 2050 5110 2100 5152
rect 9469 5184 9519 5226
rect 9677 5184 9727 5226
rect 9885 5184 9935 5226
rect 10098 5184 10148 5226
rect 6702 5089 6752 5131
rect 6915 5089 6965 5131
rect 7123 5089 7173 5131
rect 7331 5089 7381 5131
rect 3175 4971 3225 5013
rect 3383 4971 3433 5013
rect 3591 4971 3641 5013
rect 3804 4971 3854 5013
rect 359 4871 409 4913
rect 572 4871 622 4913
rect 780 4871 830 4913
rect 988 4871 1038 4913
rect 8456 4950 8506 4992
rect 8664 4950 8714 4992
rect 8872 4950 8922 4992
rect 9085 4950 9135 4992
rect 5640 4850 5690 4892
rect 5853 4850 5903 4892
rect 6061 4850 6111 4892
rect 6269 4850 6319 4892
rect 4187 4790 4237 4832
rect 4395 4790 4445 4832
rect 4603 4790 4653 4832
rect 4816 4790 4866 4832
rect 1371 4690 1421 4732
rect 1584 4690 1634 4732
rect 1792 4690 1842 4732
rect 2000 4690 2050 4732
rect 9468 4769 9518 4811
rect 9676 4769 9726 4811
rect 9884 4769 9934 4811
rect 10097 4769 10147 4811
rect 6652 4669 6702 4711
rect 6865 4669 6915 4711
rect 7073 4669 7123 4711
rect 7281 4669 7331 4711
rect 2880 4539 2930 4581
rect 3088 4539 3138 4581
rect 3296 4539 3346 4581
rect 3509 4539 3559 4581
rect 358 4456 408 4498
rect 571 4456 621 4498
rect 779 4456 829 4498
rect 987 4456 1037 4498
rect 8161 4518 8211 4560
rect 8369 4518 8419 4560
rect 8577 4518 8627 4560
rect 8790 4518 8840 4560
rect 5639 4435 5689 4477
rect 5852 4435 5902 4477
rect 6060 4435 6110 4477
rect 6268 4435 6318 4477
rect 4191 4229 4241 4271
rect 4399 4229 4449 4271
rect 4607 4229 4657 4271
rect 4820 4229 4870 4271
rect 1669 4146 1719 4188
rect 1882 4146 1932 4188
rect 2090 4146 2140 4188
rect 2298 4146 2348 4188
rect 9472 4208 9522 4250
rect 9680 4208 9730 4250
rect 9888 4208 9938 4250
rect 10101 4208 10151 4250
rect 6950 4125 7000 4167
rect 7163 4125 7213 4167
rect 7371 4125 7421 4167
rect 7579 4125 7629 4167
rect 3178 3995 3228 4037
rect 3386 3995 3436 4037
rect 3594 3995 3644 4037
rect 3807 3995 3857 4037
rect 362 3895 412 3937
rect 575 3895 625 3937
rect 783 3895 833 3937
rect 991 3895 1041 3937
rect 8459 3974 8509 4016
rect 8667 3974 8717 4016
rect 8875 3974 8925 4016
rect 9088 3974 9138 4016
rect 5643 3874 5693 3916
rect 5856 3874 5906 3916
rect 6064 3874 6114 3916
rect 6272 3874 6322 3916
rect 4190 3814 4240 3856
rect 4398 3814 4448 3856
rect 4606 3814 4656 3856
rect 4819 3814 4869 3856
rect 1374 3714 1424 3756
rect 1587 3714 1637 3756
rect 1795 3714 1845 3756
rect 2003 3714 2053 3756
rect 9471 3793 9521 3835
rect 9679 3793 9729 3835
rect 9887 3793 9937 3835
rect 10100 3793 10150 3835
rect 6655 3693 6705 3735
rect 6868 3693 6918 3735
rect 7076 3693 7126 3735
rect 7284 3693 7334 3735
rect 3128 3575 3178 3617
rect 3336 3575 3386 3617
rect 3544 3575 3594 3617
rect 3757 3575 3807 3617
rect 361 3480 411 3522
rect 574 3480 624 3522
rect 782 3480 832 3522
rect 990 3480 1040 3522
rect 8409 3554 8459 3596
rect 8617 3554 8667 3596
rect 8825 3554 8875 3596
rect 9038 3554 9088 3596
rect 5642 3459 5692 3501
rect 5855 3459 5905 3501
rect 6063 3459 6113 3501
rect 6271 3459 6321 3501
rect 4196 3248 4246 3290
rect 4404 3248 4454 3290
rect 4612 3248 4662 3290
rect 4825 3248 4875 3290
rect 1429 3153 1479 3195
rect 1642 3153 1692 3195
rect 1850 3153 1900 3195
rect 2058 3153 2108 3195
rect 9477 3227 9527 3269
rect 9685 3227 9735 3269
rect 9893 3227 9943 3269
rect 10106 3227 10156 3269
rect 6710 3132 6760 3174
rect 6923 3132 6973 3174
rect 7131 3132 7181 3174
rect 7339 3132 7389 3174
rect 3183 3014 3233 3056
rect 3391 3014 3441 3056
rect 3599 3014 3649 3056
rect 3812 3014 3862 3056
rect 367 2914 417 2956
rect 580 2914 630 2956
rect 788 2914 838 2956
rect 996 2914 1046 2956
rect 8464 2993 8514 3035
rect 8672 2993 8722 3035
rect 8880 2993 8930 3035
rect 9093 2993 9143 3035
rect 5648 2893 5698 2935
rect 5861 2893 5911 2935
rect 6069 2893 6119 2935
rect 6277 2893 6327 2935
rect 4195 2833 4245 2875
rect 4403 2833 4453 2875
rect 4611 2833 4661 2875
rect 4824 2833 4874 2875
rect 1379 2733 1429 2775
rect 1592 2733 1642 2775
rect 1800 2733 1850 2775
rect 2008 2733 2058 2775
rect 9476 2812 9526 2854
rect 9684 2812 9734 2854
rect 9892 2812 9942 2854
rect 10105 2812 10155 2854
rect 6660 2712 6710 2754
rect 6873 2712 6923 2754
rect 7081 2712 7131 2754
rect 7289 2712 7339 2754
rect 2975 2547 3025 2589
rect 3183 2547 3233 2589
rect 3391 2547 3441 2589
rect 3604 2547 3654 2589
rect 366 2499 416 2541
rect 579 2499 629 2541
rect 787 2499 837 2541
rect 995 2499 1045 2541
rect 8256 2526 8306 2568
rect 8464 2526 8514 2568
rect 8672 2526 8722 2568
rect 8885 2526 8935 2568
rect 5647 2478 5697 2520
rect 5860 2478 5910 2520
rect 6068 2478 6118 2520
rect 6276 2478 6326 2520
rect 4203 2269 4253 2311
rect 4411 2269 4461 2311
rect 4619 2269 4669 2311
rect 4832 2269 4882 2311
rect 1594 2221 1644 2263
rect 1807 2221 1857 2263
rect 2015 2221 2065 2263
rect 2223 2221 2273 2263
rect 9484 2248 9534 2290
rect 9692 2248 9742 2290
rect 9900 2248 9950 2290
rect 10113 2248 10163 2290
rect 6875 2200 6925 2242
rect 7088 2200 7138 2242
rect 7296 2200 7346 2242
rect 7504 2200 7554 2242
rect 3190 2035 3240 2077
rect 3398 2035 3448 2077
rect 3606 2035 3656 2077
rect 3819 2035 3869 2077
rect 374 1935 424 1977
rect 587 1935 637 1977
rect 795 1935 845 1977
rect 1003 1935 1053 1977
rect 8471 2014 8521 2056
rect 8679 2014 8729 2056
rect 8887 2014 8937 2056
rect 9100 2014 9150 2056
rect 5655 1914 5705 1956
rect 5868 1914 5918 1956
rect 6076 1914 6126 1956
rect 6284 1914 6334 1956
rect 4202 1854 4252 1896
rect 4410 1854 4460 1896
rect 4618 1854 4668 1896
rect 4831 1854 4881 1896
rect 1386 1754 1436 1796
rect 1599 1754 1649 1796
rect 1807 1754 1857 1796
rect 2015 1754 2065 1796
rect 9483 1833 9533 1875
rect 9691 1833 9741 1875
rect 9899 1833 9949 1875
rect 10112 1833 10162 1875
rect 6667 1733 6717 1775
rect 6880 1733 6930 1775
rect 7088 1733 7138 1775
rect 7296 1733 7346 1775
rect 3140 1615 3190 1657
rect 3348 1615 3398 1657
rect 3556 1615 3606 1657
rect 3769 1615 3819 1657
rect 373 1520 423 1562
rect 586 1520 636 1562
rect 794 1520 844 1562
rect 1002 1520 1052 1562
rect 8421 1594 8471 1636
rect 8629 1594 8679 1636
rect 8837 1594 8887 1636
rect 9050 1594 9100 1636
rect 5654 1499 5704 1541
rect 5867 1499 5917 1541
rect 6075 1499 6125 1541
rect 6283 1499 6333 1541
rect 4208 1288 4258 1330
rect 4416 1288 4466 1330
rect 4624 1288 4674 1330
rect 4837 1288 4887 1330
rect 1441 1193 1491 1235
rect 1654 1193 1704 1235
rect 1862 1193 1912 1235
rect 2070 1193 2120 1235
rect 9489 1267 9539 1309
rect 9697 1267 9747 1309
rect 9905 1267 9955 1309
rect 10118 1267 10168 1309
rect 6722 1172 6772 1214
rect 6935 1172 6985 1214
rect 7143 1172 7193 1214
rect 7351 1172 7401 1214
rect 3195 1054 3245 1096
rect 3403 1054 3453 1096
rect 3611 1054 3661 1096
rect 3824 1054 3874 1096
rect 379 954 429 996
rect 592 954 642 996
rect 800 954 850 996
rect 1008 954 1058 996
rect 8476 1033 8526 1075
rect 8684 1033 8734 1075
rect 8892 1033 8942 1075
rect 9105 1033 9155 1075
rect 5660 933 5710 975
rect 5873 933 5923 975
rect 6081 933 6131 975
rect 6289 933 6339 975
rect 4207 873 4257 915
rect 4415 873 4465 915
rect 4623 873 4673 915
rect 4836 873 4886 915
rect 1391 773 1441 815
rect 1604 773 1654 815
rect 1812 773 1862 815
rect 2020 773 2070 815
rect 9488 852 9538 894
rect 9696 852 9746 894
rect 9904 852 9954 894
rect 10117 852 10167 894
rect 6672 752 6722 794
rect 6885 752 6935 794
rect 7093 752 7143 794
rect 7301 752 7351 794
rect 378 539 428 581
rect 591 539 641 581
rect 799 539 849 581
rect 1007 539 1057 581
rect 5659 518 5709 560
rect 5872 518 5922 560
rect 6080 518 6130 560
rect 6288 518 6338 560
rect 1781 58 1831 100
rect 1994 58 2044 100
rect 2202 58 2252 100
rect 2410 58 2460 100
rect 7062 37 7112 79
rect 7275 37 7325 79
rect 7483 37 7533 79
rect 7691 37 7741 79
rect 4871 -30 4921 12
rect 5084 -30 5134 12
rect 5292 -30 5342 12
rect 5500 -30 5550 12
<< pmos >>
rect 342 7931 392 8031
rect 555 7931 605 8031
rect 763 7931 813 8031
rect 971 7931 1021 8031
rect 4171 7969 4221 8069
rect 4379 7969 4429 8069
rect 4587 7969 4637 8069
rect 4800 7969 4850 8069
rect 1354 7750 1404 7850
rect 1567 7750 1617 7850
rect 1775 7750 1825 7850
rect 1983 7750 2033 7850
rect 5623 7910 5673 8010
rect 5836 7910 5886 8010
rect 6044 7910 6094 8010
rect 6252 7910 6302 8010
rect 9452 7948 9502 8048
rect 9660 7948 9710 8048
rect 9868 7948 9918 8048
rect 10081 7948 10131 8048
rect 3158 7735 3208 7835
rect 3366 7735 3416 7835
rect 3574 7735 3624 7835
rect 3787 7735 3837 7835
rect 6635 7729 6685 7829
rect 6848 7729 6898 7829
rect 7056 7729 7106 7829
rect 7264 7729 7314 7829
rect 341 7516 391 7616
rect 554 7516 604 7616
rect 762 7516 812 7616
rect 970 7516 1020 7616
rect 4170 7554 4220 7654
rect 4378 7554 4428 7654
rect 4586 7554 4636 7654
rect 4799 7554 4849 7654
rect 8439 7714 8489 7814
rect 8647 7714 8697 7814
rect 8855 7714 8905 7814
rect 9068 7714 9118 7814
rect 5622 7495 5672 7595
rect 5835 7495 5885 7595
rect 6043 7495 6093 7595
rect 6251 7495 6301 7595
rect 9451 7533 9501 7633
rect 9659 7533 9709 7633
rect 9867 7533 9917 7633
rect 10080 7533 10130 7633
rect 3108 7315 3158 7415
rect 3316 7315 3366 7415
rect 3524 7315 3574 7415
rect 3737 7315 3787 7415
rect 8389 7294 8439 7394
rect 8597 7294 8647 7394
rect 8805 7294 8855 7394
rect 9018 7294 9068 7394
rect 1409 7189 1459 7289
rect 1622 7189 1672 7289
rect 1830 7189 1880 7289
rect 2038 7189 2088 7289
rect 6690 7168 6740 7268
rect 6903 7168 6953 7268
rect 7111 7168 7161 7268
rect 7319 7168 7369 7268
rect 347 6950 397 7050
rect 560 6950 610 7050
rect 768 6950 818 7050
rect 976 6950 1026 7050
rect 4176 6988 4226 7088
rect 4384 6988 4434 7088
rect 4592 6988 4642 7088
rect 4805 6988 4855 7088
rect 1359 6769 1409 6869
rect 1572 6769 1622 6869
rect 1780 6769 1830 6869
rect 1988 6769 2038 6869
rect 5628 6929 5678 7029
rect 5841 6929 5891 7029
rect 6049 6929 6099 7029
rect 6257 6929 6307 7029
rect 9457 6967 9507 7067
rect 9665 6967 9715 7067
rect 9873 6967 9923 7067
rect 10086 6967 10136 7067
rect 3163 6754 3213 6854
rect 3371 6754 3421 6854
rect 3579 6754 3629 6854
rect 3792 6754 3842 6854
rect 6640 6748 6690 6848
rect 6853 6748 6903 6848
rect 7061 6748 7111 6848
rect 7269 6748 7319 6848
rect 346 6535 396 6635
rect 559 6535 609 6635
rect 767 6535 817 6635
rect 975 6535 1025 6635
rect 4175 6573 4225 6673
rect 4383 6573 4433 6673
rect 4591 6573 4641 6673
rect 4804 6573 4854 6673
rect 8444 6733 8494 6833
rect 8652 6733 8702 6833
rect 8860 6733 8910 6833
rect 9073 6733 9123 6833
rect 5627 6514 5677 6614
rect 5840 6514 5890 6614
rect 6048 6514 6098 6614
rect 6256 6514 6306 6614
rect 9456 6552 9506 6652
rect 9664 6552 9714 6652
rect 9872 6552 9922 6652
rect 10085 6552 10135 6652
rect 1574 6257 1624 6357
rect 1787 6257 1837 6357
rect 1995 6257 2045 6357
rect 2203 6257 2253 6357
rect 2955 6287 3005 6387
rect 3163 6287 3213 6387
rect 3371 6287 3421 6387
rect 3584 6287 3634 6387
rect 6855 6236 6905 6336
rect 7068 6236 7118 6336
rect 7276 6236 7326 6336
rect 7484 6236 7534 6336
rect 8236 6266 8286 6366
rect 8444 6266 8494 6366
rect 8652 6266 8702 6366
rect 8865 6266 8915 6366
rect 354 5971 404 6071
rect 567 5971 617 6071
rect 775 5971 825 6071
rect 983 5971 1033 6071
rect 4183 6009 4233 6109
rect 4391 6009 4441 6109
rect 4599 6009 4649 6109
rect 4812 6009 4862 6109
rect 1366 5790 1416 5890
rect 1579 5790 1629 5890
rect 1787 5790 1837 5890
rect 1995 5790 2045 5890
rect 5635 5950 5685 6050
rect 5848 5950 5898 6050
rect 6056 5950 6106 6050
rect 6264 5950 6314 6050
rect 9464 5988 9514 6088
rect 9672 5988 9722 6088
rect 9880 5988 9930 6088
rect 10093 5988 10143 6088
rect 3170 5775 3220 5875
rect 3378 5775 3428 5875
rect 3586 5775 3636 5875
rect 3799 5775 3849 5875
rect 6647 5769 6697 5869
rect 6860 5769 6910 5869
rect 7068 5769 7118 5869
rect 7276 5769 7326 5869
rect 353 5556 403 5656
rect 566 5556 616 5656
rect 774 5556 824 5656
rect 982 5556 1032 5656
rect 4182 5594 4232 5694
rect 4390 5594 4440 5694
rect 4598 5594 4648 5694
rect 4811 5594 4861 5694
rect 8451 5754 8501 5854
rect 8659 5754 8709 5854
rect 8867 5754 8917 5854
rect 9080 5754 9130 5854
rect 5634 5535 5684 5635
rect 5847 5535 5897 5635
rect 6055 5535 6105 5635
rect 6263 5535 6313 5635
rect 9463 5573 9513 5673
rect 9671 5573 9721 5673
rect 9879 5573 9929 5673
rect 10092 5573 10142 5673
rect 3120 5355 3170 5455
rect 3328 5355 3378 5455
rect 3536 5355 3586 5455
rect 3749 5355 3799 5455
rect 8401 5334 8451 5434
rect 8609 5334 8659 5434
rect 8817 5334 8867 5434
rect 9030 5334 9080 5434
rect 1421 5229 1471 5329
rect 1634 5229 1684 5329
rect 1842 5229 1892 5329
rect 2050 5229 2100 5329
rect 6702 5208 6752 5308
rect 6915 5208 6965 5308
rect 7123 5208 7173 5308
rect 7331 5208 7381 5308
rect 359 4990 409 5090
rect 572 4990 622 5090
rect 780 4990 830 5090
rect 988 4990 1038 5090
rect 4188 5028 4238 5128
rect 4396 5028 4446 5128
rect 4604 5028 4654 5128
rect 4817 5028 4867 5128
rect 1371 4809 1421 4909
rect 1584 4809 1634 4909
rect 1792 4809 1842 4909
rect 2000 4809 2050 4909
rect 5640 4969 5690 5069
rect 5853 4969 5903 5069
rect 6061 4969 6111 5069
rect 6269 4969 6319 5069
rect 9469 5007 9519 5107
rect 9677 5007 9727 5107
rect 9885 5007 9935 5107
rect 10098 5007 10148 5107
rect 3175 4794 3225 4894
rect 3383 4794 3433 4894
rect 3591 4794 3641 4894
rect 3804 4794 3854 4894
rect 6652 4788 6702 4888
rect 6865 4788 6915 4888
rect 7073 4788 7123 4888
rect 7281 4788 7331 4888
rect 358 4575 408 4675
rect 571 4575 621 4675
rect 779 4575 829 4675
rect 987 4575 1037 4675
rect 4187 4613 4237 4713
rect 4395 4613 4445 4713
rect 4603 4613 4653 4713
rect 4816 4613 4866 4713
rect 8456 4773 8506 4873
rect 8664 4773 8714 4873
rect 8872 4773 8922 4873
rect 9085 4773 9135 4873
rect 5639 4554 5689 4654
rect 5852 4554 5902 4654
rect 6060 4554 6110 4654
rect 6268 4554 6318 4654
rect 9468 4592 9518 4692
rect 9676 4592 9726 4692
rect 9884 4592 9934 4692
rect 10097 4592 10147 4692
rect 1669 4265 1719 4365
rect 1882 4265 1932 4365
rect 2090 4265 2140 4365
rect 2298 4265 2348 4365
rect 2880 4362 2930 4462
rect 3088 4362 3138 4462
rect 3296 4362 3346 4462
rect 3509 4362 3559 4462
rect 6950 4244 7000 4344
rect 7163 4244 7213 4344
rect 7371 4244 7421 4344
rect 7579 4244 7629 4344
rect 8161 4341 8211 4441
rect 8369 4341 8419 4441
rect 8577 4341 8627 4441
rect 8790 4341 8840 4441
rect 362 4014 412 4114
rect 575 4014 625 4114
rect 783 4014 833 4114
rect 991 4014 1041 4114
rect 4191 4052 4241 4152
rect 4399 4052 4449 4152
rect 4607 4052 4657 4152
rect 4820 4052 4870 4152
rect 1374 3833 1424 3933
rect 1587 3833 1637 3933
rect 1795 3833 1845 3933
rect 2003 3833 2053 3933
rect 5643 3993 5693 4093
rect 5856 3993 5906 4093
rect 6064 3993 6114 4093
rect 6272 3993 6322 4093
rect 9472 4031 9522 4131
rect 9680 4031 9730 4131
rect 9888 4031 9938 4131
rect 10101 4031 10151 4131
rect 3178 3818 3228 3918
rect 3386 3818 3436 3918
rect 3594 3818 3644 3918
rect 3807 3818 3857 3918
rect 6655 3812 6705 3912
rect 6868 3812 6918 3912
rect 7076 3812 7126 3912
rect 7284 3812 7334 3912
rect 361 3599 411 3699
rect 574 3599 624 3699
rect 782 3599 832 3699
rect 990 3599 1040 3699
rect 4190 3637 4240 3737
rect 4398 3637 4448 3737
rect 4606 3637 4656 3737
rect 4819 3637 4869 3737
rect 8459 3797 8509 3897
rect 8667 3797 8717 3897
rect 8875 3797 8925 3897
rect 9088 3797 9138 3897
rect 5642 3578 5692 3678
rect 5855 3578 5905 3678
rect 6063 3578 6113 3678
rect 6271 3578 6321 3678
rect 9471 3616 9521 3716
rect 9679 3616 9729 3716
rect 9887 3616 9937 3716
rect 10100 3616 10150 3716
rect 3128 3398 3178 3498
rect 3336 3398 3386 3498
rect 3544 3398 3594 3498
rect 3757 3398 3807 3498
rect 8409 3377 8459 3477
rect 8617 3377 8667 3477
rect 8825 3377 8875 3477
rect 9038 3377 9088 3477
rect 1429 3272 1479 3372
rect 1642 3272 1692 3372
rect 1850 3272 1900 3372
rect 2058 3272 2108 3372
rect 6710 3251 6760 3351
rect 6923 3251 6973 3351
rect 7131 3251 7181 3351
rect 7339 3251 7389 3351
rect 367 3033 417 3133
rect 580 3033 630 3133
rect 788 3033 838 3133
rect 996 3033 1046 3133
rect 4196 3071 4246 3171
rect 4404 3071 4454 3171
rect 4612 3071 4662 3171
rect 4825 3071 4875 3171
rect 1379 2852 1429 2952
rect 1592 2852 1642 2952
rect 1800 2852 1850 2952
rect 2008 2852 2058 2952
rect 5648 3012 5698 3112
rect 5861 3012 5911 3112
rect 6069 3012 6119 3112
rect 6277 3012 6327 3112
rect 9477 3050 9527 3150
rect 9685 3050 9735 3150
rect 9893 3050 9943 3150
rect 10106 3050 10156 3150
rect 3183 2837 3233 2937
rect 3391 2837 3441 2937
rect 3599 2837 3649 2937
rect 3812 2837 3862 2937
rect 6660 2831 6710 2931
rect 6873 2831 6923 2931
rect 7081 2831 7131 2931
rect 7289 2831 7339 2931
rect 366 2618 416 2718
rect 579 2618 629 2718
rect 787 2618 837 2718
rect 995 2618 1045 2718
rect 4195 2656 4245 2756
rect 4403 2656 4453 2756
rect 4611 2656 4661 2756
rect 4824 2656 4874 2756
rect 8464 2816 8514 2916
rect 8672 2816 8722 2916
rect 8880 2816 8930 2916
rect 9093 2816 9143 2916
rect 5647 2597 5697 2697
rect 5860 2597 5910 2697
rect 6068 2597 6118 2697
rect 6276 2597 6326 2697
rect 9476 2635 9526 2735
rect 9684 2635 9734 2735
rect 9892 2635 9942 2735
rect 10105 2635 10155 2735
rect 1594 2340 1644 2440
rect 1807 2340 1857 2440
rect 2015 2340 2065 2440
rect 2223 2340 2273 2440
rect 2975 2370 3025 2470
rect 3183 2370 3233 2470
rect 3391 2370 3441 2470
rect 3604 2370 3654 2470
rect 6875 2319 6925 2419
rect 7088 2319 7138 2419
rect 7296 2319 7346 2419
rect 7504 2319 7554 2419
rect 8256 2349 8306 2449
rect 8464 2349 8514 2449
rect 8672 2349 8722 2449
rect 8885 2349 8935 2449
rect 374 2054 424 2154
rect 587 2054 637 2154
rect 795 2054 845 2154
rect 1003 2054 1053 2154
rect 4203 2092 4253 2192
rect 4411 2092 4461 2192
rect 4619 2092 4669 2192
rect 4832 2092 4882 2192
rect 1386 1873 1436 1973
rect 1599 1873 1649 1973
rect 1807 1873 1857 1973
rect 2015 1873 2065 1973
rect 5655 2033 5705 2133
rect 5868 2033 5918 2133
rect 6076 2033 6126 2133
rect 6284 2033 6334 2133
rect 9484 2071 9534 2171
rect 9692 2071 9742 2171
rect 9900 2071 9950 2171
rect 10113 2071 10163 2171
rect 3190 1858 3240 1958
rect 3398 1858 3448 1958
rect 3606 1858 3656 1958
rect 3819 1858 3869 1958
rect 6667 1852 6717 1952
rect 6880 1852 6930 1952
rect 7088 1852 7138 1952
rect 7296 1852 7346 1952
rect 373 1639 423 1739
rect 586 1639 636 1739
rect 794 1639 844 1739
rect 1002 1639 1052 1739
rect 4202 1677 4252 1777
rect 4410 1677 4460 1777
rect 4618 1677 4668 1777
rect 4831 1677 4881 1777
rect 8471 1837 8521 1937
rect 8679 1837 8729 1937
rect 8887 1837 8937 1937
rect 9100 1837 9150 1937
rect 5654 1618 5704 1718
rect 5867 1618 5917 1718
rect 6075 1618 6125 1718
rect 6283 1618 6333 1718
rect 9483 1656 9533 1756
rect 9691 1656 9741 1756
rect 9899 1656 9949 1756
rect 10112 1656 10162 1756
rect 3140 1438 3190 1538
rect 3348 1438 3398 1538
rect 3556 1438 3606 1538
rect 3769 1438 3819 1538
rect 8421 1417 8471 1517
rect 8629 1417 8679 1517
rect 8837 1417 8887 1517
rect 9050 1417 9100 1517
rect 1441 1312 1491 1412
rect 1654 1312 1704 1412
rect 1862 1312 1912 1412
rect 2070 1312 2120 1412
rect 6722 1291 6772 1391
rect 6935 1291 6985 1391
rect 7143 1291 7193 1391
rect 7351 1291 7401 1391
rect 379 1073 429 1173
rect 592 1073 642 1173
rect 800 1073 850 1173
rect 1008 1073 1058 1173
rect 4208 1111 4258 1211
rect 4416 1111 4466 1211
rect 4624 1111 4674 1211
rect 4837 1111 4887 1211
rect 1391 892 1441 992
rect 1604 892 1654 992
rect 1812 892 1862 992
rect 2020 892 2070 992
rect 5660 1052 5710 1152
rect 5873 1052 5923 1152
rect 6081 1052 6131 1152
rect 6289 1052 6339 1152
rect 9489 1090 9539 1190
rect 9697 1090 9747 1190
rect 9905 1090 9955 1190
rect 10118 1090 10168 1190
rect 3195 877 3245 977
rect 3403 877 3453 977
rect 3611 877 3661 977
rect 3824 877 3874 977
rect 6672 871 6722 971
rect 6885 871 6935 971
rect 7093 871 7143 971
rect 7301 871 7351 971
rect 378 658 428 758
rect 591 658 641 758
rect 799 658 849 758
rect 1007 658 1057 758
rect 4207 696 4257 796
rect 4415 696 4465 796
rect 4623 696 4673 796
rect 4836 696 4886 796
rect 8476 856 8526 956
rect 8684 856 8734 956
rect 8892 856 8942 956
rect 9105 856 9155 956
rect 5659 637 5709 737
rect 5872 637 5922 737
rect 6080 637 6130 737
rect 6288 637 6338 737
rect 9488 675 9538 775
rect 9696 675 9746 775
rect 9904 675 9954 775
rect 10117 675 10167 775
rect 1781 177 1831 277
rect 1994 177 2044 277
rect 2202 177 2252 277
rect 2410 177 2460 277
rect 4871 89 4921 189
rect 5084 89 5134 189
rect 5292 89 5342 189
rect 5500 89 5550 189
rect 7062 156 7112 256
rect 7275 156 7325 256
rect 7483 156 7533 256
rect 7691 156 7741 256
<< ndiff >>
rect 4122 8176 4171 8188
rect 4122 8156 4133 8176
rect 4153 8156 4171 8176
rect 4122 8146 4171 8156
rect 4221 8172 4265 8188
rect 4221 8152 4236 8172
rect 4256 8152 4265 8172
rect 4221 8146 4265 8152
rect 4335 8172 4379 8188
rect 4335 8152 4344 8172
rect 4364 8152 4379 8172
rect 4335 8146 4379 8152
rect 4429 8176 4478 8188
rect 4429 8156 4447 8176
rect 4467 8156 4478 8176
rect 4429 8146 4478 8156
rect 4543 8172 4587 8188
rect 4543 8152 4552 8172
rect 4572 8152 4587 8172
rect 4543 8146 4587 8152
rect 4637 8176 4686 8188
rect 4637 8156 4655 8176
rect 4675 8156 4686 8176
rect 4637 8146 4686 8156
rect 4756 8172 4800 8188
rect 4756 8152 4765 8172
rect 4785 8152 4800 8172
rect 4756 8146 4800 8152
rect 4850 8176 4899 8188
rect 4850 8156 4868 8176
rect 4888 8156 4899 8176
rect 4850 8146 4899 8156
rect 9403 8155 9452 8167
rect 9403 8135 9414 8155
rect 9434 8135 9452 8155
rect 9403 8125 9452 8135
rect 9502 8151 9546 8167
rect 9502 8131 9517 8151
rect 9537 8131 9546 8151
rect 9502 8125 9546 8131
rect 9616 8151 9660 8167
rect 9616 8131 9625 8151
rect 9645 8131 9660 8151
rect 9616 8125 9660 8131
rect 9710 8155 9759 8167
rect 9710 8135 9728 8155
rect 9748 8135 9759 8155
rect 9710 8125 9759 8135
rect 9824 8151 9868 8167
rect 9824 8131 9833 8151
rect 9853 8131 9868 8151
rect 9824 8125 9868 8131
rect 9918 8155 9967 8167
rect 9918 8135 9936 8155
rect 9956 8135 9967 8155
rect 9918 8125 9967 8135
rect 10037 8151 10081 8167
rect 10037 8131 10046 8151
rect 10066 8131 10081 8151
rect 10037 8125 10081 8131
rect 10131 8155 10180 8167
rect 10131 8135 10149 8155
rect 10169 8135 10180 8155
rect 10131 8125 10180 8135
rect 3109 7942 3158 7954
rect 3109 7922 3120 7942
rect 3140 7922 3158 7942
rect 3109 7912 3158 7922
rect 3208 7938 3252 7954
rect 3208 7918 3223 7938
rect 3243 7918 3252 7938
rect 3208 7912 3252 7918
rect 3322 7938 3366 7954
rect 3322 7918 3331 7938
rect 3351 7918 3366 7938
rect 3322 7912 3366 7918
rect 3416 7942 3465 7954
rect 3416 7922 3434 7942
rect 3454 7922 3465 7942
rect 3416 7912 3465 7922
rect 3530 7938 3574 7954
rect 3530 7918 3539 7938
rect 3559 7918 3574 7938
rect 3530 7912 3574 7918
rect 3624 7942 3673 7954
rect 3624 7922 3642 7942
rect 3662 7922 3673 7942
rect 3624 7912 3673 7922
rect 3743 7938 3787 7954
rect 3743 7918 3752 7938
rect 3772 7918 3787 7938
rect 3743 7912 3787 7918
rect 3837 7942 3886 7954
rect 3837 7922 3855 7942
rect 3875 7922 3886 7942
rect 3837 7912 3886 7922
rect 293 7844 342 7854
rect 293 7824 304 7844
rect 324 7824 342 7844
rect 293 7812 342 7824
rect 392 7848 436 7854
rect 392 7828 407 7848
rect 427 7828 436 7848
rect 392 7812 436 7828
rect 506 7844 555 7854
rect 506 7824 517 7844
rect 537 7824 555 7844
rect 506 7812 555 7824
rect 605 7848 649 7854
rect 605 7828 620 7848
rect 640 7828 649 7848
rect 605 7812 649 7828
rect 714 7844 763 7854
rect 714 7824 725 7844
rect 745 7824 763 7844
rect 714 7812 763 7824
rect 813 7848 857 7854
rect 813 7828 828 7848
rect 848 7828 857 7848
rect 813 7812 857 7828
rect 927 7848 971 7854
rect 927 7828 936 7848
rect 956 7828 971 7848
rect 927 7812 971 7828
rect 1021 7844 1070 7854
rect 1021 7824 1039 7844
rect 1059 7824 1070 7844
rect 1021 7812 1070 7824
rect 8390 7921 8439 7933
rect 8390 7901 8401 7921
rect 8421 7901 8439 7921
rect 8390 7891 8439 7901
rect 8489 7917 8533 7933
rect 8489 7897 8504 7917
rect 8524 7897 8533 7917
rect 8489 7891 8533 7897
rect 8603 7917 8647 7933
rect 8603 7897 8612 7917
rect 8632 7897 8647 7917
rect 8603 7891 8647 7897
rect 8697 7921 8746 7933
rect 8697 7901 8715 7921
rect 8735 7901 8746 7921
rect 8697 7891 8746 7901
rect 8811 7917 8855 7933
rect 8811 7897 8820 7917
rect 8840 7897 8855 7917
rect 8811 7891 8855 7897
rect 8905 7921 8954 7933
rect 8905 7901 8923 7921
rect 8943 7901 8954 7921
rect 8905 7891 8954 7901
rect 9024 7917 9068 7933
rect 9024 7897 9033 7917
rect 9053 7897 9068 7917
rect 9024 7891 9068 7897
rect 9118 7921 9167 7933
rect 9118 7901 9136 7921
rect 9156 7901 9167 7921
rect 9118 7891 9167 7901
rect 5574 7823 5623 7833
rect 5574 7803 5585 7823
rect 5605 7803 5623 7823
rect 5574 7791 5623 7803
rect 5673 7827 5717 7833
rect 5673 7807 5688 7827
rect 5708 7807 5717 7827
rect 5673 7791 5717 7807
rect 5787 7823 5836 7833
rect 5787 7803 5798 7823
rect 5818 7803 5836 7823
rect 5787 7791 5836 7803
rect 5886 7827 5930 7833
rect 5886 7807 5901 7827
rect 5921 7807 5930 7827
rect 5886 7791 5930 7807
rect 5995 7823 6044 7833
rect 5995 7803 6006 7823
rect 6026 7803 6044 7823
rect 5995 7791 6044 7803
rect 6094 7827 6138 7833
rect 6094 7807 6109 7827
rect 6129 7807 6138 7827
rect 6094 7791 6138 7807
rect 6208 7827 6252 7833
rect 6208 7807 6217 7827
rect 6237 7807 6252 7827
rect 6208 7791 6252 7807
rect 6302 7823 6351 7833
rect 6302 7803 6320 7823
rect 6340 7803 6351 7823
rect 6302 7791 6351 7803
rect 4121 7761 4170 7773
rect 4121 7741 4132 7761
rect 4152 7741 4170 7761
rect 4121 7731 4170 7741
rect 4220 7757 4264 7773
rect 4220 7737 4235 7757
rect 4255 7737 4264 7757
rect 4220 7731 4264 7737
rect 4334 7757 4378 7773
rect 4334 7737 4343 7757
rect 4363 7737 4378 7757
rect 4334 7731 4378 7737
rect 4428 7761 4477 7773
rect 4428 7741 4446 7761
rect 4466 7741 4477 7761
rect 4428 7731 4477 7741
rect 4542 7757 4586 7773
rect 4542 7737 4551 7757
rect 4571 7737 4586 7757
rect 4542 7731 4586 7737
rect 4636 7761 4685 7773
rect 4636 7741 4654 7761
rect 4674 7741 4685 7761
rect 4636 7731 4685 7741
rect 4755 7757 4799 7773
rect 4755 7737 4764 7757
rect 4784 7737 4799 7757
rect 4755 7731 4799 7737
rect 4849 7761 4898 7773
rect 4849 7741 4867 7761
rect 4887 7741 4898 7761
rect 4849 7731 4898 7741
rect 1305 7663 1354 7673
rect 1305 7643 1316 7663
rect 1336 7643 1354 7663
rect 1305 7631 1354 7643
rect 1404 7667 1448 7673
rect 1404 7647 1419 7667
rect 1439 7647 1448 7667
rect 1404 7631 1448 7647
rect 1518 7663 1567 7673
rect 1518 7643 1529 7663
rect 1549 7643 1567 7663
rect 1518 7631 1567 7643
rect 1617 7667 1661 7673
rect 1617 7647 1632 7667
rect 1652 7647 1661 7667
rect 1617 7631 1661 7647
rect 1726 7663 1775 7673
rect 1726 7643 1737 7663
rect 1757 7643 1775 7663
rect 1726 7631 1775 7643
rect 1825 7667 1869 7673
rect 1825 7647 1840 7667
rect 1860 7647 1869 7667
rect 1825 7631 1869 7647
rect 1939 7667 1983 7673
rect 1939 7647 1948 7667
rect 1968 7647 1983 7667
rect 1939 7631 1983 7647
rect 2033 7663 2082 7673
rect 2033 7643 2051 7663
rect 2071 7643 2082 7663
rect 2033 7631 2082 7643
rect 9402 7740 9451 7752
rect 9402 7720 9413 7740
rect 9433 7720 9451 7740
rect 9402 7710 9451 7720
rect 9501 7736 9545 7752
rect 9501 7716 9516 7736
rect 9536 7716 9545 7736
rect 9501 7710 9545 7716
rect 9615 7736 9659 7752
rect 9615 7716 9624 7736
rect 9644 7716 9659 7736
rect 9615 7710 9659 7716
rect 9709 7740 9758 7752
rect 9709 7720 9727 7740
rect 9747 7720 9758 7740
rect 9709 7710 9758 7720
rect 9823 7736 9867 7752
rect 9823 7716 9832 7736
rect 9852 7716 9867 7736
rect 9823 7710 9867 7716
rect 9917 7740 9966 7752
rect 9917 7720 9935 7740
rect 9955 7720 9966 7740
rect 9917 7710 9966 7720
rect 10036 7736 10080 7752
rect 10036 7716 10045 7736
rect 10065 7716 10080 7736
rect 10036 7710 10080 7716
rect 10130 7740 10179 7752
rect 10130 7720 10148 7740
rect 10168 7720 10179 7740
rect 10130 7710 10179 7720
rect 6586 7642 6635 7652
rect 6586 7622 6597 7642
rect 6617 7622 6635 7642
rect 6586 7610 6635 7622
rect 6685 7646 6729 7652
rect 6685 7626 6700 7646
rect 6720 7626 6729 7646
rect 6685 7610 6729 7626
rect 6799 7642 6848 7652
rect 6799 7622 6810 7642
rect 6830 7622 6848 7642
rect 6799 7610 6848 7622
rect 6898 7646 6942 7652
rect 6898 7626 6913 7646
rect 6933 7626 6942 7646
rect 6898 7610 6942 7626
rect 7007 7642 7056 7652
rect 7007 7622 7018 7642
rect 7038 7622 7056 7642
rect 7007 7610 7056 7622
rect 7106 7646 7150 7652
rect 7106 7626 7121 7646
rect 7141 7626 7150 7646
rect 7106 7610 7150 7626
rect 7220 7646 7264 7652
rect 7220 7626 7229 7646
rect 7249 7626 7264 7646
rect 7220 7610 7264 7626
rect 7314 7642 7363 7652
rect 7314 7622 7332 7642
rect 7352 7622 7363 7642
rect 7314 7610 7363 7622
rect 3059 7522 3108 7534
rect 3059 7502 3070 7522
rect 3090 7502 3108 7522
rect 3059 7492 3108 7502
rect 3158 7518 3202 7534
rect 3158 7498 3173 7518
rect 3193 7498 3202 7518
rect 3158 7492 3202 7498
rect 3272 7518 3316 7534
rect 3272 7498 3281 7518
rect 3301 7498 3316 7518
rect 3272 7492 3316 7498
rect 3366 7522 3415 7534
rect 3366 7502 3384 7522
rect 3404 7502 3415 7522
rect 3366 7492 3415 7502
rect 3480 7518 3524 7534
rect 3480 7498 3489 7518
rect 3509 7498 3524 7518
rect 3480 7492 3524 7498
rect 3574 7522 3623 7534
rect 3574 7502 3592 7522
rect 3612 7502 3623 7522
rect 3574 7492 3623 7502
rect 3693 7518 3737 7534
rect 3693 7498 3702 7518
rect 3722 7498 3737 7518
rect 3693 7492 3737 7498
rect 3787 7522 3836 7534
rect 3787 7502 3805 7522
rect 3825 7502 3836 7522
rect 3787 7492 3836 7502
rect 292 7429 341 7439
rect 292 7409 303 7429
rect 323 7409 341 7429
rect 292 7397 341 7409
rect 391 7433 435 7439
rect 391 7413 406 7433
rect 426 7413 435 7433
rect 391 7397 435 7413
rect 505 7429 554 7439
rect 505 7409 516 7429
rect 536 7409 554 7429
rect 505 7397 554 7409
rect 604 7433 648 7439
rect 604 7413 619 7433
rect 639 7413 648 7433
rect 604 7397 648 7413
rect 713 7429 762 7439
rect 713 7409 724 7429
rect 744 7409 762 7429
rect 713 7397 762 7409
rect 812 7433 856 7439
rect 812 7413 827 7433
rect 847 7413 856 7433
rect 812 7397 856 7413
rect 926 7433 970 7439
rect 926 7413 935 7433
rect 955 7413 970 7433
rect 926 7397 970 7413
rect 1020 7429 1069 7439
rect 1020 7409 1038 7429
rect 1058 7409 1069 7429
rect 8340 7501 8389 7513
rect 1020 7397 1069 7409
rect 8340 7481 8351 7501
rect 8371 7481 8389 7501
rect 8340 7471 8389 7481
rect 8439 7497 8483 7513
rect 8439 7477 8454 7497
rect 8474 7477 8483 7497
rect 8439 7471 8483 7477
rect 8553 7497 8597 7513
rect 8553 7477 8562 7497
rect 8582 7477 8597 7497
rect 8553 7471 8597 7477
rect 8647 7501 8696 7513
rect 8647 7481 8665 7501
rect 8685 7481 8696 7501
rect 8647 7471 8696 7481
rect 8761 7497 8805 7513
rect 8761 7477 8770 7497
rect 8790 7477 8805 7497
rect 8761 7471 8805 7477
rect 8855 7501 8904 7513
rect 8855 7481 8873 7501
rect 8893 7481 8904 7501
rect 8855 7471 8904 7481
rect 8974 7497 9018 7513
rect 8974 7477 8983 7497
rect 9003 7477 9018 7497
rect 8974 7471 9018 7477
rect 9068 7501 9117 7513
rect 9068 7481 9086 7501
rect 9106 7481 9117 7501
rect 9068 7471 9117 7481
rect 5573 7408 5622 7418
rect 5573 7388 5584 7408
rect 5604 7388 5622 7408
rect 5573 7376 5622 7388
rect 5672 7412 5716 7418
rect 5672 7392 5687 7412
rect 5707 7392 5716 7412
rect 5672 7376 5716 7392
rect 5786 7408 5835 7418
rect 5786 7388 5797 7408
rect 5817 7388 5835 7408
rect 5786 7376 5835 7388
rect 5885 7412 5929 7418
rect 5885 7392 5900 7412
rect 5920 7392 5929 7412
rect 5885 7376 5929 7392
rect 5994 7408 6043 7418
rect 5994 7388 6005 7408
rect 6025 7388 6043 7408
rect 5994 7376 6043 7388
rect 6093 7412 6137 7418
rect 6093 7392 6108 7412
rect 6128 7392 6137 7412
rect 6093 7376 6137 7392
rect 6207 7412 6251 7418
rect 6207 7392 6216 7412
rect 6236 7392 6251 7412
rect 6207 7376 6251 7392
rect 6301 7408 6350 7418
rect 6301 7388 6319 7408
rect 6339 7388 6350 7408
rect 6301 7376 6350 7388
rect 4127 7195 4176 7207
rect 4127 7175 4138 7195
rect 4158 7175 4176 7195
rect 4127 7165 4176 7175
rect 4226 7191 4270 7207
rect 4226 7171 4241 7191
rect 4261 7171 4270 7191
rect 4226 7165 4270 7171
rect 4340 7191 4384 7207
rect 4340 7171 4349 7191
rect 4369 7171 4384 7191
rect 4340 7165 4384 7171
rect 4434 7195 4483 7207
rect 4434 7175 4452 7195
rect 4472 7175 4483 7195
rect 4434 7165 4483 7175
rect 4548 7191 4592 7207
rect 4548 7171 4557 7191
rect 4577 7171 4592 7191
rect 4548 7165 4592 7171
rect 4642 7195 4691 7207
rect 4642 7175 4660 7195
rect 4680 7175 4691 7195
rect 4642 7165 4691 7175
rect 4761 7191 4805 7207
rect 4761 7171 4770 7191
rect 4790 7171 4805 7191
rect 4761 7165 4805 7171
rect 4855 7195 4904 7207
rect 4855 7175 4873 7195
rect 4893 7175 4904 7195
rect 4855 7165 4904 7175
rect 1360 7102 1409 7112
rect 1360 7082 1371 7102
rect 1391 7082 1409 7102
rect 1360 7070 1409 7082
rect 1459 7106 1503 7112
rect 1459 7086 1474 7106
rect 1494 7086 1503 7106
rect 1459 7070 1503 7086
rect 1573 7102 1622 7112
rect 1573 7082 1584 7102
rect 1604 7082 1622 7102
rect 1573 7070 1622 7082
rect 1672 7106 1716 7112
rect 1672 7086 1687 7106
rect 1707 7086 1716 7106
rect 1672 7070 1716 7086
rect 1781 7102 1830 7112
rect 1781 7082 1792 7102
rect 1812 7082 1830 7102
rect 1781 7070 1830 7082
rect 1880 7106 1924 7112
rect 1880 7086 1895 7106
rect 1915 7086 1924 7106
rect 1880 7070 1924 7086
rect 1994 7106 2038 7112
rect 1994 7086 2003 7106
rect 2023 7086 2038 7106
rect 1994 7070 2038 7086
rect 2088 7102 2137 7112
rect 2088 7082 2106 7102
rect 2126 7082 2137 7102
rect 9408 7174 9457 7186
rect 2088 7070 2137 7082
rect 9408 7154 9419 7174
rect 9439 7154 9457 7174
rect 9408 7144 9457 7154
rect 9507 7170 9551 7186
rect 9507 7150 9522 7170
rect 9542 7150 9551 7170
rect 9507 7144 9551 7150
rect 9621 7170 9665 7186
rect 9621 7150 9630 7170
rect 9650 7150 9665 7170
rect 9621 7144 9665 7150
rect 9715 7174 9764 7186
rect 9715 7154 9733 7174
rect 9753 7154 9764 7174
rect 9715 7144 9764 7154
rect 9829 7170 9873 7186
rect 9829 7150 9838 7170
rect 9858 7150 9873 7170
rect 9829 7144 9873 7150
rect 9923 7174 9972 7186
rect 9923 7154 9941 7174
rect 9961 7154 9972 7174
rect 9923 7144 9972 7154
rect 10042 7170 10086 7186
rect 10042 7150 10051 7170
rect 10071 7150 10086 7170
rect 10042 7144 10086 7150
rect 10136 7174 10185 7186
rect 10136 7154 10154 7174
rect 10174 7154 10185 7174
rect 10136 7144 10185 7154
rect 6641 7081 6690 7091
rect 6641 7061 6652 7081
rect 6672 7061 6690 7081
rect 6641 7049 6690 7061
rect 6740 7085 6784 7091
rect 6740 7065 6755 7085
rect 6775 7065 6784 7085
rect 6740 7049 6784 7065
rect 6854 7081 6903 7091
rect 6854 7061 6865 7081
rect 6885 7061 6903 7081
rect 6854 7049 6903 7061
rect 6953 7085 6997 7091
rect 6953 7065 6968 7085
rect 6988 7065 6997 7085
rect 6953 7049 6997 7065
rect 7062 7081 7111 7091
rect 7062 7061 7073 7081
rect 7093 7061 7111 7081
rect 7062 7049 7111 7061
rect 7161 7085 7205 7091
rect 7161 7065 7176 7085
rect 7196 7065 7205 7085
rect 7161 7049 7205 7065
rect 7275 7085 7319 7091
rect 7275 7065 7284 7085
rect 7304 7065 7319 7085
rect 7275 7049 7319 7065
rect 7369 7081 7418 7091
rect 7369 7061 7387 7081
rect 7407 7061 7418 7081
rect 7369 7049 7418 7061
rect 3114 6961 3163 6973
rect 3114 6941 3125 6961
rect 3145 6941 3163 6961
rect 3114 6931 3163 6941
rect 3213 6957 3257 6973
rect 3213 6937 3228 6957
rect 3248 6937 3257 6957
rect 3213 6931 3257 6937
rect 3327 6957 3371 6973
rect 3327 6937 3336 6957
rect 3356 6937 3371 6957
rect 3327 6931 3371 6937
rect 3421 6961 3470 6973
rect 3421 6941 3439 6961
rect 3459 6941 3470 6961
rect 3421 6931 3470 6941
rect 3535 6957 3579 6973
rect 3535 6937 3544 6957
rect 3564 6937 3579 6957
rect 3535 6931 3579 6937
rect 3629 6961 3678 6973
rect 3629 6941 3647 6961
rect 3667 6941 3678 6961
rect 3629 6931 3678 6941
rect 3748 6957 3792 6973
rect 3748 6937 3757 6957
rect 3777 6937 3792 6957
rect 3748 6931 3792 6937
rect 3842 6961 3891 6973
rect 3842 6941 3860 6961
rect 3880 6941 3891 6961
rect 3842 6931 3891 6941
rect 298 6863 347 6873
rect 298 6843 309 6863
rect 329 6843 347 6863
rect 298 6831 347 6843
rect 397 6867 441 6873
rect 397 6847 412 6867
rect 432 6847 441 6867
rect 397 6831 441 6847
rect 511 6863 560 6873
rect 511 6843 522 6863
rect 542 6843 560 6863
rect 511 6831 560 6843
rect 610 6867 654 6873
rect 610 6847 625 6867
rect 645 6847 654 6867
rect 610 6831 654 6847
rect 719 6863 768 6873
rect 719 6843 730 6863
rect 750 6843 768 6863
rect 719 6831 768 6843
rect 818 6867 862 6873
rect 818 6847 833 6867
rect 853 6847 862 6867
rect 818 6831 862 6847
rect 932 6867 976 6873
rect 932 6847 941 6867
rect 961 6847 976 6867
rect 932 6831 976 6847
rect 1026 6863 1075 6873
rect 1026 6843 1044 6863
rect 1064 6843 1075 6863
rect 1026 6831 1075 6843
rect 8395 6940 8444 6952
rect 8395 6920 8406 6940
rect 8426 6920 8444 6940
rect 8395 6910 8444 6920
rect 8494 6936 8538 6952
rect 8494 6916 8509 6936
rect 8529 6916 8538 6936
rect 8494 6910 8538 6916
rect 8608 6936 8652 6952
rect 8608 6916 8617 6936
rect 8637 6916 8652 6936
rect 8608 6910 8652 6916
rect 8702 6940 8751 6952
rect 8702 6920 8720 6940
rect 8740 6920 8751 6940
rect 8702 6910 8751 6920
rect 8816 6936 8860 6952
rect 8816 6916 8825 6936
rect 8845 6916 8860 6936
rect 8816 6910 8860 6916
rect 8910 6940 8959 6952
rect 8910 6920 8928 6940
rect 8948 6920 8959 6940
rect 8910 6910 8959 6920
rect 9029 6936 9073 6952
rect 9029 6916 9038 6936
rect 9058 6916 9073 6936
rect 9029 6910 9073 6916
rect 9123 6940 9172 6952
rect 9123 6920 9141 6940
rect 9161 6920 9172 6940
rect 9123 6910 9172 6920
rect 5579 6842 5628 6852
rect 5579 6822 5590 6842
rect 5610 6822 5628 6842
rect 5579 6810 5628 6822
rect 5678 6846 5722 6852
rect 5678 6826 5693 6846
rect 5713 6826 5722 6846
rect 5678 6810 5722 6826
rect 5792 6842 5841 6852
rect 5792 6822 5803 6842
rect 5823 6822 5841 6842
rect 5792 6810 5841 6822
rect 5891 6846 5935 6852
rect 5891 6826 5906 6846
rect 5926 6826 5935 6846
rect 5891 6810 5935 6826
rect 6000 6842 6049 6852
rect 6000 6822 6011 6842
rect 6031 6822 6049 6842
rect 6000 6810 6049 6822
rect 6099 6846 6143 6852
rect 6099 6826 6114 6846
rect 6134 6826 6143 6846
rect 6099 6810 6143 6826
rect 6213 6846 6257 6852
rect 6213 6826 6222 6846
rect 6242 6826 6257 6846
rect 6213 6810 6257 6826
rect 6307 6842 6356 6852
rect 6307 6822 6325 6842
rect 6345 6822 6356 6842
rect 6307 6810 6356 6822
rect 4126 6780 4175 6792
rect 4126 6760 4137 6780
rect 4157 6760 4175 6780
rect 4126 6750 4175 6760
rect 4225 6776 4269 6792
rect 4225 6756 4240 6776
rect 4260 6756 4269 6776
rect 4225 6750 4269 6756
rect 4339 6776 4383 6792
rect 4339 6756 4348 6776
rect 4368 6756 4383 6776
rect 4339 6750 4383 6756
rect 4433 6780 4482 6792
rect 4433 6760 4451 6780
rect 4471 6760 4482 6780
rect 4433 6750 4482 6760
rect 4547 6776 4591 6792
rect 4547 6756 4556 6776
rect 4576 6756 4591 6776
rect 4547 6750 4591 6756
rect 4641 6780 4690 6792
rect 4641 6760 4659 6780
rect 4679 6760 4690 6780
rect 4641 6750 4690 6760
rect 4760 6776 4804 6792
rect 4760 6756 4769 6776
rect 4789 6756 4804 6776
rect 4760 6750 4804 6756
rect 4854 6780 4903 6792
rect 4854 6760 4872 6780
rect 4892 6760 4903 6780
rect 4854 6750 4903 6760
rect 1310 6682 1359 6692
rect 1310 6662 1321 6682
rect 1341 6662 1359 6682
rect 1310 6650 1359 6662
rect 1409 6686 1453 6692
rect 1409 6666 1424 6686
rect 1444 6666 1453 6686
rect 1409 6650 1453 6666
rect 1523 6682 1572 6692
rect 1523 6662 1534 6682
rect 1554 6662 1572 6682
rect 1523 6650 1572 6662
rect 1622 6686 1666 6692
rect 1622 6666 1637 6686
rect 1657 6666 1666 6686
rect 1622 6650 1666 6666
rect 1731 6682 1780 6692
rect 1731 6662 1742 6682
rect 1762 6662 1780 6682
rect 1731 6650 1780 6662
rect 1830 6686 1874 6692
rect 1830 6666 1845 6686
rect 1865 6666 1874 6686
rect 1830 6650 1874 6666
rect 1944 6686 1988 6692
rect 1944 6666 1953 6686
rect 1973 6666 1988 6686
rect 1944 6650 1988 6666
rect 2038 6682 2087 6692
rect 2038 6662 2056 6682
rect 2076 6662 2087 6682
rect 2038 6650 2087 6662
rect 9407 6759 9456 6771
rect 9407 6739 9418 6759
rect 9438 6739 9456 6759
rect 9407 6729 9456 6739
rect 9506 6755 9550 6771
rect 9506 6735 9521 6755
rect 9541 6735 9550 6755
rect 9506 6729 9550 6735
rect 9620 6755 9664 6771
rect 9620 6735 9629 6755
rect 9649 6735 9664 6755
rect 9620 6729 9664 6735
rect 9714 6759 9763 6771
rect 9714 6739 9732 6759
rect 9752 6739 9763 6759
rect 9714 6729 9763 6739
rect 9828 6755 9872 6771
rect 9828 6735 9837 6755
rect 9857 6735 9872 6755
rect 9828 6729 9872 6735
rect 9922 6759 9971 6771
rect 9922 6739 9940 6759
rect 9960 6739 9971 6759
rect 9922 6729 9971 6739
rect 10041 6755 10085 6771
rect 10041 6735 10050 6755
rect 10070 6735 10085 6755
rect 10041 6729 10085 6735
rect 10135 6759 10184 6771
rect 10135 6739 10153 6759
rect 10173 6739 10184 6759
rect 10135 6729 10184 6739
rect 6591 6661 6640 6671
rect 6591 6641 6602 6661
rect 6622 6641 6640 6661
rect 6591 6629 6640 6641
rect 6690 6665 6734 6671
rect 6690 6645 6705 6665
rect 6725 6645 6734 6665
rect 6690 6629 6734 6645
rect 6804 6661 6853 6671
rect 6804 6641 6815 6661
rect 6835 6641 6853 6661
rect 6804 6629 6853 6641
rect 6903 6665 6947 6671
rect 6903 6645 6918 6665
rect 6938 6645 6947 6665
rect 6903 6629 6947 6645
rect 7012 6661 7061 6671
rect 7012 6641 7023 6661
rect 7043 6641 7061 6661
rect 7012 6629 7061 6641
rect 7111 6665 7155 6671
rect 7111 6645 7126 6665
rect 7146 6645 7155 6665
rect 7111 6629 7155 6645
rect 7225 6665 7269 6671
rect 7225 6645 7234 6665
rect 7254 6645 7269 6665
rect 7225 6629 7269 6645
rect 7319 6661 7368 6671
rect 7319 6641 7337 6661
rect 7357 6641 7368 6661
rect 7319 6629 7368 6641
rect 2906 6494 2955 6506
rect 2906 6474 2917 6494
rect 2937 6474 2955 6494
rect 2906 6464 2955 6474
rect 3005 6490 3049 6506
rect 3005 6470 3020 6490
rect 3040 6470 3049 6490
rect 3005 6464 3049 6470
rect 3119 6490 3163 6506
rect 3119 6470 3128 6490
rect 3148 6470 3163 6490
rect 3119 6464 3163 6470
rect 3213 6494 3262 6506
rect 3213 6474 3231 6494
rect 3251 6474 3262 6494
rect 3213 6464 3262 6474
rect 3327 6490 3371 6506
rect 3327 6470 3336 6490
rect 3356 6470 3371 6490
rect 3327 6464 3371 6470
rect 3421 6494 3470 6506
rect 3421 6474 3439 6494
rect 3459 6474 3470 6494
rect 3421 6464 3470 6474
rect 3540 6490 3584 6506
rect 3540 6470 3549 6490
rect 3569 6470 3584 6490
rect 3540 6464 3584 6470
rect 3634 6494 3683 6506
rect 3634 6474 3652 6494
rect 3672 6474 3683 6494
rect 3634 6464 3683 6474
rect 297 6448 346 6458
rect 297 6428 308 6448
rect 328 6428 346 6448
rect 297 6416 346 6428
rect 396 6452 440 6458
rect 396 6432 411 6452
rect 431 6432 440 6452
rect 396 6416 440 6432
rect 510 6448 559 6458
rect 510 6428 521 6448
rect 541 6428 559 6448
rect 510 6416 559 6428
rect 609 6452 653 6458
rect 609 6432 624 6452
rect 644 6432 653 6452
rect 609 6416 653 6432
rect 718 6448 767 6458
rect 718 6428 729 6448
rect 749 6428 767 6448
rect 718 6416 767 6428
rect 817 6452 861 6458
rect 817 6432 832 6452
rect 852 6432 861 6452
rect 817 6416 861 6432
rect 931 6452 975 6458
rect 931 6432 940 6452
rect 960 6432 975 6452
rect 931 6416 975 6432
rect 1025 6448 1074 6458
rect 1025 6428 1043 6448
rect 1063 6428 1074 6448
rect 1025 6416 1074 6428
rect 8187 6473 8236 6485
rect 8187 6453 8198 6473
rect 8218 6453 8236 6473
rect 8187 6443 8236 6453
rect 8286 6469 8330 6485
rect 8286 6449 8301 6469
rect 8321 6449 8330 6469
rect 8286 6443 8330 6449
rect 8400 6469 8444 6485
rect 8400 6449 8409 6469
rect 8429 6449 8444 6469
rect 8400 6443 8444 6449
rect 8494 6473 8543 6485
rect 8494 6453 8512 6473
rect 8532 6453 8543 6473
rect 8494 6443 8543 6453
rect 8608 6469 8652 6485
rect 8608 6449 8617 6469
rect 8637 6449 8652 6469
rect 8608 6443 8652 6449
rect 8702 6473 8751 6485
rect 8702 6453 8720 6473
rect 8740 6453 8751 6473
rect 8702 6443 8751 6453
rect 8821 6469 8865 6485
rect 8821 6449 8830 6469
rect 8850 6449 8865 6469
rect 8821 6443 8865 6449
rect 8915 6473 8964 6485
rect 8915 6453 8933 6473
rect 8953 6453 8964 6473
rect 8915 6443 8964 6453
rect 5578 6427 5627 6437
rect 5578 6407 5589 6427
rect 5609 6407 5627 6427
rect 5578 6395 5627 6407
rect 5677 6431 5721 6437
rect 5677 6411 5692 6431
rect 5712 6411 5721 6431
rect 5677 6395 5721 6411
rect 5791 6427 5840 6437
rect 5791 6407 5802 6427
rect 5822 6407 5840 6427
rect 5791 6395 5840 6407
rect 5890 6431 5934 6437
rect 5890 6411 5905 6431
rect 5925 6411 5934 6431
rect 5890 6395 5934 6411
rect 5999 6427 6048 6437
rect 5999 6407 6010 6427
rect 6030 6407 6048 6427
rect 5999 6395 6048 6407
rect 6098 6431 6142 6437
rect 6098 6411 6113 6431
rect 6133 6411 6142 6431
rect 6098 6395 6142 6411
rect 6212 6431 6256 6437
rect 6212 6411 6221 6431
rect 6241 6411 6256 6431
rect 6212 6395 6256 6411
rect 6306 6427 6355 6437
rect 6306 6407 6324 6427
rect 6344 6407 6355 6427
rect 6306 6395 6355 6407
rect 4134 6216 4183 6228
rect 4134 6196 4145 6216
rect 4165 6196 4183 6216
rect 4134 6186 4183 6196
rect 4233 6212 4277 6228
rect 4233 6192 4248 6212
rect 4268 6192 4277 6212
rect 4233 6186 4277 6192
rect 4347 6212 4391 6228
rect 4347 6192 4356 6212
rect 4376 6192 4391 6212
rect 4347 6186 4391 6192
rect 4441 6216 4490 6228
rect 4441 6196 4459 6216
rect 4479 6196 4490 6216
rect 4441 6186 4490 6196
rect 4555 6212 4599 6228
rect 4555 6192 4564 6212
rect 4584 6192 4599 6212
rect 4555 6186 4599 6192
rect 4649 6216 4698 6228
rect 4649 6196 4667 6216
rect 4687 6196 4698 6216
rect 4649 6186 4698 6196
rect 4768 6212 4812 6228
rect 4768 6192 4777 6212
rect 4797 6192 4812 6212
rect 4768 6186 4812 6192
rect 4862 6216 4911 6228
rect 4862 6196 4880 6216
rect 4900 6196 4911 6216
rect 4862 6186 4911 6196
rect 1525 6170 1574 6180
rect 1525 6150 1536 6170
rect 1556 6150 1574 6170
rect 1525 6138 1574 6150
rect 1624 6174 1668 6180
rect 1624 6154 1639 6174
rect 1659 6154 1668 6174
rect 1624 6138 1668 6154
rect 1738 6170 1787 6180
rect 1738 6150 1749 6170
rect 1769 6150 1787 6170
rect 1738 6138 1787 6150
rect 1837 6174 1881 6180
rect 1837 6154 1852 6174
rect 1872 6154 1881 6174
rect 1837 6138 1881 6154
rect 1946 6170 1995 6180
rect 1946 6150 1957 6170
rect 1977 6150 1995 6170
rect 1946 6138 1995 6150
rect 2045 6174 2089 6180
rect 2045 6154 2060 6174
rect 2080 6154 2089 6174
rect 2045 6138 2089 6154
rect 2159 6174 2203 6180
rect 2159 6154 2168 6174
rect 2188 6154 2203 6174
rect 2159 6138 2203 6154
rect 2253 6170 2302 6180
rect 2253 6150 2271 6170
rect 2291 6150 2302 6170
rect 2253 6138 2302 6150
rect 9415 6195 9464 6207
rect 9415 6175 9426 6195
rect 9446 6175 9464 6195
rect 9415 6165 9464 6175
rect 9514 6191 9558 6207
rect 9514 6171 9529 6191
rect 9549 6171 9558 6191
rect 9514 6165 9558 6171
rect 9628 6191 9672 6207
rect 9628 6171 9637 6191
rect 9657 6171 9672 6191
rect 9628 6165 9672 6171
rect 9722 6195 9771 6207
rect 9722 6175 9740 6195
rect 9760 6175 9771 6195
rect 9722 6165 9771 6175
rect 9836 6191 9880 6207
rect 9836 6171 9845 6191
rect 9865 6171 9880 6191
rect 9836 6165 9880 6171
rect 9930 6195 9979 6207
rect 9930 6175 9948 6195
rect 9968 6175 9979 6195
rect 9930 6165 9979 6175
rect 10049 6191 10093 6207
rect 10049 6171 10058 6191
rect 10078 6171 10093 6191
rect 10049 6165 10093 6171
rect 10143 6195 10192 6207
rect 10143 6175 10161 6195
rect 10181 6175 10192 6195
rect 10143 6165 10192 6175
rect 6806 6149 6855 6159
rect 6806 6129 6817 6149
rect 6837 6129 6855 6149
rect 6806 6117 6855 6129
rect 6905 6153 6949 6159
rect 6905 6133 6920 6153
rect 6940 6133 6949 6153
rect 6905 6117 6949 6133
rect 7019 6149 7068 6159
rect 7019 6129 7030 6149
rect 7050 6129 7068 6149
rect 7019 6117 7068 6129
rect 7118 6153 7162 6159
rect 7118 6133 7133 6153
rect 7153 6133 7162 6153
rect 7118 6117 7162 6133
rect 7227 6149 7276 6159
rect 7227 6129 7238 6149
rect 7258 6129 7276 6149
rect 7227 6117 7276 6129
rect 7326 6153 7370 6159
rect 7326 6133 7341 6153
rect 7361 6133 7370 6153
rect 7326 6117 7370 6133
rect 7440 6153 7484 6159
rect 7440 6133 7449 6153
rect 7469 6133 7484 6153
rect 7440 6117 7484 6133
rect 7534 6149 7583 6159
rect 7534 6129 7552 6149
rect 7572 6129 7583 6149
rect 7534 6117 7583 6129
rect 3121 5982 3170 5994
rect 3121 5962 3132 5982
rect 3152 5962 3170 5982
rect 3121 5952 3170 5962
rect 3220 5978 3264 5994
rect 3220 5958 3235 5978
rect 3255 5958 3264 5978
rect 3220 5952 3264 5958
rect 3334 5978 3378 5994
rect 3334 5958 3343 5978
rect 3363 5958 3378 5978
rect 3334 5952 3378 5958
rect 3428 5982 3477 5994
rect 3428 5962 3446 5982
rect 3466 5962 3477 5982
rect 3428 5952 3477 5962
rect 3542 5978 3586 5994
rect 3542 5958 3551 5978
rect 3571 5958 3586 5978
rect 3542 5952 3586 5958
rect 3636 5982 3685 5994
rect 3636 5962 3654 5982
rect 3674 5962 3685 5982
rect 3636 5952 3685 5962
rect 3755 5978 3799 5994
rect 3755 5958 3764 5978
rect 3784 5958 3799 5978
rect 3755 5952 3799 5958
rect 3849 5982 3898 5994
rect 3849 5962 3867 5982
rect 3887 5962 3898 5982
rect 3849 5952 3898 5962
rect 305 5884 354 5894
rect 305 5864 316 5884
rect 336 5864 354 5884
rect 305 5852 354 5864
rect 404 5888 448 5894
rect 404 5868 419 5888
rect 439 5868 448 5888
rect 404 5852 448 5868
rect 518 5884 567 5894
rect 518 5864 529 5884
rect 549 5864 567 5884
rect 518 5852 567 5864
rect 617 5888 661 5894
rect 617 5868 632 5888
rect 652 5868 661 5888
rect 617 5852 661 5868
rect 726 5884 775 5894
rect 726 5864 737 5884
rect 757 5864 775 5884
rect 726 5852 775 5864
rect 825 5888 869 5894
rect 825 5868 840 5888
rect 860 5868 869 5888
rect 825 5852 869 5868
rect 939 5888 983 5894
rect 939 5868 948 5888
rect 968 5868 983 5888
rect 939 5852 983 5868
rect 1033 5884 1082 5894
rect 1033 5864 1051 5884
rect 1071 5864 1082 5884
rect 1033 5852 1082 5864
rect 8402 5961 8451 5973
rect 8402 5941 8413 5961
rect 8433 5941 8451 5961
rect 8402 5931 8451 5941
rect 8501 5957 8545 5973
rect 8501 5937 8516 5957
rect 8536 5937 8545 5957
rect 8501 5931 8545 5937
rect 8615 5957 8659 5973
rect 8615 5937 8624 5957
rect 8644 5937 8659 5957
rect 8615 5931 8659 5937
rect 8709 5961 8758 5973
rect 8709 5941 8727 5961
rect 8747 5941 8758 5961
rect 8709 5931 8758 5941
rect 8823 5957 8867 5973
rect 8823 5937 8832 5957
rect 8852 5937 8867 5957
rect 8823 5931 8867 5937
rect 8917 5961 8966 5973
rect 8917 5941 8935 5961
rect 8955 5941 8966 5961
rect 8917 5931 8966 5941
rect 9036 5957 9080 5973
rect 9036 5937 9045 5957
rect 9065 5937 9080 5957
rect 9036 5931 9080 5937
rect 9130 5961 9179 5973
rect 9130 5941 9148 5961
rect 9168 5941 9179 5961
rect 9130 5931 9179 5941
rect 5586 5863 5635 5873
rect 5586 5843 5597 5863
rect 5617 5843 5635 5863
rect 5586 5831 5635 5843
rect 5685 5867 5729 5873
rect 5685 5847 5700 5867
rect 5720 5847 5729 5867
rect 5685 5831 5729 5847
rect 5799 5863 5848 5873
rect 5799 5843 5810 5863
rect 5830 5843 5848 5863
rect 5799 5831 5848 5843
rect 5898 5867 5942 5873
rect 5898 5847 5913 5867
rect 5933 5847 5942 5867
rect 5898 5831 5942 5847
rect 6007 5863 6056 5873
rect 6007 5843 6018 5863
rect 6038 5843 6056 5863
rect 6007 5831 6056 5843
rect 6106 5867 6150 5873
rect 6106 5847 6121 5867
rect 6141 5847 6150 5867
rect 6106 5831 6150 5847
rect 6220 5867 6264 5873
rect 6220 5847 6229 5867
rect 6249 5847 6264 5867
rect 6220 5831 6264 5847
rect 6314 5863 6363 5873
rect 6314 5843 6332 5863
rect 6352 5843 6363 5863
rect 6314 5831 6363 5843
rect 4133 5801 4182 5813
rect 4133 5781 4144 5801
rect 4164 5781 4182 5801
rect 4133 5771 4182 5781
rect 4232 5797 4276 5813
rect 4232 5777 4247 5797
rect 4267 5777 4276 5797
rect 4232 5771 4276 5777
rect 4346 5797 4390 5813
rect 4346 5777 4355 5797
rect 4375 5777 4390 5797
rect 4346 5771 4390 5777
rect 4440 5801 4489 5813
rect 4440 5781 4458 5801
rect 4478 5781 4489 5801
rect 4440 5771 4489 5781
rect 4554 5797 4598 5813
rect 4554 5777 4563 5797
rect 4583 5777 4598 5797
rect 4554 5771 4598 5777
rect 4648 5801 4697 5813
rect 4648 5781 4666 5801
rect 4686 5781 4697 5801
rect 4648 5771 4697 5781
rect 4767 5797 4811 5813
rect 4767 5777 4776 5797
rect 4796 5777 4811 5797
rect 4767 5771 4811 5777
rect 4861 5801 4910 5813
rect 4861 5781 4879 5801
rect 4899 5781 4910 5801
rect 4861 5771 4910 5781
rect 1317 5703 1366 5713
rect 1317 5683 1328 5703
rect 1348 5683 1366 5703
rect 1317 5671 1366 5683
rect 1416 5707 1460 5713
rect 1416 5687 1431 5707
rect 1451 5687 1460 5707
rect 1416 5671 1460 5687
rect 1530 5703 1579 5713
rect 1530 5683 1541 5703
rect 1561 5683 1579 5703
rect 1530 5671 1579 5683
rect 1629 5707 1673 5713
rect 1629 5687 1644 5707
rect 1664 5687 1673 5707
rect 1629 5671 1673 5687
rect 1738 5703 1787 5713
rect 1738 5683 1749 5703
rect 1769 5683 1787 5703
rect 1738 5671 1787 5683
rect 1837 5707 1881 5713
rect 1837 5687 1852 5707
rect 1872 5687 1881 5707
rect 1837 5671 1881 5687
rect 1951 5707 1995 5713
rect 1951 5687 1960 5707
rect 1980 5687 1995 5707
rect 1951 5671 1995 5687
rect 2045 5703 2094 5713
rect 2045 5683 2063 5703
rect 2083 5683 2094 5703
rect 2045 5671 2094 5683
rect 9414 5780 9463 5792
rect 9414 5760 9425 5780
rect 9445 5760 9463 5780
rect 9414 5750 9463 5760
rect 9513 5776 9557 5792
rect 9513 5756 9528 5776
rect 9548 5756 9557 5776
rect 9513 5750 9557 5756
rect 9627 5776 9671 5792
rect 9627 5756 9636 5776
rect 9656 5756 9671 5776
rect 9627 5750 9671 5756
rect 9721 5780 9770 5792
rect 9721 5760 9739 5780
rect 9759 5760 9770 5780
rect 9721 5750 9770 5760
rect 9835 5776 9879 5792
rect 9835 5756 9844 5776
rect 9864 5756 9879 5776
rect 9835 5750 9879 5756
rect 9929 5780 9978 5792
rect 9929 5760 9947 5780
rect 9967 5760 9978 5780
rect 9929 5750 9978 5760
rect 10048 5776 10092 5792
rect 10048 5756 10057 5776
rect 10077 5756 10092 5776
rect 10048 5750 10092 5756
rect 10142 5780 10191 5792
rect 10142 5760 10160 5780
rect 10180 5760 10191 5780
rect 10142 5750 10191 5760
rect 6598 5682 6647 5692
rect 6598 5662 6609 5682
rect 6629 5662 6647 5682
rect 6598 5650 6647 5662
rect 6697 5686 6741 5692
rect 6697 5666 6712 5686
rect 6732 5666 6741 5686
rect 6697 5650 6741 5666
rect 6811 5682 6860 5692
rect 6811 5662 6822 5682
rect 6842 5662 6860 5682
rect 6811 5650 6860 5662
rect 6910 5686 6954 5692
rect 6910 5666 6925 5686
rect 6945 5666 6954 5686
rect 6910 5650 6954 5666
rect 7019 5682 7068 5692
rect 7019 5662 7030 5682
rect 7050 5662 7068 5682
rect 7019 5650 7068 5662
rect 7118 5686 7162 5692
rect 7118 5666 7133 5686
rect 7153 5666 7162 5686
rect 7118 5650 7162 5666
rect 7232 5686 7276 5692
rect 7232 5666 7241 5686
rect 7261 5666 7276 5686
rect 7232 5650 7276 5666
rect 7326 5682 7375 5692
rect 7326 5662 7344 5682
rect 7364 5662 7375 5682
rect 7326 5650 7375 5662
rect 3071 5562 3120 5574
rect 3071 5542 3082 5562
rect 3102 5542 3120 5562
rect 3071 5532 3120 5542
rect 3170 5558 3214 5574
rect 3170 5538 3185 5558
rect 3205 5538 3214 5558
rect 3170 5532 3214 5538
rect 3284 5558 3328 5574
rect 3284 5538 3293 5558
rect 3313 5538 3328 5558
rect 3284 5532 3328 5538
rect 3378 5562 3427 5574
rect 3378 5542 3396 5562
rect 3416 5542 3427 5562
rect 3378 5532 3427 5542
rect 3492 5558 3536 5574
rect 3492 5538 3501 5558
rect 3521 5538 3536 5558
rect 3492 5532 3536 5538
rect 3586 5562 3635 5574
rect 3586 5542 3604 5562
rect 3624 5542 3635 5562
rect 3586 5532 3635 5542
rect 3705 5558 3749 5574
rect 3705 5538 3714 5558
rect 3734 5538 3749 5558
rect 3705 5532 3749 5538
rect 3799 5562 3848 5574
rect 3799 5542 3817 5562
rect 3837 5542 3848 5562
rect 3799 5532 3848 5542
rect 304 5469 353 5479
rect 304 5449 315 5469
rect 335 5449 353 5469
rect 304 5437 353 5449
rect 403 5473 447 5479
rect 403 5453 418 5473
rect 438 5453 447 5473
rect 403 5437 447 5453
rect 517 5469 566 5479
rect 517 5449 528 5469
rect 548 5449 566 5469
rect 517 5437 566 5449
rect 616 5473 660 5479
rect 616 5453 631 5473
rect 651 5453 660 5473
rect 616 5437 660 5453
rect 725 5469 774 5479
rect 725 5449 736 5469
rect 756 5449 774 5469
rect 725 5437 774 5449
rect 824 5473 868 5479
rect 824 5453 839 5473
rect 859 5453 868 5473
rect 824 5437 868 5453
rect 938 5473 982 5479
rect 938 5453 947 5473
rect 967 5453 982 5473
rect 938 5437 982 5453
rect 1032 5469 1081 5479
rect 1032 5449 1050 5469
rect 1070 5449 1081 5469
rect 8352 5541 8401 5553
rect 1032 5437 1081 5449
rect 8352 5521 8363 5541
rect 8383 5521 8401 5541
rect 8352 5511 8401 5521
rect 8451 5537 8495 5553
rect 8451 5517 8466 5537
rect 8486 5517 8495 5537
rect 8451 5511 8495 5517
rect 8565 5537 8609 5553
rect 8565 5517 8574 5537
rect 8594 5517 8609 5537
rect 8565 5511 8609 5517
rect 8659 5541 8708 5553
rect 8659 5521 8677 5541
rect 8697 5521 8708 5541
rect 8659 5511 8708 5521
rect 8773 5537 8817 5553
rect 8773 5517 8782 5537
rect 8802 5517 8817 5537
rect 8773 5511 8817 5517
rect 8867 5541 8916 5553
rect 8867 5521 8885 5541
rect 8905 5521 8916 5541
rect 8867 5511 8916 5521
rect 8986 5537 9030 5553
rect 8986 5517 8995 5537
rect 9015 5517 9030 5537
rect 8986 5511 9030 5517
rect 9080 5541 9129 5553
rect 9080 5521 9098 5541
rect 9118 5521 9129 5541
rect 9080 5511 9129 5521
rect 5585 5448 5634 5458
rect 5585 5428 5596 5448
rect 5616 5428 5634 5448
rect 5585 5416 5634 5428
rect 5684 5452 5728 5458
rect 5684 5432 5699 5452
rect 5719 5432 5728 5452
rect 5684 5416 5728 5432
rect 5798 5448 5847 5458
rect 5798 5428 5809 5448
rect 5829 5428 5847 5448
rect 5798 5416 5847 5428
rect 5897 5452 5941 5458
rect 5897 5432 5912 5452
rect 5932 5432 5941 5452
rect 5897 5416 5941 5432
rect 6006 5448 6055 5458
rect 6006 5428 6017 5448
rect 6037 5428 6055 5448
rect 6006 5416 6055 5428
rect 6105 5452 6149 5458
rect 6105 5432 6120 5452
rect 6140 5432 6149 5452
rect 6105 5416 6149 5432
rect 6219 5452 6263 5458
rect 6219 5432 6228 5452
rect 6248 5432 6263 5452
rect 6219 5416 6263 5432
rect 6313 5448 6362 5458
rect 6313 5428 6331 5448
rect 6351 5428 6362 5448
rect 6313 5416 6362 5428
rect 4139 5235 4188 5247
rect 4139 5215 4150 5235
rect 4170 5215 4188 5235
rect 4139 5205 4188 5215
rect 4238 5231 4282 5247
rect 4238 5211 4253 5231
rect 4273 5211 4282 5231
rect 4238 5205 4282 5211
rect 4352 5231 4396 5247
rect 4352 5211 4361 5231
rect 4381 5211 4396 5231
rect 4352 5205 4396 5211
rect 4446 5235 4495 5247
rect 4446 5215 4464 5235
rect 4484 5215 4495 5235
rect 4446 5205 4495 5215
rect 4560 5231 4604 5247
rect 4560 5211 4569 5231
rect 4589 5211 4604 5231
rect 4560 5205 4604 5211
rect 4654 5235 4703 5247
rect 4654 5215 4672 5235
rect 4692 5215 4703 5235
rect 4654 5205 4703 5215
rect 4773 5231 4817 5247
rect 4773 5211 4782 5231
rect 4802 5211 4817 5231
rect 4773 5205 4817 5211
rect 4867 5235 4916 5247
rect 4867 5215 4885 5235
rect 4905 5215 4916 5235
rect 4867 5205 4916 5215
rect 1372 5142 1421 5152
rect 1372 5122 1383 5142
rect 1403 5122 1421 5142
rect 1372 5110 1421 5122
rect 1471 5146 1515 5152
rect 1471 5126 1486 5146
rect 1506 5126 1515 5146
rect 1471 5110 1515 5126
rect 1585 5142 1634 5152
rect 1585 5122 1596 5142
rect 1616 5122 1634 5142
rect 1585 5110 1634 5122
rect 1684 5146 1728 5152
rect 1684 5126 1699 5146
rect 1719 5126 1728 5146
rect 1684 5110 1728 5126
rect 1793 5142 1842 5152
rect 1793 5122 1804 5142
rect 1824 5122 1842 5142
rect 1793 5110 1842 5122
rect 1892 5146 1936 5152
rect 1892 5126 1907 5146
rect 1927 5126 1936 5146
rect 1892 5110 1936 5126
rect 2006 5146 2050 5152
rect 2006 5126 2015 5146
rect 2035 5126 2050 5146
rect 2006 5110 2050 5126
rect 2100 5142 2149 5152
rect 2100 5122 2118 5142
rect 2138 5122 2149 5142
rect 9420 5214 9469 5226
rect 2100 5110 2149 5122
rect 9420 5194 9431 5214
rect 9451 5194 9469 5214
rect 9420 5184 9469 5194
rect 9519 5210 9563 5226
rect 9519 5190 9534 5210
rect 9554 5190 9563 5210
rect 9519 5184 9563 5190
rect 9633 5210 9677 5226
rect 9633 5190 9642 5210
rect 9662 5190 9677 5210
rect 9633 5184 9677 5190
rect 9727 5214 9776 5226
rect 9727 5194 9745 5214
rect 9765 5194 9776 5214
rect 9727 5184 9776 5194
rect 9841 5210 9885 5226
rect 9841 5190 9850 5210
rect 9870 5190 9885 5210
rect 9841 5184 9885 5190
rect 9935 5214 9984 5226
rect 9935 5194 9953 5214
rect 9973 5194 9984 5214
rect 9935 5184 9984 5194
rect 10054 5210 10098 5226
rect 10054 5190 10063 5210
rect 10083 5190 10098 5210
rect 10054 5184 10098 5190
rect 10148 5214 10197 5226
rect 10148 5194 10166 5214
rect 10186 5194 10197 5214
rect 10148 5184 10197 5194
rect 6653 5121 6702 5131
rect 6653 5101 6664 5121
rect 6684 5101 6702 5121
rect 6653 5089 6702 5101
rect 6752 5125 6796 5131
rect 6752 5105 6767 5125
rect 6787 5105 6796 5125
rect 6752 5089 6796 5105
rect 6866 5121 6915 5131
rect 6866 5101 6877 5121
rect 6897 5101 6915 5121
rect 6866 5089 6915 5101
rect 6965 5125 7009 5131
rect 6965 5105 6980 5125
rect 7000 5105 7009 5125
rect 6965 5089 7009 5105
rect 7074 5121 7123 5131
rect 7074 5101 7085 5121
rect 7105 5101 7123 5121
rect 7074 5089 7123 5101
rect 7173 5125 7217 5131
rect 7173 5105 7188 5125
rect 7208 5105 7217 5125
rect 7173 5089 7217 5105
rect 7287 5125 7331 5131
rect 7287 5105 7296 5125
rect 7316 5105 7331 5125
rect 7287 5089 7331 5105
rect 7381 5121 7430 5131
rect 7381 5101 7399 5121
rect 7419 5101 7430 5121
rect 7381 5089 7430 5101
rect 3126 5001 3175 5013
rect 3126 4981 3137 5001
rect 3157 4981 3175 5001
rect 3126 4971 3175 4981
rect 3225 4997 3269 5013
rect 3225 4977 3240 4997
rect 3260 4977 3269 4997
rect 3225 4971 3269 4977
rect 3339 4997 3383 5013
rect 3339 4977 3348 4997
rect 3368 4977 3383 4997
rect 3339 4971 3383 4977
rect 3433 5001 3482 5013
rect 3433 4981 3451 5001
rect 3471 4981 3482 5001
rect 3433 4971 3482 4981
rect 3547 4997 3591 5013
rect 3547 4977 3556 4997
rect 3576 4977 3591 4997
rect 3547 4971 3591 4977
rect 3641 5001 3690 5013
rect 3641 4981 3659 5001
rect 3679 4981 3690 5001
rect 3641 4971 3690 4981
rect 3760 4997 3804 5013
rect 3760 4977 3769 4997
rect 3789 4977 3804 4997
rect 3760 4971 3804 4977
rect 3854 5001 3903 5013
rect 3854 4981 3872 5001
rect 3892 4981 3903 5001
rect 3854 4971 3903 4981
rect 310 4903 359 4913
rect 310 4883 321 4903
rect 341 4883 359 4903
rect 310 4871 359 4883
rect 409 4907 453 4913
rect 409 4887 424 4907
rect 444 4887 453 4907
rect 409 4871 453 4887
rect 523 4903 572 4913
rect 523 4883 534 4903
rect 554 4883 572 4903
rect 523 4871 572 4883
rect 622 4907 666 4913
rect 622 4887 637 4907
rect 657 4887 666 4907
rect 622 4871 666 4887
rect 731 4903 780 4913
rect 731 4883 742 4903
rect 762 4883 780 4903
rect 731 4871 780 4883
rect 830 4907 874 4913
rect 830 4887 845 4907
rect 865 4887 874 4907
rect 830 4871 874 4887
rect 944 4907 988 4913
rect 944 4887 953 4907
rect 973 4887 988 4907
rect 944 4871 988 4887
rect 1038 4903 1087 4913
rect 1038 4883 1056 4903
rect 1076 4883 1087 4903
rect 1038 4871 1087 4883
rect 8407 4980 8456 4992
rect 8407 4960 8418 4980
rect 8438 4960 8456 4980
rect 8407 4950 8456 4960
rect 8506 4976 8550 4992
rect 8506 4956 8521 4976
rect 8541 4956 8550 4976
rect 8506 4950 8550 4956
rect 8620 4976 8664 4992
rect 8620 4956 8629 4976
rect 8649 4956 8664 4976
rect 8620 4950 8664 4956
rect 8714 4980 8763 4992
rect 8714 4960 8732 4980
rect 8752 4960 8763 4980
rect 8714 4950 8763 4960
rect 8828 4976 8872 4992
rect 8828 4956 8837 4976
rect 8857 4956 8872 4976
rect 8828 4950 8872 4956
rect 8922 4980 8971 4992
rect 8922 4960 8940 4980
rect 8960 4960 8971 4980
rect 8922 4950 8971 4960
rect 9041 4976 9085 4992
rect 9041 4956 9050 4976
rect 9070 4956 9085 4976
rect 9041 4950 9085 4956
rect 9135 4980 9184 4992
rect 9135 4960 9153 4980
rect 9173 4960 9184 4980
rect 9135 4950 9184 4960
rect 5591 4882 5640 4892
rect 5591 4862 5602 4882
rect 5622 4862 5640 4882
rect 5591 4850 5640 4862
rect 5690 4886 5734 4892
rect 5690 4866 5705 4886
rect 5725 4866 5734 4886
rect 5690 4850 5734 4866
rect 5804 4882 5853 4892
rect 5804 4862 5815 4882
rect 5835 4862 5853 4882
rect 5804 4850 5853 4862
rect 5903 4886 5947 4892
rect 5903 4866 5918 4886
rect 5938 4866 5947 4886
rect 5903 4850 5947 4866
rect 6012 4882 6061 4892
rect 6012 4862 6023 4882
rect 6043 4862 6061 4882
rect 6012 4850 6061 4862
rect 6111 4886 6155 4892
rect 6111 4866 6126 4886
rect 6146 4866 6155 4886
rect 6111 4850 6155 4866
rect 6225 4886 6269 4892
rect 6225 4866 6234 4886
rect 6254 4866 6269 4886
rect 6225 4850 6269 4866
rect 6319 4882 6368 4892
rect 6319 4862 6337 4882
rect 6357 4862 6368 4882
rect 6319 4850 6368 4862
rect 4138 4820 4187 4832
rect 4138 4800 4149 4820
rect 4169 4800 4187 4820
rect 4138 4790 4187 4800
rect 4237 4816 4281 4832
rect 4237 4796 4252 4816
rect 4272 4796 4281 4816
rect 4237 4790 4281 4796
rect 4351 4816 4395 4832
rect 4351 4796 4360 4816
rect 4380 4796 4395 4816
rect 4351 4790 4395 4796
rect 4445 4820 4494 4832
rect 4445 4800 4463 4820
rect 4483 4800 4494 4820
rect 4445 4790 4494 4800
rect 4559 4816 4603 4832
rect 4559 4796 4568 4816
rect 4588 4796 4603 4816
rect 4559 4790 4603 4796
rect 4653 4820 4702 4832
rect 4653 4800 4671 4820
rect 4691 4800 4702 4820
rect 4653 4790 4702 4800
rect 4772 4816 4816 4832
rect 4772 4796 4781 4816
rect 4801 4796 4816 4816
rect 4772 4790 4816 4796
rect 4866 4820 4915 4832
rect 4866 4800 4884 4820
rect 4904 4800 4915 4820
rect 4866 4790 4915 4800
rect 1322 4722 1371 4732
rect 1322 4702 1333 4722
rect 1353 4702 1371 4722
rect 1322 4690 1371 4702
rect 1421 4726 1465 4732
rect 1421 4706 1436 4726
rect 1456 4706 1465 4726
rect 1421 4690 1465 4706
rect 1535 4722 1584 4732
rect 1535 4702 1546 4722
rect 1566 4702 1584 4722
rect 1535 4690 1584 4702
rect 1634 4726 1678 4732
rect 1634 4706 1649 4726
rect 1669 4706 1678 4726
rect 1634 4690 1678 4706
rect 1743 4722 1792 4732
rect 1743 4702 1754 4722
rect 1774 4702 1792 4722
rect 1743 4690 1792 4702
rect 1842 4726 1886 4732
rect 1842 4706 1857 4726
rect 1877 4706 1886 4726
rect 1842 4690 1886 4706
rect 1956 4726 2000 4732
rect 1956 4706 1965 4726
rect 1985 4706 2000 4726
rect 1956 4690 2000 4706
rect 2050 4722 2099 4732
rect 2050 4702 2068 4722
rect 2088 4702 2099 4722
rect 2050 4690 2099 4702
rect 9419 4799 9468 4811
rect 9419 4779 9430 4799
rect 9450 4779 9468 4799
rect 9419 4769 9468 4779
rect 9518 4795 9562 4811
rect 9518 4775 9533 4795
rect 9553 4775 9562 4795
rect 9518 4769 9562 4775
rect 9632 4795 9676 4811
rect 9632 4775 9641 4795
rect 9661 4775 9676 4795
rect 9632 4769 9676 4775
rect 9726 4799 9775 4811
rect 9726 4779 9744 4799
rect 9764 4779 9775 4799
rect 9726 4769 9775 4779
rect 9840 4795 9884 4811
rect 9840 4775 9849 4795
rect 9869 4775 9884 4795
rect 9840 4769 9884 4775
rect 9934 4799 9983 4811
rect 9934 4779 9952 4799
rect 9972 4779 9983 4799
rect 9934 4769 9983 4779
rect 10053 4795 10097 4811
rect 10053 4775 10062 4795
rect 10082 4775 10097 4795
rect 10053 4769 10097 4775
rect 10147 4799 10196 4811
rect 10147 4779 10165 4799
rect 10185 4779 10196 4799
rect 10147 4769 10196 4779
rect 6603 4701 6652 4711
rect 6603 4681 6614 4701
rect 6634 4681 6652 4701
rect 6603 4669 6652 4681
rect 6702 4705 6746 4711
rect 6702 4685 6717 4705
rect 6737 4685 6746 4705
rect 6702 4669 6746 4685
rect 6816 4701 6865 4711
rect 6816 4681 6827 4701
rect 6847 4681 6865 4701
rect 6816 4669 6865 4681
rect 6915 4705 6959 4711
rect 6915 4685 6930 4705
rect 6950 4685 6959 4705
rect 6915 4669 6959 4685
rect 7024 4701 7073 4711
rect 7024 4681 7035 4701
rect 7055 4681 7073 4701
rect 7024 4669 7073 4681
rect 7123 4705 7167 4711
rect 7123 4685 7138 4705
rect 7158 4685 7167 4705
rect 7123 4669 7167 4685
rect 7237 4705 7281 4711
rect 7237 4685 7246 4705
rect 7266 4685 7281 4705
rect 7237 4669 7281 4685
rect 7331 4701 7380 4711
rect 7331 4681 7349 4701
rect 7369 4681 7380 4701
rect 7331 4669 7380 4681
rect 2831 4569 2880 4581
rect 2831 4549 2842 4569
rect 2862 4549 2880 4569
rect 2831 4539 2880 4549
rect 2930 4565 2974 4581
rect 2930 4545 2945 4565
rect 2965 4545 2974 4565
rect 2930 4539 2974 4545
rect 3044 4565 3088 4581
rect 3044 4545 3053 4565
rect 3073 4545 3088 4565
rect 3044 4539 3088 4545
rect 3138 4569 3187 4581
rect 3138 4549 3156 4569
rect 3176 4549 3187 4569
rect 3138 4539 3187 4549
rect 3252 4565 3296 4581
rect 3252 4545 3261 4565
rect 3281 4545 3296 4565
rect 3252 4539 3296 4545
rect 3346 4569 3395 4581
rect 3346 4549 3364 4569
rect 3384 4549 3395 4569
rect 3346 4539 3395 4549
rect 3465 4565 3509 4581
rect 3465 4545 3474 4565
rect 3494 4545 3509 4565
rect 3465 4539 3509 4545
rect 3559 4569 3608 4581
rect 3559 4549 3577 4569
rect 3597 4549 3608 4569
rect 3559 4539 3608 4549
rect 309 4488 358 4498
rect 309 4468 320 4488
rect 340 4468 358 4488
rect 309 4456 358 4468
rect 408 4492 452 4498
rect 408 4472 423 4492
rect 443 4472 452 4492
rect 408 4456 452 4472
rect 522 4488 571 4498
rect 522 4468 533 4488
rect 553 4468 571 4488
rect 522 4456 571 4468
rect 621 4492 665 4498
rect 621 4472 636 4492
rect 656 4472 665 4492
rect 621 4456 665 4472
rect 730 4488 779 4498
rect 730 4468 741 4488
rect 761 4468 779 4488
rect 730 4456 779 4468
rect 829 4492 873 4498
rect 829 4472 844 4492
rect 864 4472 873 4492
rect 829 4456 873 4472
rect 943 4492 987 4498
rect 943 4472 952 4492
rect 972 4472 987 4492
rect 943 4456 987 4472
rect 1037 4488 1086 4498
rect 1037 4468 1055 4488
rect 1075 4468 1086 4488
rect 1037 4456 1086 4468
rect 8112 4548 8161 4560
rect 8112 4528 8123 4548
rect 8143 4528 8161 4548
rect 8112 4518 8161 4528
rect 8211 4544 8255 4560
rect 8211 4524 8226 4544
rect 8246 4524 8255 4544
rect 8211 4518 8255 4524
rect 8325 4544 8369 4560
rect 8325 4524 8334 4544
rect 8354 4524 8369 4544
rect 8325 4518 8369 4524
rect 8419 4548 8468 4560
rect 8419 4528 8437 4548
rect 8457 4528 8468 4548
rect 8419 4518 8468 4528
rect 8533 4544 8577 4560
rect 8533 4524 8542 4544
rect 8562 4524 8577 4544
rect 8533 4518 8577 4524
rect 8627 4548 8676 4560
rect 8627 4528 8645 4548
rect 8665 4528 8676 4548
rect 8627 4518 8676 4528
rect 8746 4544 8790 4560
rect 8746 4524 8755 4544
rect 8775 4524 8790 4544
rect 8746 4518 8790 4524
rect 8840 4548 8889 4560
rect 8840 4528 8858 4548
rect 8878 4528 8889 4548
rect 8840 4518 8889 4528
rect 5590 4467 5639 4477
rect 5590 4447 5601 4467
rect 5621 4447 5639 4467
rect 5590 4435 5639 4447
rect 5689 4471 5733 4477
rect 5689 4451 5704 4471
rect 5724 4451 5733 4471
rect 5689 4435 5733 4451
rect 5803 4467 5852 4477
rect 5803 4447 5814 4467
rect 5834 4447 5852 4467
rect 5803 4435 5852 4447
rect 5902 4471 5946 4477
rect 5902 4451 5917 4471
rect 5937 4451 5946 4471
rect 5902 4435 5946 4451
rect 6011 4467 6060 4477
rect 6011 4447 6022 4467
rect 6042 4447 6060 4467
rect 6011 4435 6060 4447
rect 6110 4471 6154 4477
rect 6110 4451 6125 4471
rect 6145 4451 6154 4471
rect 6110 4435 6154 4451
rect 6224 4471 6268 4477
rect 6224 4451 6233 4471
rect 6253 4451 6268 4471
rect 6224 4435 6268 4451
rect 6318 4467 6367 4477
rect 6318 4447 6336 4467
rect 6356 4447 6367 4467
rect 6318 4435 6367 4447
rect 4142 4259 4191 4271
rect 4142 4239 4153 4259
rect 4173 4239 4191 4259
rect 4142 4229 4191 4239
rect 4241 4255 4285 4271
rect 4241 4235 4256 4255
rect 4276 4235 4285 4255
rect 4241 4229 4285 4235
rect 4355 4255 4399 4271
rect 4355 4235 4364 4255
rect 4384 4235 4399 4255
rect 4355 4229 4399 4235
rect 4449 4259 4498 4271
rect 4449 4239 4467 4259
rect 4487 4239 4498 4259
rect 4449 4229 4498 4239
rect 4563 4255 4607 4271
rect 4563 4235 4572 4255
rect 4592 4235 4607 4255
rect 4563 4229 4607 4235
rect 4657 4259 4706 4271
rect 4657 4239 4675 4259
rect 4695 4239 4706 4259
rect 4657 4229 4706 4239
rect 4776 4255 4820 4271
rect 4776 4235 4785 4255
rect 4805 4235 4820 4255
rect 4776 4229 4820 4235
rect 4870 4259 4919 4271
rect 4870 4239 4888 4259
rect 4908 4239 4919 4259
rect 4870 4229 4919 4239
rect 1620 4178 1669 4188
rect 1620 4158 1631 4178
rect 1651 4158 1669 4178
rect 1620 4146 1669 4158
rect 1719 4182 1763 4188
rect 1719 4162 1734 4182
rect 1754 4162 1763 4182
rect 1719 4146 1763 4162
rect 1833 4178 1882 4188
rect 1833 4158 1844 4178
rect 1864 4158 1882 4178
rect 1833 4146 1882 4158
rect 1932 4182 1976 4188
rect 1932 4162 1947 4182
rect 1967 4162 1976 4182
rect 1932 4146 1976 4162
rect 2041 4178 2090 4188
rect 2041 4158 2052 4178
rect 2072 4158 2090 4178
rect 2041 4146 2090 4158
rect 2140 4182 2184 4188
rect 2140 4162 2155 4182
rect 2175 4162 2184 4182
rect 2140 4146 2184 4162
rect 2254 4182 2298 4188
rect 2254 4162 2263 4182
rect 2283 4162 2298 4182
rect 2254 4146 2298 4162
rect 2348 4178 2397 4188
rect 2348 4158 2366 4178
rect 2386 4158 2397 4178
rect 2348 4146 2397 4158
rect 9423 4238 9472 4250
rect 9423 4218 9434 4238
rect 9454 4218 9472 4238
rect 9423 4208 9472 4218
rect 9522 4234 9566 4250
rect 9522 4214 9537 4234
rect 9557 4214 9566 4234
rect 9522 4208 9566 4214
rect 9636 4234 9680 4250
rect 9636 4214 9645 4234
rect 9665 4214 9680 4234
rect 9636 4208 9680 4214
rect 9730 4238 9779 4250
rect 9730 4218 9748 4238
rect 9768 4218 9779 4238
rect 9730 4208 9779 4218
rect 9844 4234 9888 4250
rect 9844 4214 9853 4234
rect 9873 4214 9888 4234
rect 9844 4208 9888 4214
rect 9938 4238 9987 4250
rect 9938 4218 9956 4238
rect 9976 4218 9987 4238
rect 9938 4208 9987 4218
rect 10057 4234 10101 4250
rect 10057 4214 10066 4234
rect 10086 4214 10101 4234
rect 10057 4208 10101 4214
rect 10151 4238 10200 4250
rect 10151 4218 10169 4238
rect 10189 4218 10200 4238
rect 10151 4208 10200 4218
rect 6901 4157 6950 4167
rect 6901 4137 6912 4157
rect 6932 4137 6950 4157
rect 6901 4125 6950 4137
rect 7000 4161 7044 4167
rect 7000 4141 7015 4161
rect 7035 4141 7044 4161
rect 7000 4125 7044 4141
rect 7114 4157 7163 4167
rect 7114 4137 7125 4157
rect 7145 4137 7163 4157
rect 7114 4125 7163 4137
rect 7213 4161 7257 4167
rect 7213 4141 7228 4161
rect 7248 4141 7257 4161
rect 7213 4125 7257 4141
rect 7322 4157 7371 4167
rect 7322 4137 7333 4157
rect 7353 4137 7371 4157
rect 7322 4125 7371 4137
rect 7421 4161 7465 4167
rect 7421 4141 7436 4161
rect 7456 4141 7465 4161
rect 7421 4125 7465 4141
rect 7535 4161 7579 4167
rect 7535 4141 7544 4161
rect 7564 4141 7579 4161
rect 7535 4125 7579 4141
rect 7629 4157 7678 4167
rect 7629 4137 7647 4157
rect 7667 4137 7678 4157
rect 7629 4125 7678 4137
rect 3129 4025 3178 4037
rect 3129 4005 3140 4025
rect 3160 4005 3178 4025
rect 3129 3995 3178 4005
rect 3228 4021 3272 4037
rect 3228 4001 3243 4021
rect 3263 4001 3272 4021
rect 3228 3995 3272 4001
rect 3342 4021 3386 4037
rect 3342 4001 3351 4021
rect 3371 4001 3386 4021
rect 3342 3995 3386 4001
rect 3436 4025 3485 4037
rect 3436 4005 3454 4025
rect 3474 4005 3485 4025
rect 3436 3995 3485 4005
rect 3550 4021 3594 4037
rect 3550 4001 3559 4021
rect 3579 4001 3594 4021
rect 3550 3995 3594 4001
rect 3644 4025 3693 4037
rect 3644 4005 3662 4025
rect 3682 4005 3693 4025
rect 3644 3995 3693 4005
rect 3763 4021 3807 4037
rect 3763 4001 3772 4021
rect 3792 4001 3807 4021
rect 3763 3995 3807 4001
rect 3857 4025 3906 4037
rect 3857 4005 3875 4025
rect 3895 4005 3906 4025
rect 3857 3995 3906 4005
rect 313 3927 362 3937
rect 313 3907 324 3927
rect 344 3907 362 3927
rect 313 3895 362 3907
rect 412 3931 456 3937
rect 412 3911 427 3931
rect 447 3911 456 3931
rect 412 3895 456 3911
rect 526 3927 575 3937
rect 526 3907 537 3927
rect 557 3907 575 3927
rect 526 3895 575 3907
rect 625 3931 669 3937
rect 625 3911 640 3931
rect 660 3911 669 3931
rect 625 3895 669 3911
rect 734 3927 783 3937
rect 734 3907 745 3927
rect 765 3907 783 3927
rect 734 3895 783 3907
rect 833 3931 877 3937
rect 833 3911 848 3931
rect 868 3911 877 3931
rect 833 3895 877 3911
rect 947 3931 991 3937
rect 947 3911 956 3931
rect 976 3911 991 3931
rect 947 3895 991 3911
rect 1041 3927 1090 3937
rect 1041 3907 1059 3927
rect 1079 3907 1090 3927
rect 1041 3895 1090 3907
rect 8410 4004 8459 4016
rect 8410 3984 8421 4004
rect 8441 3984 8459 4004
rect 8410 3974 8459 3984
rect 8509 4000 8553 4016
rect 8509 3980 8524 4000
rect 8544 3980 8553 4000
rect 8509 3974 8553 3980
rect 8623 4000 8667 4016
rect 8623 3980 8632 4000
rect 8652 3980 8667 4000
rect 8623 3974 8667 3980
rect 8717 4004 8766 4016
rect 8717 3984 8735 4004
rect 8755 3984 8766 4004
rect 8717 3974 8766 3984
rect 8831 4000 8875 4016
rect 8831 3980 8840 4000
rect 8860 3980 8875 4000
rect 8831 3974 8875 3980
rect 8925 4004 8974 4016
rect 8925 3984 8943 4004
rect 8963 3984 8974 4004
rect 8925 3974 8974 3984
rect 9044 4000 9088 4016
rect 9044 3980 9053 4000
rect 9073 3980 9088 4000
rect 9044 3974 9088 3980
rect 9138 4004 9187 4016
rect 9138 3984 9156 4004
rect 9176 3984 9187 4004
rect 9138 3974 9187 3984
rect 5594 3906 5643 3916
rect 5594 3886 5605 3906
rect 5625 3886 5643 3906
rect 5594 3874 5643 3886
rect 5693 3910 5737 3916
rect 5693 3890 5708 3910
rect 5728 3890 5737 3910
rect 5693 3874 5737 3890
rect 5807 3906 5856 3916
rect 5807 3886 5818 3906
rect 5838 3886 5856 3906
rect 5807 3874 5856 3886
rect 5906 3910 5950 3916
rect 5906 3890 5921 3910
rect 5941 3890 5950 3910
rect 5906 3874 5950 3890
rect 6015 3906 6064 3916
rect 6015 3886 6026 3906
rect 6046 3886 6064 3906
rect 6015 3874 6064 3886
rect 6114 3910 6158 3916
rect 6114 3890 6129 3910
rect 6149 3890 6158 3910
rect 6114 3874 6158 3890
rect 6228 3910 6272 3916
rect 6228 3890 6237 3910
rect 6257 3890 6272 3910
rect 6228 3874 6272 3890
rect 6322 3906 6371 3916
rect 6322 3886 6340 3906
rect 6360 3886 6371 3906
rect 6322 3874 6371 3886
rect 4141 3844 4190 3856
rect 4141 3824 4152 3844
rect 4172 3824 4190 3844
rect 4141 3814 4190 3824
rect 4240 3840 4284 3856
rect 4240 3820 4255 3840
rect 4275 3820 4284 3840
rect 4240 3814 4284 3820
rect 4354 3840 4398 3856
rect 4354 3820 4363 3840
rect 4383 3820 4398 3840
rect 4354 3814 4398 3820
rect 4448 3844 4497 3856
rect 4448 3824 4466 3844
rect 4486 3824 4497 3844
rect 4448 3814 4497 3824
rect 4562 3840 4606 3856
rect 4562 3820 4571 3840
rect 4591 3820 4606 3840
rect 4562 3814 4606 3820
rect 4656 3844 4705 3856
rect 4656 3824 4674 3844
rect 4694 3824 4705 3844
rect 4656 3814 4705 3824
rect 4775 3840 4819 3856
rect 4775 3820 4784 3840
rect 4804 3820 4819 3840
rect 4775 3814 4819 3820
rect 4869 3844 4918 3856
rect 4869 3824 4887 3844
rect 4907 3824 4918 3844
rect 4869 3814 4918 3824
rect 1325 3746 1374 3756
rect 1325 3726 1336 3746
rect 1356 3726 1374 3746
rect 1325 3714 1374 3726
rect 1424 3750 1468 3756
rect 1424 3730 1439 3750
rect 1459 3730 1468 3750
rect 1424 3714 1468 3730
rect 1538 3746 1587 3756
rect 1538 3726 1549 3746
rect 1569 3726 1587 3746
rect 1538 3714 1587 3726
rect 1637 3750 1681 3756
rect 1637 3730 1652 3750
rect 1672 3730 1681 3750
rect 1637 3714 1681 3730
rect 1746 3746 1795 3756
rect 1746 3726 1757 3746
rect 1777 3726 1795 3746
rect 1746 3714 1795 3726
rect 1845 3750 1889 3756
rect 1845 3730 1860 3750
rect 1880 3730 1889 3750
rect 1845 3714 1889 3730
rect 1959 3750 2003 3756
rect 1959 3730 1968 3750
rect 1988 3730 2003 3750
rect 1959 3714 2003 3730
rect 2053 3746 2102 3756
rect 2053 3726 2071 3746
rect 2091 3726 2102 3746
rect 2053 3714 2102 3726
rect 9422 3823 9471 3835
rect 9422 3803 9433 3823
rect 9453 3803 9471 3823
rect 9422 3793 9471 3803
rect 9521 3819 9565 3835
rect 9521 3799 9536 3819
rect 9556 3799 9565 3819
rect 9521 3793 9565 3799
rect 9635 3819 9679 3835
rect 9635 3799 9644 3819
rect 9664 3799 9679 3819
rect 9635 3793 9679 3799
rect 9729 3823 9778 3835
rect 9729 3803 9747 3823
rect 9767 3803 9778 3823
rect 9729 3793 9778 3803
rect 9843 3819 9887 3835
rect 9843 3799 9852 3819
rect 9872 3799 9887 3819
rect 9843 3793 9887 3799
rect 9937 3823 9986 3835
rect 9937 3803 9955 3823
rect 9975 3803 9986 3823
rect 9937 3793 9986 3803
rect 10056 3819 10100 3835
rect 10056 3799 10065 3819
rect 10085 3799 10100 3819
rect 10056 3793 10100 3799
rect 10150 3823 10199 3835
rect 10150 3803 10168 3823
rect 10188 3803 10199 3823
rect 10150 3793 10199 3803
rect 6606 3725 6655 3735
rect 6606 3705 6617 3725
rect 6637 3705 6655 3725
rect 6606 3693 6655 3705
rect 6705 3729 6749 3735
rect 6705 3709 6720 3729
rect 6740 3709 6749 3729
rect 6705 3693 6749 3709
rect 6819 3725 6868 3735
rect 6819 3705 6830 3725
rect 6850 3705 6868 3725
rect 6819 3693 6868 3705
rect 6918 3729 6962 3735
rect 6918 3709 6933 3729
rect 6953 3709 6962 3729
rect 6918 3693 6962 3709
rect 7027 3725 7076 3735
rect 7027 3705 7038 3725
rect 7058 3705 7076 3725
rect 7027 3693 7076 3705
rect 7126 3729 7170 3735
rect 7126 3709 7141 3729
rect 7161 3709 7170 3729
rect 7126 3693 7170 3709
rect 7240 3729 7284 3735
rect 7240 3709 7249 3729
rect 7269 3709 7284 3729
rect 7240 3693 7284 3709
rect 7334 3725 7383 3735
rect 7334 3705 7352 3725
rect 7372 3705 7383 3725
rect 7334 3693 7383 3705
rect 3079 3605 3128 3617
rect 3079 3585 3090 3605
rect 3110 3585 3128 3605
rect 3079 3575 3128 3585
rect 3178 3601 3222 3617
rect 3178 3581 3193 3601
rect 3213 3581 3222 3601
rect 3178 3575 3222 3581
rect 3292 3601 3336 3617
rect 3292 3581 3301 3601
rect 3321 3581 3336 3601
rect 3292 3575 3336 3581
rect 3386 3605 3435 3617
rect 3386 3585 3404 3605
rect 3424 3585 3435 3605
rect 3386 3575 3435 3585
rect 3500 3601 3544 3617
rect 3500 3581 3509 3601
rect 3529 3581 3544 3601
rect 3500 3575 3544 3581
rect 3594 3605 3643 3617
rect 3594 3585 3612 3605
rect 3632 3585 3643 3605
rect 3594 3575 3643 3585
rect 3713 3601 3757 3617
rect 3713 3581 3722 3601
rect 3742 3581 3757 3601
rect 3713 3575 3757 3581
rect 3807 3605 3856 3617
rect 3807 3585 3825 3605
rect 3845 3585 3856 3605
rect 3807 3575 3856 3585
rect 312 3512 361 3522
rect 312 3492 323 3512
rect 343 3492 361 3512
rect 312 3480 361 3492
rect 411 3516 455 3522
rect 411 3496 426 3516
rect 446 3496 455 3516
rect 411 3480 455 3496
rect 525 3512 574 3522
rect 525 3492 536 3512
rect 556 3492 574 3512
rect 525 3480 574 3492
rect 624 3516 668 3522
rect 624 3496 639 3516
rect 659 3496 668 3516
rect 624 3480 668 3496
rect 733 3512 782 3522
rect 733 3492 744 3512
rect 764 3492 782 3512
rect 733 3480 782 3492
rect 832 3516 876 3522
rect 832 3496 847 3516
rect 867 3496 876 3516
rect 832 3480 876 3496
rect 946 3516 990 3522
rect 946 3496 955 3516
rect 975 3496 990 3516
rect 946 3480 990 3496
rect 1040 3512 1089 3522
rect 1040 3492 1058 3512
rect 1078 3492 1089 3512
rect 8360 3584 8409 3596
rect 1040 3480 1089 3492
rect 8360 3564 8371 3584
rect 8391 3564 8409 3584
rect 8360 3554 8409 3564
rect 8459 3580 8503 3596
rect 8459 3560 8474 3580
rect 8494 3560 8503 3580
rect 8459 3554 8503 3560
rect 8573 3580 8617 3596
rect 8573 3560 8582 3580
rect 8602 3560 8617 3580
rect 8573 3554 8617 3560
rect 8667 3584 8716 3596
rect 8667 3564 8685 3584
rect 8705 3564 8716 3584
rect 8667 3554 8716 3564
rect 8781 3580 8825 3596
rect 8781 3560 8790 3580
rect 8810 3560 8825 3580
rect 8781 3554 8825 3560
rect 8875 3584 8924 3596
rect 8875 3564 8893 3584
rect 8913 3564 8924 3584
rect 8875 3554 8924 3564
rect 8994 3580 9038 3596
rect 8994 3560 9003 3580
rect 9023 3560 9038 3580
rect 8994 3554 9038 3560
rect 9088 3584 9137 3596
rect 9088 3564 9106 3584
rect 9126 3564 9137 3584
rect 9088 3554 9137 3564
rect 5593 3491 5642 3501
rect 5593 3471 5604 3491
rect 5624 3471 5642 3491
rect 5593 3459 5642 3471
rect 5692 3495 5736 3501
rect 5692 3475 5707 3495
rect 5727 3475 5736 3495
rect 5692 3459 5736 3475
rect 5806 3491 5855 3501
rect 5806 3471 5817 3491
rect 5837 3471 5855 3491
rect 5806 3459 5855 3471
rect 5905 3495 5949 3501
rect 5905 3475 5920 3495
rect 5940 3475 5949 3495
rect 5905 3459 5949 3475
rect 6014 3491 6063 3501
rect 6014 3471 6025 3491
rect 6045 3471 6063 3491
rect 6014 3459 6063 3471
rect 6113 3495 6157 3501
rect 6113 3475 6128 3495
rect 6148 3475 6157 3495
rect 6113 3459 6157 3475
rect 6227 3495 6271 3501
rect 6227 3475 6236 3495
rect 6256 3475 6271 3495
rect 6227 3459 6271 3475
rect 6321 3491 6370 3501
rect 6321 3471 6339 3491
rect 6359 3471 6370 3491
rect 6321 3459 6370 3471
rect 4147 3278 4196 3290
rect 4147 3258 4158 3278
rect 4178 3258 4196 3278
rect 4147 3248 4196 3258
rect 4246 3274 4290 3290
rect 4246 3254 4261 3274
rect 4281 3254 4290 3274
rect 4246 3248 4290 3254
rect 4360 3274 4404 3290
rect 4360 3254 4369 3274
rect 4389 3254 4404 3274
rect 4360 3248 4404 3254
rect 4454 3278 4503 3290
rect 4454 3258 4472 3278
rect 4492 3258 4503 3278
rect 4454 3248 4503 3258
rect 4568 3274 4612 3290
rect 4568 3254 4577 3274
rect 4597 3254 4612 3274
rect 4568 3248 4612 3254
rect 4662 3278 4711 3290
rect 4662 3258 4680 3278
rect 4700 3258 4711 3278
rect 4662 3248 4711 3258
rect 4781 3274 4825 3290
rect 4781 3254 4790 3274
rect 4810 3254 4825 3274
rect 4781 3248 4825 3254
rect 4875 3278 4924 3290
rect 4875 3258 4893 3278
rect 4913 3258 4924 3278
rect 4875 3248 4924 3258
rect 1380 3185 1429 3195
rect 1380 3165 1391 3185
rect 1411 3165 1429 3185
rect 1380 3153 1429 3165
rect 1479 3189 1523 3195
rect 1479 3169 1494 3189
rect 1514 3169 1523 3189
rect 1479 3153 1523 3169
rect 1593 3185 1642 3195
rect 1593 3165 1604 3185
rect 1624 3165 1642 3185
rect 1593 3153 1642 3165
rect 1692 3189 1736 3195
rect 1692 3169 1707 3189
rect 1727 3169 1736 3189
rect 1692 3153 1736 3169
rect 1801 3185 1850 3195
rect 1801 3165 1812 3185
rect 1832 3165 1850 3185
rect 1801 3153 1850 3165
rect 1900 3189 1944 3195
rect 1900 3169 1915 3189
rect 1935 3169 1944 3189
rect 1900 3153 1944 3169
rect 2014 3189 2058 3195
rect 2014 3169 2023 3189
rect 2043 3169 2058 3189
rect 2014 3153 2058 3169
rect 2108 3185 2157 3195
rect 2108 3165 2126 3185
rect 2146 3165 2157 3185
rect 9428 3257 9477 3269
rect 2108 3153 2157 3165
rect 9428 3237 9439 3257
rect 9459 3237 9477 3257
rect 9428 3227 9477 3237
rect 9527 3253 9571 3269
rect 9527 3233 9542 3253
rect 9562 3233 9571 3253
rect 9527 3227 9571 3233
rect 9641 3253 9685 3269
rect 9641 3233 9650 3253
rect 9670 3233 9685 3253
rect 9641 3227 9685 3233
rect 9735 3257 9784 3269
rect 9735 3237 9753 3257
rect 9773 3237 9784 3257
rect 9735 3227 9784 3237
rect 9849 3253 9893 3269
rect 9849 3233 9858 3253
rect 9878 3233 9893 3253
rect 9849 3227 9893 3233
rect 9943 3257 9992 3269
rect 9943 3237 9961 3257
rect 9981 3237 9992 3257
rect 9943 3227 9992 3237
rect 10062 3253 10106 3269
rect 10062 3233 10071 3253
rect 10091 3233 10106 3253
rect 10062 3227 10106 3233
rect 10156 3257 10205 3269
rect 10156 3237 10174 3257
rect 10194 3237 10205 3257
rect 10156 3227 10205 3237
rect 6661 3164 6710 3174
rect 6661 3144 6672 3164
rect 6692 3144 6710 3164
rect 6661 3132 6710 3144
rect 6760 3168 6804 3174
rect 6760 3148 6775 3168
rect 6795 3148 6804 3168
rect 6760 3132 6804 3148
rect 6874 3164 6923 3174
rect 6874 3144 6885 3164
rect 6905 3144 6923 3164
rect 6874 3132 6923 3144
rect 6973 3168 7017 3174
rect 6973 3148 6988 3168
rect 7008 3148 7017 3168
rect 6973 3132 7017 3148
rect 7082 3164 7131 3174
rect 7082 3144 7093 3164
rect 7113 3144 7131 3164
rect 7082 3132 7131 3144
rect 7181 3168 7225 3174
rect 7181 3148 7196 3168
rect 7216 3148 7225 3168
rect 7181 3132 7225 3148
rect 7295 3168 7339 3174
rect 7295 3148 7304 3168
rect 7324 3148 7339 3168
rect 7295 3132 7339 3148
rect 7389 3164 7438 3174
rect 7389 3144 7407 3164
rect 7427 3144 7438 3164
rect 7389 3132 7438 3144
rect 3134 3044 3183 3056
rect 3134 3024 3145 3044
rect 3165 3024 3183 3044
rect 3134 3014 3183 3024
rect 3233 3040 3277 3056
rect 3233 3020 3248 3040
rect 3268 3020 3277 3040
rect 3233 3014 3277 3020
rect 3347 3040 3391 3056
rect 3347 3020 3356 3040
rect 3376 3020 3391 3040
rect 3347 3014 3391 3020
rect 3441 3044 3490 3056
rect 3441 3024 3459 3044
rect 3479 3024 3490 3044
rect 3441 3014 3490 3024
rect 3555 3040 3599 3056
rect 3555 3020 3564 3040
rect 3584 3020 3599 3040
rect 3555 3014 3599 3020
rect 3649 3044 3698 3056
rect 3649 3024 3667 3044
rect 3687 3024 3698 3044
rect 3649 3014 3698 3024
rect 3768 3040 3812 3056
rect 3768 3020 3777 3040
rect 3797 3020 3812 3040
rect 3768 3014 3812 3020
rect 3862 3044 3911 3056
rect 3862 3024 3880 3044
rect 3900 3024 3911 3044
rect 3862 3014 3911 3024
rect 318 2946 367 2956
rect 318 2926 329 2946
rect 349 2926 367 2946
rect 318 2914 367 2926
rect 417 2950 461 2956
rect 417 2930 432 2950
rect 452 2930 461 2950
rect 417 2914 461 2930
rect 531 2946 580 2956
rect 531 2926 542 2946
rect 562 2926 580 2946
rect 531 2914 580 2926
rect 630 2950 674 2956
rect 630 2930 645 2950
rect 665 2930 674 2950
rect 630 2914 674 2930
rect 739 2946 788 2956
rect 739 2926 750 2946
rect 770 2926 788 2946
rect 739 2914 788 2926
rect 838 2950 882 2956
rect 838 2930 853 2950
rect 873 2930 882 2950
rect 838 2914 882 2930
rect 952 2950 996 2956
rect 952 2930 961 2950
rect 981 2930 996 2950
rect 952 2914 996 2930
rect 1046 2946 1095 2956
rect 1046 2926 1064 2946
rect 1084 2926 1095 2946
rect 1046 2914 1095 2926
rect 8415 3023 8464 3035
rect 8415 3003 8426 3023
rect 8446 3003 8464 3023
rect 8415 2993 8464 3003
rect 8514 3019 8558 3035
rect 8514 2999 8529 3019
rect 8549 2999 8558 3019
rect 8514 2993 8558 2999
rect 8628 3019 8672 3035
rect 8628 2999 8637 3019
rect 8657 2999 8672 3019
rect 8628 2993 8672 2999
rect 8722 3023 8771 3035
rect 8722 3003 8740 3023
rect 8760 3003 8771 3023
rect 8722 2993 8771 3003
rect 8836 3019 8880 3035
rect 8836 2999 8845 3019
rect 8865 2999 8880 3019
rect 8836 2993 8880 2999
rect 8930 3023 8979 3035
rect 8930 3003 8948 3023
rect 8968 3003 8979 3023
rect 8930 2993 8979 3003
rect 9049 3019 9093 3035
rect 9049 2999 9058 3019
rect 9078 2999 9093 3019
rect 9049 2993 9093 2999
rect 9143 3023 9192 3035
rect 9143 3003 9161 3023
rect 9181 3003 9192 3023
rect 9143 2993 9192 3003
rect 5599 2925 5648 2935
rect 5599 2905 5610 2925
rect 5630 2905 5648 2925
rect 5599 2893 5648 2905
rect 5698 2929 5742 2935
rect 5698 2909 5713 2929
rect 5733 2909 5742 2929
rect 5698 2893 5742 2909
rect 5812 2925 5861 2935
rect 5812 2905 5823 2925
rect 5843 2905 5861 2925
rect 5812 2893 5861 2905
rect 5911 2929 5955 2935
rect 5911 2909 5926 2929
rect 5946 2909 5955 2929
rect 5911 2893 5955 2909
rect 6020 2925 6069 2935
rect 6020 2905 6031 2925
rect 6051 2905 6069 2925
rect 6020 2893 6069 2905
rect 6119 2929 6163 2935
rect 6119 2909 6134 2929
rect 6154 2909 6163 2929
rect 6119 2893 6163 2909
rect 6233 2929 6277 2935
rect 6233 2909 6242 2929
rect 6262 2909 6277 2929
rect 6233 2893 6277 2909
rect 6327 2925 6376 2935
rect 6327 2905 6345 2925
rect 6365 2905 6376 2925
rect 6327 2893 6376 2905
rect 4146 2863 4195 2875
rect 4146 2843 4157 2863
rect 4177 2843 4195 2863
rect 4146 2833 4195 2843
rect 4245 2859 4289 2875
rect 4245 2839 4260 2859
rect 4280 2839 4289 2859
rect 4245 2833 4289 2839
rect 4359 2859 4403 2875
rect 4359 2839 4368 2859
rect 4388 2839 4403 2859
rect 4359 2833 4403 2839
rect 4453 2863 4502 2875
rect 4453 2843 4471 2863
rect 4491 2843 4502 2863
rect 4453 2833 4502 2843
rect 4567 2859 4611 2875
rect 4567 2839 4576 2859
rect 4596 2839 4611 2859
rect 4567 2833 4611 2839
rect 4661 2863 4710 2875
rect 4661 2843 4679 2863
rect 4699 2843 4710 2863
rect 4661 2833 4710 2843
rect 4780 2859 4824 2875
rect 4780 2839 4789 2859
rect 4809 2839 4824 2859
rect 4780 2833 4824 2839
rect 4874 2863 4923 2875
rect 4874 2843 4892 2863
rect 4912 2843 4923 2863
rect 4874 2833 4923 2843
rect 1330 2765 1379 2775
rect 1330 2745 1341 2765
rect 1361 2745 1379 2765
rect 1330 2733 1379 2745
rect 1429 2769 1473 2775
rect 1429 2749 1444 2769
rect 1464 2749 1473 2769
rect 1429 2733 1473 2749
rect 1543 2765 1592 2775
rect 1543 2745 1554 2765
rect 1574 2745 1592 2765
rect 1543 2733 1592 2745
rect 1642 2769 1686 2775
rect 1642 2749 1657 2769
rect 1677 2749 1686 2769
rect 1642 2733 1686 2749
rect 1751 2765 1800 2775
rect 1751 2745 1762 2765
rect 1782 2745 1800 2765
rect 1751 2733 1800 2745
rect 1850 2769 1894 2775
rect 1850 2749 1865 2769
rect 1885 2749 1894 2769
rect 1850 2733 1894 2749
rect 1964 2769 2008 2775
rect 1964 2749 1973 2769
rect 1993 2749 2008 2769
rect 1964 2733 2008 2749
rect 2058 2765 2107 2775
rect 2058 2745 2076 2765
rect 2096 2745 2107 2765
rect 2058 2733 2107 2745
rect 9427 2842 9476 2854
rect 9427 2822 9438 2842
rect 9458 2822 9476 2842
rect 9427 2812 9476 2822
rect 9526 2838 9570 2854
rect 9526 2818 9541 2838
rect 9561 2818 9570 2838
rect 9526 2812 9570 2818
rect 9640 2838 9684 2854
rect 9640 2818 9649 2838
rect 9669 2818 9684 2838
rect 9640 2812 9684 2818
rect 9734 2842 9783 2854
rect 9734 2822 9752 2842
rect 9772 2822 9783 2842
rect 9734 2812 9783 2822
rect 9848 2838 9892 2854
rect 9848 2818 9857 2838
rect 9877 2818 9892 2838
rect 9848 2812 9892 2818
rect 9942 2842 9991 2854
rect 9942 2822 9960 2842
rect 9980 2822 9991 2842
rect 9942 2812 9991 2822
rect 10061 2838 10105 2854
rect 10061 2818 10070 2838
rect 10090 2818 10105 2838
rect 10061 2812 10105 2818
rect 10155 2842 10204 2854
rect 10155 2822 10173 2842
rect 10193 2822 10204 2842
rect 10155 2812 10204 2822
rect 6611 2744 6660 2754
rect 6611 2724 6622 2744
rect 6642 2724 6660 2744
rect 6611 2712 6660 2724
rect 6710 2748 6754 2754
rect 6710 2728 6725 2748
rect 6745 2728 6754 2748
rect 6710 2712 6754 2728
rect 6824 2744 6873 2754
rect 6824 2724 6835 2744
rect 6855 2724 6873 2744
rect 6824 2712 6873 2724
rect 6923 2748 6967 2754
rect 6923 2728 6938 2748
rect 6958 2728 6967 2748
rect 6923 2712 6967 2728
rect 7032 2744 7081 2754
rect 7032 2724 7043 2744
rect 7063 2724 7081 2744
rect 7032 2712 7081 2724
rect 7131 2748 7175 2754
rect 7131 2728 7146 2748
rect 7166 2728 7175 2748
rect 7131 2712 7175 2728
rect 7245 2748 7289 2754
rect 7245 2728 7254 2748
rect 7274 2728 7289 2748
rect 7245 2712 7289 2728
rect 7339 2744 7388 2754
rect 7339 2724 7357 2744
rect 7377 2724 7388 2744
rect 7339 2712 7388 2724
rect 2926 2577 2975 2589
rect 2926 2557 2937 2577
rect 2957 2557 2975 2577
rect 2926 2547 2975 2557
rect 3025 2573 3069 2589
rect 3025 2553 3040 2573
rect 3060 2553 3069 2573
rect 3025 2547 3069 2553
rect 3139 2573 3183 2589
rect 3139 2553 3148 2573
rect 3168 2553 3183 2573
rect 3139 2547 3183 2553
rect 3233 2577 3282 2589
rect 3233 2557 3251 2577
rect 3271 2557 3282 2577
rect 3233 2547 3282 2557
rect 3347 2573 3391 2589
rect 3347 2553 3356 2573
rect 3376 2553 3391 2573
rect 3347 2547 3391 2553
rect 3441 2577 3490 2589
rect 3441 2557 3459 2577
rect 3479 2557 3490 2577
rect 3441 2547 3490 2557
rect 3560 2573 3604 2589
rect 3560 2553 3569 2573
rect 3589 2553 3604 2573
rect 3560 2547 3604 2553
rect 3654 2577 3703 2589
rect 3654 2557 3672 2577
rect 3692 2557 3703 2577
rect 3654 2547 3703 2557
rect 317 2531 366 2541
rect 317 2511 328 2531
rect 348 2511 366 2531
rect 317 2499 366 2511
rect 416 2535 460 2541
rect 416 2515 431 2535
rect 451 2515 460 2535
rect 416 2499 460 2515
rect 530 2531 579 2541
rect 530 2511 541 2531
rect 561 2511 579 2531
rect 530 2499 579 2511
rect 629 2535 673 2541
rect 629 2515 644 2535
rect 664 2515 673 2535
rect 629 2499 673 2515
rect 738 2531 787 2541
rect 738 2511 749 2531
rect 769 2511 787 2531
rect 738 2499 787 2511
rect 837 2535 881 2541
rect 837 2515 852 2535
rect 872 2515 881 2535
rect 837 2499 881 2515
rect 951 2535 995 2541
rect 951 2515 960 2535
rect 980 2515 995 2535
rect 951 2499 995 2515
rect 1045 2531 1094 2541
rect 1045 2511 1063 2531
rect 1083 2511 1094 2531
rect 1045 2499 1094 2511
rect 8207 2556 8256 2568
rect 8207 2536 8218 2556
rect 8238 2536 8256 2556
rect 8207 2526 8256 2536
rect 8306 2552 8350 2568
rect 8306 2532 8321 2552
rect 8341 2532 8350 2552
rect 8306 2526 8350 2532
rect 8420 2552 8464 2568
rect 8420 2532 8429 2552
rect 8449 2532 8464 2552
rect 8420 2526 8464 2532
rect 8514 2556 8563 2568
rect 8514 2536 8532 2556
rect 8552 2536 8563 2556
rect 8514 2526 8563 2536
rect 8628 2552 8672 2568
rect 8628 2532 8637 2552
rect 8657 2532 8672 2552
rect 8628 2526 8672 2532
rect 8722 2556 8771 2568
rect 8722 2536 8740 2556
rect 8760 2536 8771 2556
rect 8722 2526 8771 2536
rect 8841 2552 8885 2568
rect 8841 2532 8850 2552
rect 8870 2532 8885 2552
rect 8841 2526 8885 2532
rect 8935 2556 8984 2568
rect 8935 2536 8953 2556
rect 8973 2536 8984 2556
rect 8935 2526 8984 2536
rect 5598 2510 5647 2520
rect 5598 2490 5609 2510
rect 5629 2490 5647 2510
rect 5598 2478 5647 2490
rect 5697 2514 5741 2520
rect 5697 2494 5712 2514
rect 5732 2494 5741 2514
rect 5697 2478 5741 2494
rect 5811 2510 5860 2520
rect 5811 2490 5822 2510
rect 5842 2490 5860 2510
rect 5811 2478 5860 2490
rect 5910 2514 5954 2520
rect 5910 2494 5925 2514
rect 5945 2494 5954 2514
rect 5910 2478 5954 2494
rect 6019 2510 6068 2520
rect 6019 2490 6030 2510
rect 6050 2490 6068 2510
rect 6019 2478 6068 2490
rect 6118 2514 6162 2520
rect 6118 2494 6133 2514
rect 6153 2494 6162 2514
rect 6118 2478 6162 2494
rect 6232 2514 6276 2520
rect 6232 2494 6241 2514
rect 6261 2494 6276 2514
rect 6232 2478 6276 2494
rect 6326 2510 6375 2520
rect 6326 2490 6344 2510
rect 6364 2490 6375 2510
rect 6326 2478 6375 2490
rect 4154 2299 4203 2311
rect 4154 2279 4165 2299
rect 4185 2279 4203 2299
rect 4154 2269 4203 2279
rect 4253 2295 4297 2311
rect 4253 2275 4268 2295
rect 4288 2275 4297 2295
rect 4253 2269 4297 2275
rect 4367 2295 4411 2311
rect 4367 2275 4376 2295
rect 4396 2275 4411 2295
rect 4367 2269 4411 2275
rect 4461 2299 4510 2311
rect 4461 2279 4479 2299
rect 4499 2279 4510 2299
rect 4461 2269 4510 2279
rect 4575 2295 4619 2311
rect 4575 2275 4584 2295
rect 4604 2275 4619 2295
rect 4575 2269 4619 2275
rect 4669 2299 4718 2311
rect 4669 2279 4687 2299
rect 4707 2279 4718 2299
rect 4669 2269 4718 2279
rect 4788 2295 4832 2311
rect 4788 2275 4797 2295
rect 4817 2275 4832 2295
rect 4788 2269 4832 2275
rect 4882 2299 4931 2311
rect 4882 2279 4900 2299
rect 4920 2279 4931 2299
rect 4882 2269 4931 2279
rect 1545 2253 1594 2263
rect 1545 2233 1556 2253
rect 1576 2233 1594 2253
rect 1545 2221 1594 2233
rect 1644 2257 1688 2263
rect 1644 2237 1659 2257
rect 1679 2237 1688 2257
rect 1644 2221 1688 2237
rect 1758 2253 1807 2263
rect 1758 2233 1769 2253
rect 1789 2233 1807 2253
rect 1758 2221 1807 2233
rect 1857 2257 1901 2263
rect 1857 2237 1872 2257
rect 1892 2237 1901 2257
rect 1857 2221 1901 2237
rect 1966 2253 2015 2263
rect 1966 2233 1977 2253
rect 1997 2233 2015 2253
rect 1966 2221 2015 2233
rect 2065 2257 2109 2263
rect 2065 2237 2080 2257
rect 2100 2237 2109 2257
rect 2065 2221 2109 2237
rect 2179 2257 2223 2263
rect 2179 2237 2188 2257
rect 2208 2237 2223 2257
rect 2179 2221 2223 2237
rect 2273 2253 2322 2263
rect 2273 2233 2291 2253
rect 2311 2233 2322 2253
rect 2273 2221 2322 2233
rect 9435 2278 9484 2290
rect 9435 2258 9446 2278
rect 9466 2258 9484 2278
rect 9435 2248 9484 2258
rect 9534 2274 9578 2290
rect 9534 2254 9549 2274
rect 9569 2254 9578 2274
rect 9534 2248 9578 2254
rect 9648 2274 9692 2290
rect 9648 2254 9657 2274
rect 9677 2254 9692 2274
rect 9648 2248 9692 2254
rect 9742 2278 9791 2290
rect 9742 2258 9760 2278
rect 9780 2258 9791 2278
rect 9742 2248 9791 2258
rect 9856 2274 9900 2290
rect 9856 2254 9865 2274
rect 9885 2254 9900 2274
rect 9856 2248 9900 2254
rect 9950 2278 9999 2290
rect 9950 2258 9968 2278
rect 9988 2258 9999 2278
rect 9950 2248 9999 2258
rect 10069 2274 10113 2290
rect 10069 2254 10078 2274
rect 10098 2254 10113 2274
rect 10069 2248 10113 2254
rect 10163 2278 10212 2290
rect 10163 2258 10181 2278
rect 10201 2258 10212 2278
rect 10163 2248 10212 2258
rect 6826 2232 6875 2242
rect 6826 2212 6837 2232
rect 6857 2212 6875 2232
rect 6826 2200 6875 2212
rect 6925 2236 6969 2242
rect 6925 2216 6940 2236
rect 6960 2216 6969 2236
rect 6925 2200 6969 2216
rect 7039 2232 7088 2242
rect 7039 2212 7050 2232
rect 7070 2212 7088 2232
rect 7039 2200 7088 2212
rect 7138 2236 7182 2242
rect 7138 2216 7153 2236
rect 7173 2216 7182 2236
rect 7138 2200 7182 2216
rect 7247 2232 7296 2242
rect 7247 2212 7258 2232
rect 7278 2212 7296 2232
rect 7247 2200 7296 2212
rect 7346 2236 7390 2242
rect 7346 2216 7361 2236
rect 7381 2216 7390 2236
rect 7346 2200 7390 2216
rect 7460 2236 7504 2242
rect 7460 2216 7469 2236
rect 7489 2216 7504 2236
rect 7460 2200 7504 2216
rect 7554 2232 7603 2242
rect 7554 2212 7572 2232
rect 7592 2212 7603 2232
rect 7554 2200 7603 2212
rect 3141 2065 3190 2077
rect 3141 2045 3152 2065
rect 3172 2045 3190 2065
rect 3141 2035 3190 2045
rect 3240 2061 3284 2077
rect 3240 2041 3255 2061
rect 3275 2041 3284 2061
rect 3240 2035 3284 2041
rect 3354 2061 3398 2077
rect 3354 2041 3363 2061
rect 3383 2041 3398 2061
rect 3354 2035 3398 2041
rect 3448 2065 3497 2077
rect 3448 2045 3466 2065
rect 3486 2045 3497 2065
rect 3448 2035 3497 2045
rect 3562 2061 3606 2077
rect 3562 2041 3571 2061
rect 3591 2041 3606 2061
rect 3562 2035 3606 2041
rect 3656 2065 3705 2077
rect 3656 2045 3674 2065
rect 3694 2045 3705 2065
rect 3656 2035 3705 2045
rect 3775 2061 3819 2077
rect 3775 2041 3784 2061
rect 3804 2041 3819 2061
rect 3775 2035 3819 2041
rect 3869 2065 3918 2077
rect 3869 2045 3887 2065
rect 3907 2045 3918 2065
rect 3869 2035 3918 2045
rect 325 1967 374 1977
rect 325 1947 336 1967
rect 356 1947 374 1967
rect 325 1935 374 1947
rect 424 1971 468 1977
rect 424 1951 439 1971
rect 459 1951 468 1971
rect 424 1935 468 1951
rect 538 1967 587 1977
rect 538 1947 549 1967
rect 569 1947 587 1967
rect 538 1935 587 1947
rect 637 1971 681 1977
rect 637 1951 652 1971
rect 672 1951 681 1971
rect 637 1935 681 1951
rect 746 1967 795 1977
rect 746 1947 757 1967
rect 777 1947 795 1967
rect 746 1935 795 1947
rect 845 1971 889 1977
rect 845 1951 860 1971
rect 880 1951 889 1971
rect 845 1935 889 1951
rect 959 1971 1003 1977
rect 959 1951 968 1971
rect 988 1951 1003 1971
rect 959 1935 1003 1951
rect 1053 1967 1102 1977
rect 1053 1947 1071 1967
rect 1091 1947 1102 1967
rect 1053 1935 1102 1947
rect 8422 2044 8471 2056
rect 8422 2024 8433 2044
rect 8453 2024 8471 2044
rect 8422 2014 8471 2024
rect 8521 2040 8565 2056
rect 8521 2020 8536 2040
rect 8556 2020 8565 2040
rect 8521 2014 8565 2020
rect 8635 2040 8679 2056
rect 8635 2020 8644 2040
rect 8664 2020 8679 2040
rect 8635 2014 8679 2020
rect 8729 2044 8778 2056
rect 8729 2024 8747 2044
rect 8767 2024 8778 2044
rect 8729 2014 8778 2024
rect 8843 2040 8887 2056
rect 8843 2020 8852 2040
rect 8872 2020 8887 2040
rect 8843 2014 8887 2020
rect 8937 2044 8986 2056
rect 8937 2024 8955 2044
rect 8975 2024 8986 2044
rect 8937 2014 8986 2024
rect 9056 2040 9100 2056
rect 9056 2020 9065 2040
rect 9085 2020 9100 2040
rect 9056 2014 9100 2020
rect 9150 2044 9199 2056
rect 9150 2024 9168 2044
rect 9188 2024 9199 2044
rect 9150 2014 9199 2024
rect 5606 1946 5655 1956
rect 5606 1926 5617 1946
rect 5637 1926 5655 1946
rect 5606 1914 5655 1926
rect 5705 1950 5749 1956
rect 5705 1930 5720 1950
rect 5740 1930 5749 1950
rect 5705 1914 5749 1930
rect 5819 1946 5868 1956
rect 5819 1926 5830 1946
rect 5850 1926 5868 1946
rect 5819 1914 5868 1926
rect 5918 1950 5962 1956
rect 5918 1930 5933 1950
rect 5953 1930 5962 1950
rect 5918 1914 5962 1930
rect 6027 1946 6076 1956
rect 6027 1926 6038 1946
rect 6058 1926 6076 1946
rect 6027 1914 6076 1926
rect 6126 1950 6170 1956
rect 6126 1930 6141 1950
rect 6161 1930 6170 1950
rect 6126 1914 6170 1930
rect 6240 1950 6284 1956
rect 6240 1930 6249 1950
rect 6269 1930 6284 1950
rect 6240 1914 6284 1930
rect 6334 1946 6383 1956
rect 6334 1926 6352 1946
rect 6372 1926 6383 1946
rect 6334 1914 6383 1926
rect 4153 1884 4202 1896
rect 4153 1864 4164 1884
rect 4184 1864 4202 1884
rect 4153 1854 4202 1864
rect 4252 1880 4296 1896
rect 4252 1860 4267 1880
rect 4287 1860 4296 1880
rect 4252 1854 4296 1860
rect 4366 1880 4410 1896
rect 4366 1860 4375 1880
rect 4395 1860 4410 1880
rect 4366 1854 4410 1860
rect 4460 1884 4509 1896
rect 4460 1864 4478 1884
rect 4498 1864 4509 1884
rect 4460 1854 4509 1864
rect 4574 1880 4618 1896
rect 4574 1860 4583 1880
rect 4603 1860 4618 1880
rect 4574 1854 4618 1860
rect 4668 1884 4717 1896
rect 4668 1864 4686 1884
rect 4706 1864 4717 1884
rect 4668 1854 4717 1864
rect 4787 1880 4831 1896
rect 4787 1860 4796 1880
rect 4816 1860 4831 1880
rect 4787 1854 4831 1860
rect 4881 1884 4930 1896
rect 4881 1864 4899 1884
rect 4919 1864 4930 1884
rect 4881 1854 4930 1864
rect 1337 1786 1386 1796
rect 1337 1766 1348 1786
rect 1368 1766 1386 1786
rect 1337 1754 1386 1766
rect 1436 1790 1480 1796
rect 1436 1770 1451 1790
rect 1471 1770 1480 1790
rect 1436 1754 1480 1770
rect 1550 1786 1599 1796
rect 1550 1766 1561 1786
rect 1581 1766 1599 1786
rect 1550 1754 1599 1766
rect 1649 1790 1693 1796
rect 1649 1770 1664 1790
rect 1684 1770 1693 1790
rect 1649 1754 1693 1770
rect 1758 1786 1807 1796
rect 1758 1766 1769 1786
rect 1789 1766 1807 1786
rect 1758 1754 1807 1766
rect 1857 1790 1901 1796
rect 1857 1770 1872 1790
rect 1892 1770 1901 1790
rect 1857 1754 1901 1770
rect 1971 1790 2015 1796
rect 1971 1770 1980 1790
rect 2000 1770 2015 1790
rect 1971 1754 2015 1770
rect 2065 1786 2114 1796
rect 2065 1766 2083 1786
rect 2103 1766 2114 1786
rect 2065 1754 2114 1766
rect 9434 1863 9483 1875
rect 9434 1843 9445 1863
rect 9465 1843 9483 1863
rect 9434 1833 9483 1843
rect 9533 1859 9577 1875
rect 9533 1839 9548 1859
rect 9568 1839 9577 1859
rect 9533 1833 9577 1839
rect 9647 1859 9691 1875
rect 9647 1839 9656 1859
rect 9676 1839 9691 1859
rect 9647 1833 9691 1839
rect 9741 1863 9790 1875
rect 9741 1843 9759 1863
rect 9779 1843 9790 1863
rect 9741 1833 9790 1843
rect 9855 1859 9899 1875
rect 9855 1839 9864 1859
rect 9884 1839 9899 1859
rect 9855 1833 9899 1839
rect 9949 1863 9998 1875
rect 9949 1843 9967 1863
rect 9987 1843 9998 1863
rect 9949 1833 9998 1843
rect 10068 1859 10112 1875
rect 10068 1839 10077 1859
rect 10097 1839 10112 1859
rect 10068 1833 10112 1839
rect 10162 1863 10211 1875
rect 10162 1843 10180 1863
rect 10200 1843 10211 1863
rect 10162 1833 10211 1843
rect 6618 1765 6667 1775
rect 6618 1745 6629 1765
rect 6649 1745 6667 1765
rect 6618 1733 6667 1745
rect 6717 1769 6761 1775
rect 6717 1749 6732 1769
rect 6752 1749 6761 1769
rect 6717 1733 6761 1749
rect 6831 1765 6880 1775
rect 6831 1745 6842 1765
rect 6862 1745 6880 1765
rect 6831 1733 6880 1745
rect 6930 1769 6974 1775
rect 6930 1749 6945 1769
rect 6965 1749 6974 1769
rect 6930 1733 6974 1749
rect 7039 1765 7088 1775
rect 7039 1745 7050 1765
rect 7070 1745 7088 1765
rect 7039 1733 7088 1745
rect 7138 1769 7182 1775
rect 7138 1749 7153 1769
rect 7173 1749 7182 1769
rect 7138 1733 7182 1749
rect 7252 1769 7296 1775
rect 7252 1749 7261 1769
rect 7281 1749 7296 1769
rect 7252 1733 7296 1749
rect 7346 1765 7395 1775
rect 7346 1745 7364 1765
rect 7384 1745 7395 1765
rect 7346 1733 7395 1745
rect 3091 1645 3140 1657
rect 3091 1625 3102 1645
rect 3122 1625 3140 1645
rect 3091 1615 3140 1625
rect 3190 1641 3234 1657
rect 3190 1621 3205 1641
rect 3225 1621 3234 1641
rect 3190 1615 3234 1621
rect 3304 1641 3348 1657
rect 3304 1621 3313 1641
rect 3333 1621 3348 1641
rect 3304 1615 3348 1621
rect 3398 1645 3447 1657
rect 3398 1625 3416 1645
rect 3436 1625 3447 1645
rect 3398 1615 3447 1625
rect 3512 1641 3556 1657
rect 3512 1621 3521 1641
rect 3541 1621 3556 1641
rect 3512 1615 3556 1621
rect 3606 1645 3655 1657
rect 3606 1625 3624 1645
rect 3644 1625 3655 1645
rect 3606 1615 3655 1625
rect 3725 1641 3769 1657
rect 3725 1621 3734 1641
rect 3754 1621 3769 1641
rect 3725 1615 3769 1621
rect 3819 1645 3868 1657
rect 3819 1625 3837 1645
rect 3857 1625 3868 1645
rect 3819 1615 3868 1625
rect 324 1552 373 1562
rect 324 1532 335 1552
rect 355 1532 373 1552
rect 324 1520 373 1532
rect 423 1556 467 1562
rect 423 1536 438 1556
rect 458 1536 467 1556
rect 423 1520 467 1536
rect 537 1552 586 1562
rect 537 1532 548 1552
rect 568 1532 586 1552
rect 537 1520 586 1532
rect 636 1556 680 1562
rect 636 1536 651 1556
rect 671 1536 680 1556
rect 636 1520 680 1536
rect 745 1552 794 1562
rect 745 1532 756 1552
rect 776 1532 794 1552
rect 745 1520 794 1532
rect 844 1556 888 1562
rect 844 1536 859 1556
rect 879 1536 888 1556
rect 844 1520 888 1536
rect 958 1556 1002 1562
rect 958 1536 967 1556
rect 987 1536 1002 1556
rect 958 1520 1002 1536
rect 1052 1552 1101 1562
rect 1052 1532 1070 1552
rect 1090 1532 1101 1552
rect 8372 1624 8421 1636
rect 1052 1520 1101 1532
rect 8372 1604 8383 1624
rect 8403 1604 8421 1624
rect 8372 1594 8421 1604
rect 8471 1620 8515 1636
rect 8471 1600 8486 1620
rect 8506 1600 8515 1620
rect 8471 1594 8515 1600
rect 8585 1620 8629 1636
rect 8585 1600 8594 1620
rect 8614 1600 8629 1620
rect 8585 1594 8629 1600
rect 8679 1624 8728 1636
rect 8679 1604 8697 1624
rect 8717 1604 8728 1624
rect 8679 1594 8728 1604
rect 8793 1620 8837 1636
rect 8793 1600 8802 1620
rect 8822 1600 8837 1620
rect 8793 1594 8837 1600
rect 8887 1624 8936 1636
rect 8887 1604 8905 1624
rect 8925 1604 8936 1624
rect 8887 1594 8936 1604
rect 9006 1620 9050 1636
rect 9006 1600 9015 1620
rect 9035 1600 9050 1620
rect 9006 1594 9050 1600
rect 9100 1624 9149 1636
rect 9100 1604 9118 1624
rect 9138 1604 9149 1624
rect 9100 1594 9149 1604
rect 5605 1531 5654 1541
rect 5605 1511 5616 1531
rect 5636 1511 5654 1531
rect 5605 1499 5654 1511
rect 5704 1535 5748 1541
rect 5704 1515 5719 1535
rect 5739 1515 5748 1535
rect 5704 1499 5748 1515
rect 5818 1531 5867 1541
rect 5818 1511 5829 1531
rect 5849 1511 5867 1531
rect 5818 1499 5867 1511
rect 5917 1535 5961 1541
rect 5917 1515 5932 1535
rect 5952 1515 5961 1535
rect 5917 1499 5961 1515
rect 6026 1531 6075 1541
rect 6026 1511 6037 1531
rect 6057 1511 6075 1531
rect 6026 1499 6075 1511
rect 6125 1535 6169 1541
rect 6125 1515 6140 1535
rect 6160 1515 6169 1535
rect 6125 1499 6169 1515
rect 6239 1535 6283 1541
rect 6239 1515 6248 1535
rect 6268 1515 6283 1535
rect 6239 1499 6283 1515
rect 6333 1531 6382 1541
rect 6333 1511 6351 1531
rect 6371 1511 6382 1531
rect 6333 1499 6382 1511
rect 4159 1318 4208 1330
rect 4159 1298 4170 1318
rect 4190 1298 4208 1318
rect 4159 1288 4208 1298
rect 4258 1314 4302 1330
rect 4258 1294 4273 1314
rect 4293 1294 4302 1314
rect 4258 1288 4302 1294
rect 4372 1314 4416 1330
rect 4372 1294 4381 1314
rect 4401 1294 4416 1314
rect 4372 1288 4416 1294
rect 4466 1318 4515 1330
rect 4466 1298 4484 1318
rect 4504 1298 4515 1318
rect 4466 1288 4515 1298
rect 4580 1314 4624 1330
rect 4580 1294 4589 1314
rect 4609 1294 4624 1314
rect 4580 1288 4624 1294
rect 4674 1318 4723 1330
rect 4674 1298 4692 1318
rect 4712 1298 4723 1318
rect 4674 1288 4723 1298
rect 4793 1314 4837 1330
rect 4793 1294 4802 1314
rect 4822 1294 4837 1314
rect 4793 1288 4837 1294
rect 4887 1318 4936 1330
rect 4887 1298 4905 1318
rect 4925 1298 4936 1318
rect 4887 1288 4936 1298
rect 1392 1225 1441 1235
rect 1392 1205 1403 1225
rect 1423 1205 1441 1225
rect 1392 1193 1441 1205
rect 1491 1229 1535 1235
rect 1491 1209 1506 1229
rect 1526 1209 1535 1229
rect 1491 1193 1535 1209
rect 1605 1225 1654 1235
rect 1605 1205 1616 1225
rect 1636 1205 1654 1225
rect 1605 1193 1654 1205
rect 1704 1229 1748 1235
rect 1704 1209 1719 1229
rect 1739 1209 1748 1229
rect 1704 1193 1748 1209
rect 1813 1225 1862 1235
rect 1813 1205 1824 1225
rect 1844 1205 1862 1225
rect 1813 1193 1862 1205
rect 1912 1229 1956 1235
rect 1912 1209 1927 1229
rect 1947 1209 1956 1229
rect 1912 1193 1956 1209
rect 2026 1229 2070 1235
rect 2026 1209 2035 1229
rect 2055 1209 2070 1229
rect 2026 1193 2070 1209
rect 2120 1225 2169 1235
rect 2120 1205 2138 1225
rect 2158 1205 2169 1225
rect 9440 1297 9489 1309
rect 2120 1193 2169 1205
rect 9440 1277 9451 1297
rect 9471 1277 9489 1297
rect 9440 1267 9489 1277
rect 9539 1293 9583 1309
rect 9539 1273 9554 1293
rect 9574 1273 9583 1293
rect 9539 1267 9583 1273
rect 9653 1293 9697 1309
rect 9653 1273 9662 1293
rect 9682 1273 9697 1293
rect 9653 1267 9697 1273
rect 9747 1297 9796 1309
rect 9747 1277 9765 1297
rect 9785 1277 9796 1297
rect 9747 1267 9796 1277
rect 9861 1293 9905 1309
rect 9861 1273 9870 1293
rect 9890 1273 9905 1293
rect 9861 1267 9905 1273
rect 9955 1297 10004 1309
rect 9955 1277 9973 1297
rect 9993 1277 10004 1297
rect 9955 1267 10004 1277
rect 10074 1293 10118 1309
rect 10074 1273 10083 1293
rect 10103 1273 10118 1293
rect 10074 1267 10118 1273
rect 10168 1297 10217 1309
rect 10168 1277 10186 1297
rect 10206 1277 10217 1297
rect 10168 1267 10217 1277
rect 6673 1204 6722 1214
rect 6673 1184 6684 1204
rect 6704 1184 6722 1204
rect 6673 1172 6722 1184
rect 6772 1208 6816 1214
rect 6772 1188 6787 1208
rect 6807 1188 6816 1208
rect 6772 1172 6816 1188
rect 6886 1204 6935 1214
rect 6886 1184 6897 1204
rect 6917 1184 6935 1204
rect 6886 1172 6935 1184
rect 6985 1208 7029 1214
rect 6985 1188 7000 1208
rect 7020 1188 7029 1208
rect 6985 1172 7029 1188
rect 7094 1204 7143 1214
rect 7094 1184 7105 1204
rect 7125 1184 7143 1204
rect 7094 1172 7143 1184
rect 7193 1208 7237 1214
rect 7193 1188 7208 1208
rect 7228 1188 7237 1208
rect 7193 1172 7237 1188
rect 7307 1208 7351 1214
rect 7307 1188 7316 1208
rect 7336 1188 7351 1208
rect 7307 1172 7351 1188
rect 7401 1204 7450 1214
rect 7401 1184 7419 1204
rect 7439 1184 7450 1204
rect 7401 1172 7450 1184
rect 3146 1084 3195 1096
rect 3146 1064 3157 1084
rect 3177 1064 3195 1084
rect 3146 1054 3195 1064
rect 3245 1080 3289 1096
rect 3245 1060 3260 1080
rect 3280 1060 3289 1080
rect 3245 1054 3289 1060
rect 3359 1080 3403 1096
rect 3359 1060 3368 1080
rect 3388 1060 3403 1080
rect 3359 1054 3403 1060
rect 3453 1084 3502 1096
rect 3453 1064 3471 1084
rect 3491 1064 3502 1084
rect 3453 1054 3502 1064
rect 3567 1080 3611 1096
rect 3567 1060 3576 1080
rect 3596 1060 3611 1080
rect 3567 1054 3611 1060
rect 3661 1084 3710 1096
rect 3661 1064 3679 1084
rect 3699 1064 3710 1084
rect 3661 1054 3710 1064
rect 3780 1080 3824 1096
rect 3780 1060 3789 1080
rect 3809 1060 3824 1080
rect 3780 1054 3824 1060
rect 3874 1084 3923 1096
rect 3874 1064 3892 1084
rect 3912 1064 3923 1084
rect 3874 1054 3923 1064
rect 330 986 379 996
rect 330 966 341 986
rect 361 966 379 986
rect 330 954 379 966
rect 429 990 473 996
rect 429 970 444 990
rect 464 970 473 990
rect 429 954 473 970
rect 543 986 592 996
rect 543 966 554 986
rect 574 966 592 986
rect 543 954 592 966
rect 642 990 686 996
rect 642 970 657 990
rect 677 970 686 990
rect 642 954 686 970
rect 751 986 800 996
rect 751 966 762 986
rect 782 966 800 986
rect 751 954 800 966
rect 850 990 894 996
rect 850 970 865 990
rect 885 970 894 990
rect 850 954 894 970
rect 964 990 1008 996
rect 964 970 973 990
rect 993 970 1008 990
rect 964 954 1008 970
rect 1058 986 1107 996
rect 1058 966 1076 986
rect 1096 966 1107 986
rect 1058 954 1107 966
rect 8427 1063 8476 1075
rect 8427 1043 8438 1063
rect 8458 1043 8476 1063
rect 8427 1033 8476 1043
rect 8526 1059 8570 1075
rect 8526 1039 8541 1059
rect 8561 1039 8570 1059
rect 8526 1033 8570 1039
rect 8640 1059 8684 1075
rect 8640 1039 8649 1059
rect 8669 1039 8684 1059
rect 8640 1033 8684 1039
rect 8734 1063 8783 1075
rect 8734 1043 8752 1063
rect 8772 1043 8783 1063
rect 8734 1033 8783 1043
rect 8848 1059 8892 1075
rect 8848 1039 8857 1059
rect 8877 1039 8892 1059
rect 8848 1033 8892 1039
rect 8942 1063 8991 1075
rect 8942 1043 8960 1063
rect 8980 1043 8991 1063
rect 8942 1033 8991 1043
rect 9061 1059 9105 1075
rect 9061 1039 9070 1059
rect 9090 1039 9105 1059
rect 9061 1033 9105 1039
rect 9155 1063 9204 1075
rect 9155 1043 9173 1063
rect 9193 1043 9204 1063
rect 9155 1033 9204 1043
rect 5611 965 5660 975
rect 5611 945 5622 965
rect 5642 945 5660 965
rect 5611 933 5660 945
rect 5710 969 5754 975
rect 5710 949 5725 969
rect 5745 949 5754 969
rect 5710 933 5754 949
rect 5824 965 5873 975
rect 5824 945 5835 965
rect 5855 945 5873 965
rect 5824 933 5873 945
rect 5923 969 5967 975
rect 5923 949 5938 969
rect 5958 949 5967 969
rect 5923 933 5967 949
rect 6032 965 6081 975
rect 6032 945 6043 965
rect 6063 945 6081 965
rect 6032 933 6081 945
rect 6131 969 6175 975
rect 6131 949 6146 969
rect 6166 949 6175 969
rect 6131 933 6175 949
rect 6245 969 6289 975
rect 6245 949 6254 969
rect 6274 949 6289 969
rect 6245 933 6289 949
rect 6339 965 6388 975
rect 6339 945 6357 965
rect 6377 945 6388 965
rect 6339 933 6388 945
rect 4158 903 4207 915
rect 4158 883 4169 903
rect 4189 883 4207 903
rect 4158 873 4207 883
rect 4257 899 4301 915
rect 4257 879 4272 899
rect 4292 879 4301 899
rect 4257 873 4301 879
rect 4371 899 4415 915
rect 4371 879 4380 899
rect 4400 879 4415 899
rect 4371 873 4415 879
rect 4465 903 4514 915
rect 4465 883 4483 903
rect 4503 883 4514 903
rect 4465 873 4514 883
rect 4579 899 4623 915
rect 4579 879 4588 899
rect 4608 879 4623 899
rect 4579 873 4623 879
rect 4673 903 4722 915
rect 4673 883 4691 903
rect 4711 883 4722 903
rect 4673 873 4722 883
rect 4792 899 4836 915
rect 4792 879 4801 899
rect 4821 879 4836 899
rect 4792 873 4836 879
rect 4886 903 4935 915
rect 4886 883 4904 903
rect 4924 883 4935 903
rect 4886 873 4935 883
rect 1342 805 1391 815
rect 1342 785 1353 805
rect 1373 785 1391 805
rect 1342 773 1391 785
rect 1441 809 1485 815
rect 1441 789 1456 809
rect 1476 789 1485 809
rect 1441 773 1485 789
rect 1555 805 1604 815
rect 1555 785 1566 805
rect 1586 785 1604 805
rect 1555 773 1604 785
rect 1654 809 1698 815
rect 1654 789 1669 809
rect 1689 789 1698 809
rect 1654 773 1698 789
rect 1763 805 1812 815
rect 1763 785 1774 805
rect 1794 785 1812 805
rect 1763 773 1812 785
rect 1862 809 1906 815
rect 1862 789 1877 809
rect 1897 789 1906 809
rect 1862 773 1906 789
rect 1976 809 2020 815
rect 1976 789 1985 809
rect 2005 789 2020 809
rect 1976 773 2020 789
rect 2070 805 2119 815
rect 2070 785 2088 805
rect 2108 785 2119 805
rect 2070 773 2119 785
rect 9439 882 9488 894
rect 9439 862 9450 882
rect 9470 862 9488 882
rect 9439 852 9488 862
rect 9538 878 9582 894
rect 9538 858 9553 878
rect 9573 858 9582 878
rect 9538 852 9582 858
rect 9652 878 9696 894
rect 9652 858 9661 878
rect 9681 858 9696 878
rect 9652 852 9696 858
rect 9746 882 9795 894
rect 9746 862 9764 882
rect 9784 862 9795 882
rect 9746 852 9795 862
rect 9860 878 9904 894
rect 9860 858 9869 878
rect 9889 858 9904 878
rect 9860 852 9904 858
rect 9954 882 10003 894
rect 9954 862 9972 882
rect 9992 862 10003 882
rect 9954 852 10003 862
rect 10073 878 10117 894
rect 10073 858 10082 878
rect 10102 858 10117 878
rect 10073 852 10117 858
rect 10167 882 10216 894
rect 10167 862 10185 882
rect 10205 862 10216 882
rect 10167 852 10216 862
rect 6623 784 6672 794
rect 6623 764 6634 784
rect 6654 764 6672 784
rect 6623 752 6672 764
rect 6722 788 6766 794
rect 6722 768 6737 788
rect 6757 768 6766 788
rect 6722 752 6766 768
rect 6836 784 6885 794
rect 6836 764 6847 784
rect 6867 764 6885 784
rect 6836 752 6885 764
rect 6935 788 6979 794
rect 6935 768 6950 788
rect 6970 768 6979 788
rect 6935 752 6979 768
rect 7044 784 7093 794
rect 7044 764 7055 784
rect 7075 764 7093 784
rect 7044 752 7093 764
rect 7143 788 7187 794
rect 7143 768 7158 788
rect 7178 768 7187 788
rect 7143 752 7187 768
rect 7257 788 7301 794
rect 7257 768 7266 788
rect 7286 768 7301 788
rect 7257 752 7301 768
rect 7351 784 7400 794
rect 7351 764 7369 784
rect 7389 764 7400 784
rect 7351 752 7400 764
rect 329 571 378 581
rect 329 551 340 571
rect 360 551 378 571
rect 329 539 378 551
rect 428 575 472 581
rect 428 555 443 575
rect 463 555 472 575
rect 428 539 472 555
rect 542 571 591 581
rect 542 551 553 571
rect 573 551 591 571
rect 542 539 591 551
rect 641 575 685 581
rect 641 555 656 575
rect 676 555 685 575
rect 641 539 685 555
rect 750 571 799 581
rect 750 551 761 571
rect 781 551 799 571
rect 750 539 799 551
rect 849 575 893 581
rect 849 555 864 575
rect 884 555 893 575
rect 849 539 893 555
rect 963 575 1007 581
rect 963 555 972 575
rect 992 555 1007 575
rect 963 539 1007 555
rect 1057 571 1106 581
rect 1057 551 1075 571
rect 1095 551 1106 571
rect 1057 539 1106 551
rect 5610 550 5659 560
rect 5610 530 5621 550
rect 5641 530 5659 550
rect 5610 518 5659 530
rect 5709 554 5753 560
rect 5709 534 5724 554
rect 5744 534 5753 554
rect 5709 518 5753 534
rect 5823 550 5872 560
rect 5823 530 5834 550
rect 5854 530 5872 550
rect 5823 518 5872 530
rect 5922 554 5966 560
rect 5922 534 5937 554
rect 5957 534 5966 554
rect 5922 518 5966 534
rect 6031 550 6080 560
rect 6031 530 6042 550
rect 6062 530 6080 550
rect 6031 518 6080 530
rect 6130 554 6174 560
rect 6130 534 6145 554
rect 6165 534 6174 554
rect 6130 518 6174 534
rect 6244 554 6288 560
rect 6244 534 6253 554
rect 6273 534 6288 554
rect 6244 518 6288 534
rect 6338 550 6387 560
rect 6338 530 6356 550
rect 6376 530 6387 550
rect 6338 518 6387 530
rect 1732 90 1781 100
rect 1732 70 1743 90
rect 1763 70 1781 90
rect 1732 58 1781 70
rect 1831 94 1875 100
rect 1831 74 1846 94
rect 1866 74 1875 94
rect 1831 58 1875 74
rect 1945 90 1994 100
rect 1945 70 1956 90
rect 1976 70 1994 90
rect 1945 58 1994 70
rect 2044 94 2088 100
rect 2044 74 2059 94
rect 2079 74 2088 94
rect 2044 58 2088 74
rect 2153 90 2202 100
rect 2153 70 2164 90
rect 2184 70 2202 90
rect 2153 58 2202 70
rect 2252 94 2296 100
rect 2252 74 2267 94
rect 2287 74 2296 94
rect 2252 58 2296 74
rect 2366 94 2410 100
rect 2366 74 2375 94
rect 2395 74 2410 94
rect 2366 58 2410 74
rect 2460 90 2509 100
rect 2460 70 2478 90
rect 2498 70 2509 90
rect 2460 58 2509 70
rect 7013 69 7062 79
rect 7013 49 7024 69
rect 7044 49 7062 69
rect 7013 37 7062 49
rect 7112 73 7156 79
rect 7112 53 7127 73
rect 7147 53 7156 73
rect 7112 37 7156 53
rect 7226 69 7275 79
rect 7226 49 7237 69
rect 7257 49 7275 69
rect 7226 37 7275 49
rect 7325 73 7369 79
rect 7325 53 7340 73
rect 7360 53 7369 73
rect 7325 37 7369 53
rect 7434 69 7483 79
rect 7434 49 7445 69
rect 7465 49 7483 69
rect 7434 37 7483 49
rect 7533 73 7577 79
rect 7533 53 7548 73
rect 7568 53 7577 73
rect 7533 37 7577 53
rect 7647 73 7691 79
rect 7647 53 7656 73
rect 7676 53 7691 73
rect 7647 37 7691 53
rect 7741 69 7790 79
rect 7741 49 7759 69
rect 7779 49 7790 69
rect 7741 37 7790 49
rect 4822 2 4871 12
rect 4822 -18 4833 2
rect 4853 -18 4871 2
rect 4822 -30 4871 -18
rect 4921 6 4965 12
rect 4921 -14 4936 6
rect 4956 -14 4965 6
rect 4921 -30 4965 -14
rect 5035 2 5084 12
rect 5035 -18 5046 2
rect 5066 -18 5084 2
rect 5035 -30 5084 -18
rect 5134 6 5178 12
rect 5134 -14 5149 6
rect 5169 -14 5178 6
rect 5134 -30 5178 -14
rect 5243 2 5292 12
rect 5243 -18 5254 2
rect 5274 -18 5292 2
rect 5243 -30 5292 -18
rect 5342 6 5386 12
rect 5342 -14 5357 6
rect 5377 -14 5386 6
rect 5342 -30 5386 -14
rect 5456 6 5500 12
rect 5456 -14 5465 6
rect 5485 -14 5500 6
rect 5456 -30 5500 -14
rect 5550 2 5599 12
rect 5550 -18 5568 2
rect 5588 -18 5599 2
rect 5550 -30 5599 -18
<< pdiff >>
rect 298 7993 342 8031
rect 298 7973 310 7993
rect 330 7973 342 7993
rect 298 7931 342 7973
rect 392 7993 434 8031
rect 392 7973 406 7993
rect 426 7973 434 7993
rect 392 7931 434 7973
rect 511 7993 555 8031
rect 511 7973 523 7993
rect 543 7973 555 7993
rect 511 7931 555 7973
rect 605 7993 647 8031
rect 605 7973 619 7993
rect 639 7973 647 7993
rect 605 7931 647 7973
rect 719 7993 763 8031
rect 719 7973 731 7993
rect 751 7973 763 7993
rect 719 7931 763 7973
rect 813 7993 855 8031
rect 813 7973 827 7993
rect 847 7973 855 7993
rect 813 7931 855 7973
rect 929 7993 971 8031
rect 929 7973 937 7993
rect 957 7973 971 7993
rect 929 7931 971 7973
rect 1021 8000 1066 8031
rect 4127 8027 4171 8069
rect 4127 8007 4139 8027
rect 4159 8007 4171 8027
rect 4127 8000 4171 8007
rect 1021 7993 1065 8000
rect 1021 7973 1033 7993
rect 1053 7973 1065 7993
rect 1021 7931 1065 7973
rect 4126 7969 4171 8000
rect 4221 8027 4263 8069
rect 4221 8007 4235 8027
rect 4255 8007 4263 8027
rect 4221 7969 4263 8007
rect 4337 8027 4379 8069
rect 4337 8007 4345 8027
rect 4365 8007 4379 8027
rect 4337 7969 4379 8007
rect 4429 8027 4473 8069
rect 4429 8007 4441 8027
rect 4461 8007 4473 8027
rect 4429 7969 4473 8007
rect 4545 8027 4587 8069
rect 4545 8007 4553 8027
rect 4573 8007 4587 8027
rect 4545 7969 4587 8007
rect 4637 8027 4681 8069
rect 4637 8007 4649 8027
rect 4669 8007 4681 8027
rect 4637 7969 4681 8007
rect 4758 8027 4800 8069
rect 4758 8007 4766 8027
rect 4786 8007 4800 8027
rect 4758 7969 4800 8007
rect 4850 8027 4894 8069
rect 4850 8007 4862 8027
rect 4882 8007 4894 8027
rect 4850 7969 4894 8007
rect 5579 7972 5623 8010
rect 5579 7952 5591 7972
rect 5611 7952 5623 7972
rect 1310 7812 1354 7850
rect 1310 7792 1322 7812
rect 1342 7792 1354 7812
rect 1310 7750 1354 7792
rect 1404 7812 1446 7850
rect 1404 7792 1418 7812
rect 1438 7792 1446 7812
rect 1404 7750 1446 7792
rect 1523 7812 1567 7850
rect 1523 7792 1535 7812
rect 1555 7792 1567 7812
rect 1523 7750 1567 7792
rect 1617 7812 1659 7850
rect 1617 7792 1631 7812
rect 1651 7792 1659 7812
rect 1617 7750 1659 7792
rect 1731 7812 1775 7850
rect 1731 7792 1743 7812
rect 1763 7792 1775 7812
rect 1731 7750 1775 7792
rect 1825 7812 1867 7850
rect 1825 7792 1839 7812
rect 1859 7792 1867 7812
rect 1825 7750 1867 7792
rect 1941 7812 1983 7850
rect 1941 7792 1949 7812
rect 1969 7792 1983 7812
rect 1941 7750 1983 7792
rect 2033 7819 2078 7850
rect 5579 7910 5623 7952
rect 5673 7972 5715 8010
rect 5673 7952 5687 7972
rect 5707 7952 5715 7972
rect 5673 7910 5715 7952
rect 5792 7972 5836 8010
rect 5792 7952 5804 7972
rect 5824 7952 5836 7972
rect 5792 7910 5836 7952
rect 5886 7972 5928 8010
rect 5886 7952 5900 7972
rect 5920 7952 5928 7972
rect 5886 7910 5928 7952
rect 6000 7972 6044 8010
rect 6000 7952 6012 7972
rect 6032 7952 6044 7972
rect 6000 7910 6044 7952
rect 6094 7972 6136 8010
rect 6094 7952 6108 7972
rect 6128 7952 6136 7972
rect 6094 7910 6136 7952
rect 6210 7972 6252 8010
rect 6210 7952 6218 7972
rect 6238 7952 6252 7972
rect 6210 7910 6252 7952
rect 6302 7979 6347 8010
rect 9408 8006 9452 8048
rect 9408 7986 9420 8006
rect 9440 7986 9452 8006
rect 9408 7979 9452 7986
rect 6302 7972 6346 7979
rect 6302 7952 6314 7972
rect 6334 7952 6346 7972
rect 6302 7910 6346 7952
rect 9407 7948 9452 7979
rect 9502 8006 9544 8048
rect 9502 7986 9516 8006
rect 9536 7986 9544 8006
rect 9502 7948 9544 7986
rect 9618 8006 9660 8048
rect 9618 7986 9626 8006
rect 9646 7986 9660 8006
rect 9618 7948 9660 7986
rect 9710 8006 9754 8048
rect 9710 7986 9722 8006
rect 9742 7986 9754 8006
rect 9710 7948 9754 7986
rect 9826 8006 9868 8048
rect 9826 7986 9834 8006
rect 9854 7986 9868 8006
rect 9826 7948 9868 7986
rect 9918 8006 9962 8048
rect 9918 7986 9930 8006
rect 9950 7986 9962 8006
rect 9918 7948 9962 7986
rect 10039 8006 10081 8048
rect 10039 7986 10047 8006
rect 10067 7986 10081 8006
rect 10039 7948 10081 7986
rect 10131 8006 10175 8048
rect 10131 7986 10143 8006
rect 10163 7986 10175 8006
rect 10131 7948 10175 7986
rect 2033 7812 2077 7819
rect 2033 7792 2045 7812
rect 2065 7792 2077 7812
rect 2033 7750 2077 7792
rect 3114 7793 3158 7835
rect 3114 7773 3126 7793
rect 3146 7773 3158 7793
rect 3114 7766 3158 7773
rect 3113 7735 3158 7766
rect 3208 7793 3250 7835
rect 3208 7773 3222 7793
rect 3242 7773 3250 7793
rect 3208 7735 3250 7773
rect 3324 7793 3366 7835
rect 3324 7773 3332 7793
rect 3352 7773 3366 7793
rect 3324 7735 3366 7773
rect 3416 7793 3460 7835
rect 3416 7773 3428 7793
rect 3448 7773 3460 7793
rect 3416 7735 3460 7773
rect 3532 7793 3574 7835
rect 3532 7773 3540 7793
rect 3560 7773 3574 7793
rect 3532 7735 3574 7773
rect 3624 7793 3668 7835
rect 3624 7773 3636 7793
rect 3656 7773 3668 7793
rect 3624 7735 3668 7773
rect 3745 7793 3787 7835
rect 3745 7773 3753 7793
rect 3773 7773 3787 7793
rect 3745 7735 3787 7773
rect 3837 7793 3881 7835
rect 3837 7773 3849 7793
rect 3869 7773 3881 7793
rect 6591 7791 6635 7829
rect 3837 7735 3881 7773
rect 6591 7771 6603 7791
rect 6623 7771 6635 7791
rect 6591 7729 6635 7771
rect 6685 7791 6727 7829
rect 6685 7771 6699 7791
rect 6719 7771 6727 7791
rect 6685 7729 6727 7771
rect 6804 7791 6848 7829
rect 6804 7771 6816 7791
rect 6836 7771 6848 7791
rect 6804 7729 6848 7771
rect 6898 7791 6940 7829
rect 6898 7771 6912 7791
rect 6932 7771 6940 7791
rect 6898 7729 6940 7771
rect 7012 7791 7056 7829
rect 7012 7771 7024 7791
rect 7044 7771 7056 7791
rect 7012 7729 7056 7771
rect 7106 7791 7148 7829
rect 7106 7771 7120 7791
rect 7140 7771 7148 7791
rect 7106 7729 7148 7771
rect 7222 7791 7264 7829
rect 7222 7771 7230 7791
rect 7250 7771 7264 7791
rect 7222 7729 7264 7771
rect 7314 7798 7359 7829
rect 7314 7791 7358 7798
rect 7314 7771 7326 7791
rect 7346 7771 7358 7791
rect 7314 7729 7358 7771
rect 8395 7772 8439 7814
rect 8395 7752 8407 7772
rect 8427 7752 8439 7772
rect 8395 7745 8439 7752
rect 297 7578 341 7616
rect 297 7558 309 7578
rect 329 7558 341 7578
rect 297 7516 341 7558
rect 391 7578 433 7616
rect 391 7558 405 7578
rect 425 7558 433 7578
rect 391 7516 433 7558
rect 510 7578 554 7616
rect 510 7558 522 7578
rect 542 7558 554 7578
rect 510 7516 554 7558
rect 604 7578 646 7616
rect 604 7558 618 7578
rect 638 7558 646 7578
rect 604 7516 646 7558
rect 718 7578 762 7616
rect 718 7558 730 7578
rect 750 7558 762 7578
rect 718 7516 762 7558
rect 812 7578 854 7616
rect 812 7558 826 7578
rect 846 7558 854 7578
rect 812 7516 854 7558
rect 928 7578 970 7616
rect 928 7558 936 7578
rect 956 7558 970 7578
rect 928 7516 970 7558
rect 1020 7585 1065 7616
rect 4126 7612 4170 7654
rect 4126 7592 4138 7612
rect 4158 7592 4170 7612
rect 4126 7585 4170 7592
rect 1020 7578 1064 7585
rect 1020 7558 1032 7578
rect 1052 7558 1064 7578
rect 1020 7516 1064 7558
rect 4125 7554 4170 7585
rect 4220 7612 4262 7654
rect 4220 7592 4234 7612
rect 4254 7592 4262 7612
rect 4220 7554 4262 7592
rect 4336 7612 4378 7654
rect 4336 7592 4344 7612
rect 4364 7592 4378 7612
rect 4336 7554 4378 7592
rect 4428 7612 4472 7654
rect 4428 7592 4440 7612
rect 4460 7592 4472 7612
rect 4428 7554 4472 7592
rect 4544 7612 4586 7654
rect 4544 7592 4552 7612
rect 4572 7592 4586 7612
rect 4544 7554 4586 7592
rect 4636 7612 4680 7654
rect 4636 7592 4648 7612
rect 4668 7592 4680 7612
rect 4636 7554 4680 7592
rect 4757 7612 4799 7654
rect 4757 7592 4765 7612
rect 4785 7592 4799 7612
rect 4757 7554 4799 7592
rect 4849 7612 4893 7654
rect 8394 7714 8439 7745
rect 8489 7772 8531 7814
rect 8489 7752 8503 7772
rect 8523 7752 8531 7772
rect 8489 7714 8531 7752
rect 8605 7772 8647 7814
rect 8605 7752 8613 7772
rect 8633 7752 8647 7772
rect 8605 7714 8647 7752
rect 8697 7772 8741 7814
rect 8697 7752 8709 7772
rect 8729 7752 8741 7772
rect 8697 7714 8741 7752
rect 8813 7772 8855 7814
rect 8813 7752 8821 7772
rect 8841 7752 8855 7772
rect 8813 7714 8855 7752
rect 8905 7772 8949 7814
rect 8905 7752 8917 7772
rect 8937 7752 8949 7772
rect 8905 7714 8949 7752
rect 9026 7772 9068 7814
rect 9026 7752 9034 7772
rect 9054 7752 9068 7772
rect 9026 7714 9068 7752
rect 9118 7772 9162 7814
rect 9118 7752 9130 7772
rect 9150 7752 9162 7772
rect 9118 7714 9162 7752
rect 4849 7592 4861 7612
rect 4881 7592 4893 7612
rect 4849 7554 4893 7592
rect 5578 7557 5622 7595
rect 5578 7537 5590 7557
rect 5610 7537 5622 7557
rect 5578 7495 5622 7537
rect 5672 7557 5714 7595
rect 5672 7537 5686 7557
rect 5706 7537 5714 7557
rect 5672 7495 5714 7537
rect 5791 7557 5835 7595
rect 5791 7537 5803 7557
rect 5823 7537 5835 7557
rect 5791 7495 5835 7537
rect 5885 7557 5927 7595
rect 5885 7537 5899 7557
rect 5919 7537 5927 7557
rect 5885 7495 5927 7537
rect 5999 7557 6043 7595
rect 5999 7537 6011 7557
rect 6031 7537 6043 7557
rect 5999 7495 6043 7537
rect 6093 7557 6135 7595
rect 6093 7537 6107 7557
rect 6127 7537 6135 7557
rect 6093 7495 6135 7537
rect 6209 7557 6251 7595
rect 6209 7537 6217 7557
rect 6237 7537 6251 7557
rect 6209 7495 6251 7537
rect 6301 7564 6346 7595
rect 9407 7591 9451 7633
rect 9407 7571 9419 7591
rect 9439 7571 9451 7591
rect 9407 7564 9451 7571
rect 6301 7557 6345 7564
rect 6301 7537 6313 7557
rect 6333 7537 6345 7557
rect 6301 7495 6345 7537
rect 9406 7533 9451 7564
rect 9501 7591 9543 7633
rect 9501 7571 9515 7591
rect 9535 7571 9543 7591
rect 9501 7533 9543 7571
rect 9617 7591 9659 7633
rect 9617 7571 9625 7591
rect 9645 7571 9659 7591
rect 9617 7533 9659 7571
rect 9709 7591 9753 7633
rect 9709 7571 9721 7591
rect 9741 7571 9753 7591
rect 9709 7533 9753 7571
rect 9825 7591 9867 7633
rect 9825 7571 9833 7591
rect 9853 7571 9867 7591
rect 9825 7533 9867 7571
rect 9917 7591 9961 7633
rect 9917 7571 9929 7591
rect 9949 7571 9961 7591
rect 9917 7533 9961 7571
rect 10038 7591 10080 7633
rect 10038 7571 10046 7591
rect 10066 7571 10080 7591
rect 10038 7533 10080 7571
rect 10130 7591 10174 7633
rect 10130 7571 10142 7591
rect 10162 7571 10174 7591
rect 10130 7533 10174 7571
rect 3064 7373 3108 7415
rect 3064 7353 3076 7373
rect 3096 7353 3108 7373
rect 3064 7346 3108 7353
rect 3063 7315 3108 7346
rect 3158 7373 3200 7415
rect 3158 7353 3172 7373
rect 3192 7353 3200 7373
rect 3158 7315 3200 7353
rect 3274 7373 3316 7415
rect 3274 7353 3282 7373
rect 3302 7353 3316 7373
rect 3274 7315 3316 7353
rect 3366 7373 3410 7415
rect 3366 7353 3378 7373
rect 3398 7353 3410 7373
rect 3366 7315 3410 7353
rect 3482 7373 3524 7415
rect 3482 7353 3490 7373
rect 3510 7353 3524 7373
rect 3482 7315 3524 7353
rect 3574 7373 3618 7415
rect 3574 7353 3586 7373
rect 3606 7353 3618 7373
rect 3574 7315 3618 7353
rect 3695 7373 3737 7415
rect 3695 7353 3703 7373
rect 3723 7353 3737 7373
rect 3695 7315 3737 7353
rect 3787 7373 3831 7415
rect 3787 7353 3799 7373
rect 3819 7353 3831 7373
rect 3787 7315 3831 7353
rect 8345 7352 8389 7394
rect 8345 7332 8357 7352
rect 8377 7332 8389 7352
rect 8345 7325 8389 7332
rect 8344 7294 8389 7325
rect 8439 7352 8481 7394
rect 8439 7332 8453 7352
rect 8473 7332 8481 7352
rect 8439 7294 8481 7332
rect 8555 7352 8597 7394
rect 8555 7332 8563 7352
rect 8583 7332 8597 7352
rect 8555 7294 8597 7332
rect 8647 7352 8691 7394
rect 8647 7332 8659 7352
rect 8679 7332 8691 7352
rect 8647 7294 8691 7332
rect 8763 7352 8805 7394
rect 8763 7332 8771 7352
rect 8791 7332 8805 7352
rect 8763 7294 8805 7332
rect 8855 7352 8899 7394
rect 8855 7332 8867 7352
rect 8887 7332 8899 7352
rect 8855 7294 8899 7332
rect 8976 7352 9018 7394
rect 8976 7332 8984 7352
rect 9004 7332 9018 7352
rect 8976 7294 9018 7332
rect 9068 7352 9112 7394
rect 9068 7332 9080 7352
rect 9100 7332 9112 7352
rect 9068 7294 9112 7332
rect 1365 7251 1409 7289
rect 1365 7231 1377 7251
rect 1397 7231 1409 7251
rect 1365 7189 1409 7231
rect 1459 7251 1501 7289
rect 1459 7231 1473 7251
rect 1493 7231 1501 7251
rect 1459 7189 1501 7231
rect 1578 7251 1622 7289
rect 1578 7231 1590 7251
rect 1610 7231 1622 7251
rect 1578 7189 1622 7231
rect 1672 7251 1714 7289
rect 1672 7231 1686 7251
rect 1706 7231 1714 7251
rect 1672 7189 1714 7231
rect 1786 7251 1830 7289
rect 1786 7231 1798 7251
rect 1818 7231 1830 7251
rect 1786 7189 1830 7231
rect 1880 7251 1922 7289
rect 1880 7231 1894 7251
rect 1914 7231 1922 7251
rect 1880 7189 1922 7231
rect 1996 7251 2038 7289
rect 1996 7231 2004 7251
rect 2024 7231 2038 7251
rect 1996 7189 2038 7231
rect 2088 7258 2133 7289
rect 2088 7251 2132 7258
rect 2088 7231 2100 7251
rect 2120 7231 2132 7251
rect 2088 7189 2132 7231
rect 6646 7230 6690 7268
rect 6646 7210 6658 7230
rect 6678 7210 6690 7230
rect 6646 7168 6690 7210
rect 6740 7230 6782 7268
rect 6740 7210 6754 7230
rect 6774 7210 6782 7230
rect 6740 7168 6782 7210
rect 6859 7230 6903 7268
rect 6859 7210 6871 7230
rect 6891 7210 6903 7230
rect 6859 7168 6903 7210
rect 6953 7230 6995 7268
rect 6953 7210 6967 7230
rect 6987 7210 6995 7230
rect 6953 7168 6995 7210
rect 7067 7230 7111 7268
rect 7067 7210 7079 7230
rect 7099 7210 7111 7230
rect 7067 7168 7111 7210
rect 7161 7230 7203 7268
rect 7161 7210 7175 7230
rect 7195 7210 7203 7230
rect 7161 7168 7203 7210
rect 7277 7230 7319 7268
rect 7277 7210 7285 7230
rect 7305 7210 7319 7230
rect 7277 7168 7319 7210
rect 7369 7237 7414 7268
rect 7369 7230 7413 7237
rect 7369 7210 7381 7230
rect 7401 7210 7413 7230
rect 7369 7168 7413 7210
rect 303 7012 347 7050
rect 303 6992 315 7012
rect 335 6992 347 7012
rect 303 6950 347 6992
rect 397 7012 439 7050
rect 397 6992 411 7012
rect 431 6992 439 7012
rect 397 6950 439 6992
rect 516 7012 560 7050
rect 516 6992 528 7012
rect 548 6992 560 7012
rect 516 6950 560 6992
rect 610 7012 652 7050
rect 610 6992 624 7012
rect 644 6992 652 7012
rect 610 6950 652 6992
rect 724 7012 768 7050
rect 724 6992 736 7012
rect 756 6992 768 7012
rect 724 6950 768 6992
rect 818 7012 860 7050
rect 818 6992 832 7012
rect 852 6992 860 7012
rect 818 6950 860 6992
rect 934 7012 976 7050
rect 934 6992 942 7012
rect 962 6992 976 7012
rect 934 6950 976 6992
rect 1026 7019 1071 7050
rect 4132 7046 4176 7088
rect 4132 7026 4144 7046
rect 4164 7026 4176 7046
rect 4132 7019 4176 7026
rect 1026 7012 1070 7019
rect 1026 6992 1038 7012
rect 1058 6992 1070 7012
rect 1026 6950 1070 6992
rect 4131 6988 4176 7019
rect 4226 7046 4268 7088
rect 4226 7026 4240 7046
rect 4260 7026 4268 7046
rect 4226 6988 4268 7026
rect 4342 7046 4384 7088
rect 4342 7026 4350 7046
rect 4370 7026 4384 7046
rect 4342 6988 4384 7026
rect 4434 7046 4478 7088
rect 4434 7026 4446 7046
rect 4466 7026 4478 7046
rect 4434 6988 4478 7026
rect 4550 7046 4592 7088
rect 4550 7026 4558 7046
rect 4578 7026 4592 7046
rect 4550 6988 4592 7026
rect 4642 7046 4686 7088
rect 4642 7026 4654 7046
rect 4674 7026 4686 7046
rect 4642 6988 4686 7026
rect 4763 7046 4805 7088
rect 4763 7026 4771 7046
rect 4791 7026 4805 7046
rect 4763 6988 4805 7026
rect 4855 7046 4899 7088
rect 4855 7026 4867 7046
rect 4887 7026 4899 7046
rect 4855 6988 4899 7026
rect 5584 6991 5628 7029
rect 5584 6971 5596 6991
rect 5616 6971 5628 6991
rect 1315 6831 1359 6869
rect 1315 6811 1327 6831
rect 1347 6811 1359 6831
rect 1315 6769 1359 6811
rect 1409 6831 1451 6869
rect 1409 6811 1423 6831
rect 1443 6811 1451 6831
rect 1409 6769 1451 6811
rect 1528 6831 1572 6869
rect 1528 6811 1540 6831
rect 1560 6811 1572 6831
rect 1528 6769 1572 6811
rect 1622 6831 1664 6869
rect 1622 6811 1636 6831
rect 1656 6811 1664 6831
rect 1622 6769 1664 6811
rect 1736 6831 1780 6869
rect 1736 6811 1748 6831
rect 1768 6811 1780 6831
rect 1736 6769 1780 6811
rect 1830 6831 1872 6869
rect 1830 6811 1844 6831
rect 1864 6811 1872 6831
rect 1830 6769 1872 6811
rect 1946 6831 1988 6869
rect 1946 6811 1954 6831
rect 1974 6811 1988 6831
rect 1946 6769 1988 6811
rect 2038 6838 2083 6869
rect 5584 6929 5628 6971
rect 5678 6991 5720 7029
rect 5678 6971 5692 6991
rect 5712 6971 5720 6991
rect 5678 6929 5720 6971
rect 5797 6991 5841 7029
rect 5797 6971 5809 6991
rect 5829 6971 5841 6991
rect 5797 6929 5841 6971
rect 5891 6991 5933 7029
rect 5891 6971 5905 6991
rect 5925 6971 5933 6991
rect 5891 6929 5933 6971
rect 6005 6991 6049 7029
rect 6005 6971 6017 6991
rect 6037 6971 6049 6991
rect 6005 6929 6049 6971
rect 6099 6991 6141 7029
rect 6099 6971 6113 6991
rect 6133 6971 6141 6991
rect 6099 6929 6141 6971
rect 6215 6991 6257 7029
rect 6215 6971 6223 6991
rect 6243 6971 6257 6991
rect 6215 6929 6257 6971
rect 6307 6998 6352 7029
rect 9413 7025 9457 7067
rect 9413 7005 9425 7025
rect 9445 7005 9457 7025
rect 9413 6998 9457 7005
rect 6307 6991 6351 6998
rect 6307 6971 6319 6991
rect 6339 6971 6351 6991
rect 6307 6929 6351 6971
rect 9412 6967 9457 6998
rect 9507 7025 9549 7067
rect 9507 7005 9521 7025
rect 9541 7005 9549 7025
rect 9507 6967 9549 7005
rect 9623 7025 9665 7067
rect 9623 7005 9631 7025
rect 9651 7005 9665 7025
rect 9623 6967 9665 7005
rect 9715 7025 9759 7067
rect 9715 7005 9727 7025
rect 9747 7005 9759 7025
rect 9715 6967 9759 7005
rect 9831 7025 9873 7067
rect 9831 7005 9839 7025
rect 9859 7005 9873 7025
rect 9831 6967 9873 7005
rect 9923 7025 9967 7067
rect 9923 7005 9935 7025
rect 9955 7005 9967 7025
rect 9923 6967 9967 7005
rect 10044 7025 10086 7067
rect 10044 7005 10052 7025
rect 10072 7005 10086 7025
rect 10044 6967 10086 7005
rect 10136 7025 10180 7067
rect 10136 7005 10148 7025
rect 10168 7005 10180 7025
rect 10136 6967 10180 7005
rect 2038 6831 2082 6838
rect 2038 6811 2050 6831
rect 2070 6811 2082 6831
rect 2038 6769 2082 6811
rect 3119 6812 3163 6854
rect 3119 6792 3131 6812
rect 3151 6792 3163 6812
rect 3119 6785 3163 6792
rect 3118 6754 3163 6785
rect 3213 6812 3255 6854
rect 3213 6792 3227 6812
rect 3247 6792 3255 6812
rect 3213 6754 3255 6792
rect 3329 6812 3371 6854
rect 3329 6792 3337 6812
rect 3357 6792 3371 6812
rect 3329 6754 3371 6792
rect 3421 6812 3465 6854
rect 3421 6792 3433 6812
rect 3453 6792 3465 6812
rect 3421 6754 3465 6792
rect 3537 6812 3579 6854
rect 3537 6792 3545 6812
rect 3565 6792 3579 6812
rect 3537 6754 3579 6792
rect 3629 6812 3673 6854
rect 3629 6792 3641 6812
rect 3661 6792 3673 6812
rect 3629 6754 3673 6792
rect 3750 6812 3792 6854
rect 3750 6792 3758 6812
rect 3778 6792 3792 6812
rect 3750 6754 3792 6792
rect 3842 6812 3886 6854
rect 3842 6792 3854 6812
rect 3874 6792 3886 6812
rect 6596 6810 6640 6848
rect 3842 6754 3886 6792
rect 6596 6790 6608 6810
rect 6628 6790 6640 6810
rect 6596 6748 6640 6790
rect 6690 6810 6732 6848
rect 6690 6790 6704 6810
rect 6724 6790 6732 6810
rect 6690 6748 6732 6790
rect 6809 6810 6853 6848
rect 6809 6790 6821 6810
rect 6841 6790 6853 6810
rect 6809 6748 6853 6790
rect 6903 6810 6945 6848
rect 6903 6790 6917 6810
rect 6937 6790 6945 6810
rect 6903 6748 6945 6790
rect 7017 6810 7061 6848
rect 7017 6790 7029 6810
rect 7049 6790 7061 6810
rect 7017 6748 7061 6790
rect 7111 6810 7153 6848
rect 7111 6790 7125 6810
rect 7145 6790 7153 6810
rect 7111 6748 7153 6790
rect 7227 6810 7269 6848
rect 7227 6790 7235 6810
rect 7255 6790 7269 6810
rect 7227 6748 7269 6790
rect 7319 6817 7364 6848
rect 7319 6810 7363 6817
rect 7319 6790 7331 6810
rect 7351 6790 7363 6810
rect 7319 6748 7363 6790
rect 8400 6791 8444 6833
rect 8400 6771 8412 6791
rect 8432 6771 8444 6791
rect 8400 6764 8444 6771
rect 302 6597 346 6635
rect 302 6577 314 6597
rect 334 6577 346 6597
rect 302 6535 346 6577
rect 396 6597 438 6635
rect 396 6577 410 6597
rect 430 6577 438 6597
rect 396 6535 438 6577
rect 515 6597 559 6635
rect 515 6577 527 6597
rect 547 6577 559 6597
rect 515 6535 559 6577
rect 609 6597 651 6635
rect 609 6577 623 6597
rect 643 6577 651 6597
rect 609 6535 651 6577
rect 723 6597 767 6635
rect 723 6577 735 6597
rect 755 6577 767 6597
rect 723 6535 767 6577
rect 817 6597 859 6635
rect 817 6577 831 6597
rect 851 6577 859 6597
rect 817 6535 859 6577
rect 933 6597 975 6635
rect 933 6577 941 6597
rect 961 6577 975 6597
rect 933 6535 975 6577
rect 1025 6604 1070 6635
rect 4131 6631 4175 6673
rect 4131 6611 4143 6631
rect 4163 6611 4175 6631
rect 4131 6604 4175 6611
rect 1025 6597 1069 6604
rect 1025 6577 1037 6597
rect 1057 6577 1069 6597
rect 1025 6535 1069 6577
rect 4130 6573 4175 6604
rect 4225 6631 4267 6673
rect 4225 6611 4239 6631
rect 4259 6611 4267 6631
rect 4225 6573 4267 6611
rect 4341 6631 4383 6673
rect 4341 6611 4349 6631
rect 4369 6611 4383 6631
rect 4341 6573 4383 6611
rect 4433 6631 4477 6673
rect 4433 6611 4445 6631
rect 4465 6611 4477 6631
rect 4433 6573 4477 6611
rect 4549 6631 4591 6673
rect 4549 6611 4557 6631
rect 4577 6611 4591 6631
rect 4549 6573 4591 6611
rect 4641 6631 4685 6673
rect 4641 6611 4653 6631
rect 4673 6611 4685 6631
rect 4641 6573 4685 6611
rect 4762 6631 4804 6673
rect 4762 6611 4770 6631
rect 4790 6611 4804 6631
rect 4762 6573 4804 6611
rect 4854 6631 4898 6673
rect 8399 6733 8444 6764
rect 8494 6791 8536 6833
rect 8494 6771 8508 6791
rect 8528 6771 8536 6791
rect 8494 6733 8536 6771
rect 8610 6791 8652 6833
rect 8610 6771 8618 6791
rect 8638 6771 8652 6791
rect 8610 6733 8652 6771
rect 8702 6791 8746 6833
rect 8702 6771 8714 6791
rect 8734 6771 8746 6791
rect 8702 6733 8746 6771
rect 8818 6791 8860 6833
rect 8818 6771 8826 6791
rect 8846 6771 8860 6791
rect 8818 6733 8860 6771
rect 8910 6791 8954 6833
rect 8910 6771 8922 6791
rect 8942 6771 8954 6791
rect 8910 6733 8954 6771
rect 9031 6791 9073 6833
rect 9031 6771 9039 6791
rect 9059 6771 9073 6791
rect 9031 6733 9073 6771
rect 9123 6791 9167 6833
rect 9123 6771 9135 6791
rect 9155 6771 9167 6791
rect 9123 6733 9167 6771
rect 4854 6611 4866 6631
rect 4886 6611 4898 6631
rect 4854 6573 4898 6611
rect 5583 6576 5627 6614
rect 5583 6556 5595 6576
rect 5615 6556 5627 6576
rect 5583 6514 5627 6556
rect 5677 6576 5719 6614
rect 5677 6556 5691 6576
rect 5711 6556 5719 6576
rect 5677 6514 5719 6556
rect 5796 6576 5840 6614
rect 5796 6556 5808 6576
rect 5828 6556 5840 6576
rect 5796 6514 5840 6556
rect 5890 6576 5932 6614
rect 5890 6556 5904 6576
rect 5924 6556 5932 6576
rect 5890 6514 5932 6556
rect 6004 6576 6048 6614
rect 6004 6556 6016 6576
rect 6036 6556 6048 6576
rect 6004 6514 6048 6556
rect 6098 6576 6140 6614
rect 6098 6556 6112 6576
rect 6132 6556 6140 6576
rect 6098 6514 6140 6556
rect 6214 6576 6256 6614
rect 6214 6556 6222 6576
rect 6242 6556 6256 6576
rect 6214 6514 6256 6556
rect 6306 6583 6351 6614
rect 9412 6610 9456 6652
rect 9412 6590 9424 6610
rect 9444 6590 9456 6610
rect 9412 6583 9456 6590
rect 6306 6576 6350 6583
rect 6306 6556 6318 6576
rect 6338 6556 6350 6576
rect 6306 6514 6350 6556
rect 9411 6552 9456 6583
rect 9506 6610 9548 6652
rect 9506 6590 9520 6610
rect 9540 6590 9548 6610
rect 9506 6552 9548 6590
rect 9622 6610 9664 6652
rect 9622 6590 9630 6610
rect 9650 6590 9664 6610
rect 9622 6552 9664 6590
rect 9714 6610 9758 6652
rect 9714 6590 9726 6610
rect 9746 6590 9758 6610
rect 9714 6552 9758 6590
rect 9830 6610 9872 6652
rect 9830 6590 9838 6610
rect 9858 6590 9872 6610
rect 9830 6552 9872 6590
rect 9922 6610 9966 6652
rect 9922 6590 9934 6610
rect 9954 6590 9966 6610
rect 9922 6552 9966 6590
rect 10043 6610 10085 6652
rect 10043 6590 10051 6610
rect 10071 6590 10085 6610
rect 10043 6552 10085 6590
rect 10135 6610 10179 6652
rect 10135 6590 10147 6610
rect 10167 6590 10179 6610
rect 10135 6552 10179 6590
rect 1530 6319 1574 6357
rect 1530 6299 1542 6319
rect 1562 6299 1574 6319
rect 1530 6257 1574 6299
rect 1624 6319 1666 6357
rect 1624 6299 1638 6319
rect 1658 6299 1666 6319
rect 1624 6257 1666 6299
rect 1743 6319 1787 6357
rect 1743 6299 1755 6319
rect 1775 6299 1787 6319
rect 1743 6257 1787 6299
rect 1837 6319 1879 6357
rect 1837 6299 1851 6319
rect 1871 6299 1879 6319
rect 1837 6257 1879 6299
rect 1951 6319 1995 6357
rect 1951 6299 1963 6319
rect 1983 6299 1995 6319
rect 1951 6257 1995 6299
rect 2045 6319 2087 6357
rect 2045 6299 2059 6319
rect 2079 6299 2087 6319
rect 2045 6257 2087 6299
rect 2161 6319 2203 6357
rect 2161 6299 2169 6319
rect 2189 6299 2203 6319
rect 2161 6257 2203 6299
rect 2253 6326 2298 6357
rect 2911 6345 2955 6387
rect 2253 6319 2297 6326
rect 2253 6299 2265 6319
rect 2285 6299 2297 6319
rect 2911 6325 2923 6345
rect 2943 6325 2955 6345
rect 2911 6318 2955 6325
rect 2253 6257 2297 6299
rect 2910 6287 2955 6318
rect 3005 6345 3047 6387
rect 3005 6325 3019 6345
rect 3039 6325 3047 6345
rect 3005 6287 3047 6325
rect 3121 6345 3163 6387
rect 3121 6325 3129 6345
rect 3149 6325 3163 6345
rect 3121 6287 3163 6325
rect 3213 6345 3257 6387
rect 3213 6325 3225 6345
rect 3245 6325 3257 6345
rect 3213 6287 3257 6325
rect 3329 6345 3371 6387
rect 3329 6325 3337 6345
rect 3357 6325 3371 6345
rect 3329 6287 3371 6325
rect 3421 6345 3465 6387
rect 3421 6325 3433 6345
rect 3453 6325 3465 6345
rect 3421 6287 3465 6325
rect 3542 6345 3584 6387
rect 3542 6325 3550 6345
rect 3570 6325 3584 6345
rect 3542 6287 3584 6325
rect 3634 6345 3678 6387
rect 3634 6325 3646 6345
rect 3666 6325 3678 6345
rect 3634 6287 3678 6325
rect 6811 6298 6855 6336
rect 6811 6278 6823 6298
rect 6843 6278 6855 6298
rect 6811 6236 6855 6278
rect 6905 6298 6947 6336
rect 6905 6278 6919 6298
rect 6939 6278 6947 6298
rect 6905 6236 6947 6278
rect 7024 6298 7068 6336
rect 7024 6278 7036 6298
rect 7056 6278 7068 6298
rect 7024 6236 7068 6278
rect 7118 6298 7160 6336
rect 7118 6278 7132 6298
rect 7152 6278 7160 6298
rect 7118 6236 7160 6278
rect 7232 6298 7276 6336
rect 7232 6278 7244 6298
rect 7264 6278 7276 6298
rect 7232 6236 7276 6278
rect 7326 6298 7368 6336
rect 7326 6278 7340 6298
rect 7360 6278 7368 6298
rect 7326 6236 7368 6278
rect 7442 6298 7484 6336
rect 7442 6278 7450 6298
rect 7470 6278 7484 6298
rect 7442 6236 7484 6278
rect 7534 6305 7579 6336
rect 8192 6324 8236 6366
rect 7534 6298 7578 6305
rect 7534 6278 7546 6298
rect 7566 6278 7578 6298
rect 8192 6304 8204 6324
rect 8224 6304 8236 6324
rect 8192 6297 8236 6304
rect 7534 6236 7578 6278
rect 8191 6266 8236 6297
rect 8286 6324 8328 6366
rect 8286 6304 8300 6324
rect 8320 6304 8328 6324
rect 8286 6266 8328 6304
rect 8402 6324 8444 6366
rect 8402 6304 8410 6324
rect 8430 6304 8444 6324
rect 8402 6266 8444 6304
rect 8494 6324 8538 6366
rect 8494 6304 8506 6324
rect 8526 6304 8538 6324
rect 8494 6266 8538 6304
rect 8610 6324 8652 6366
rect 8610 6304 8618 6324
rect 8638 6304 8652 6324
rect 8610 6266 8652 6304
rect 8702 6324 8746 6366
rect 8702 6304 8714 6324
rect 8734 6304 8746 6324
rect 8702 6266 8746 6304
rect 8823 6324 8865 6366
rect 8823 6304 8831 6324
rect 8851 6304 8865 6324
rect 8823 6266 8865 6304
rect 8915 6324 8959 6366
rect 8915 6304 8927 6324
rect 8947 6304 8959 6324
rect 8915 6266 8959 6304
rect 310 6033 354 6071
rect 310 6013 322 6033
rect 342 6013 354 6033
rect 310 5971 354 6013
rect 404 6033 446 6071
rect 404 6013 418 6033
rect 438 6013 446 6033
rect 404 5971 446 6013
rect 523 6033 567 6071
rect 523 6013 535 6033
rect 555 6013 567 6033
rect 523 5971 567 6013
rect 617 6033 659 6071
rect 617 6013 631 6033
rect 651 6013 659 6033
rect 617 5971 659 6013
rect 731 6033 775 6071
rect 731 6013 743 6033
rect 763 6013 775 6033
rect 731 5971 775 6013
rect 825 6033 867 6071
rect 825 6013 839 6033
rect 859 6013 867 6033
rect 825 5971 867 6013
rect 941 6033 983 6071
rect 941 6013 949 6033
rect 969 6013 983 6033
rect 941 5971 983 6013
rect 1033 6040 1078 6071
rect 4139 6067 4183 6109
rect 4139 6047 4151 6067
rect 4171 6047 4183 6067
rect 4139 6040 4183 6047
rect 1033 6033 1077 6040
rect 1033 6013 1045 6033
rect 1065 6013 1077 6033
rect 1033 5971 1077 6013
rect 4138 6009 4183 6040
rect 4233 6067 4275 6109
rect 4233 6047 4247 6067
rect 4267 6047 4275 6067
rect 4233 6009 4275 6047
rect 4349 6067 4391 6109
rect 4349 6047 4357 6067
rect 4377 6047 4391 6067
rect 4349 6009 4391 6047
rect 4441 6067 4485 6109
rect 4441 6047 4453 6067
rect 4473 6047 4485 6067
rect 4441 6009 4485 6047
rect 4557 6067 4599 6109
rect 4557 6047 4565 6067
rect 4585 6047 4599 6067
rect 4557 6009 4599 6047
rect 4649 6067 4693 6109
rect 4649 6047 4661 6067
rect 4681 6047 4693 6067
rect 4649 6009 4693 6047
rect 4770 6067 4812 6109
rect 4770 6047 4778 6067
rect 4798 6047 4812 6067
rect 4770 6009 4812 6047
rect 4862 6067 4906 6109
rect 4862 6047 4874 6067
rect 4894 6047 4906 6067
rect 4862 6009 4906 6047
rect 5591 6012 5635 6050
rect 5591 5992 5603 6012
rect 5623 5992 5635 6012
rect 1322 5852 1366 5890
rect 1322 5832 1334 5852
rect 1354 5832 1366 5852
rect 1322 5790 1366 5832
rect 1416 5852 1458 5890
rect 1416 5832 1430 5852
rect 1450 5832 1458 5852
rect 1416 5790 1458 5832
rect 1535 5852 1579 5890
rect 1535 5832 1547 5852
rect 1567 5832 1579 5852
rect 1535 5790 1579 5832
rect 1629 5852 1671 5890
rect 1629 5832 1643 5852
rect 1663 5832 1671 5852
rect 1629 5790 1671 5832
rect 1743 5852 1787 5890
rect 1743 5832 1755 5852
rect 1775 5832 1787 5852
rect 1743 5790 1787 5832
rect 1837 5852 1879 5890
rect 1837 5832 1851 5852
rect 1871 5832 1879 5852
rect 1837 5790 1879 5832
rect 1953 5852 1995 5890
rect 1953 5832 1961 5852
rect 1981 5832 1995 5852
rect 1953 5790 1995 5832
rect 2045 5859 2090 5890
rect 5591 5950 5635 5992
rect 5685 6012 5727 6050
rect 5685 5992 5699 6012
rect 5719 5992 5727 6012
rect 5685 5950 5727 5992
rect 5804 6012 5848 6050
rect 5804 5992 5816 6012
rect 5836 5992 5848 6012
rect 5804 5950 5848 5992
rect 5898 6012 5940 6050
rect 5898 5992 5912 6012
rect 5932 5992 5940 6012
rect 5898 5950 5940 5992
rect 6012 6012 6056 6050
rect 6012 5992 6024 6012
rect 6044 5992 6056 6012
rect 6012 5950 6056 5992
rect 6106 6012 6148 6050
rect 6106 5992 6120 6012
rect 6140 5992 6148 6012
rect 6106 5950 6148 5992
rect 6222 6012 6264 6050
rect 6222 5992 6230 6012
rect 6250 5992 6264 6012
rect 6222 5950 6264 5992
rect 6314 6019 6359 6050
rect 9420 6046 9464 6088
rect 9420 6026 9432 6046
rect 9452 6026 9464 6046
rect 9420 6019 9464 6026
rect 6314 6012 6358 6019
rect 6314 5992 6326 6012
rect 6346 5992 6358 6012
rect 6314 5950 6358 5992
rect 9419 5988 9464 6019
rect 9514 6046 9556 6088
rect 9514 6026 9528 6046
rect 9548 6026 9556 6046
rect 9514 5988 9556 6026
rect 9630 6046 9672 6088
rect 9630 6026 9638 6046
rect 9658 6026 9672 6046
rect 9630 5988 9672 6026
rect 9722 6046 9766 6088
rect 9722 6026 9734 6046
rect 9754 6026 9766 6046
rect 9722 5988 9766 6026
rect 9838 6046 9880 6088
rect 9838 6026 9846 6046
rect 9866 6026 9880 6046
rect 9838 5988 9880 6026
rect 9930 6046 9974 6088
rect 9930 6026 9942 6046
rect 9962 6026 9974 6046
rect 9930 5988 9974 6026
rect 10051 6046 10093 6088
rect 10051 6026 10059 6046
rect 10079 6026 10093 6046
rect 10051 5988 10093 6026
rect 10143 6046 10187 6088
rect 10143 6026 10155 6046
rect 10175 6026 10187 6046
rect 10143 5988 10187 6026
rect 2045 5852 2089 5859
rect 2045 5832 2057 5852
rect 2077 5832 2089 5852
rect 2045 5790 2089 5832
rect 3126 5833 3170 5875
rect 3126 5813 3138 5833
rect 3158 5813 3170 5833
rect 3126 5806 3170 5813
rect 3125 5775 3170 5806
rect 3220 5833 3262 5875
rect 3220 5813 3234 5833
rect 3254 5813 3262 5833
rect 3220 5775 3262 5813
rect 3336 5833 3378 5875
rect 3336 5813 3344 5833
rect 3364 5813 3378 5833
rect 3336 5775 3378 5813
rect 3428 5833 3472 5875
rect 3428 5813 3440 5833
rect 3460 5813 3472 5833
rect 3428 5775 3472 5813
rect 3544 5833 3586 5875
rect 3544 5813 3552 5833
rect 3572 5813 3586 5833
rect 3544 5775 3586 5813
rect 3636 5833 3680 5875
rect 3636 5813 3648 5833
rect 3668 5813 3680 5833
rect 3636 5775 3680 5813
rect 3757 5833 3799 5875
rect 3757 5813 3765 5833
rect 3785 5813 3799 5833
rect 3757 5775 3799 5813
rect 3849 5833 3893 5875
rect 3849 5813 3861 5833
rect 3881 5813 3893 5833
rect 6603 5831 6647 5869
rect 3849 5775 3893 5813
rect 6603 5811 6615 5831
rect 6635 5811 6647 5831
rect 6603 5769 6647 5811
rect 6697 5831 6739 5869
rect 6697 5811 6711 5831
rect 6731 5811 6739 5831
rect 6697 5769 6739 5811
rect 6816 5831 6860 5869
rect 6816 5811 6828 5831
rect 6848 5811 6860 5831
rect 6816 5769 6860 5811
rect 6910 5831 6952 5869
rect 6910 5811 6924 5831
rect 6944 5811 6952 5831
rect 6910 5769 6952 5811
rect 7024 5831 7068 5869
rect 7024 5811 7036 5831
rect 7056 5811 7068 5831
rect 7024 5769 7068 5811
rect 7118 5831 7160 5869
rect 7118 5811 7132 5831
rect 7152 5811 7160 5831
rect 7118 5769 7160 5811
rect 7234 5831 7276 5869
rect 7234 5811 7242 5831
rect 7262 5811 7276 5831
rect 7234 5769 7276 5811
rect 7326 5838 7371 5869
rect 7326 5831 7370 5838
rect 7326 5811 7338 5831
rect 7358 5811 7370 5831
rect 7326 5769 7370 5811
rect 8407 5812 8451 5854
rect 8407 5792 8419 5812
rect 8439 5792 8451 5812
rect 8407 5785 8451 5792
rect 309 5618 353 5656
rect 309 5598 321 5618
rect 341 5598 353 5618
rect 309 5556 353 5598
rect 403 5618 445 5656
rect 403 5598 417 5618
rect 437 5598 445 5618
rect 403 5556 445 5598
rect 522 5618 566 5656
rect 522 5598 534 5618
rect 554 5598 566 5618
rect 522 5556 566 5598
rect 616 5618 658 5656
rect 616 5598 630 5618
rect 650 5598 658 5618
rect 616 5556 658 5598
rect 730 5618 774 5656
rect 730 5598 742 5618
rect 762 5598 774 5618
rect 730 5556 774 5598
rect 824 5618 866 5656
rect 824 5598 838 5618
rect 858 5598 866 5618
rect 824 5556 866 5598
rect 940 5618 982 5656
rect 940 5598 948 5618
rect 968 5598 982 5618
rect 940 5556 982 5598
rect 1032 5625 1077 5656
rect 4138 5652 4182 5694
rect 4138 5632 4150 5652
rect 4170 5632 4182 5652
rect 4138 5625 4182 5632
rect 1032 5618 1076 5625
rect 1032 5598 1044 5618
rect 1064 5598 1076 5618
rect 1032 5556 1076 5598
rect 4137 5594 4182 5625
rect 4232 5652 4274 5694
rect 4232 5632 4246 5652
rect 4266 5632 4274 5652
rect 4232 5594 4274 5632
rect 4348 5652 4390 5694
rect 4348 5632 4356 5652
rect 4376 5632 4390 5652
rect 4348 5594 4390 5632
rect 4440 5652 4484 5694
rect 4440 5632 4452 5652
rect 4472 5632 4484 5652
rect 4440 5594 4484 5632
rect 4556 5652 4598 5694
rect 4556 5632 4564 5652
rect 4584 5632 4598 5652
rect 4556 5594 4598 5632
rect 4648 5652 4692 5694
rect 4648 5632 4660 5652
rect 4680 5632 4692 5652
rect 4648 5594 4692 5632
rect 4769 5652 4811 5694
rect 4769 5632 4777 5652
rect 4797 5632 4811 5652
rect 4769 5594 4811 5632
rect 4861 5652 4905 5694
rect 8406 5754 8451 5785
rect 8501 5812 8543 5854
rect 8501 5792 8515 5812
rect 8535 5792 8543 5812
rect 8501 5754 8543 5792
rect 8617 5812 8659 5854
rect 8617 5792 8625 5812
rect 8645 5792 8659 5812
rect 8617 5754 8659 5792
rect 8709 5812 8753 5854
rect 8709 5792 8721 5812
rect 8741 5792 8753 5812
rect 8709 5754 8753 5792
rect 8825 5812 8867 5854
rect 8825 5792 8833 5812
rect 8853 5792 8867 5812
rect 8825 5754 8867 5792
rect 8917 5812 8961 5854
rect 8917 5792 8929 5812
rect 8949 5792 8961 5812
rect 8917 5754 8961 5792
rect 9038 5812 9080 5854
rect 9038 5792 9046 5812
rect 9066 5792 9080 5812
rect 9038 5754 9080 5792
rect 9130 5812 9174 5854
rect 9130 5792 9142 5812
rect 9162 5792 9174 5812
rect 9130 5754 9174 5792
rect 4861 5632 4873 5652
rect 4893 5632 4905 5652
rect 4861 5594 4905 5632
rect 5590 5597 5634 5635
rect 5590 5577 5602 5597
rect 5622 5577 5634 5597
rect 5590 5535 5634 5577
rect 5684 5597 5726 5635
rect 5684 5577 5698 5597
rect 5718 5577 5726 5597
rect 5684 5535 5726 5577
rect 5803 5597 5847 5635
rect 5803 5577 5815 5597
rect 5835 5577 5847 5597
rect 5803 5535 5847 5577
rect 5897 5597 5939 5635
rect 5897 5577 5911 5597
rect 5931 5577 5939 5597
rect 5897 5535 5939 5577
rect 6011 5597 6055 5635
rect 6011 5577 6023 5597
rect 6043 5577 6055 5597
rect 6011 5535 6055 5577
rect 6105 5597 6147 5635
rect 6105 5577 6119 5597
rect 6139 5577 6147 5597
rect 6105 5535 6147 5577
rect 6221 5597 6263 5635
rect 6221 5577 6229 5597
rect 6249 5577 6263 5597
rect 6221 5535 6263 5577
rect 6313 5604 6358 5635
rect 9419 5631 9463 5673
rect 9419 5611 9431 5631
rect 9451 5611 9463 5631
rect 9419 5604 9463 5611
rect 6313 5597 6357 5604
rect 6313 5577 6325 5597
rect 6345 5577 6357 5597
rect 6313 5535 6357 5577
rect 9418 5573 9463 5604
rect 9513 5631 9555 5673
rect 9513 5611 9527 5631
rect 9547 5611 9555 5631
rect 9513 5573 9555 5611
rect 9629 5631 9671 5673
rect 9629 5611 9637 5631
rect 9657 5611 9671 5631
rect 9629 5573 9671 5611
rect 9721 5631 9765 5673
rect 9721 5611 9733 5631
rect 9753 5611 9765 5631
rect 9721 5573 9765 5611
rect 9837 5631 9879 5673
rect 9837 5611 9845 5631
rect 9865 5611 9879 5631
rect 9837 5573 9879 5611
rect 9929 5631 9973 5673
rect 9929 5611 9941 5631
rect 9961 5611 9973 5631
rect 9929 5573 9973 5611
rect 10050 5631 10092 5673
rect 10050 5611 10058 5631
rect 10078 5611 10092 5631
rect 10050 5573 10092 5611
rect 10142 5631 10186 5673
rect 10142 5611 10154 5631
rect 10174 5611 10186 5631
rect 10142 5573 10186 5611
rect 3076 5413 3120 5455
rect 3076 5393 3088 5413
rect 3108 5393 3120 5413
rect 3076 5386 3120 5393
rect 3075 5355 3120 5386
rect 3170 5413 3212 5455
rect 3170 5393 3184 5413
rect 3204 5393 3212 5413
rect 3170 5355 3212 5393
rect 3286 5413 3328 5455
rect 3286 5393 3294 5413
rect 3314 5393 3328 5413
rect 3286 5355 3328 5393
rect 3378 5413 3422 5455
rect 3378 5393 3390 5413
rect 3410 5393 3422 5413
rect 3378 5355 3422 5393
rect 3494 5413 3536 5455
rect 3494 5393 3502 5413
rect 3522 5393 3536 5413
rect 3494 5355 3536 5393
rect 3586 5413 3630 5455
rect 3586 5393 3598 5413
rect 3618 5393 3630 5413
rect 3586 5355 3630 5393
rect 3707 5413 3749 5455
rect 3707 5393 3715 5413
rect 3735 5393 3749 5413
rect 3707 5355 3749 5393
rect 3799 5413 3843 5455
rect 3799 5393 3811 5413
rect 3831 5393 3843 5413
rect 3799 5355 3843 5393
rect 8357 5392 8401 5434
rect 8357 5372 8369 5392
rect 8389 5372 8401 5392
rect 8357 5365 8401 5372
rect 8356 5334 8401 5365
rect 8451 5392 8493 5434
rect 8451 5372 8465 5392
rect 8485 5372 8493 5392
rect 8451 5334 8493 5372
rect 8567 5392 8609 5434
rect 8567 5372 8575 5392
rect 8595 5372 8609 5392
rect 8567 5334 8609 5372
rect 8659 5392 8703 5434
rect 8659 5372 8671 5392
rect 8691 5372 8703 5392
rect 8659 5334 8703 5372
rect 8775 5392 8817 5434
rect 8775 5372 8783 5392
rect 8803 5372 8817 5392
rect 8775 5334 8817 5372
rect 8867 5392 8911 5434
rect 8867 5372 8879 5392
rect 8899 5372 8911 5392
rect 8867 5334 8911 5372
rect 8988 5392 9030 5434
rect 8988 5372 8996 5392
rect 9016 5372 9030 5392
rect 8988 5334 9030 5372
rect 9080 5392 9124 5434
rect 9080 5372 9092 5392
rect 9112 5372 9124 5392
rect 9080 5334 9124 5372
rect 1377 5291 1421 5329
rect 1377 5271 1389 5291
rect 1409 5271 1421 5291
rect 1377 5229 1421 5271
rect 1471 5291 1513 5329
rect 1471 5271 1485 5291
rect 1505 5271 1513 5291
rect 1471 5229 1513 5271
rect 1590 5291 1634 5329
rect 1590 5271 1602 5291
rect 1622 5271 1634 5291
rect 1590 5229 1634 5271
rect 1684 5291 1726 5329
rect 1684 5271 1698 5291
rect 1718 5271 1726 5291
rect 1684 5229 1726 5271
rect 1798 5291 1842 5329
rect 1798 5271 1810 5291
rect 1830 5271 1842 5291
rect 1798 5229 1842 5271
rect 1892 5291 1934 5329
rect 1892 5271 1906 5291
rect 1926 5271 1934 5291
rect 1892 5229 1934 5271
rect 2008 5291 2050 5329
rect 2008 5271 2016 5291
rect 2036 5271 2050 5291
rect 2008 5229 2050 5271
rect 2100 5298 2145 5329
rect 2100 5291 2144 5298
rect 2100 5271 2112 5291
rect 2132 5271 2144 5291
rect 2100 5229 2144 5271
rect 6658 5270 6702 5308
rect 6658 5250 6670 5270
rect 6690 5250 6702 5270
rect 6658 5208 6702 5250
rect 6752 5270 6794 5308
rect 6752 5250 6766 5270
rect 6786 5250 6794 5270
rect 6752 5208 6794 5250
rect 6871 5270 6915 5308
rect 6871 5250 6883 5270
rect 6903 5250 6915 5270
rect 6871 5208 6915 5250
rect 6965 5270 7007 5308
rect 6965 5250 6979 5270
rect 6999 5250 7007 5270
rect 6965 5208 7007 5250
rect 7079 5270 7123 5308
rect 7079 5250 7091 5270
rect 7111 5250 7123 5270
rect 7079 5208 7123 5250
rect 7173 5270 7215 5308
rect 7173 5250 7187 5270
rect 7207 5250 7215 5270
rect 7173 5208 7215 5250
rect 7289 5270 7331 5308
rect 7289 5250 7297 5270
rect 7317 5250 7331 5270
rect 7289 5208 7331 5250
rect 7381 5277 7426 5308
rect 7381 5270 7425 5277
rect 7381 5250 7393 5270
rect 7413 5250 7425 5270
rect 7381 5208 7425 5250
rect 315 5052 359 5090
rect 315 5032 327 5052
rect 347 5032 359 5052
rect 315 4990 359 5032
rect 409 5052 451 5090
rect 409 5032 423 5052
rect 443 5032 451 5052
rect 409 4990 451 5032
rect 528 5052 572 5090
rect 528 5032 540 5052
rect 560 5032 572 5052
rect 528 4990 572 5032
rect 622 5052 664 5090
rect 622 5032 636 5052
rect 656 5032 664 5052
rect 622 4990 664 5032
rect 736 5052 780 5090
rect 736 5032 748 5052
rect 768 5032 780 5052
rect 736 4990 780 5032
rect 830 5052 872 5090
rect 830 5032 844 5052
rect 864 5032 872 5052
rect 830 4990 872 5032
rect 946 5052 988 5090
rect 946 5032 954 5052
rect 974 5032 988 5052
rect 946 4990 988 5032
rect 1038 5059 1083 5090
rect 4144 5086 4188 5128
rect 4144 5066 4156 5086
rect 4176 5066 4188 5086
rect 4144 5059 4188 5066
rect 1038 5052 1082 5059
rect 1038 5032 1050 5052
rect 1070 5032 1082 5052
rect 1038 4990 1082 5032
rect 4143 5028 4188 5059
rect 4238 5086 4280 5128
rect 4238 5066 4252 5086
rect 4272 5066 4280 5086
rect 4238 5028 4280 5066
rect 4354 5086 4396 5128
rect 4354 5066 4362 5086
rect 4382 5066 4396 5086
rect 4354 5028 4396 5066
rect 4446 5086 4490 5128
rect 4446 5066 4458 5086
rect 4478 5066 4490 5086
rect 4446 5028 4490 5066
rect 4562 5086 4604 5128
rect 4562 5066 4570 5086
rect 4590 5066 4604 5086
rect 4562 5028 4604 5066
rect 4654 5086 4698 5128
rect 4654 5066 4666 5086
rect 4686 5066 4698 5086
rect 4654 5028 4698 5066
rect 4775 5086 4817 5128
rect 4775 5066 4783 5086
rect 4803 5066 4817 5086
rect 4775 5028 4817 5066
rect 4867 5086 4911 5128
rect 4867 5066 4879 5086
rect 4899 5066 4911 5086
rect 4867 5028 4911 5066
rect 5596 5031 5640 5069
rect 5596 5011 5608 5031
rect 5628 5011 5640 5031
rect 1327 4871 1371 4909
rect 1327 4851 1339 4871
rect 1359 4851 1371 4871
rect 1327 4809 1371 4851
rect 1421 4871 1463 4909
rect 1421 4851 1435 4871
rect 1455 4851 1463 4871
rect 1421 4809 1463 4851
rect 1540 4871 1584 4909
rect 1540 4851 1552 4871
rect 1572 4851 1584 4871
rect 1540 4809 1584 4851
rect 1634 4871 1676 4909
rect 1634 4851 1648 4871
rect 1668 4851 1676 4871
rect 1634 4809 1676 4851
rect 1748 4871 1792 4909
rect 1748 4851 1760 4871
rect 1780 4851 1792 4871
rect 1748 4809 1792 4851
rect 1842 4871 1884 4909
rect 1842 4851 1856 4871
rect 1876 4851 1884 4871
rect 1842 4809 1884 4851
rect 1958 4871 2000 4909
rect 1958 4851 1966 4871
rect 1986 4851 2000 4871
rect 1958 4809 2000 4851
rect 2050 4878 2095 4909
rect 5596 4969 5640 5011
rect 5690 5031 5732 5069
rect 5690 5011 5704 5031
rect 5724 5011 5732 5031
rect 5690 4969 5732 5011
rect 5809 5031 5853 5069
rect 5809 5011 5821 5031
rect 5841 5011 5853 5031
rect 5809 4969 5853 5011
rect 5903 5031 5945 5069
rect 5903 5011 5917 5031
rect 5937 5011 5945 5031
rect 5903 4969 5945 5011
rect 6017 5031 6061 5069
rect 6017 5011 6029 5031
rect 6049 5011 6061 5031
rect 6017 4969 6061 5011
rect 6111 5031 6153 5069
rect 6111 5011 6125 5031
rect 6145 5011 6153 5031
rect 6111 4969 6153 5011
rect 6227 5031 6269 5069
rect 6227 5011 6235 5031
rect 6255 5011 6269 5031
rect 6227 4969 6269 5011
rect 6319 5038 6364 5069
rect 9425 5065 9469 5107
rect 9425 5045 9437 5065
rect 9457 5045 9469 5065
rect 9425 5038 9469 5045
rect 6319 5031 6363 5038
rect 6319 5011 6331 5031
rect 6351 5011 6363 5031
rect 6319 4969 6363 5011
rect 9424 5007 9469 5038
rect 9519 5065 9561 5107
rect 9519 5045 9533 5065
rect 9553 5045 9561 5065
rect 9519 5007 9561 5045
rect 9635 5065 9677 5107
rect 9635 5045 9643 5065
rect 9663 5045 9677 5065
rect 9635 5007 9677 5045
rect 9727 5065 9771 5107
rect 9727 5045 9739 5065
rect 9759 5045 9771 5065
rect 9727 5007 9771 5045
rect 9843 5065 9885 5107
rect 9843 5045 9851 5065
rect 9871 5045 9885 5065
rect 9843 5007 9885 5045
rect 9935 5065 9979 5107
rect 9935 5045 9947 5065
rect 9967 5045 9979 5065
rect 9935 5007 9979 5045
rect 10056 5065 10098 5107
rect 10056 5045 10064 5065
rect 10084 5045 10098 5065
rect 10056 5007 10098 5045
rect 10148 5065 10192 5107
rect 10148 5045 10160 5065
rect 10180 5045 10192 5065
rect 10148 5007 10192 5045
rect 2050 4871 2094 4878
rect 2050 4851 2062 4871
rect 2082 4851 2094 4871
rect 2050 4809 2094 4851
rect 3131 4852 3175 4894
rect 3131 4832 3143 4852
rect 3163 4832 3175 4852
rect 3131 4825 3175 4832
rect 3130 4794 3175 4825
rect 3225 4852 3267 4894
rect 3225 4832 3239 4852
rect 3259 4832 3267 4852
rect 3225 4794 3267 4832
rect 3341 4852 3383 4894
rect 3341 4832 3349 4852
rect 3369 4832 3383 4852
rect 3341 4794 3383 4832
rect 3433 4852 3477 4894
rect 3433 4832 3445 4852
rect 3465 4832 3477 4852
rect 3433 4794 3477 4832
rect 3549 4852 3591 4894
rect 3549 4832 3557 4852
rect 3577 4832 3591 4852
rect 3549 4794 3591 4832
rect 3641 4852 3685 4894
rect 3641 4832 3653 4852
rect 3673 4832 3685 4852
rect 3641 4794 3685 4832
rect 3762 4852 3804 4894
rect 3762 4832 3770 4852
rect 3790 4832 3804 4852
rect 3762 4794 3804 4832
rect 3854 4852 3898 4894
rect 3854 4832 3866 4852
rect 3886 4832 3898 4852
rect 6608 4850 6652 4888
rect 3854 4794 3898 4832
rect 6608 4830 6620 4850
rect 6640 4830 6652 4850
rect 6608 4788 6652 4830
rect 6702 4850 6744 4888
rect 6702 4830 6716 4850
rect 6736 4830 6744 4850
rect 6702 4788 6744 4830
rect 6821 4850 6865 4888
rect 6821 4830 6833 4850
rect 6853 4830 6865 4850
rect 6821 4788 6865 4830
rect 6915 4850 6957 4888
rect 6915 4830 6929 4850
rect 6949 4830 6957 4850
rect 6915 4788 6957 4830
rect 7029 4850 7073 4888
rect 7029 4830 7041 4850
rect 7061 4830 7073 4850
rect 7029 4788 7073 4830
rect 7123 4850 7165 4888
rect 7123 4830 7137 4850
rect 7157 4830 7165 4850
rect 7123 4788 7165 4830
rect 7239 4850 7281 4888
rect 7239 4830 7247 4850
rect 7267 4830 7281 4850
rect 7239 4788 7281 4830
rect 7331 4857 7376 4888
rect 7331 4850 7375 4857
rect 7331 4830 7343 4850
rect 7363 4830 7375 4850
rect 7331 4788 7375 4830
rect 8412 4831 8456 4873
rect 8412 4811 8424 4831
rect 8444 4811 8456 4831
rect 8412 4804 8456 4811
rect 314 4637 358 4675
rect 314 4617 326 4637
rect 346 4617 358 4637
rect 314 4575 358 4617
rect 408 4637 450 4675
rect 408 4617 422 4637
rect 442 4617 450 4637
rect 408 4575 450 4617
rect 527 4637 571 4675
rect 527 4617 539 4637
rect 559 4617 571 4637
rect 527 4575 571 4617
rect 621 4637 663 4675
rect 621 4617 635 4637
rect 655 4617 663 4637
rect 621 4575 663 4617
rect 735 4637 779 4675
rect 735 4617 747 4637
rect 767 4617 779 4637
rect 735 4575 779 4617
rect 829 4637 871 4675
rect 829 4617 843 4637
rect 863 4617 871 4637
rect 829 4575 871 4617
rect 945 4637 987 4675
rect 945 4617 953 4637
rect 973 4617 987 4637
rect 945 4575 987 4617
rect 1037 4644 1082 4675
rect 4143 4671 4187 4713
rect 4143 4651 4155 4671
rect 4175 4651 4187 4671
rect 4143 4644 4187 4651
rect 1037 4637 1081 4644
rect 1037 4617 1049 4637
rect 1069 4617 1081 4637
rect 1037 4575 1081 4617
rect 4142 4613 4187 4644
rect 4237 4671 4279 4713
rect 4237 4651 4251 4671
rect 4271 4651 4279 4671
rect 4237 4613 4279 4651
rect 4353 4671 4395 4713
rect 4353 4651 4361 4671
rect 4381 4651 4395 4671
rect 4353 4613 4395 4651
rect 4445 4671 4489 4713
rect 4445 4651 4457 4671
rect 4477 4651 4489 4671
rect 4445 4613 4489 4651
rect 4561 4671 4603 4713
rect 4561 4651 4569 4671
rect 4589 4651 4603 4671
rect 4561 4613 4603 4651
rect 4653 4671 4697 4713
rect 4653 4651 4665 4671
rect 4685 4651 4697 4671
rect 4653 4613 4697 4651
rect 4774 4671 4816 4713
rect 4774 4651 4782 4671
rect 4802 4651 4816 4671
rect 4774 4613 4816 4651
rect 4866 4671 4910 4713
rect 8411 4773 8456 4804
rect 8506 4831 8548 4873
rect 8506 4811 8520 4831
rect 8540 4811 8548 4831
rect 8506 4773 8548 4811
rect 8622 4831 8664 4873
rect 8622 4811 8630 4831
rect 8650 4811 8664 4831
rect 8622 4773 8664 4811
rect 8714 4831 8758 4873
rect 8714 4811 8726 4831
rect 8746 4811 8758 4831
rect 8714 4773 8758 4811
rect 8830 4831 8872 4873
rect 8830 4811 8838 4831
rect 8858 4811 8872 4831
rect 8830 4773 8872 4811
rect 8922 4831 8966 4873
rect 8922 4811 8934 4831
rect 8954 4811 8966 4831
rect 8922 4773 8966 4811
rect 9043 4831 9085 4873
rect 9043 4811 9051 4831
rect 9071 4811 9085 4831
rect 9043 4773 9085 4811
rect 9135 4831 9179 4873
rect 9135 4811 9147 4831
rect 9167 4811 9179 4831
rect 9135 4773 9179 4811
rect 4866 4651 4878 4671
rect 4898 4651 4910 4671
rect 4866 4613 4910 4651
rect 5595 4616 5639 4654
rect 5595 4596 5607 4616
rect 5627 4596 5639 4616
rect 5595 4554 5639 4596
rect 5689 4616 5731 4654
rect 5689 4596 5703 4616
rect 5723 4596 5731 4616
rect 5689 4554 5731 4596
rect 5808 4616 5852 4654
rect 5808 4596 5820 4616
rect 5840 4596 5852 4616
rect 5808 4554 5852 4596
rect 5902 4616 5944 4654
rect 5902 4596 5916 4616
rect 5936 4596 5944 4616
rect 5902 4554 5944 4596
rect 6016 4616 6060 4654
rect 6016 4596 6028 4616
rect 6048 4596 6060 4616
rect 6016 4554 6060 4596
rect 6110 4616 6152 4654
rect 6110 4596 6124 4616
rect 6144 4596 6152 4616
rect 6110 4554 6152 4596
rect 6226 4616 6268 4654
rect 6226 4596 6234 4616
rect 6254 4596 6268 4616
rect 6226 4554 6268 4596
rect 6318 4623 6363 4654
rect 9424 4650 9468 4692
rect 9424 4630 9436 4650
rect 9456 4630 9468 4650
rect 9424 4623 9468 4630
rect 6318 4616 6362 4623
rect 6318 4596 6330 4616
rect 6350 4596 6362 4616
rect 6318 4554 6362 4596
rect 9423 4592 9468 4623
rect 9518 4650 9560 4692
rect 9518 4630 9532 4650
rect 9552 4630 9560 4650
rect 9518 4592 9560 4630
rect 9634 4650 9676 4692
rect 9634 4630 9642 4650
rect 9662 4630 9676 4650
rect 9634 4592 9676 4630
rect 9726 4650 9770 4692
rect 9726 4630 9738 4650
rect 9758 4630 9770 4650
rect 9726 4592 9770 4630
rect 9842 4650 9884 4692
rect 9842 4630 9850 4650
rect 9870 4630 9884 4650
rect 9842 4592 9884 4630
rect 9934 4650 9978 4692
rect 9934 4630 9946 4650
rect 9966 4630 9978 4650
rect 9934 4592 9978 4630
rect 10055 4650 10097 4692
rect 10055 4630 10063 4650
rect 10083 4630 10097 4650
rect 10055 4592 10097 4630
rect 10147 4650 10191 4692
rect 10147 4630 10159 4650
rect 10179 4630 10191 4650
rect 10147 4592 10191 4630
rect 2836 4420 2880 4462
rect 2836 4400 2848 4420
rect 2868 4400 2880 4420
rect 2836 4393 2880 4400
rect 1625 4327 1669 4365
rect 1625 4307 1637 4327
rect 1657 4307 1669 4327
rect 1625 4265 1669 4307
rect 1719 4327 1761 4365
rect 1719 4307 1733 4327
rect 1753 4307 1761 4327
rect 1719 4265 1761 4307
rect 1838 4327 1882 4365
rect 1838 4307 1850 4327
rect 1870 4307 1882 4327
rect 1838 4265 1882 4307
rect 1932 4327 1974 4365
rect 1932 4307 1946 4327
rect 1966 4307 1974 4327
rect 1932 4265 1974 4307
rect 2046 4327 2090 4365
rect 2046 4307 2058 4327
rect 2078 4307 2090 4327
rect 2046 4265 2090 4307
rect 2140 4327 2182 4365
rect 2140 4307 2154 4327
rect 2174 4307 2182 4327
rect 2140 4265 2182 4307
rect 2256 4327 2298 4365
rect 2256 4307 2264 4327
rect 2284 4307 2298 4327
rect 2256 4265 2298 4307
rect 2348 4334 2393 4365
rect 2835 4362 2880 4393
rect 2930 4420 2972 4462
rect 2930 4400 2944 4420
rect 2964 4400 2972 4420
rect 2930 4362 2972 4400
rect 3046 4420 3088 4462
rect 3046 4400 3054 4420
rect 3074 4400 3088 4420
rect 3046 4362 3088 4400
rect 3138 4420 3182 4462
rect 3138 4400 3150 4420
rect 3170 4400 3182 4420
rect 3138 4362 3182 4400
rect 3254 4420 3296 4462
rect 3254 4400 3262 4420
rect 3282 4400 3296 4420
rect 3254 4362 3296 4400
rect 3346 4420 3390 4462
rect 3346 4400 3358 4420
rect 3378 4400 3390 4420
rect 3346 4362 3390 4400
rect 3467 4420 3509 4462
rect 3467 4400 3475 4420
rect 3495 4400 3509 4420
rect 3467 4362 3509 4400
rect 3559 4420 3603 4462
rect 3559 4400 3571 4420
rect 3591 4400 3603 4420
rect 3559 4362 3603 4400
rect 8117 4399 8161 4441
rect 8117 4379 8129 4399
rect 8149 4379 8161 4399
rect 8117 4372 8161 4379
rect 2348 4327 2392 4334
rect 2348 4307 2360 4327
rect 2380 4307 2392 4327
rect 2348 4265 2392 4307
rect 6906 4306 6950 4344
rect 6906 4286 6918 4306
rect 6938 4286 6950 4306
rect 6906 4244 6950 4286
rect 7000 4306 7042 4344
rect 7000 4286 7014 4306
rect 7034 4286 7042 4306
rect 7000 4244 7042 4286
rect 7119 4306 7163 4344
rect 7119 4286 7131 4306
rect 7151 4286 7163 4306
rect 7119 4244 7163 4286
rect 7213 4306 7255 4344
rect 7213 4286 7227 4306
rect 7247 4286 7255 4306
rect 7213 4244 7255 4286
rect 7327 4306 7371 4344
rect 7327 4286 7339 4306
rect 7359 4286 7371 4306
rect 7327 4244 7371 4286
rect 7421 4306 7463 4344
rect 7421 4286 7435 4306
rect 7455 4286 7463 4306
rect 7421 4244 7463 4286
rect 7537 4306 7579 4344
rect 7537 4286 7545 4306
rect 7565 4286 7579 4306
rect 7537 4244 7579 4286
rect 7629 4313 7674 4344
rect 8116 4341 8161 4372
rect 8211 4399 8253 4441
rect 8211 4379 8225 4399
rect 8245 4379 8253 4399
rect 8211 4341 8253 4379
rect 8327 4399 8369 4441
rect 8327 4379 8335 4399
rect 8355 4379 8369 4399
rect 8327 4341 8369 4379
rect 8419 4399 8463 4441
rect 8419 4379 8431 4399
rect 8451 4379 8463 4399
rect 8419 4341 8463 4379
rect 8535 4399 8577 4441
rect 8535 4379 8543 4399
rect 8563 4379 8577 4399
rect 8535 4341 8577 4379
rect 8627 4399 8671 4441
rect 8627 4379 8639 4399
rect 8659 4379 8671 4399
rect 8627 4341 8671 4379
rect 8748 4399 8790 4441
rect 8748 4379 8756 4399
rect 8776 4379 8790 4399
rect 8748 4341 8790 4379
rect 8840 4399 8884 4441
rect 8840 4379 8852 4399
rect 8872 4379 8884 4399
rect 8840 4341 8884 4379
rect 7629 4306 7673 4313
rect 7629 4286 7641 4306
rect 7661 4286 7673 4306
rect 7629 4244 7673 4286
rect 318 4076 362 4114
rect 318 4056 330 4076
rect 350 4056 362 4076
rect 318 4014 362 4056
rect 412 4076 454 4114
rect 412 4056 426 4076
rect 446 4056 454 4076
rect 412 4014 454 4056
rect 531 4076 575 4114
rect 531 4056 543 4076
rect 563 4056 575 4076
rect 531 4014 575 4056
rect 625 4076 667 4114
rect 625 4056 639 4076
rect 659 4056 667 4076
rect 625 4014 667 4056
rect 739 4076 783 4114
rect 739 4056 751 4076
rect 771 4056 783 4076
rect 739 4014 783 4056
rect 833 4076 875 4114
rect 833 4056 847 4076
rect 867 4056 875 4076
rect 833 4014 875 4056
rect 949 4076 991 4114
rect 949 4056 957 4076
rect 977 4056 991 4076
rect 949 4014 991 4056
rect 1041 4083 1086 4114
rect 4147 4110 4191 4152
rect 4147 4090 4159 4110
rect 4179 4090 4191 4110
rect 4147 4083 4191 4090
rect 1041 4076 1085 4083
rect 1041 4056 1053 4076
rect 1073 4056 1085 4076
rect 1041 4014 1085 4056
rect 4146 4052 4191 4083
rect 4241 4110 4283 4152
rect 4241 4090 4255 4110
rect 4275 4090 4283 4110
rect 4241 4052 4283 4090
rect 4357 4110 4399 4152
rect 4357 4090 4365 4110
rect 4385 4090 4399 4110
rect 4357 4052 4399 4090
rect 4449 4110 4493 4152
rect 4449 4090 4461 4110
rect 4481 4090 4493 4110
rect 4449 4052 4493 4090
rect 4565 4110 4607 4152
rect 4565 4090 4573 4110
rect 4593 4090 4607 4110
rect 4565 4052 4607 4090
rect 4657 4110 4701 4152
rect 4657 4090 4669 4110
rect 4689 4090 4701 4110
rect 4657 4052 4701 4090
rect 4778 4110 4820 4152
rect 4778 4090 4786 4110
rect 4806 4090 4820 4110
rect 4778 4052 4820 4090
rect 4870 4110 4914 4152
rect 4870 4090 4882 4110
rect 4902 4090 4914 4110
rect 4870 4052 4914 4090
rect 5599 4055 5643 4093
rect 5599 4035 5611 4055
rect 5631 4035 5643 4055
rect 1330 3895 1374 3933
rect 1330 3875 1342 3895
rect 1362 3875 1374 3895
rect 1330 3833 1374 3875
rect 1424 3895 1466 3933
rect 1424 3875 1438 3895
rect 1458 3875 1466 3895
rect 1424 3833 1466 3875
rect 1543 3895 1587 3933
rect 1543 3875 1555 3895
rect 1575 3875 1587 3895
rect 1543 3833 1587 3875
rect 1637 3895 1679 3933
rect 1637 3875 1651 3895
rect 1671 3875 1679 3895
rect 1637 3833 1679 3875
rect 1751 3895 1795 3933
rect 1751 3875 1763 3895
rect 1783 3875 1795 3895
rect 1751 3833 1795 3875
rect 1845 3895 1887 3933
rect 1845 3875 1859 3895
rect 1879 3875 1887 3895
rect 1845 3833 1887 3875
rect 1961 3895 2003 3933
rect 1961 3875 1969 3895
rect 1989 3875 2003 3895
rect 1961 3833 2003 3875
rect 2053 3902 2098 3933
rect 5599 3993 5643 4035
rect 5693 4055 5735 4093
rect 5693 4035 5707 4055
rect 5727 4035 5735 4055
rect 5693 3993 5735 4035
rect 5812 4055 5856 4093
rect 5812 4035 5824 4055
rect 5844 4035 5856 4055
rect 5812 3993 5856 4035
rect 5906 4055 5948 4093
rect 5906 4035 5920 4055
rect 5940 4035 5948 4055
rect 5906 3993 5948 4035
rect 6020 4055 6064 4093
rect 6020 4035 6032 4055
rect 6052 4035 6064 4055
rect 6020 3993 6064 4035
rect 6114 4055 6156 4093
rect 6114 4035 6128 4055
rect 6148 4035 6156 4055
rect 6114 3993 6156 4035
rect 6230 4055 6272 4093
rect 6230 4035 6238 4055
rect 6258 4035 6272 4055
rect 6230 3993 6272 4035
rect 6322 4062 6367 4093
rect 9428 4089 9472 4131
rect 9428 4069 9440 4089
rect 9460 4069 9472 4089
rect 9428 4062 9472 4069
rect 6322 4055 6366 4062
rect 6322 4035 6334 4055
rect 6354 4035 6366 4055
rect 6322 3993 6366 4035
rect 9427 4031 9472 4062
rect 9522 4089 9564 4131
rect 9522 4069 9536 4089
rect 9556 4069 9564 4089
rect 9522 4031 9564 4069
rect 9638 4089 9680 4131
rect 9638 4069 9646 4089
rect 9666 4069 9680 4089
rect 9638 4031 9680 4069
rect 9730 4089 9774 4131
rect 9730 4069 9742 4089
rect 9762 4069 9774 4089
rect 9730 4031 9774 4069
rect 9846 4089 9888 4131
rect 9846 4069 9854 4089
rect 9874 4069 9888 4089
rect 9846 4031 9888 4069
rect 9938 4089 9982 4131
rect 9938 4069 9950 4089
rect 9970 4069 9982 4089
rect 9938 4031 9982 4069
rect 10059 4089 10101 4131
rect 10059 4069 10067 4089
rect 10087 4069 10101 4089
rect 10059 4031 10101 4069
rect 10151 4089 10195 4131
rect 10151 4069 10163 4089
rect 10183 4069 10195 4089
rect 10151 4031 10195 4069
rect 2053 3895 2097 3902
rect 2053 3875 2065 3895
rect 2085 3875 2097 3895
rect 2053 3833 2097 3875
rect 3134 3876 3178 3918
rect 3134 3856 3146 3876
rect 3166 3856 3178 3876
rect 3134 3849 3178 3856
rect 3133 3818 3178 3849
rect 3228 3876 3270 3918
rect 3228 3856 3242 3876
rect 3262 3856 3270 3876
rect 3228 3818 3270 3856
rect 3344 3876 3386 3918
rect 3344 3856 3352 3876
rect 3372 3856 3386 3876
rect 3344 3818 3386 3856
rect 3436 3876 3480 3918
rect 3436 3856 3448 3876
rect 3468 3856 3480 3876
rect 3436 3818 3480 3856
rect 3552 3876 3594 3918
rect 3552 3856 3560 3876
rect 3580 3856 3594 3876
rect 3552 3818 3594 3856
rect 3644 3876 3688 3918
rect 3644 3856 3656 3876
rect 3676 3856 3688 3876
rect 3644 3818 3688 3856
rect 3765 3876 3807 3918
rect 3765 3856 3773 3876
rect 3793 3856 3807 3876
rect 3765 3818 3807 3856
rect 3857 3876 3901 3918
rect 3857 3856 3869 3876
rect 3889 3856 3901 3876
rect 6611 3874 6655 3912
rect 3857 3818 3901 3856
rect 6611 3854 6623 3874
rect 6643 3854 6655 3874
rect 6611 3812 6655 3854
rect 6705 3874 6747 3912
rect 6705 3854 6719 3874
rect 6739 3854 6747 3874
rect 6705 3812 6747 3854
rect 6824 3874 6868 3912
rect 6824 3854 6836 3874
rect 6856 3854 6868 3874
rect 6824 3812 6868 3854
rect 6918 3874 6960 3912
rect 6918 3854 6932 3874
rect 6952 3854 6960 3874
rect 6918 3812 6960 3854
rect 7032 3874 7076 3912
rect 7032 3854 7044 3874
rect 7064 3854 7076 3874
rect 7032 3812 7076 3854
rect 7126 3874 7168 3912
rect 7126 3854 7140 3874
rect 7160 3854 7168 3874
rect 7126 3812 7168 3854
rect 7242 3874 7284 3912
rect 7242 3854 7250 3874
rect 7270 3854 7284 3874
rect 7242 3812 7284 3854
rect 7334 3881 7379 3912
rect 7334 3874 7378 3881
rect 7334 3854 7346 3874
rect 7366 3854 7378 3874
rect 7334 3812 7378 3854
rect 8415 3855 8459 3897
rect 8415 3835 8427 3855
rect 8447 3835 8459 3855
rect 8415 3828 8459 3835
rect 317 3661 361 3699
rect 317 3641 329 3661
rect 349 3641 361 3661
rect 317 3599 361 3641
rect 411 3661 453 3699
rect 411 3641 425 3661
rect 445 3641 453 3661
rect 411 3599 453 3641
rect 530 3661 574 3699
rect 530 3641 542 3661
rect 562 3641 574 3661
rect 530 3599 574 3641
rect 624 3661 666 3699
rect 624 3641 638 3661
rect 658 3641 666 3661
rect 624 3599 666 3641
rect 738 3661 782 3699
rect 738 3641 750 3661
rect 770 3641 782 3661
rect 738 3599 782 3641
rect 832 3661 874 3699
rect 832 3641 846 3661
rect 866 3641 874 3661
rect 832 3599 874 3641
rect 948 3661 990 3699
rect 948 3641 956 3661
rect 976 3641 990 3661
rect 948 3599 990 3641
rect 1040 3668 1085 3699
rect 4146 3695 4190 3737
rect 4146 3675 4158 3695
rect 4178 3675 4190 3695
rect 4146 3668 4190 3675
rect 1040 3661 1084 3668
rect 1040 3641 1052 3661
rect 1072 3641 1084 3661
rect 1040 3599 1084 3641
rect 4145 3637 4190 3668
rect 4240 3695 4282 3737
rect 4240 3675 4254 3695
rect 4274 3675 4282 3695
rect 4240 3637 4282 3675
rect 4356 3695 4398 3737
rect 4356 3675 4364 3695
rect 4384 3675 4398 3695
rect 4356 3637 4398 3675
rect 4448 3695 4492 3737
rect 4448 3675 4460 3695
rect 4480 3675 4492 3695
rect 4448 3637 4492 3675
rect 4564 3695 4606 3737
rect 4564 3675 4572 3695
rect 4592 3675 4606 3695
rect 4564 3637 4606 3675
rect 4656 3695 4700 3737
rect 4656 3675 4668 3695
rect 4688 3675 4700 3695
rect 4656 3637 4700 3675
rect 4777 3695 4819 3737
rect 4777 3675 4785 3695
rect 4805 3675 4819 3695
rect 4777 3637 4819 3675
rect 4869 3695 4913 3737
rect 8414 3797 8459 3828
rect 8509 3855 8551 3897
rect 8509 3835 8523 3855
rect 8543 3835 8551 3855
rect 8509 3797 8551 3835
rect 8625 3855 8667 3897
rect 8625 3835 8633 3855
rect 8653 3835 8667 3855
rect 8625 3797 8667 3835
rect 8717 3855 8761 3897
rect 8717 3835 8729 3855
rect 8749 3835 8761 3855
rect 8717 3797 8761 3835
rect 8833 3855 8875 3897
rect 8833 3835 8841 3855
rect 8861 3835 8875 3855
rect 8833 3797 8875 3835
rect 8925 3855 8969 3897
rect 8925 3835 8937 3855
rect 8957 3835 8969 3855
rect 8925 3797 8969 3835
rect 9046 3855 9088 3897
rect 9046 3835 9054 3855
rect 9074 3835 9088 3855
rect 9046 3797 9088 3835
rect 9138 3855 9182 3897
rect 9138 3835 9150 3855
rect 9170 3835 9182 3855
rect 9138 3797 9182 3835
rect 4869 3675 4881 3695
rect 4901 3675 4913 3695
rect 4869 3637 4913 3675
rect 5598 3640 5642 3678
rect 5598 3620 5610 3640
rect 5630 3620 5642 3640
rect 5598 3578 5642 3620
rect 5692 3640 5734 3678
rect 5692 3620 5706 3640
rect 5726 3620 5734 3640
rect 5692 3578 5734 3620
rect 5811 3640 5855 3678
rect 5811 3620 5823 3640
rect 5843 3620 5855 3640
rect 5811 3578 5855 3620
rect 5905 3640 5947 3678
rect 5905 3620 5919 3640
rect 5939 3620 5947 3640
rect 5905 3578 5947 3620
rect 6019 3640 6063 3678
rect 6019 3620 6031 3640
rect 6051 3620 6063 3640
rect 6019 3578 6063 3620
rect 6113 3640 6155 3678
rect 6113 3620 6127 3640
rect 6147 3620 6155 3640
rect 6113 3578 6155 3620
rect 6229 3640 6271 3678
rect 6229 3620 6237 3640
rect 6257 3620 6271 3640
rect 6229 3578 6271 3620
rect 6321 3647 6366 3678
rect 9427 3674 9471 3716
rect 9427 3654 9439 3674
rect 9459 3654 9471 3674
rect 9427 3647 9471 3654
rect 6321 3640 6365 3647
rect 6321 3620 6333 3640
rect 6353 3620 6365 3640
rect 6321 3578 6365 3620
rect 9426 3616 9471 3647
rect 9521 3674 9563 3716
rect 9521 3654 9535 3674
rect 9555 3654 9563 3674
rect 9521 3616 9563 3654
rect 9637 3674 9679 3716
rect 9637 3654 9645 3674
rect 9665 3654 9679 3674
rect 9637 3616 9679 3654
rect 9729 3674 9773 3716
rect 9729 3654 9741 3674
rect 9761 3654 9773 3674
rect 9729 3616 9773 3654
rect 9845 3674 9887 3716
rect 9845 3654 9853 3674
rect 9873 3654 9887 3674
rect 9845 3616 9887 3654
rect 9937 3674 9981 3716
rect 9937 3654 9949 3674
rect 9969 3654 9981 3674
rect 9937 3616 9981 3654
rect 10058 3674 10100 3716
rect 10058 3654 10066 3674
rect 10086 3654 10100 3674
rect 10058 3616 10100 3654
rect 10150 3674 10194 3716
rect 10150 3654 10162 3674
rect 10182 3654 10194 3674
rect 10150 3616 10194 3654
rect 3084 3456 3128 3498
rect 3084 3436 3096 3456
rect 3116 3436 3128 3456
rect 3084 3429 3128 3436
rect 3083 3398 3128 3429
rect 3178 3456 3220 3498
rect 3178 3436 3192 3456
rect 3212 3436 3220 3456
rect 3178 3398 3220 3436
rect 3294 3456 3336 3498
rect 3294 3436 3302 3456
rect 3322 3436 3336 3456
rect 3294 3398 3336 3436
rect 3386 3456 3430 3498
rect 3386 3436 3398 3456
rect 3418 3436 3430 3456
rect 3386 3398 3430 3436
rect 3502 3456 3544 3498
rect 3502 3436 3510 3456
rect 3530 3436 3544 3456
rect 3502 3398 3544 3436
rect 3594 3456 3638 3498
rect 3594 3436 3606 3456
rect 3626 3436 3638 3456
rect 3594 3398 3638 3436
rect 3715 3456 3757 3498
rect 3715 3436 3723 3456
rect 3743 3436 3757 3456
rect 3715 3398 3757 3436
rect 3807 3456 3851 3498
rect 3807 3436 3819 3456
rect 3839 3436 3851 3456
rect 3807 3398 3851 3436
rect 8365 3435 8409 3477
rect 8365 3415 8377 3435
rect 8397 3415 8409 3435
rect 8365 3408 8409 3415
rect 8364 3377 8409 3408
rect 8459 3435 8501 3477
rect 8459 3415 8473 3435
rect 8493 3415 8501 3435
rect 8459 3377 8501 3415
rect 8575 3435 8617 3477
rect 8575 3415 8583 3435
rect 8603 3415 8617 3435
rect 8575 3377 8617 3415
rect 8667 3435 8711 3477
rect 8667 3415 8679 3435
rect 8699 3415 8711 3435
rect 8667 3377 8711 3415
rect 8783 3435 8825 3477
rect 8783 3415 8791 3435
rect 8811 3415 8825 3435
rect 8783 3377 8825 3415
rect 8875 3435 8919 3477
rect 8875 3415 8887 3435
rect 8907 3415 8919 3435
rect 8875 3377 8919 3415
rect 8996 3435 9038 3477
rect 8996 3415 9004 3435
rect 9024 3415 9038 3435
rect 8996 3377 9038 3415
rect 9088 3435 9132 3477
rect 9088 3415 9100 3435
rect 9120 3415 9132 3435
rect 9088 3377 9132 3415
rect 1385 3334 1429 3372
rect 1385 3314 1397 3334
rect 1417 3314 1429 3334
rect 1385 3272 1429 3314
rect 1479 3334 1521 3372
rect 1479 3314 1493 3334
rect 1513 3314 1521 3334
rect 1479 3272 1521 3314
rect 1598 3334 1642 3372
rect 1598 3314 1610 3334
rect 1630 3314 1642 3334
rect 1598 3272 1642 3314
rect 1692 3334 1734 3372
rect 1692 3314 1706 3334
rect 1726 3314 1734 3334
rect 1692 3272 1734 3314
rect 1806 3334 1850 3372
rect 1806 3314 1818 3334
rect 1838 3314 1850 3334
rect 1806 3272 1850 3314
rect 1900 3334 1942 3372
rect 1900 3314 1914 3334
rect 1934 3314 1942 3334
rect 1900 3272 1942 3314
rect 2016 3334 2058 3372
rect 2016 3314 2024 3334
rect 2044 3314 2058 3334
rect 2016 3272 2058 3314
rect 2108 3341 2153 3372
rect 2108 3334 2152 3341
rect 2108 3314 2120 3334
rect 2140 3314 2152 3334
rect 2108 3272 2152 3314
rect 6666 3313 6710 3351
rect 6666 3293 6678 3313
rect 6698 3293 6710 3313
rect 6666 3251 6710 3293
rect 6760 3313 6802 3351
rect 6760 3293 6774 3313
rect 6794 3293 6802 3313
rect 6760 3251 6802 3293
rect 6879 3313 6923 3351
rect 6879 3293 6891 3313
rect 6911 3293 6923 3313
rect 6879 3251 6923 3293
rect 6973 3313 7015 3351
rect 6973 3293 6987 3313
rect 7007 3293 7015 3313
rect 6973 3251 7015 3293
rect 7087 3313 7131 3351
rect 7087 3293 7099 3313
rect 7119 3293 7131 3313
rect 7087 3251 7131 3293
rect 7181 3313 7223 3351
rect 7181 3293 7195 3313
rect 7215 3293 7223 3313
rect 7181 3251 7223 3293
rect 7297 3313 7339 3351
rect 7297 3293 7305 3313
rect 7325 3293 7339 3313
rect 7297 3251 7339 3293
rect 7389 3320 7434 3351
rect 7389 3313 7433 3320
rect 7389 3293 7401 3313
rect 7421 3293 7433 3313
rect 7389 3251 7433 3293
rect 323 3095 367 3133
rect 323 3075 335 3095
rect 355 3075 367 3095
rect 323 3033 367 3075
rect 417 3095 459 3133
rect 417 3075 431 3095
rect 451 3075 459 3095
rect 417 3033 459 3075
rect 536 3095 580 3133
rect 536 3075 548 3095
rect 568 3075 580 3095
rect 536 3033 580 3075
rect 630 3095 672 3133
rect 630 3075 644 3095
rect 664 3075 672 3095
rect 630 3033 672 3075
rect 744 3095 788 3133
rect 744 3075 756 3095
rect 776 3075 788 3095
rect 744 3033 788 3075
rect 838 3095 880 3133
rect 838 3075 852 3095
rect 872 3075 880 3095
rect 838 3033 880 3075
rect 954 3095 996 3133
rect 954 3075 962 3095
rect 982 3075 996 3095
rect 954 3033 996 3075
rect 1046 3102 1091 3133
rect 4152 3129 4196 3171
rect 4152 3109 4164 3129
rect 4184 3109 4196 3129
rect 4152 3102 4196 3109
rect 1046 3095 1090 3102
rect 1046 3075 1058 3095
rect 1078 3075 1090 3095
rect 1046 3033 1090 3075
rect 4151 3071 4196 3102
rect 4246 3129 4288 3171
rect 4246 3109 4260 3129
rect 4280 3109 4288 3129
rect 4246 3071 4288 3109
rect 4362 3129 4404 3171
rect 4362 3109 4370 3129
rect 4390 3109 4404 3129
rect 4362 3071 4404 3109
rect 4454 3129 4498 3171
rect 4454 3109 4466 3129
rect 4486 3109 4498 3129
rect 4454 3071 4498 3109
rect 4570 3129 4612 3171
rect 4570 3109 4578 3129
rect 4598 3109 4612 3129
rect 4570 3071 4612 3109
rect 4662 3129 4706 3171
rect 4662 3109 4674 3129
rect 4694 3109 4706 3129
rect 4662 3071 4706 3109
rect 4783 3129 4825 3171
rect 4783 3109 4791 3129
rect 4811 3109 4825 3129
rect 4783 3071 4825 3109
rect 4875 3129 4919 3171
rect 4875 3109 4887 3129
rect 4907 3109 4919 3129
rect 4875 3071 4919 3109
rect 5604 3074 5648 3112
rect 5604 3054 5616 3074
rect 5636 3054 5648 3074
rect 1335 2914 1379 2952
rect 1335 2894 1347 2914
rect 1367 2894 1379 2914
rect 1335 2852 1379 2894
rect 1429 2914 1471 2952
rect 1429 2894 1443 2914
rect 1463 2894 1471 2914
rect 1429 2852 1471 2894
rect 1548 2914 1592 2952
rect 1548 2894 1560 2914
rect 1580 2894 1592 2914
rect 1548 2852 1592 2894
rect 1642 2914 1684 2952
rect 1642 2894 1656 2914
rect 1676 2894 1684 2914
rect 1642 2852 1684 2894
rect 1756 2914 1800 2952
rect 1756 2894 1768 2914
rect 1788 2894 1800 2914
rect 1756 2852 1800 2894
rect 1850 2914 1892 2952
rect 1850 2894 1864 2914
rect 1884 2894 1892 2914
rect 1850 2852 1892 2894
rect 1966 2914 2008 2952
rect 1966 2894 1974 2914
rect 1994 2894 2008 2914
rect 1966 2852 2008 2894
rect 2058 2921 2103 2952
rect 5604 3012 5648 3054
rect 5698 3074 5740 3112
rect 5698 3054 5712 3074
rect 5732 3054 5740 3074
rect 5698 3012 5740 3054
rect 5817 3074 5861 3112
rect 5817 3054 5829 3074
rect 5849 3054 5861 3074
rect 5817 3012 5861 3054
rect 5911 3074 5953 3112
rect 5911 3054 5925 3074
rect 5945 3054 5953 3074
rect 5911 3012 5953 3054
rect 6025 3074 6069 3112
rect 6025 3054 6037 3074
rect 6057 3054 6069 3074
rect 6025 3012 6069 3054
rect 6119 3074 6161 3112
rect 6119 3054 6133 3074
rect 6153 3054 6161 3074
rect 6119 3012 6161 3054
rect 6235 3074 6277 3112
rect 6235 3054 6243 3074
rect 6263 3054 6277 3074
rect 6235 3012 6277 3054
rect 6327 3081 6372 3112
rect 9433 3108 9477 3150
rect 9433 3088 9445 3108
rect 9465 3088 9477 3108
rect 9433 3081 9477 3088
rect 6327 3074 6371 3081
rect 6327 3054 6339 3074
rect 6359 3054 6371 3074
rect 6327 3012 6371 3054
rect 9432 3050 9477 3081
rect 9527 3108 9569 3150
rect 9527 3088 9541 3108
rect 9561 3088 9569 3108
rect 9527 3050 9569 3088
rect 9643 3108 9685 3150
rect 9643 3088 9651 3108
rect 9671 3088 9685 3108
rect 9643 3050 9685 3088
rect 9735 3108 9779 3150
rect 9735 3088 9747 3108
rect 9767 3088 9779 3108
rect 9735 3050 9779 3088
rect 9851 3108 9893 3150
rect 9851 3088 9859 3108
rect 9879 3088 9893 3108
rect 9851 3050 9893 3088
rect 9943 3108 9987 3150
rect 9943 3088 9955 3108
rect 9975 3088 9987 3108
rect 9943 3050 9987 3088
rect 10064 3108 10106 3150
rect 10064 3088 10072 3108
rect 10092 3088 10106 3108
rect 10064 3050 10106 3088
rect 10156 3108 10200 3150
rect 10156 3088 10168 3108
rect 10188 3088 10200 3108
rect 10156 3050 10200 3088
rect 2058 2914 2102 2921
rect 2058 2894 2070 2914
rect 2090 2894 2102 2914
rect 2058 2852 2102 2894
rect 3139 2895 3183 2937
rect 3139 2875 3151 2895
rect 3171 2875 3183 2895
rect 3139 2868 3183 2875
rect 3138 2837 3183 2868
rect 3233 2895 3275 2937
rect 3233 2875 3247 2895
rect 3267 2875 3275 2895
rect 3233 2837 3275 2875
rect 3349 2895 3391 2937
rect 3349 2875 3357 2895
rect 3377 2875 3391 2895
rect 3349 2837 3391 2875
rect 3441 2895 3485 2937
rect 3441 2875 3453 2895
rect 3473 2875 3485 2895
rect 3441 2837 3485 2875
rect 3557 2895 3599 2937
rect 3557 2875 3565 2895
rect 3585 2875 3599 2895
rect 3557 2837 3599 2875
rect 3649 2895 3693 2937
rect 3649 2875 3661 2895
rect 3681 2875 3693 2895
rect 3649 2837 3693 2875
rect 3770 2895 3812 2937
rect 3770 2875 3778 2895
rect 3798 2875 3812 2895
rect 3770 2837 3812 2875
rect 3862 2895 3906 2937
rect 3862 2875 3874 2895
rect 3894 2875 3906 2895
rect 6616 2893 6660 2931
rect 3862 2837 3906 2875
rect 6616 2873 6628 2893
rect 6648 2873 6660 2893
rect 6616 2831 6660 2873
rect 6710 2893 6752 2931
rect 6710 2873 6724 2893
rect 6744 2873 6752 2893
rect 6710 2831 6752 2873
rect 6829 2893 6873 2931
rect 6829 2873 6841 2893
rect 6861 2873 6873 2893
rect 6829 2831 6873 2873
rect 6923 2893 6965 2931
rect 6923 2873 6937 2893
rect 6957 2873 6965 2893
rect 6923 2831 6965 2873
rect 7037 2893 7081 2931
rect 7037 2873 7049 2893
rect 7069 2873 7081 2893
rect 7037 2831 7081 2873
rect 7131 2893 7173 2931
rect 7131 2873 7145 2893
rect 7165 2873 7173 2893
rect 7131 2831 7173 2873
rect 7247 2893 7289 2931
rect 7247 2873 7255 2893
rect 7275 2873 7289 2893
rect 7247 2831 7289 2873
rect 7339 2900 7384 2931
rect 7339 2893 7383 2900
rect 7339 2873 7351 2893
rect 7371 2873 7383 2893
rect 7339 2831 7383 2873
rect 8420 2874 8464 2916
rect 8420 2854 8432 2874
rect 8452 2854 8464 2874
rect 8420 2847 8464 2854
rect 322 2680 366 2718
rect 322 2660 334 2680
rect 354 2660 366 2680
rect 322 2618 366 2660
rect 416 2680 458 2718
rect 416 2660 430 2680
rect 450 2660 458 2680
rect 416 2618 458 2660
rect 535 2680 579 2718
rect 535 2660 547 2680
rect 567 2660 579 2680
rect 535 2618 579 2660
rect 629 2680 671 2718
rect 629 2660 643 2680
rect 663 2660 671 2680
rect 629 2618 671 2660
rect 743 2680 787 2718
rect 743 2660 755 2680
rect 775 2660 787 2680
rect 743 2618 787 2660
rect 837 2680 879 2718
rect 837 2660 851 2680
rect 871 2660 879 2680
rect 837 2618 879 2660
rect 953 2680 995 2718
rect 953 2660 961 2680
rect 981 2660 995 2680
rect 953 2618 995 2660
rect 1045 2687 1090 2718
rect 4151 2714 4195 2756
rect 4151 2694 4163 2714
rect 4183 2694 4195 2714
rect 4151 2687 4195 2694
rect 1045 2680 1089 2687
rect 1045 2660 1057 2680
rect 1077 2660 1089 2680
rect 1045 2618 1089 2660
rect 4150 2656 4195 2687
rect 4245 2714 4287 2756
rect 4245 2694 4259 2714
rect 4279 2694 4287 2714
rect 4245 2656 4287 2694
rect 4361 2714 4403 2756
rect 4361 2694 4369 2714
rect 4389 2694 4403 2714
rect 4361 2656 4403 2694
rect 4453 2714 4497 2756
rect 4453 2694 4465 2714
rect 4485 2694 4497 2714
rect 4453 2656 4497 2694
rect 4569 2714 4611 2756
rect 4569 2694 4577 2714
rect 4597 2694 4611 2714
rect 4569 2656 4611 2694
rect 4661 2714 4705 2756
rect 4661 2694 4673 2714
rect 4693 2694 4705 2714
rect 4661 2656 4705 2694
rect 4782 2714 4824 2756
rect 4782 2694 4790 2714
rect 4810 2694 4824 2714
rect 4782 2656 4824 2694
rect 4874 2714 4918 2756
rect 8419 2816 8464 2847
rect 8514 2874 8556 2916
rect 8514 2854 8528 2874
rect 8548 2854 8556 2874
rect 8514 2816 8556 2854
rect 8630 2874 8672 2916
rect 8630 2854 8638 2874
rect 8658 2854 8672 2874
rect 8630 2816 8672 2854
rect 8722 2874 8766 2916
rect 8722 2854 8734 2874
rect 8754 2854 8766 2874
rect 8722 2816 8766 2854
rect 8838 2874 8880 2916
rect 8838 2854 8846 2874
rect 8866 2854 8880 2874
rect 8838 2816 8880 2854
rect 8930 2874 8974 2916
rect 8930 2854 8942 2874
rect 8962 2854 8974 2874
rect 8930 2816 8974 2854
rect 9051 2874 9093 2916
rect 9051 2854 9059 2874
rect 9079 2854 9093 2874
rect 9051 2816 9093 2854
rect 9143 2874 9187 2916
rect 9143 2854 9155 2874
rect 9175 2854 9187 2874
rect 9143 2816 9187 2854
rect 4874 2694 4886 2714
rect 4906 2694 4918 2714
rect 4874 2656 4918 2694
rect 5603 2659 5647 2697
rect 5603 2639 5615 2659
rect 5635 2639 5647 2659
rect 5603 2597 5647 2639
rect 5697 2659 5739 2697
rect 5697 2639 5711 2659
rect 5731 2639 5739 2659
rect 5697 2597 5739 2639
rect 5816 2659 5860 2697
rect 5816 2639 5828 2659
rect 5848 2639 5860 2659
rect 5816 2597 5860 2639
rect 5910 2659 5952 2697
rect 5910 2639 5924 2659
rect 5944 2639 5952 2659
rect 5910 2597 5952 2639
rect 6024 2659 6068 2697
rect 6024 2639 6036 2659
rect 6056 2639 6068 2659
rect 6024 2597 6068 2639
rect 6118 2659 6160 2697
rect 6118 2639 6132 2659
rect 6152 2639 6160 2659
rect 6118 2597 6160 2639
rect 6234 2659 6276 2697
rect 6234 2639 6242 2659
rect 6262 2639 6276 2659
rect 6234 2597 6276 2639
rect 6326 2666 6371 2697
rect 9432 2693 9476 2735
rect 9432 2673 9444 2693
rect 9464 2673 9476 2693
rect 9432 2666 9476 2673
rect 6326 2659 6370 2666
rect 6326 2639 6338 2659
rect 6358 2639 6370 2659
rect 6326 2597 6370 2639
rect 9431 2635 9476 2666
rect 9526 2693 9568 2735
rect 9526 2673 9540 2693
rect 9560 2673 9568 2693
rect 9526 2635 9568 2673
rect 9642 2693 9684 2735
rect 9642 2673 9650 2693
rect 9670 2673 9684 2693
rect 9642 2635 9684 2673
rect 9734 2693 9778 2735
rect 9734 2673 9746 2693
rect 9766 2673 9778 2693
rect 9734 2635 9778 2673
rect 9850 2693 9892 2735
rect 9850 2673 9858 2693
rect 9878 2673 9892 2693
rect 9850 2635 9892 2673
rect 9942 2693 9986 2735
rect 9942 2673 9954 2693
rect 9974 2673 9986 2693
rect 9942 2635 9986 2673
rect 10063 2693 10105 2735
rect 10063 2673 10071 2693
rect 10091 2673 10105 2693
rect 10063 2635 10105 2673
rect 10155 2693 10199 2735
rect 10155 2673 10167 2693
rect 10187 2673 10199 2693
rect 10155 2635 10199 2673
rect 1550 2402 1594 2440
rect 1550 2382 1562 2402
rect 1582 2382 1594 2402
rect 1550 2340 1594 2382
rect 1644 2402 1686 2440
rect 1644 2382 1658 2402
rect 1678 2382 1686 2402
rect 1644 2340 1686 2382
rect 1763 2402 1807 2440
rect 1763 2382 1775 2402
rect 1795 2382 1807 2402
rect 1763 2340 1807 2382
rect 1857 2402 1899 2440
rect 1857 2382 1871 2402
rect 1891 2382 1899 2402
rect 1857 2340 1899 2382
rect 1971 2402 2015 2440
rect 1971 2382 1983 2402
rect 2003 2382 2015 2402
rect 1971 2340 2015 2382
rect 2065 2402 2107 2440
rect 2065 2382 2079 2402
rect 2099 2382 2107 2402
rect 2065 2340 2107 2382
rect 2181 2402 2223 2440
rect 2181 2382 2189 2402
rect 2209 2382 2223 2402
rect 2181 2340 2223 2382
rect 2273 2409 2318 2440
rect 2931 2428 2975 2470
rect 2273 2402 2317 2409
rect 2273 2382 2285 2402
rect 2305 2382 2317 2402
rect 2931 2408 2943 2428
rect 2963 2408 2975 2428
rect 2931 2401 2975 2408
rect 2273 2340 2317 2382
rect 2930 2370 2975 2401
rect 3025 2428 3067 2470
rect 3025 2408 3039 2428
rect 3059 2408 3067 2428
rect 3025 2370 3067 2408
rect 3141 2428 3183 2470
rect 3141 2408 3149 2428
rect 3169 2408 3183 2428
rect 3141 2370 3183 2408
rect 3233 2428 3277 2470
rect 3233 2408 3245 2428
rect 3265 2408 3277 2428
rect 3233 2370 3277 2408
rect 3349 2428 3391 2470
rect 3349 2408 3357 2428
rect 3377 2408 3391 2428
rect 3349 2370 3391 2408
rect 3441 2428 3485 2470
rect 3441 2408 3453 2428
rect 3473 2408 3485 2428
rect 3441 2370 3485 2408
rect 3562 2428 3604 2470
rect 3562 2408 3570 2428
rect 3590 2408 3604 2428
rect 3562 2370 3604 2408
rect 3654 2428 3698 2470
rect 3654 2408 3666 2428
rect 3686 2408 3698 2428
rect 3654 2370 3698 2408
rect 6831 2381 6875 2419
rect 6831 2361 6843 2381
rect 6863 2361 6875 2381
rect 6831 2319 6875 2361
rect 6925 2381 6967 2419
rect 6925 2361 6939 2381
rect 6959 2361 6967 2381
rect 6925 2319 6967 2361
rect 7044 2381 7088 2419
rect 7044 2361 7056 2381
rect 7076 2361 7088 2381
rect 7044 2319 7088 2361
rect 7138 2381 7180 2419
rect 7138 2361 7152 2381
rect 7172 2361 7180 2381
rect 7138 2319 7180 2361
rect 7252 2381 7296 2419
rect 7252 2361 7264 2381
rect 7284 2361 7296 2381
rect 7252 2319 7296 2361
rect 7346 2381 7388 2419
rect 7346 2361 7360 2381
rect 7380 2361 7388 2381
rect 7346 2319 7388 2361
rect 7462 2381 7504 2419
rect 7462 2361 7470 2381
rect 7490 2361 7504 2381
rect 7462 2319 7504 2361
rect 7554 2388 7599 2419
rect 8212 2407 8256 2449
rect 7554 2381 7598 2388
rect 7554 2361 7566 2381
rect 7586 2361 7598 2381
rect 8212 2387 8224 2407
rect 8244 2387 8256 2407
rect 8212 2380 8256 2387
rect 7554 2319 7598 2361
rect 8211 2349 8256 2380
rect 8306 2407 8348 2449
rect 8306 2387 8320 2407
rect 8340 2387 8348 2407
rect 8306 2349 8348 2387
rect 8422 2407 8464 2449
rect 8422 2387 8430 2407
rect 8450 2387 8464 2407
rect 8422 2349 8464 2387
rect 8514 2407 8558 2449
rect 8514 2387 8526 2407
rect 8546 2387 8558 2407
rect 8514 2349 8558 2387
rect 8630 2407 8672 2449
rect 8630 2387 8638 2407
rect 8658 2387 8672 2407
rect 8630 2349 8672 2387
rect 8722 2407 8766 2449
rect 8722 2387 8734 2407
rect 8754 2387 8766 2407
rect 8722 2349 8766 2387
rect 8843 2407 8885 2449
rect 8843 2387 8851 2407
rect 8871 2387 8885 2407
rect 8843 2349 8885 2387
rect 8935 2407 8979 2449
rect 8935 2387 8947 2407
rect 8967 2387 8979 2407
rect 8935 2349 8979 2387
rect 330 2116 374 2154
rect 330 2096 342 2116
rect 362 2096 374 2116
rect 330 2054 374 2096
rect 424 2116 466 2154
rect 424 2096 438 2116
rect 458 2096 466 2116
rect 424 2054 466 2096
rect 543 2116 587 2154
rect 543 2096 555 2116
rect 575 2096 587 2116
rect 543 2054 587 2096
rect 637 2116 679 2154
rect 637 2096 651 2116
rect 671 2096 679 2116
rect 637 2054 679 2096
rect 751 2116 795 2154
rect 751 2096 763 2116
rect 783 2096 795 2116
rect 751 2054 795 2096
rect 845 2116 887 2154
rect 845 2096 859 2116
rect 879 2096 887 2116
rect 845 2054 887 2096
rect 961 2116 1003 2154
rect 961 2096 969 2116
rect 989 2096 1003 2116
rect 961 2054 1003 2096
rect 1053 2123 1098 2154
rect 4159 2150 4203 2192
rect 4159 2130 4171 2150
rect 4191 2130 4203 2150
rect 4159 2123 4203 2130
rect 1053 2116 1097 2123
rect 1053 2096 1065 2116
rect 1085 2096 1097 2116
rect 1053 2054 1097 2096
rect 4158 2092 4203 2123
rect 4253 2150 4295 2192
rect 4253 2130 4267 2150
rect 4287 2130 4295 2150
rect 4253 2092 4295 2130
rect 4369 2150 4411 2192
rect 4369 2130 4377 2150
rect 4397 2130 4411 2150
rect 4369 2092 4411 2130
rect 4461 2150 4505 2192
rect 4461 2130 4473 2150
rect 4493 2130 4505 2150
rect 4461 2092 4505 2130
rect 4577 2150 4619 2192
rect 4577 2130 4585 2150
rect 4605 2130 4619 2150
rect 4577 2092 4619 2130
rect 4669 2150 4713 2192
rect 4669 2130 4681 2150
rect 4701 2130 4713 2150
rect 4669 2092 4713 2130
rect 4790 2150 4832 2192
rect 4790 2130 4798 2150
rect 4818 2130 4832 2150
rect 4790 2092 4832 2130
rect 4882 2150 4926 2192
rect 4882 2130 4894 2150
rect 4914 2130 4926 2150
rect 4882 2092 4926 2130
rect 5611 2095 5655 2133
rect 5611 2075 5623 2095
rect 5643 2075 5655 2095
rect 1342 1935 1386 1973
rect 1342 1915 1354 1935
rect 1374 1915 1386 1935
rect 1342 1873 1386 1915
rect 1436 1935 1478 1973
rect 1436 1915 1450 1935
rect 1470 1915 1478 1935
rect 1436 1873 1478 1915
rect 1555 1935 1599 1973
rect 1555 1915 1567 1935
rect 1587 1915 1599 1935
rect 1555 1873 1599 1915
rect 1649 1935 1691 1973
rect 1649 1915 1663 1935
rect 1683 1915 1691 1935
rect 1649 1873 1691 1915
rect 1763 1935 1807 1973
rect 1763 1915 1775 1935
rect 1795 1915 1807 1935
rect 1763 1873 1807 1915
rect 1857 1935 1899 1973
rect 1857 1915 1871 1935
rect 1891 1915 1899 1935
rect 1857 1873 1899 1915
rect 1973 1935 2015 1973
rect 1973 1915 1981 1935
rect 2001 1915 2015 1935
rect 1973 1873 2015 1915
rect 2065 1942 2110 1973
rect 5611 2033 5655 2075
rect 5705 2095 5747 2133
rect 5705 2075 5719 2095
rect 5739 2075 5747 2095
rect 5705 2033 5747 2075
rect 5824 2095 5868 2133
rect 5824 2075 5836 2095
rect 5856 2075 5868 2095
rect 5824 2033 5868 2075
rect 5918 2095 5960 2133
rect 5918 2075 5932 2095
rect 5952 2075 5960 2095
rect 5918 2033 5960 2075
rect 6032 2095 6076 2133
rect 6032 2075 6044 2095
rect 6064 2075 6076 2095
rect 6032 2033 6076 2075
rect 6126 2095 6168 2133
rect 6126 2075 6140 2095
rect 6160 2075 6168 2095
rect 6126 2033 6168 2075
rect 6242 2095 6284 2133
rect 6242 2075 6250 2095
rect 6270 2075 6284 2095
rect 6242 2033 6284 2075
rect 6334 2102 6379 2133
rect 9440 2129 9484 2171
rect 9440 2109 9452 2129
rect 9472 2109 9484 2129
rect 9440 2102 9484 2109
rect 6334 2095 6378 2102
rect 6334 2075 6346 2095
rect 6366 2075 6378 2095
rect 6334 2033 6378 2075
rect 9439 2071 9484 2102
rect 9534 2129 9576 2171
rect 9534 2109 9548 2129
rect 9568 2109 9576 2129
rect 9534 2071 9576 2109
rect 9650 2129 9692 2171
rect 9650 2109 9658 2129
rect 9678 2109 9692 2129
rect 9650 2071 9692 2109
rect 9742 2129 9786 2171
rect 9742 2109 9754 2129
rect 9774 2109 9786 2129
rect 9742 2071 9786 2109
rect 9858 2129 9900 2171
rect 9858 2109 9866 2129
rect 9886 2109 9900 2129
rect 9858 2071 9900 2109
rect 9950 2129 9994 2171
rect 9950 2109 9962 2129
rect 9982 2109 9994 2129
rect 9950 2071 9994 2109
rect 10071 2129 10113 2171
rect 10071 2109 10079 2129
rect 10099 2109 10113 2129
rect 10071 2071 10113 2109
rect 10163 2129 10207 2171
rect 10163 2109 10175 2129
rect 10195 2109 10207 2129
rect 10163 2071 10207 2109
rect 2065 1935 2109 1942
rect 2065 1915 2077 1935
rect 2097 1915 2109 1935
rect 2065 1873 2109 1915
rect 3146 1916 3190 1958
rect 3146 1896 3158 1916
rect 3178 1896 3190 1916
rect 3146 1889 3190 1896
rect 3145 1858 3190 1889
rect 3240 1916 3282 1958
rect 3240 1896 3254 1916
rect 3274 1896 3282 1916
rect 3240 1858 3282 1896
rect 3356 1916 3398 1958
rect 3356 1896 3364 1916
rect 3384 1896 3398 1916
rect 3356 1858 3398 1896
rect 3448 1916 3492 1958
rect 3448 1896 3460 1916
rect 3480 1896 3492 1916
rect 3448 1858 3492 1896
rect 3564 1916 3606 1958
rect 3564 1896 3572 1916
rect 3592 1896 3606 1916
rect 3564 1858 3606 1896
rect 3656 1916 3700 1958
rect 3656 1896 3668 1916
rect 3688 1896 3700 1916
rect 3656 1858 3700 1896
rect 3777 1916 3819 1958
rect 3777 1896 3785 1916
rect 3805 1896 3819 1916
rect 3777 1858 3819 1896
rect 3869 1916 3913 1958
rect 3869 1896 3881 1916
rect 3901 1896 3913 1916
rect 6623 1914 6667 1952
rect 3869 1858 3913 1896
rect 6623 1894 6635 1914
rect 6655 1894 6667 1914
rect 6623 1852 6667 1894
rect 6717 1914 6759 1952
rect 6717 1894 6731 1914
rect 6751 1894 6759 1914
rect 6717 1852 6759 1894
rect 6836 1914 6880 1952
rect 6836 1894 6848 1914
rect 6868 1894 6880 1914
rect 6836 1852 6880 1894
rect 6930 1914 6972 1952
rect 6930 1894 6944 1914
rect 6964 1894 6972 1914
rect 6930 1852 6972 1894
rect 7044 1914 7088 1952
rect 7044 1894 7056 1914
rect 7076 1894 7088 1914
rect 7044 1852 7088 1894
rect 7138 1914 7180 1952
rect 7138 1894 7152 1914
rect 7172 1894 7180 1914
rect 7138 1852 7180 1894
rect 7254 1914 7296 1952
rect 7254 1894 7262 1914
rect 7282 1894 7296 1914
rect 7254 1852 7296 1894
rect 7346 1921 7391 1952
rect 7346 1914 7390 1921
rect 7346 1894 7358 1914
rect 7378 1894 7390 1914
rect 7346 1852 7390 1894
rect 8427 1895 8471 1937
rect 8427 1875 8439 1895
rect 8459 1875 8471 1895
rect 8427 1868 8471 1875
rect 329 1701 373 1739
rect 329 1681 341 1701
rect 361 1681 373 1701
rect 329 1639 373 1681
rect 423 1701 465 1739
rect 423 1681 437 1701
rect 457 1681 465 1701
rect 423 1639 465 1681
rect 542 1701 586 1739
rect 542 1681 554 1701
rect 574 1681 586 1701
rect 542 1639 586 1681
rect 636 1701 678 1739
rect 636 1681 650 1701
rect 670 1681 678 1701
rect 636 1639 678 1681
rect 750 1701 794 1739
rect 750 1681 762 1701
rect 782 1681 794 1701
rect 750 1639 794 1681
rect 844 1701 886 1739
rect 844 1681 858 1701
rect 878 1681 886 1701
rect 844 1639 886 1681
rect 960 1701 1002 1739
rect 960 1681 968 1701
rect 988 1681 1002 1701
rect 960 1639 1002 1681
rect 1052 1708 1097 1739
rect 4158 1735 4202 1777
rect 4158 1715 4170 1735
rect 4190 1715 4202 1735
rect 4158 1708 4202 1715
rect 1052 1701 1096 1708
rect 1052 1681 1064 1701
rect 1084 1681 1096 1701
rect 1052 1639 1096 1681
rect 4157 1677 4202 1708
rect 4252 1735 4294 1777
rect 4252 1715 4266 1735
rect 4286 1715 4294 1735
rect 4252 1677 4294 1715
rect 4368 1735 4410 1777
rect 4368 1715 4376 1735
rect 4396 1715 4410 1735
rect 4368 1677 4410 1715
rect 4460 1735 4504 1777
rect 4460 1715 4472 1735
rect 4492 1715 4504 1735
rect 4460 1677 4504 1715
rect 4576 1735 4618 1777
rect 4576 1715 4584 1735
rect 4604 1715 4618 1735
rect 4576 1677 4618 1715
rect 4668 1735 4712 1777
rect 4668 1715 4680 1735
rect 4700 1715 4712 1735
rect 4668 1677 4712 1715
rect 4789 1735 4831 1777
rect 4789 1715 4797 1735
rect 4817 1715 4831 1735
rect 4789 1677 4831 1715
rect 4881 1735 4925 1777
rect 8426 1837 8471 1868
rect 8521 1895 8563 1937
rect 8521 1875 8535 1895
rect 8555 1875 8563 1895
rect 8521 1837 8563 1875
rect 8637 1895 8679 1937
rect 8637 1875 8645 1895
rect 8665 1875 8679 1895
rect 8637 1837 8679 1875
rect 8729 1895 8773 1937
rect 8729 1875 8741 1895
rect 8761 1875 8773 1895
rect 8729 1837 8773 1875
rect 8845 1895 8887 1937
rect 8845 1875 8853 1895
rect 8873 1875 8887 1895
rect 8845 1837 8887 1875
rect 8937 1895 8981 1937
rect 8937 1875 8949 1895
rect 8969 1875 8981 1895
rect 8937 1837 8981 1875
rect 9058 1895 9100 1937
rect 9058 1875 9066 1895
rect 9086 1875 9100 1895
rect 9058 1837 9100 1875
rect 9150 1895 9194 1937
rect 9150 1875 9162 1895
rect 9182 1875 9194 1895
rect 9150 1837 9194 1875
rect 4881 1715 4893 1735
rect 4913 1715 4925 1735
rect 4881 1677 4925 1715
rect 5610 1680 5654 1718
rect 5610 1660 5622 1680
rect 5642 1660 5654 1680
rect 5610 1618 5654 1660
rect 5704 1680 5746 1718
rect 5704 1660 5718 1680
rect 5738 1660 5746 1680
rect 5704 1618 5746 1660
rect 5823 1680 5867 1718
rect 5823 1660 5835 1680
rect 5855 1660 5867 1680
rect 5823 1618 5867 1660
rect 5917 1680 5959 1718
rect 5917 1660 5931 1680
rect 5951 1660 5959 1680
rect 5917 1618 5959 1660
rect 6031 1680 6075 1718
rect 6031 1660 6043 1680
rect 6063 1660 6075 1680
rect 6031 1618 6075 1660
rect 6125 1680 6167 1718
rect 6125 1660 6139 1680
rect 6159 1660 6167 1680
rect 6125 1618 6167 1660
rect 6241 1680 6283 1718
rect 6241 1660 6249 1680
rect 6269 1660 6283 1680
rect 6241 1618 6283 1660
rect 6333 1687 6378 1718
rect 9439 1714 9483 1756
rect 9439 1694 9451 1714
rect 9471 1694 9483 1714
rect 9439 1687 9483 1694
rect 6333 1680 6377 1687
rect 6333 1660 6345 1680
rect 6365 1660 6377 1680
rect 6333 1618 6377 1660
rect 9438 1656 9483 1687
rect 9533 1714 9575 1756
rect 9533 1694 9547 1714
rect 9567 1694 9575 1714
rect 9533 1656 9575 1694
rect 9649 1714 9691 1756
rect 9649 1694 9657 1714
rect 9677 1694 9691 1714
rect 9649 1656 9691 1694
rect 9741 1714 9785 1756
rect 9741 1694 9753 1714
rect 9773 1694 9785 1714
rect 9741 1656 9785 1694
rect 9857 1714 9899 1756
rect 9857 1694 9865 1714
rect 9885 1694 9899 1714
rect 9857 1656 9899 1694
rect 9949 1714 9993 1756
rect 9949 1694 9961 1714
rect 9981 1694 9993 1714
rect 9949 1656 9993 1694
rect 10070 1714 10112 1756
rect 10070 1694 10078 1714
rect 10098 1694 10112 1714
rect 10070 1656 10112 1694
rect 10162 1714 10206 1756
rect 10162 1694 10174 1714
rect 10194 1694 10206 1714
rect 10162 1656 10206 1694
rect 3096 1496 3140 1538
rect 3096 1476 3108 1496
rect 3128 1476 3140 1496
rect 3096 1469 3140 1476
rect 3095 1438 3140 1469
rect 3190 1496 3232 1538
rect 3190 1476 3204 1496
rect 3224 1476 3232 1496
rect 3190 1438 3232 1476
rect 3306 1496 3348 1538
rect 3306 1476 3314 1496
rect 3334 1476 3348 1496
rect 3306 1438 3348 1476
rect 3398 1496 3442 1538
rect 3398 1476 3410 1496
rect 3430 1476 3442 1496
rect 3398 1438 3442 1476
rect 3514 1496 3556 1538
rect 3514 1476 3522 1496
rect 3542 1476 3556 1496
rect 3514 1438 3556 1476
rect 3606 1496 3650 1538
rect 3606 1476 3618 1496
rect 3638 1476 3650 1496
rect 3606 1438 3650 1476
rect 3727 1496 3769 1538
rect 3727 1476 3735 1496
rect 3755 1476 3769 1496
rect 3727 1438 3769 1476
rect 3819 1496 3863 1538
rect 3819 1476 3831 1496
rect 3851 1476 3863 1496
rect 3819 1438 3863 1476
rect 8377 1475 8421 1517
rect 8377 1455 8389 1475
rect 8409 1455 8421 1475
rect 8377 1448 8421 1455
rect 8376 1417 8421 1448
rect 8471 1475 8513 1517
rect 8471 1455 8485 1475
rect 8505 1455 8513 1475
rect 8471 1417 8513 1455
rect 8587 1475 8629 1517
rect 8587 1455 8595 1475
rect 8615 1455 8629 1475
rect 8587 1417 8629 1455
rect 8679 1475 8723 1517
rect 8679 1455 8691 1475
rect 8711 1455 8723 1475
rect 8679 1417 8723 1455
rect 8795 1475 8837 1517
rect 8795 1455 8803 1475
rect 8823 1455 8837 1475
rect 8795 1417 8837 1455
rect 8887 1475 8931 1517
rect 8887 1455 8899 1475
rect 8919 1455 8931 1475
rect 8887 1417 8931 1455
rect 9008 1475 9050 1517
rect 9008 1455 9016 1475
rect 9036 1455 9050 1475
rect 9008 1417 9050 1455
rect 9100 1475 9144 1517
rect 9100 1455 9112 1475
rect 9132 1455 9144 1475
rect 9100 1417 9144 1455
rect 1397 1374 1441 1412
rect 1397 1354 1409 1374
rect 1429 1354 1441 1374
rect 1397 1312 1441 1354
rect 1491 1374 1533 1412
rect 1491 1354 1505 1374
rect 1525 1354 1533 1374
rect 1491 1312 1533 1354
rect 1610 1374 1654 1412
rect 1610 1354 1622 1374
rect 1642 1354 1654 1374
rect 1610 1312 1654 1354
rect 1704 1374 1746 1412
rect 1704 1354 1718 1374
rect 1738 1354 1746 1374
rect 1704 1312 1746 1354
rect 1818 1374 1862 1412
rect 1818 1354 1830 1374
rect 1850 1354 1862 1374
rect 1818 1312 1862 1354
rect 1912 1374 1954 1412
rect 1912 1354 1926 1374
rect 1946 1354 1954 1374
rect 1912 1312 1954 1354
rect 2028 1374 2070 1412
rect 2028 1354 2036 1374
rect 2056 1354 2070 1374
rect 2028 1312 2070 1354
rect 2120 1381 2165 1412
rect 2120 1374 2164 1381
rect 2120 1354 2132 1374
rect 2152 1354 2164 1374
rect 2120 1312 2164 1354
rect 6678 1353 6722 1391
rect 6678 1333 6690 1353
rect 6710 1333 6722 1353
rect 6678 1291 6722 1333
rect 6772 1353 6814 1391
rect 6772 1333 6786 1353
rect 6806 1333 6814 1353
rect 6772 1291 6814 1333
rect 6891 1353 6935 1391
rect 6891 1333 6903 1353
rect 6923 1333 6935 1353
rect 6891 1291 6935 1333
rect 6985 1353 7027 1391
rect 6985 1333 6999 1353
rect 7019 1333 7027 1353
rect 6985 1291 7027 1333
rect 7099 1353 7143 1391
rect 7099 1333 7111 1353
rect 7131 1333 7143 1353
rect 7099 1291 7143 1333
rect 7193 1353 7235 1391
rect 7193 1333 7207 1353
rect 7227 1333 7235 1353
rect 7193 1291 7235 1333
rect 7309 1353 7351 1391
rect 7309 1333 7317 1353
rect 7337 1333 7351 1353
rect 7309 1291 7351 1333
rect 7401 1360 7446 1391
rect 7401 1353 7445 1360
rect 7401 1333 7413 1353
rect 7433 1333 7445 1353
rect 7401 1291 7445 1333
rect 335 1135 379 1173
rect 335 1115 347 1135
rect 367 1115 379 1135
rect 335 1073 379 1115
rect 429 1135 471 1173
rect 429 1115 443 1135
rect 463 1115 471 1135
rect 429 1073 471 1115
rect 548 1135 592 1173
rect 548 1115 560 1135
rect 580 1115 592 1135
rect 548 1073 592 1115
rect 642 1135 684 1173
rect 642 1115 656 1135
rect 676 1115 684 1135
rect 642 1073 684 1115
rect 756 1135 800 1173
rect 756 1115 768 1135
rect 788 1115 800 1135
rect 756 1073 800 1115
rect 850 1135 892 1173
rect 850 1115 864 1135
rect 884 1115 892 1135
rect 850 1073 892 1115
rect 966 1135 1008 1173
rect 966 1115 974 1135
rect 994 1115 1008 1135
rect 966 1073 1008 1115
rect 1058 1142 1103 1173
rect 4164 1169 4208 1211
rect 4164 1149 4176 1169
rect 4196 1149 4208 1169
rect 4164 1142 4208 1149
rect 1058 1135 1102 1142
rect 1058 1115 1070 1135
rect 1090 1115 1102 1135
rect 1058 1073 1102 1115
rect 4163 1111 4208 1142
rect 4258 1169 4300 1211
rect 4258 1149 4272 1169
rect 4292 1149 4300 1169
rect 4258 1111 4300 1149
rect 4374 1169 4416 1211
rect 4374 1149 4382 1169
rect 4402 1149 4416 1169
rect 4374 1111 4416 1149
rect 4466 1169 4510 1211
rect 4466 1149 4478 1169
rect 4498 1149 4510 1169
rect 4466 1111 4510 1149
rect 4582 1169 4624 1211
rect 4582 1149 4590 1169
rect 4610 1149 4624 1169
rect 4582 1111 4624 1149
rect 4674 1169 4718 1211
rect 4674 1149 4686 1169
rect 4706 1149 4718 1169
rect 4674 1111 4718 1149
rect 4795 1169 4837 1211
rect 4795 1149 4803 1169
rect 4823 1149 4837 1169
rect 4795 1111 4837 1149
rect 4887 1169 4931 1211
rect 4887 1149 4899 1169
rect 4919 1149 4931 1169
rect 4887 1111 4931 1149
rect 5616 1114 5660 1152
rect 5616 1094 5628 1114
rect 5648 1094 5660 1114
rect 1347 954 1391 992
rect 1347 934 1359 954
rect 1379 934 1391 954
rect 1347 892 1391 934
rect 1441 954 1483 992
rect 1441 934 1455 954
rect 1475 934 1483 954
rect 1441 892 1483 934
rect 1560 954 1604 992
rect 1560 934 1572 954
rect 1592 934 1604 954
rect 1560 892 1604 934
rect 1654 954 1696 992
rect 1654 934 1668 954
rect 1688 934 1696 954
rect 1654 892 1696 934
rect 1768 954 1812 992
rect 1768 934 1780 954
rect 1800 934 1812 954
rect 1768 892 1812 934
rect 1862 954 1904 992
rect 1862 934 1876 954
rect 1896 934 1904 954
rect 1862 892 1904 934
rect 1978 954 2020 992
rect 1978 934 1986 954
rect 2006 934 2020 954
rect 1978 892 2020 934
rect 2070 961 2115 992
rect 5616 1052 5660 1094
rect 5710 1114 5752 1152
rect 5710 1094 5724 1114
rect 5744 1094 5752 1114
rect 5710 1052 5752 1094
rect 5829 1114 5873 1152
rect 5829 1094 5841 1114
rect 5861 1094 5873 1114
rect 5829 1052 5873 1094
rect 5923 1114 5965 1152
rect 5923 1094 5937 1114
rect 5957 1094 5965 1114
rect 5923 1052 5965 1094
rect 6037 1114 6081 1152
rect 6037 1094 6049 1114
rect 6069 1094 6081 1114
rect 6037 1052 6081 1094
rect 6131 1114 6173 1152
rect 6131 1094 6145 1114
rect 6165 1094 6173 1114
rect 6131 1052 6173 1094
rect 6247 1114 6289 1152
rect 6247 1094 6255 1114
rect 6275 1094 6289 1114
rect 6247 1052 6289 1094
rect 6339 1121 6384 1152
rect 9445 1148 9489 1190
rect 9445 1128 9457 1148
rect 9477 1128 9489 1148
rect 9445 1121 9489 1128
rect 6339 1114 6383 1121
rect 6339 1094 6351 1114
rect 6371 1094 6383 1114
rect 6339 1052 6383 1094
rect 9444 1090 9489 1121
rect 9539 1148 9581 1190
rect 9539 1128 9553 1148
rect 9573 1128 9581 1148
rect 9539 1090 9581 1128
rect 9655 1148 9697 1190
rect 9655 1128 9663 1148
rect 9683 1128 9697 1148
rect 9655 1090 9697 1128
rect 9747 1148 9791 1190
rect 9747 1128 9759 1148
rect 9779 1128 9791 1148
rect 9747 1090 9791 1128
rect 9863 1148 9905 1190
rect 9863 1128 9871 1148
rect 9891 1128 9905 1148
rect 9863 1090 9905 1128
rect 9955 1148 9999 1190
rect 9955 1128 9967 1148
rect 9987 1128 9999 1148
rect 9955 1090 9999 1128
rect 10076 1148 10118 1190
rect 10076 1128 10084 1148
rect 10104 1128 10118 1148
rect 10076 1090 10118 1128
rect 10168 1148 10212 1190
rect 10168 1128 10180 1148
rect 10200 1128 10212 1148
rect 10168 1090 10212 1128
rect 2070 954 2114 961
rect 2070 934 2082 954
rect 2102 934 2114 954
rect 2070 892 2114 934
rect 3151 935 3195 977
rect 3151 915 3163 935
rect 3183 915 3195 935
rect 3151 908 3195 915
rect 3150 877 3195 908
rect 3245 935 3287 977
rect 3245 915 3259 935
rect 3279 915 3287 935
rect 3245 877 3287 915
rect 3361 935 3403 977
rect 3361 915 3369 935
rect 3389 915 3403 935
rect 3361 877 3403 915
rect 3453 935 3497 977
rect 3453 915 3465 935
rect 3485 915 3497 935
rect 3453 877 3497 915
rect 3569 935 3611 977
rect 3569 915 3577 935
rect 3597 915 3611 935
rect 3569 877 3611 915
rect 3661 935 3705 977
rect 3661 915 3673 935
rect 3693 915 3705 935
rect 3661 877 3705 915
rect 3782 935 3824 977
rect 3782 915 3790 935
rect 3810 915 3824 935
rect 3782 877 3824 915
rect 3874 935 3918 977
rect 3874 915 3886 935
rect 3906 915 3918 935
rect 6628 933 6672 971
rect 3874 877 3918 915
rect 6628 913 6640 933
rect 6660 913 6672 933
rect 6628 871 6672 913
rect 6722 933 6764 971
rect 6722 913 6736 933
rect 6756 913 6764 933
rect 6722 871 6764 913
rect 6841 933 6885 971
rect 6841 913 6853 933
rect 6873 913 6885 933
rect 6841 871 6885 913
rect 6935 933 6977 971
rect 6935 913 6949 933
rect 6969 913 6977 933
rect 6935 871 6977 913
rect 7049 933 7093 971
rect 7049 913 7061 933
rect 7081 913 7093 933
rect 7049 871 7093 913
rect 7143 933 7185 971
rect 7143 913 7157 933
rect 7177 913 7185 933
rect 7143 871 7185 913
rect 7259 933 7301 971
rect 7259 913 7267 933
rect 7287 913 7301 933
rect 7259 871 7301 913
rect 7351 940 7396 971
rect 7351 933 7395 940
rect 7351 913 7363 933
rect 7383 913 7395 933
rect 7351 871 7395 913
rect 8432 914 8476 956
rect 8432 894 8444 914
rect 8464 894 8476 914
rect 8432 887 8476 894
rect 334 720 378 758
rect 334 700 346 720
rect 366 700 378 720
rect 334 658 378 700
rect 428 720 470 758
rect 428 700 442 720
rect 462 700 470 720
rect 428 658 470 700
rect 547 720 591 758
rect 547 700 559 720
rect 579 700 591 720
rect 547 658 591 700
rect 641 720 683 758
rect 641 700 655 720
rect 675 700 683 720
rect 641 658 683 700
rect 755 720 799 758
rect 755 700 767 720
rect 787 700 799 720
rect 755 658 799 700
rect 849 720 891 758
rect 849 700 863 720
rect 883 700 891 720
rect 849 658 891 700
rect 965 720 1007 758
rect 965 700 973 720
rect 993 700 1007 720
rect 965 658 1007 700
rect 1057 727 1102 758
rect 4163 754 4207 796
rect 4163 734 4175 754
rect 4195 734 4207 754
rect 4163 727 4207 734
rect 1057 720 1101 727
rect 1057 700 1069 720
rect 1089 700 1101 720
rect 1057 658 1101 700
rect 4162 696 4207 727
rect 4257 754 4299 796
rect 4257 734 4271 754
rect 4291 734 4299 754
rect 4257 696 4299 734
rect 4373 754 4415 796
rect 4373 734 4381 754
rect 4401 734 4415 754
rect 4373 696 4415 734
rect 4465 754 4509 796
rect 4465 734 4477 754
rect 4497 734 4509 754
rect 4465 696 4509 734
rect 4581 754 4623 796
rect 4581 734 4589 754
rect 4609 734 4623 754
rect 4581 696 4623 734
rect 4673 754 4717 796
rect 4673 734 4685 754
rect 4705 734 4717 754
rect 4673 696 4717 734
rect 4794 754 4836 796
rect 4794 734 4802 754
rect 4822 734 4836 754
rect 4794 696 4836 734
rect 4886 754 4930 796
rect 8431 856 8476 887
rect 8526 914 8568 956
rect 8526 894 8540 914
rect 8560 894 8568 914
rect 8526 856 8568 894
rect 8642 914 8684 956
rect 8642 894 8650 914
rect 8670 894 8684 914
rect 8642 856 8684 894
rect 8734 914 8778 956
rect 8734 894 8746 914
rect 8766 894 8778 914
rect 8734 856 8778 894
rect 8850 914 8892 956
rect 8850 894 8858 914
rect 8878 894 8892 914
rect 8850 856 8892 894
rect 8942 914 8986 956
rect 8942 894 8954 914
rect 8974 894 8986 914
rect 8942 856 8986 894
rect 9063 914 9105 956
rect 9063 894 9071 914
rect 9091 894 9105 914
rect 9063 856 9105 894
rect 9155 914 9199 956
rect 9155 894 9167 914
rect 9187 894 9199 914
rect 9155 856 9199 894
rect 4886 734 4898 754
rect 4918 734 4930 754
rect 4886 696 4930 734
rect 5615 699 5659 737
rect 5615 679 5627 699
rect 5647 679 5659 699
rect 5615 637 5659 679
rect 5709 699 5751 737
rect 5709 679 5723 699
rect 5743 679 5751 699
rect 5709 637 5751 679
rect 5828 699 5872 737
rect 5828 679 5840 699
rect 5860 679 5872 699
rect 5828 637 5872 679
rect 5922 699 5964 737
rect 5922 679 5936 699
rect 5956 679 5964 699
rect 5922 637 5964 679
rect 6036 699 6080 737
rect 6036 679 6048 699
rect 6068 679 6080 699
rect 6036 637 6080 679
rect 6130 699 6172 737
rect 6130 679 6144 699
rect 6164 679 6172 699
rect 6130 637 6172 679
rect 6246 699 6288 737
rect 6246 679 6254 699
rect 6274 679 6288 699
rect 6246 637 6288 679
rect 6338 706 6383 737
rect 9444 733 9488 775
rect 9444 713 9456 733
rect 9476 713 9488 733
rect 9444 706 9488 713
rect 6338 699 6382 706
rect 6338 679 6350 699
rect 6370 679 6382 699
rect 6338 637 6382 679
rect 9443 675 9488 706
rect 9538 733 9580 775
rect 9538 713 9552 733
rect 9572 713 9580 733
rect 9538 675 9580 713
rect 9654 733 9696 775
rect 9654 713 9662 733
rect 9682 713 9696 733
rect 9654 675 9696 713
rect 9746 733 9790 775
rect 9746 713 9758 733
rect 9778 713 9790 733
rect 9746 675 9790 713
rect 9862 733 9904 775
rect 9862 713 9870 733
rect 9890 713 9904 733
rect 9862 675 9904 713
rect 9954 733 9998 775
rect 9954 713 9966 733
rect 9986 713 9998 733
rect 9954 675 9998 713
rect 10075 733 10117 775
rect 10075 713 10083 733
rect 10103 713 10117 733
rect 10075 675 10117 713
rect 10167 733 10211 775
rect 10167 713 10179 733
rect 10199 713 10211 733
rect 10167 675 10211 713
rect 1737 239 1781 277
rect 1737 219 1749 239
rect 1769 219 1781 239
rect 1737 177 1781 219
rect 1831 239 1873 277
rect 1831 219 1845 239
rect 1865 219 1873 239
rect 1831 177 1873 219
rect 1950 239 1994 277
rect 1950 219 1962 239
rect 1982 219 1994 239
rect 1950 177 1994 219
rect 2044 239 2086 277
rect 2044 219 2058 239
rect 2078 219 2086 239
rect 2044 177 2086 219
rect 2158 239 2202 277
rect 2158 219 2170 239
rect 2190 219 2202 239
rect 2158 177 2202 219
rect 2252 239 2294 277
rect 2252 219 2266 239
rect 2286 219 2294 239
rect 2252 177 2294 219
rect 2368 239 2410 277
rect 2368 219 2376 239
rect 2396 219 2410 239
rect 2368 177 2410 219
rect 2460 246 2505 277
rect 2460 239 2504 246
rect 2460 219 2472 239
rect 2492 219 2504 239
rect 2460 177 2504 219
rect 7018 218 7062 256
rect 7018 198 7030 218
rect 7050 198 7062 218
rect 4827 151 4871 189
rect 4827 131 4839 151
rect 4859 131 4871 151
rect 4827 89 4871 131
rect 4921 151 4963 189
rect 4921 131 4935 151
rect 4955 131 4963 151
rect 4921 89 4963 131
rect 5040 151 5084 189
rect 5040 131 5052 151
rect 5072 131 5084 151
rect 5040 89 5084 131
rect 5134 151 5176 189
rect 5134 131 5148 151
rect 5168 131 5176 151
rect 5134 89 5176 131
rect 5248 151 5292 189
rect 5248 131 5260 151
rect 5280 131 5292 151
rect 5248 89 5292 131
rect 5342 151 5384 189
rect 5342 131 5356 151
rect 5376 131 5384 151
rect 5342 89 5384 131
rect 5458 151 5500 189
rect 5458 131 5466 151
rect 5486 131 5500 151
rect 5458 89 5500 131
rect 5550 158 5595 189
rect 5550 151 5594 158
rect 7018 156 7062 198
rect 7112 218 7154 256
rect 7112 198 7126 218
rect 7146 198 7154 218
rect 7112 156 7154 198
rect 7231 218 7275 256
rect 7231 198 7243 218
rect 7263 198 7275 218
rect 7231 156 7275 198
rect 7325 218 7367 256
rect 7325 198 7339 218
rect 7359 198 7367 218
rect 7325 156 7367 198
rect 7439 218 7483 256
rect 7439 198 7451 218
rect 7471 198 7483 218
rect 7439 156 7483 198
rect 7533 218 7575 256
rect 7533 198 7547 218
rect 7567 198 7575 218
rect 7533 156 7575 198
rect 7649 218 7691 256
rect 7649 198 7657 218
rect 7677 198 7691 218
rect 7649 156 7691 198
rect 7741 225 7786 256
rect 7741 218 7785 225
rect 7741 198 7753 218
rect 7773 198 7785 218
rect 7741 156 7785 198
rect 5550 131 5562 151
rect 5582 131 5594 151
rect 5550 89 5594 131
<< ndiffc >>
rect 118 8208 136 8226
rect 4133 8156 4153 8176
rect 4236 8152 4256 8172
rect 4344 8152 4364 8172
rect 4447 8156 4467 8176
rect 4552 8152 4572 8172
rect 4655 8156 4675 8176
rect 4765 8152 4785 8172
rect 4868 8156 4888 8176
rect 5399 8187 5417 8205
rect 5048 8155 5066 8173
rect 120 8109 138 8127
rect 9414 8135 9434 8155
rect 9517 8131 9537 8151
rect 9625 8131 9645 8151
rect 9728 8135 9748 8155
rect 9833 8131 9853 8151
rect 9936 8135 9956 8155
rect 10046 8131 10066 8151
rect 10149 8135 10169 8155
rect 10329 8134 10347 8152
rect 5401 8088 5419 8106
rect 116 7994 134 8012
rect 5050 8056 5068 8074
rect 5055 7954 5073 7972
rect 118 7895 136 7913
rect 3120 7922 3140 7942
rect 3223 7918 3243 7938
rect 3331 7918 3351 7938
rect 3434 7922 3454 7942
rect 3539 7918 3559 7938
rect 3642 7922 3662 7942
rect 3752 7918 3772 7938
rect 3855 7922 3875 7942
rect 5397 7973 5415 7991
rect 304 7824 324 7844
rect 407 7828 427 7848
rect 517 7824 537 7844
rect 620 7828 640 7848
rect 725 7824 745 7844
rect 828 7828 848 7848
rect 936 7828 956 7848
rect 1039 7824 1059 7844
rect 5057 7855 5075 7873
rect 10331 8035 10349 8053
rect 10336 7933 10354 7951
rect 5399 7874 5417 7892
rect 116 7712 134 7730
rect 8401 7901 8421 7921
rect 8504 7897 8524 7917
rect 8612 7897 8632 7917
rect 8715 7901 8735 7921
rect 8820 7897 8840 7917
rect 8923 7901 8943 7921
rect 9033 7897 9053 7917
rect 9136 7901 9156 7921
rect 5585 7803 5605 7823
rect 5688 7807 5708 7827
rect 5798 7803 5818 7823
rect 5901 7807 5921 7827
rect 6006 7803 6026 7823
rect 6109 7807 6129 7827
rect 6217 7807 6237 7827
rect 6320 7803 6340 7823
rect 4132 7741 4152 7761
rect 4235 7737 4255 7757
rect 4343 7737 4363 7757
rect 4446 7741 4466 7761
rect 4551 7737 4571 7757
rect 4654 7741 4674 7761
rect 4764 7737 4784 7757
rect 4867 7741 4887 7761
rect 1316 7643 1336 7663
rect 1419 7647 1439 7667
rect 1529 7643 1549 7663
rect 1632 7647 1652 7667
rect 1737 7643 1757 7663
rect 1840 7647 1860 7667
rect 1948 7647 1968 7667
rect 2051 7643 2071 7663
rect 10338 7834 10356 7852
rect 5055 7672 5073 7690
rect 118 7613 136 7631
rect 123 7511 141 7529
rect 5397 7691 5415 7709
rect 9413 7720 9433 7740
rect 9516 7716 9536 7736
rect 9624 7716 9644 7736
rect 9727 7720 9747 7740
rect 9832 7716 9852 7736
rect 9935 7720 9955 7740
rect 10045 7716 10065 7736
rect 10148 7720 10168 7740
rect 5057 7573 5075 7591
rect 6597 7622 6617 7642
rect 6700 7626 6720 7646
rect 6810 7622 6830 7642
rect 6913 7626 6933 7646
rect 7018 7622 7038 7642
rect 7121 7626 7141 7646
rect 7229 7626 7249 7646
rect 7332 7622 7352 7642
rect 10336 7651 10354 7669
rect 5399 7592 5417 7610
rect 3070 7502 3090 7522
rect 3173 7498 3193 7518
rect 3281 7498 3301 7518
rect 3384 7502 3404 7522
rect 3489 7498 3509 7518
rect 3592 7502 3612 7522
rect 3702 7498 3722 7518
rect 3805 7502 3825 7522
rect 125 7412 143 7430
rect 303 7409 323 7429
rect 406 7413 426 7433
rect 516 7409 536 7429
rect 619 7413 639 7433
rect 724 7409 744 7429
rect 827 7413 847 7433
rect 935 7413 955 7433
rect 1038 7409 1058 7429
rect 5404 7490 5422 7508
rect 10338 7552 10356 7570
rect 5053 7458 5071 7476
rect 8351 7481 8371 7501
rect 8454 7477 8474 7497
rect 8562 7477 8582 7497
rect 8665 7481 8685 7501
rect 8770 7477 8790 7497
rect 8873 7481 8893 7501
rect 8983 7477 9003 7497
rect 9086 7481 9106 7501
rect 5406 7391 5424 7409
rect 5055 7359 5073 7377
rect 5584 7388 5604 7408
rect 5687 7392 5707 7412
rect 5797 7388 5817 7408
rect 5900 7392 5920 7412
rect 6005 7388 6025 7408
rect 6108 7392 6128 7412
rect 6216 7392 6236 7412
rect 6319 7388 6339 7408
rect 10334 7437 10352 7455
rect 10336 7338 10354 7356
rect 123 7227 141 7245
rect 125 7128 143 7146
rect 4138 7175 4158 7195
rect 4241 7171 4261 7191
rect 4349 7171 4369 7191
rect 4452 7175 4472 7195
rect 4557 7171 4577 7191
rect 4660 7175 4680 7195
rect 4770 7171 4790 7191
rect 4873 7175 4893 7195
rect 5404 7206 5422 7224
rect 5053 7174 5071 7192
rect 1371 7082 1391 7102
rect 1474 7086 1494 7106
rect 1584 7082 1604 7102
rect 1687 7086 1707 7106
rect 1792 7082 1812 7102
rect 1895 7086 1915 7106
rect 2003 7086 2023 7106
rect 2106 7082 2126 7102
rect 5406 7107 5424 7125
rect 121 7013 139 7031
rect 5055 7075 5073 7093
rect 9419 7154 9439 7174
rect 9522 7150 9542 7170
rect 9630 7150 9650 7170
rect 9733 7154 9753 7174
rect 9838 7150 9858 7170
rect 9941 7154 9961 7174
rect 10051 7150 10071 7170
rect 10154 7154 10174 7174
rect 10334 7153 10352 7171
rect 6652 7061 6672 7081
rect 6755 7065 6775 7085
rect 6865 7061 6885 7081
rect 6968 7065 6988 7085
rect 7073 7061 7093 7081
rect 7176 7065 7196 7085
rect 7284 7065 7304 7085
rect 7387 7061 7407 7081
rect 5060 6973 5078 6991
rect 123 6914 141 6932
rect 3125 6941 3145 6961
rect 3228 6937 3248 6957
rect 3336 6937 3356 6957
rect 3439 6941 3459 6961
rect 3544 6937 3564 6957
rect 3647 6941 3667 6961
rect 3757 6937 3777 6957
rect 3860 6941 3880 6961
rect 5402 6992 5420 7010
rect 309 6843 329 6863
rect 412 6847 432 6867
rect 522 6843 542 6863
rect 625 6847 645 6867
rect 730 6843 750 6863
rect 833 6847 853 6867
rect 941 6847 961 6867
rect 1044 6843 1064 6863
rect 5062 6874 5080 6892
rect 10336 7054 10354 7072
rect 10341 6952 10359 6970
rect 5404 6893 5422 6911
rect 121 6731 139 6749
rect 8406 6920 8426 6940
rect 8509 6916 8529 6936
rect 8617 6916 8637 6936
rect 8720 6920 8740 6940
rect 8825 6916 8845 6936
rect 8928 6920 8948 6940
rect 9038 6916 9058 6936
rect 9141 6920 9161 6940
rect 5590 6822 5610 6842
rect 5693 6826 5713 6846
rect 5803 6822 5823 6842
rect 5906 6826 5926 6846
rect 6011 6822 6031 6842
rect 6114 6826 6134 6846
rect 6222 6826 6242 6846
rect 6325 6822 6345 6842
rect 4137 6760 4157 6780
rect 4240 6756 4260 6776
rect 4348 6756 4368 6776
rect 4451 6760 4471 6780
rect 4556 6756 4576 6776
rect 4659 6760 4679 6780
rect 4769 6756 4789 6776
rect 4872 6760 4892 6780
rect 1321 6662 1341 6682
rect 1424 6666 1444 6686
rect 1534 6662 1554 6682
rect 1637 6666 1657 6686
rect 1742 6662 1762 6682
rect 1845 6666 1865 6686
rect 1953 6666 1973 6686
rect 2056 6662 2076 6682
rect 10343 6853 10361 6871
rect 5060 6691 5078 6709
rect 123 6632 141 6650
rect 128 6530 146 6548
rect 5402 6710 5420 6728
rect 9418 6739 9438 6759
rect 9521 6735 9541 6755
rect 9629 6735 9649 6755
rect 9732 6739 9752 6759
rect 9837 6735 9857 6755
rect 9940 6739 9960 6759
rect 10050 6735 10070 6755
rect 10153 6739 10173 6759
rect 5062 6592 5080 6610
rect 6602 6641 6622 6661
rect 6705 6645 6725 6665
rect 6815 6641 6835 6661
rect 6918 6645 6938 6665
rect 7023 6641 7043 6661
rect 7126 6645 7146 6665
rect 7234 6645 7254 6665
rect 7337 6641 7357 6661
rect 10341 6670 10359 6688
rect 5404 6611 5422 6629
rect 2917 6474 2937 6494
rect 3020 6470 3040 6490
rect 3128 6470 3148 6490
rect 3231 6474 3251 6494
rect 3336 6470 3356 6490
rect 3439 6474 3459 6494
rect 3549 6470 3569 6490
rect 3652 6474 3672 6494
rect 5409 6509 5427 6527
rect 10343 6571 10361 6589
rect 5058 6477 5076 6495
rect 130 6431 148 6449
rect 308 6428 328 6448
rect 411 6432 431 6452
rect 521 6428 541 6448
rect 624 6432 644 6452
rect 729 6428 749 6448
rect 832 6432 852 6452
rect 940 6432 960 6452
rect 1043 6428 1063 6448
rect 8198 6453 8218 6473
rect 8301 6449 8321 6469
rect 8409 6449 8429 6469
rect 8512 6453 8532 6473
rect 8617 6449 8637 6469
rect 8720 6453 8740 6473
rect 8830 6449 8850 6469
rect 8933 6453 8953 6473
rect 10339 6456 10357 6474
rect 5411 6410 5429 6428
rect 130 6248 148 6266
rect 5060 6378 5078 6396
rect 5589 6407 5609 6427
rect 5692 6411 5712 6431
rect 5802 6407 5822 6427
rect 5905 6411 5925 6431
rect 6010 6407 6030 6427
rect 6113 6411 6133 6431
rect 6221 6411 6241 6431
rect 6324 6407 6344 6427
rect 4145 6196 4165 6216
rect 4248 6192 4268 6212
rect 4356 6192 4376 6212
rect 4459 6196 4479 6216
rect 4564 6192 4584 6212
rect 4667 6196 4687 6216
rect 4777 6192 4797 6212
rect 4880 6196 4900 6216
rect 5411 6227 5429 6245
rect 10341 6357 10359 6375
rect 5060 6195 5078 6213
rect 132 6149 150 6167
rect 1536 6150 1556 6170
rect 1639 6154 1659 6174
rect 1749 6150 1769 6170
rect 1852 6154 1872 6174
rect 1957 6150 1977 6170
rect 2060 6154 2080 6174
rect 2168 6154 2188 6174
rect 2271 6150 2291 6170
rect 9426 6175 9446 6195
rect 9529 6171 9549 6191
rect 9637 6171 9657 6191
rect 9740 6175 9760 6195
rect 9845 6171 9865 6191
rect 9948 6175 9968 6195
rect 10058 6171 10078 6191
rect 10161 6175 10181 6195
rect 10341 6174 10359 6192
rect 5413 6128 5431 6146
rect 128 6034 146 6052
rect 5062 6096 5080 6114
rect 6817 6129 6837 6149
rect 6920 6133 6940 6153
rect 7030 6129 7050 6149
rect 7133 6133 7153 6153
rect 7238 6129 7258 6149
rect 7341 6133 7361 6153
rect 7449 6133 7469 6153
rect 7552 6129 7572 6149
rect 5067 5994 5085 6012
rect 130 5935 148 5953
rect 3132 5962 3152 5982
rect 3235 5958 3255 5978
rect 3343 5958 3363 5978
rect 3446 5962 3466 5982
rect 3551 5958 3571 5978
rect 3654 5962 3674 5982
rect 3764 5958 3784 5978
rect 3867 5962 3887 5982
rect 5409 6013 5427 6031
rect 316 5864 336 5884
rect 419 5868 439 5888
rect 529 5864 549 5884
rect 632 5868 652 5888
rect 737 5864 757 5884
rect 840 5868 860 5888
rect 948 5868 968 5888
rect 1051 5864 1071 5884
rect 5069 5895 5087 5913
rect 10343 6075 10361 6093
rect 10348 5973 10366 5991
rect 5411 5914 5429 5932
rect 128 5752 146 5770
rect 8413 5941 8433 5961
rect 8516 5937 8536 5957
rect 8624 5937 8644 5957
rect 8727 5941 8747 5961
rect 8832 5937 8852 5957
rect 8935 5941 8955 5961
rect 9045 5937 9065 5957
rect 9148 5941 9168 5961
rect 5597 5843 5617 5863
rect 5700 5847 5720 5867
rect 5810 5843 5830 5863
rect 5913 5847 5933 5867
rect 6018 5843 6038 5863
rect 6121 5847 6141 5867
rect 6229 5847 6249 5867
rect 6332 5843 6352 5863
rect 4144 5781 4164 5801
rect 4247 5777 4267 5797
rect 4355 5777 4375 5797
rect 4458 5781 4478 5801
rect 4563 5777 4583 5797
rect 4666 5781 4686 5801
rect 4776 5777 4796 5797
rect 4879 5781 4899 5801
rect 1328 5683 1348 5703
rect 1431 5687 1451 5707
rect 1541 5683 1561 5703
rect 1644 5687 1664 5707
rect 1749 5683 1769 5703
rect 1852 5687 1872 5707
rect 1960 5687 1980 5707
rect 2063 5683 2083 5703
rect 10350 5874 10368 5892
rect 5067 5712 5085 5730
rect 130 5653 148 5671
rect 135 5551 153 5569
rect 5409 5731 5427 5749
rect 9425 5760 9445 5780
rect 9528 5756 9548 5776
rect 9636 5756 9656 5776
rect 9739 5760 9759 5780
rect 9844 5756 9864 5776
rect 9947 5760 9967 5780
rect 10057 5756 10077 5776
rect 10160 5760 10180 5780
rect 5069 5613 5087 5631
rect 6609 5662 6629 5682
rect 6712 5666 6732 5686
rect 6822 5662 6842 5682
rect 6925 5666 6945 5686
rect 7030 5662 7050 5682
rect 7133 5666 7153 5686
rect 7241 5666 7261 5686
rect 7344 5662 7364 5682
rect 10348 5691 10366 5709
rect 5411 5632 5429 5650
rect 3082 5542 3102 5562
rect 3185 5538 3205 5558
rect 3293 5538 3313 5558
rect 3396 5542 3416 5562
rect 3501 5538 3521 5558
rect 3604 5542 3624 5562
rect 3714 5538 3734 5558
rect 3817 5542 3837 5562
rect 137 5452 155 5470
rect 315 5449 335 5469
rect 418 5453 438 5473
rect 528 5449 548 5469
rect 631 5453 651 5473
rect 736 5449 756 5469
rect 839 5453 859 5473
rect 947 5453 967 5473
rect 1050 5449 1070 5469
rect 5416 5530 5434 5548
rect 10350 5592 10368 5610
rect 5065 5498 5083 5516
rect 8363 5521 8383 5541
rect 8466 5517 8486 5537
rect 8574 5517 8594 5537
rect 8677 5521 8697 5541
rect 8782 5517 8802 5537
rect 8885 5521 8905 5541
rect 8995 5517 9015 5537
rect 9098 5521 9118 5541
rect 5418 5431 5436 5449
rect 5067 5399 5085 5417
rect 5596 5428 5616 5448
rect 5699 5432 5719 5452
rect 5809 5428 5829 5448
rect 5912 5432 5932 5452
rect 6017 5428 6037 5448
rect 6120 5432 6140 5452
rect 6228 5432 6248 5452
rect 6331 5428 6351 5448
rect 10346 5477 10364 5495
rect 10348 5378 10366 5396
rect 135 5267 153 5285
rect 137 5168 155 5186
rect 4150 5215 4170 5235
rect 4253 5211 4273 5231
rect 4361 5211 4381 5231
rect 4464 5215 4484 5235
rect 4569 5211 4589 5231
rect 4672 5215 4692 5235
rect 4782 5211 4802 5231
rect 4885 5215 4905 5235
rect 5416 5246 5434 5264
rect 5065 5214 5083 5232
rect 1383 5122 1403 5142
rect 1486 5126 1506 5146
rect 1596 5122 1616 5142
rect 1699 5126 1719 5146
rect 1804 5122 1824 5142
rect 1907 5126 1927 5146
rect 2015 5126 2035 5146
rect 2118 5122 2138 5142
rect 5418 5147 5436 5165
rect 133 5053 151 5071
rect 5067 5115 5085 5133
rect 9431 5194 9451 5214
rect 9534 5190 9554 5210
rect 9642 5190 9662 5210
rect 9745 5194 9765 5214
rect 9850 5190 9870 5210
rect 9953 5194 9973 5214
rect 10063 5190 10083 5210
rect 10166 5194 10186 5214
rect 10346 5193 10364 5211
rect 6664 5101 6684 5121
rect 6767 5105 6787 5125
rect 6877 5101 6897 5121
rect 6980 5105 7000 5125
rect 7085 5101 7105 5121
rect 7188 5105 7208 5125
rect 7296 5105 7316 5125
rect 7399 5101 7419 5121
rect 5072 5013 5090 5031
rect 135 4954 153 4972
rect 3137 4981 3157 5001
rect 3240 4977 3260 4997
rect 3348 4977 3368 4997
rect 3451 4981 3471 5001
rect 3556 4977 3576 4997
rect 3659 4981 3679 5001
rect 3769 4977 3789 4997
rect 3872 4981 3892 5001
rect 5414 5032 5432 5050
rect 321 4883 341 4903
rect 424 4887 444 4907
rect 534 4883 554 4903
rect 637 4887 657 4907
rect 742 4883 762 4903
rect 845 4887 865 4907
rect 953 4887 973 4907
rect 1056 4883 1076 4903
rect 5074 4914 5092 4932
rect 10348 5094 10366 5112
rect 10353 4992 10371 5010
rect 5416 4933 5434 4951
rect 133 4771 151 4789
rect 8418 4960 8438 4980
rect 8521 4956 8541 4976
rect 8629 4956 8649 4976
rect 8732 4960 8752 4980
rect 8837 4956 8857 4976
rect 8940 4960 8960 4980
rect 9050 4956 9070 4976
rect 9153 4960 9173 4980
rect 5602 4862 5622 4882
rect 5705 4866 5725 4886
rect 5815 4862 5835 4882
rect 5918 4866 5938 4886
rect 6023 4862 6043 4882
rect 6126 4866 6146 4886
rect 6234 4866 6254 4886
rect 6337 4862 6357 4882
rect 4149 4800 4169 4820
rect 4252 4796 4272 4816
rect 4360 4796 4380 4816
rect 4463 4800 4483 4820
rect 4568 4796 4588 4816
rect 4671 4800 4691 4820
rect 4781 4796 4801 4816
rect 4884 4800 4904 4820
rect 1333 4702 1353 4722
rect 1436 4706 1456 4726
rect 1546 4702 1566 4722
rect 1649 4706 1669 4726
rect 1754 4702 1774 4722
rect 1857 4706 1877 4726
rect 1965 4706 1985 4726
rect 2068 4702 2088 4722
rect 10355 4893 10373 4911
rect 5072 4731 5090 4749
rect 135 4672 153 4690
rect 140 4570 158 4588
rect 5414 4750 5432 4768
rect 9430 4779 9450 4799
rect 9533 4775 9553 4795
rect 9641 4775 9661 4795
rect 9744 4779 9764 4799
rect 9849 4775 9869 4795
rect 9952 4779 9972 4799
rect 10062 4775 10082 4795
rect 10165 4779 10185 4799
rect 5074 4632 5092 4650
rect 6614 4681 6634 4701
rect 6717 4685 6737 4705
rect 6827 4681 6847 4701
rect 6930 4685 6950 4705
rect 7035 4681 7055 4701
rect 7138 4685 7158 4705
rect 7246 4685 7266 4705
rect 7349 4681 7369 4701
rect 10353 4710 10371 4728
rect 5416 4651 5434 4669
rect 2842 4549 2862 4569
rect 2945 4545 2965 4565
rect 3053 4545 3073 4565
rect 3156 4549 3176 4569
rect 3261 4545 3281 4565
rect 3364 4549 3384 4569
rect 3474 4545 3494 4565
rect 3577 4549 3597 4569
rect 5421 4549 5439 4567
rect 10355 4611 10373 4629
rect 142 4471 160 4489
rect 320 4468 340 4488
rect 423 4472 443 4492
rect 533 4468 553 4488
rect 636 4472 656 4492
rect 741 4468 761 4488
rect 844 4472 864 4492
rect 952 4472 972 4492
rect 1055 4468 1075 4488
rect 5070 4517 5088 4535
rect 138 4291 156 4309
rect 8123 4528 8143 4548
rect 8226 4524 8246 4544
rect 8334 4524 8354 4544
rect 8437 4528 8457 4548
rect 8542 4524 8562 4544
rect 8645 4528 8665 4548
rect 8755 4524 8775 4544
rect 8858 4528 8878 4548
rect 5423 4450 5441 4468
rect 5072 4418 5090 4436
rect 5601 4447 5621 4467
rect 5704 4451 5724 4471
rect 5814 4447 5834 4467
rect 5917 4451 5937 4471
rect 6022 4447 6042 4467
rect 6125 4451 6145 4471
rect 6233 4451 6253 4471
rect 6336 4447 6356 4467
rect 10351 4496 10369 4514
rect 140 4192 158 4210
rect 4153 4239 4173 4259
rect 4256 4235 4276 4255
rect 4364 4235 4384 4255
rect 4467 4239 4487 4259
rect 4572 4235 4592 4255
rect 4675 4239 4695 4259
rect 4785 4235 4805 4255
rect 4888 4239 4908 4259
rect 5419 4270 5437 4288
rect 5068 4238 5086 4256
rect 1631 4158 1651 4178
rect 1734 4162 1754 4182
rect 1844 4158 1864 4178
rect 1947 4162 1967 4182
rect 2052 4158 2072 4178
rect 2155 4162 2175 4182
rect 2263 4162 2283 4182
rect 2366 4158 2386 4178
rect 10353 4397 10371 4415
rect 5421 4171 5439 4189
rect 9434 4218 9454 4238
rect 9537 4214 9557 4234
rect 9645 4214 9665 4234
rect 9748 4218 9768 4238
rect 9853 4214 9873 4234
rect 9956 4218 9976 4238
rect 10066 4214 10086 4234
rect 10169 4218 10189 4238
rect 10349 4217 10367 4235
rect 136 4077 154 4095
rect 5070 4139 5088 4157
rect 6912 4137 6932 4157
rect 7015 4141 7035 4161
rect 7125 4137 7145 4157
rect 7228 4141 7248 4161
rect 7333 4137 7353 4157
rect 7436 4141 7456 4161
rect 7544 4141 7564 4161
rect 7647 4137 7667 4157
rect 5075 4037 5093 4055
rect 138 3978 156 3996
rect 3140 4005 3160 4025
rect 3243 4001 3263 4021
rect 3351 4001 3371 4021
rect 3454 4005 3474 4025
rect 3559 4001 3579 4021
rect 3662 4005 3682 4025
rect 3772 4001 3792 4021
rect 3875 4005 3895 4025
rect 5417 4056 5435 4074
rect 324 3907 344 3927
rect 427 3911 447 3931
rect 537 3907 557 3927
rect 640 3911 660 3931
rect 745 3907 765 3927
rect 848 3911 868 3931
rect 956 3911 976 3931
rect 1059 3907 1079 3927
rect 5077 3938 5095 3956
rect 10351 4118 10369 4136
rect 10356 4016 10374 4034
rect 5419 3957 5437 3975
rect 136 3795 154 3813
rect 8421 3984 8441 4004
rect 8524 3980 8544 4000
rect 8632 3980 8652 4000
rect 8735 3984 8755 4004
rect 8840 3980 8860 4000
rect 8943 3984 8963 4004
rect 9053 3980 9073 4000
rect 9156 3984 9176 4004
rect 5605 3886 5625 3906
rect 5708 3890 5728 3910
rect 5818 3886 5838 3906
rect 5921 3890 5941 3910
rect 6026 3886 6046 3906
rect 6129 3890 6149 3910
rect 6237 3890 6257 3910
rect 6340 3886 6360 3906
rect 4152 3824 4172 3844
rect 4255 3820 4275 3840
rect 4363 3820 4383 3840
rect 4466 3824 4486 3844
rect 4571 3820 4591 3840
rect 4674 3824 4694 3844
rect 4784 3820 4804 3840
rect 4887 3824 4907 3844
rect 1336 3726 1356 3746
rect 1439 3730 1459 3750
rect 1549 3726 1569 3746
rect 1652 3730 1672 3750
rect 1757 3726 1777 3746
rect 1860 3730 1880 3750
rect 1968 3730 1988 3750
rect 2071 3726 2091 3746
rect 10358 3917 10376 3935
rect 5075 3755 5093 3773
rect 138 3696 156 3714
rect 143 3594 161 3612
rect 5417 3774 5435 3792
rect 9433 3803 9453 3823
rect 9536 3799 9556 3819
rect 9644 3799 9664 3819
rect 9747 3803 9767 3823
rect 9852 3799 9872 3819
rect 9955 3803 9975 3823
rect 10065 3799 10085 3819
rect 10168 3803 10188 3823
rect 5077 3656 5095 3674
rect 6617 3705 6637 3725
rect 6720 3709 6740 3729
rect 6830 3705 6850 3725
rect 6933 3709 6953 3729
rect 7038 3705 7058 3725
rect 7141 3709 7161 3729
rect 7249 3709 7269 3729
rect 7352 3705 7372 3725
rect 10356 3734 10374 3752
rect 5419 3675 5437 3693
rect 3090 3585 3110 3605
rect 3193 3581 3213 3601
rect 3301 3581 3321 3601
rect 3404 3585 3424 3605
rect 3509 3581 3529 3601
rect 3612 3585 3632 3605
rect 3722 3581 3742 3601
rect 3825 3585 3845 3605
rect 145 3495 163 3513
rect 323 3492 343 3512
rect 426 3496 446 3516
rect 536 3492 556 3512
rect 639 3496 659 3516
rect 744 3492 764 3512
rect 847 3496 867 3516
rect 955 3496 975 3516
rect 1058 3492 1078 3512
rect 5424 3573 5442 3591
rect 10358 3635 10376 3653
rect 5073 3541 5091 3559
rect 8371 3564 8391 3584
rect 8474 3560 8494 3580
rect 8582 3560 8602 3580
rect 8685 3564 8705 3584
rect 8790 3560 8810 3580
rect 8893 3564 8913 3584
rect 9003 3560 9023 3580
rect 9106 3564 9126 3584
rect 5426 3474 5444 3492
rect 5075 3442 5093 3460
rect 5604 3471 5624 3491
rect 5707 3475 5727 3495
rect 5817 3471 5837 3491
rect 5920 3475 5940 3495
rect 6025 3471 6045 3491
rect 6128 3475 6148 3495
rect 6236 3475 6256 3495
rect 6339 3471 6359 3491
rect 10354 3520 10372 3538
rect 10356 3421 10374 3439
rect 143 3310 161 3328
rect 145 3211 163 3229
rect 4158 3258 4178 3278
rect 4261 3254 4281 3274
rect 4369 3254 4389 3274
rect 4472 3258 4492 3278
rect 4577 3254 4597 3274
rect 4680 3258 4700 3278
rect 4790 3254 4810 3274
rect 4893 3258 4913 3278
rect 5424 3289 5442 3307
rect 5073 3257 5091 3275
rect 1391 3165 1411 3185
rect 1494 3169 1514 3189
rect 1604 3165 1624 3185
rect 1707 3169 1727 3189
rect 1812 3165 1832 3185
rect 1915 3169 1935 3189
rect 2023 3169 2043 3189
rect 2126 3165 2146 3185
rect 5426 3190 5444 3208
rect 141 3096 159 3114
rect 5075 3158 5093 3176
rect 9439 3237 9459 3257
rect 9542 3233 9562 3253
rect 9650 3233 9670 3253
rect 9753 3237 9773 3257
rect 9858 3233 9878 3253
rect 9961 3237 9981 3257
rect 10071 3233 10091 3253
rect 10174 3237 10194 3257
rect 10354 3236 10372 3254
rect 6672 3144 6692 3164
rect 6775 3148 6795 3168
rect 6885 3144 6905 3164
rect 6988 3148 7008 3168
rect 7093 3144 7113 3164
rect 7196 3148 7216 3168
rect 7304 3148 7324 3168
rect 7407 3144 7427 3164
rect 5080 3056 5098 3074
rect 143 2997 161 3015
rect 3145 3024 3165 3044
rect 3248 3020 3268 3040
rect 3356 3020 3376 3040
rect 3459 3024 3479 3044
rect 3564 3020 3584 3040
rect 3667 3024 3687 3044
rect 3777 3020 3797 3040
rect 3880 3024 3900 3044
rect 5422 3075 5440 3093
rect 329 2926 349 2946
rect 432 2930 452 2950
rect 542 2926 562 2946
rect 645 2930 665 2950
rect 750 2926 770 2946
rect 853 2930 873 2950
rect 961 2930 981 2950
rect 1064 2926 1084 2946
rect 5082 2957 5100 2975
rect 10356 3137 10374 3155
rect 10361 3035 10379 3053
rect 5424 2976 5442 2994
rect 141 2814 159 2832
rect 8426 3003 8446 3023
rect 8529 2999 8549 3019
rect 8637 2999 8657 3019
rect 8740 3003 8760 3023
rect 8845 2999 8865 3019
rect 8948 3003 8968 3023
rect 9058 2999 9078 3019
rect 9161 3003 9181 3023
rect 5610 2905 5630 2925
rect 5713 2909 5733 2929
rect 5823 2905 5843 2925
rect 5926 2909 5946 2929
rect 6031 2905 6051 2925
rect 6134 2909 6154 2929
rect 6242 2909 6262 2929
rect 6345 2905 6365 2925
rect 4157 2843 4177 2863
rect 4260 2839 4280 2859
rect 4368 2839 4388 2859
rect 4471 2843 4491 2863
rect 4576 2839 4596 2859
rect 4679 2843 4699 2863
rect 4789 2839 4809 2859
rect 4892 2843 4912 2863
rect 1341 2745 1361 2765
rect 1444 2749 1464 2769
rect 1554 2745 1574 2765
rect 1657 2749 1677 2769
rect 1762 2745 1782 2765
rect 1865 2749 1885 2769
rect 1973 2749 1993 2769
rect 2076 2745 2096 2765
rect 10363 2936 10381 2954
rect 5080 2774 5098 2792
rect 143 2715 161 2733
rect 148 2613 166 2631
rect 5422 2793 5440 2811
rect 9438 2822 9458 2842
rect 9541 2818 9561 2838
rect 9649 2818 9669 2838
rect 9752 2822 9772 2842
rect 9857 2818 9877 2838
rect 9960 2822 9980 2842
rect 10070 2818 10090 2838
rect 10173 2822 10193 2842
rect 5082 2675 5100 2693
rect 6622 2724 6642 2744
rect 6725 2728 6745 2748
rect 6835 2724 6855 2744
rect 6938 2728 6958 2748
rect 7043 2724 7063 2744
rect 7146 2728 7166 2748
rect 7254 2728 7274 2748
rect 7357 2724 7377 2744
rect 10361 2753 10379 2771
rect 5424 2694 5442 2712
rect 2937 2557 2957 2577
rect 3040 2553 3060 2573
rect 3148 2553 3168 2573
rect 3251 2557 3271 2577
rect 3356 2553 3376 2573
rect 3459 2557 3479 2577
rect 3569 2553 3589 2573
rect 3672 2557 3692 2577
rect 5429 2592 5447 2610
rect 10363 2654 10381 2672
rect 5078 2560 5096 2578
rect 150 2514 168 2532
rect 328 2511 348 2531
rect 431 2515 451 2535
rect 541 2511 561 2531
rect 644 2515 664 2535
rect 749 2511 769 2531
rect 852 2515 872 2535
rect 960 2515 980 2535
rect 1063 2511 1083 2531
rect 8218 2536 8238 2556
rect 8321 2532 8341 2552
rect 8429 2532 8449 2552
rect 8532 2536 8552 2556
rect 8637 2532 8657 2552
rect 8740 2536 8760 2556
rect 8850 2532 8870 2552
rect 8953 2536 8973 2556
rect 10359 2539 10377 2557
rect 5431 2493 5449 2511
rect 150 2331 168 2349
rect 5080 2461 5098 2479
rect 5609 2490 5629 2510
rect 5712 2494 5732 2514
rect 5822 2490 5842 2510
rect 5925 2494 5945 2514
rect 6030 2490 6050 2510
rect 6133 2494 6153 2514
rect 6241 2494 6261 2514
rect 6344 2490 6364 2510
rect 4165 2279 4185 2299
rect 4268 2275 4288 2295
rect 4376 2275 4396 2295
rect 4479 2279 4499 2299
rect 4584 2275 4604 2295
rect 4687 2279 4707 2299
rect 4797 2275 4817 2295
rect 4900 2279 4920 2299
rect 5431 2310 5449 2328
rect 10361 2440 10379 2458
rect 5080 2278 5098 2296
rect 152 2232 170 2250
rect 1556 2233 1576 2253
rect 1659 2237 1679 2257
rect 1769 2233 1789 2253
rect 1872 2237 1892 2257
rect 1977 2233 1997 2253
rect 2080 2237 2100 2257
rect 2188 2237 2208 2257
rect 2291 2233 2311 2253
rect 9446 2258 9466 2278
rect 9549 2254 9569 2274
rect 9657 2254 9677 2274
rect 9760 2258 9780 2278
rect 9865 2254 9885 2274
rect 9968 2258 9988 2278
rect 10078 2254 10098 2274
rect 10181 2258 10201 2278
rect 10361 2257 10379 2275
rect 5433 2211 5451 2229
rect 148 2117 166 2135
rect 5082 2179 5100 2197
rect 6837 2212 6857 2232
rect 6940 2216 6960 2236
rect 7050 2212 7070 2232
rect 7153 2216 7173 2236
rect 7258 2212 7278 2232
rect 7361 2216 7381 2236
rect 7469 2216 7489 2236
rect 7572 2212 7592 2232
rect 5087 2077 5105 2095
rect 150 2018 168 2036
rect 3152 2045 3172 2065
rect 3255 2041 3275 2061
rect 3363 2041 3383 2061
rect 3466 2045 3486 2065
rect 3571 2041 3591 2061
rect 3674 2045 3694 2065
rect 3784 2041 3804 2061
rect 3887 2045 3907 2065
rect 5429 2096 5447 2114
rect 336 1947 356 1967
rect 439 1951 459 1971
rect 549 1947 569 1967
rect 652 1951 672 1971
rect 757 1947 777 1967
rect 860 1951 880 1971
rect 968 1951 988 1971
rect 1071 1947 1091 1967
rect 5089 1978 5107 1996
rect 10363 2158 10381 2176
rect 10368 2056 10386 2074
rect 5431 1997 5449 2015
rect 148 1835 166 1853
rect 8433 2024 8453 2044
rect 8536 2020 8556 2040
rect 8644 2020 8664 2040
rect 8747 2024 8767 2044
rect 8852 2020 8872 2040
rect 8955 2024 8975 2044
rect 9065 2020 9085 2040
rect 9168 2024 9188 2044
rect 5617 1926 5637 1946
rect 5720 1930 5740 1950
rect 5830 1926 5850 1946
rect 5933 1930 5953 1950
rect 6038 1926 6058 1946
rect 6141 1930 6161 1950
rect 6249 1930 6269 1950
rect 6352 1926 6372 1946
rect 4164 1864 4184 1884
rect 4267 1860 4287 1880
rect 4375 1860 4395 1880
rect 4478 1864 4498 1884
rect 4583 1860 4603 1880
rect 4686 1864 4706 1884
rect 4796 1860 4816 1880
rect 4899 1864 4919 1884
rect 1348 1766 1368 1786
rect 1451 1770 1471 1790
rect 1561 1766 1581 1786
rect 1664 1770 1684 1790
rect 1769 1766 1789 1786
rect 1872 1770 1892 1790
rect 1980 1770 2000 1790
rect 2083 1766 2103 1786
rect 10370 1957 10388 1975
rect 5087 1795 5105 1813
rect 150 1736 168 1754
rect 155 1634 173 1652
rect 5429 1814 5447 1832
rect 9445 1843 9465 1863
rect 9548 1839 9568 1859
rect 9656 1839 9676 1859
rect 9759 1843 9779 1863
rect 9864 1839 9884 1859
rect 9967 1843 9987 1863
rect 10077 1839 10097 1859
rect 10180 1843 10200 1863
rect 5089 1696 5107 1714
rect 6629 1745 6649 1765
rect 6732 1749 6752 1769
rect 6842 1745 6862 1765
rect 6945 1749 6965 1769
rect 7050 1745 7070 1765
rect 7153 1749 7173 1769
rect 7261 1749 7281 1769
rect 7364 1745 7384 1765
rect 10368 1774 10386 1792
rect 5431 1715 5449 1733
rect 3102 1625 3122 1645
rect 3205 1621 3225 1641
rect 3313 1621 3333 1641
rect 3416 1625 3436 1645
rect 3521 1621 3541 1641
rect 3624 1625 3644 1645
rect 3734 1621 3754 1641
rect 3837 1625 3857 1645
rect 157 1535 175 1553
rect 335 1532 355 1552
rect 438 1536 458 1556
rect 548 1532 568 1552
rect 651 1536 671 1556
rect 756 1532 776 1552
rect 859 1536 879 1556
rect 967 1536 987 1556
rect 1070 1532 1090 1552
rect 5436 1613 5454 1631
rect 10370 1675 10388 1693
rect 5085 1581 5103 1599
rect 8383 1604 8403 1624
rect 8486 1600 8506 1620
rect 8594 1600 8614 1620
rect 8697 1604 8717 1624
rect 8802 1600 8822 1620
rect 8905 1604 8925 1624
rect 9015 1600 9035 1620
rect 9118 1604 9138 1624
rect 5438 1514 5456 1532
rect 5087 1482 5105 1500
rect 5616 1511 5636 1531
rect 5719 1515 5739 1535
rect 5829 1511 5849 1531
rect 5932 1515 5952 1535
rect 6037 1511 6057 1531
rect 6140 1515 6160 1535
rect 6248 1515 6268 1535
rect 6351 1511 6371 1531
rect 10366 1560 10384 1578
rect 10368 1461 10386 1479
rect 155 1350 173 1368
rect 157 1251 175 1269
rect 4170 1298 4190 1318
rect 4273 1294 4293 1314
rect 4381 1294 4401 1314
rect 4484 1298 4504 1318
rect 4589 1294 4609 1314
rect 4692 1298 4712 1318
rect 4802 1294 4822 1314
rect 4905 1298 4925 1318
rect 5436 1329 5454 1347
rect 5085 1297 5103 1315
rect 1403 1205 1423 1225
rect 1506 1209 1526 1229
rect 1616 1205 1636 1225
rect 1719 1209 1739 1229
rect 1824 1205 1844 1225
rect 1927 1209 1947 1229
rect 2035 1209 2055 1229
rect 2138 1205 2158 1225
rect 5438 1230 5456 1248
rect 153 1136 171 1154
rect 5087 1198 5105 1216
rect 9451 1277 9471 1297
rect 9554 1273 9574 1293
rect 9662 1273 9682 1293
rect 9765 1277 9785 1297
rect 9870 1273 9890 1293
rect 9973 1277 9993 1297
rect 10083 1273 10103 1293
rect 10186 1277 10206 1297
rect 10366 1276 10384 1294
rect 6684 1184 6704 1204
rect 6787 1188 6807 1208
rect 6897 1184 6917 1204
rect 7000 1188 7020 1208
rect 7105 1184 7125 1204
rect 7208 1188 7228 1208
rect 7316 1188 7336 1208
rect 7419 1184 7439 1204
rect 5092 1096 5110 1114
rect 155 1037 173 1055
rect 3157 1064 3177 1084
rect 3260 1060 3280 1080
rect 3368 1060 3388 1080
rect 3471 1064 3491 1084
rect 3576 1060 3596 1080
rect 3679 1064 3699 1084
rect 3789 1060 3809 1080
rect 3892 1064 3912 1084
rect 5434 1115 5452 1133
rect 341 966 361 986
rect 444 970 464 990
rect 554 966 574 986
rect 657 970 677 990
rect 762 966 782 986
rect 865 970 885 990
rect 973 970 993 990
rect 1076 966 1096 986
rect 5094 997 5112 1015
rect 10368 1177 10386 1195
rect 10373 1075 10391 1093
rect 5436 1016 5454 1034
rect 153 854 171 872
rect 8438 1043 8458 1063
rect 8541 1039 8561 1059
rect 8649 1039 8669 1059
rect 8752 1043 8772 1063
rect 8857 1039 8877 1059
rect 8960 1043 8980 1063
rect 9070 1039 9090 1059
rect 9173 1043 9193 1063
rect 5622 945 5642 965
rect 5725 949 5745 969
rect 5835 945 5855 965
rect 5938 949 5958 969
rect 6043 945 6063 965
rect 6146 949 6166 969
rect 6254 949 6274 969
rect 6357 945 6377 965
rect 4169 883 4189 903
rect 4272 879 4292 899
rect 4380 879 4400 899
rect 4483 883 4503 903
rect 4588 879 4608 899
rect 4691 883 4711 903
rect 4801 879 4821 899
rect 4904 883 4924 903
rect 1353 785 1373 805
rect 1456 789 1476 809
rect 1566 785 1586 805
rect 1669 789 1689 809
rect 1774 785 1794 805
rect 1877 789 1897 809
rect 1985 789 2005 809
rect 2088 785 2108 805
rect 10375 976 10393 994
rect 5092 814 5110 832
rect 155 755 173 773
rect 160 653 178 671
rect 5434 833 5452 851
rect 9450 862 9470 882
rect 9553 858 9573 878
rect 9661 858 9681 878
rect 9764 862 9784 882
rect 9869 858 9889 878
rect 9972 862 9992 882
rect 10082 858 10102 878
rect 10185 862 10205 882
rect 5094 715 5112 733
rect 6634 764 6654 784
rect 6737 768 6757 788
rect 6847 764 6867 784
rect 6950 768 6970 788
rect 7055 764 7075 784
rect 7158 768 7178 788
rect 7266 768 7286 788
rect 7369 764 7389 784
rect 10373 793 10391 811
rect 5436 734 5454 752
rect 5441 632 5459 650
rect 10375 694 10393 712
rect 5090 600 5108 618
rect 162 554 180 572
rect 340 551 360 571
rect 443 555 463 575
rect 553 551 573 571
rect 656 555 676 575
rect 761 551 781 571
rect 864 555 884 575
rect 972 555 992 575
rect 1075 551 1095 571
rect 10371 579 10389 597
rect 5443 533 5461 551
rect 5092 501 5110 519
rect 5621 530 5641 550
rect 5724 534 5744 554
rect 5834 530 5854 550
rect 5937 534 5957 554
rect 6042 530 6062 550
rect 6145 534 6165 554
rect 6253 534 6273 554
rect 6356 530 6376 550
rect 10373 480 10391 498
rect 1743 70 1763 90
rect 1846 74 1866 94
rect 1956 70 1976 90
rect 2059 74 2079 94
rect 2164 70 2184 90
rect 2267 74 2287 94
rect 2375 74 2395 94
rect 2478 70 2498 90
rect 7024 49 7044 69
rect 7127 53 7147 73
rect 7237 49 7257 69
rect 7340 53 7360 73
rect 7445 49 7465 69
rect 7548 53 7568 73
rect 7656 53 7676 73
rect 7759 49 7779 69
rect 4833 -18 4853 2
rect 4936 -14 4956 6
rect 5046 -18 5066 2
rect 5149 -14 5169 6
rect 5254 -18 5274 2
rect 5357 -14 5377 6
rect 5465 -14 5485 6
rect 5568 -18 5588 2
<< pdiffc >>
rect 310 7973 330 7993
rect 406 7973 426 7993
rect 523 7973 543 7993
rect 619 7973 639 7993
rect 731 7973 751 7993
rect 827 7973 847 7993
rect 937 7973 957 7993
rect 4139 8007 4159 8027
rect 1033 7973 1053 7993
rect 4235 8007 4255 8027
rect 4345 8007 4365 8027
rect 4441 8007 4461 8027
rect 4553 8007 4573 8027
rect 4649 8007 4669 8027
rect 4766 8007 4786 8027
rect 4862 8007 4882 8027
rect 5591 7952 5611 7972
rect 1322 7792 1342 7812
rect 1418 7792 1438 7812
rect 1535 7792 1555 7812
rect 1631 7792 1651 7812
rect 1743 7792 1763 7812
rect 1839 7792 1859 7812
rect 1949 7792 1969 7812
rect 5687 7952 5707 7972
rect 5804 7952 5824 7972
rect 5900 7952 5920 7972
rect 6012 7952 6032 7972
rect 6108 7952 6128 7972
rect 6218 7952 6238 7972
rect 9420 7986 9440 8006
rect 6314 7952 6334 7972
rect 9516 7986 9536 8006
rect 9626 7986 9646 8006
rect 9722 7986 9742 8006
rect 9834 7986 9854 8006
rect 9930 7986 9950 8006
rect 10047 7986 10067 8006
rect 10143 7986 10163 8006
rect 2045 7792 2065 7812
rect 3126 7773 3146 7793
rect 3222 7773 3242 7793
rect 3332 7773 3352 7793
rect 3428 7773 3448 7793
rect 3540 7773 3560 7793
rect 3636 7773 3656 7793
rect 3753 7773 3773 7793
rect 3849 7773 3869 7793
rect 6603 7771 6623 7791
rect 6699 7771 6719 7791
rect 6816 7771 6836 7791
rect 6912 7771 6932 7791
rect 7024 7771 7044 7791
rect 7120 7771 7140 7791
rect 7230 7771 7250 7791
rect 7326 7771 7346 7791
rect 8407 7752 8427 7772
rect 309 7558 329 7578
rect 405 7558 425 7578
rect 522 7558 542 7578
rect 618 7558 638 7578
rect 730 7558 750 7578
rect 826 7558 846 7578
rect 936 7558 956 7578
rect 4138 7592 4158 7612
rect 1032 7558 1052 7578
rect 4234 7592 4254 7612
rect 4344 7592 4364 7612
rect 4440 7592 4460 7612
rect 4552 7592 4572 7612
rect 4648 7592 4668 7612
rect 4765 7592 4785 7612
rect 8503 7752 8523 7772
rect 8613 7752 8633 7772
rect 8709 7752 8729 7772
rect 8821 7752 8841 7772
rect 8917 7752 8937 7772
rect 9034 7752 9054 7772
rect 9130 7752 9150 7772
rect 4861 7592 4881 7612
rect 5590 7537 5610 7557
rect 5686 7537 5706 7557
rect 5803 7537 5823 7557
rect 5899 7537 5919 7557
rect 6011 7537 6031 7557
rect 6107 7537 6127 7557
rect 6217 7537 6237 7557
rect 9419 7571 9439 7591
rect 6313 7537 6333 7557
rect 9515 7571 9535 7591
rect 9625 7571 9645 7591
rect 9721 7571 9741 7591
rect 9833 7571 9853 7591
rect 9929 7571 9949 7591
rect 10046 7571 10066 7591
rect 10142 7571 10162 7591
rect 3076 7353 3096 7373
rect 3172 7353 3192 7373
rect 3282 7353 3302 7373
rect 3378 7353 3398 7373
rect 3490 7353 3510 7373
rect 3586 7353 3606 7373
rect 3703 7353 3723 7373
rect 3799 7353 3819 7373
rect 8357 7332 8377 7352
rect 8453 7332 8473 7352
rect 8563 7332 8583 7352
rect 8659 7332 8679 7352
rect 8771 7332 8791 7352
rect 8867 7332 8887 7352
rect 8984 7332 9004 7352
rect 9080 7332 9100 7352
rect 1377 7231 1397 7251
rect 1473 7231 1493 7251
rect 1590 7231 1610 7251
rect 1686 7231 1706 7251
rect 1798 7231 1818 7251
rect 1894 7231 1914 7251
rect 2004 7231 2024 7251
rect 2100 7231 2120 7251
rect 6658 7210 6678 7230
rect 6754 7210 6774 7230
rect 6871 7210 6891 7230
rect 6967 7210 6987 7230
rect 7079 7210 7099 7230
rect 7175 7210 7195 7230
rect 7285 7210 7305 7230
rect 7381 7210 7401 7230
rect 315 6992 335 7012
rect 411 6992 431 7012
rect 528 6992 548 7012
rect 624 6992 644 7012
rect 736 6992 756 7012
rect 832 6992 852 7012
rect 942 6992 962 7012
rect 4144 7026 4164 7046
rect 1038 6992 1058 7012
rect 4240 7026 4260 7046
rect 4350 7026 4370 7046
rect 4446 7026 4466 7046
rect 4558 7026 4578 7046
rect 4654 7026 4674 7046
rect 4771 7026 4791 7046
rect 4867 7026 4887 7046
rect 5596 6971 5616 6991
rect 1327 6811 1347 6831
rect 1423 6811 1443 6831
rect 1540 6811 1560 6831
rect 1636 6811 1656 6831
rect 1748 6811 1768 6831
rect 1844 6811 1864 6831
rect 1954 6811 1974 6831
rect 5692 6971 5712 6991
rect 5809 6971 5829 6991
rect 5905 6971 5925 6991
rect 6017 6971 6037 6991
rect 6113 6971 6133 6991
rect 6223 6971 6243 6991
rect 9425 7005 9445 7025
rect 6319 6971 6339 6991
rect 9521 7005 9541 7025
rect 9631 7005 9651 7025
rect 9727 7005 9747 7025
rect 9839 7005 9859 7025
rect 9935 7005 9955 7025
rect 10052 7005 10072 7025
rect 10148 7005 10168 7025
rect 2050 6811 2070 6831
rect 3131 6792 3151 6812
rect 3227 6792 3247 6812
rect 3337 6792 3357 6812
rect 3433 6792 3453 6812
rect 3545 6792 3565 6812
rect 3641 6792 3661 6812
rect 3758 6792 3778 6812
rect 3854 6792 3874 6812
rect 6608 6790 6628 6810
rect 6704 6790 6724 6810
rect 6821 6790 6841 6810
rect 6917 6790 6937 6810
rect 7029 6790 7049 6810
rect 7125 6790 7145 6810
rect 7235 6790 7255 6810
rect 7331 6790 7351 6810
rect 8412 6771 8432 6791
rect 314 6577 334 6597
rect 410 6577 430 6597
rect 527 6577 547 6597
rect 623 6577 643 6597
rect 735 6577 755 6597
rect 831 6577 851 6597
rect 941 6577 961 6597
rect 4143 6611 4163 6631
rect 1037 6577 1057 6597
rect 4239 6611 4259 6631
rect 4349 6611 4369 6631
rect 4445 6611 4465 6631
rect 4557 6611 4577 6631
rect 4653 6611 4673 6631
rect 4770 6611 4790 6631
rect 8508 6771 8528 6791
rect 8618 6771 8638 6791
rect 8714 6771 8734 6791
rect 8826 6771 8846 6791
rect 8922 6771 8942 6791
rect 9039 6771 9059 6791
rect 9135 6771 9155 6791
rect 4866 6611 4886 6631
rect 5595 6556 5615 6576
rect 5691 6556 5711 6576
rect 5808 6556 5828 6576
rect 5904 6556 5924 6576
rect 6016 6556 6036 6576
rect 6112 6556 6132 6576
rect 6222 6556 6242 6576
rect 9424 6590 9444 6610
rect 6318 6556 6338 6576
rect 9520 6590 9540 6610
rect 9630 6590 9650 6610
rect 9726 6590 9746 6610
rect 9838 6590 9858 6610
rect 9934 6590 9954 6610
rect 10051 6590 10071 6610
rect 10147 6590 10167 6610
rect 1542 6299 1562 6319
rect 1638 6299 1658 6319
rect 1755 6299 1775 6319
rect 1851 6299 1871 6319
rect 1963 6299 1983 6319
rect 2059 6299 2079 6319
rect 2169 6299 2189 6319
rect 2265 6299 2285 6319
rect 2923 6325 2943 6345
rect 3019 6325 3039 6345
rect 3129 6325 3149 6345
rect 3225 6325 3245 6345
rect 3337 6325 3357 6345
rect 3433 6325 3453 6345
rect 3550 6325 3570 6345
rect 3646 6325 3666 6345
rect 6823 6278 6843 6298
rect 6919 6278 6939 6298
rect 7036 6278 7056 6298
rect 7132 6278 7152 6298
rect 7244 6278 7264 6298
rect 7340 6278 7360 6298
rect 7450 6278 7470 6298
rect 7546 6278 7566 6298
rect 8204 6304 8224 6324
rect 8300 6304 8320 6324
rect 8410 6304 8430 6324
rect 8506 6304 8526 6324
rect 8618 6304 8638 6324
rect 8714 6304 8734 6324
rect 8831 6304 8851 6324
rect 8927 6304 8947 6324
rect 322 6013 342 6033
rect 418 6013 438 6033
rect 535 6013 555 6033
rect 631 6013 651 6033
rect 743 6013 763 6033
rect 839 6013 859 6033
rect 949 6013 969 6033
rect 4151 6047 4171 6067
rect 1045 6013 1065 6033
rect 4247 6047 4267 6067
rect 4357 6047 4377 6067
rect 4453 6047 4473 6067
rect 4565 6047 4585 6067
rect 4661 6047 4681 6067
rect 4778 6047 4798 6067
rect 4874 6047 4894 6067
rect 5603 5992 5623 6012
rect 1334 5832 1354 5852
rect 1430 5832 1450 5852
rect 1547 5832 1567 5852
rect 1643 5832 1663 5852
rect 1755 5832 1775 5852
rect 1851 5832 1871 5852
rect 1961 5832 1981 5852
rect 5699 5992 5719 6012
rect 5816 5992 5836 6012
rect 5912 5992 5932 6012
rect 6024 5992 6044 6012
rect 6120 5992 6140 6012
rect 6230 5992 6250 6012
rect 9432 6026 9452 6046
rect 6326 5992 6346 6012
rect 9528 6026 9548 6046
rect 9638 6026 9658 6046
rect 9734 6026 9754 6046
rect 9846 6026 9866 6046
rect 9942 6026 9962 6046
rect 10059 6026 10079 6046
rect 10155 6026 10175 6046
rect 2057 5832 2077 5852
rect 3138 5813 3158 5833
rect 3234 5813 3254 5833
rect 3344 5813 3364 5833
rect 3440 5813 3460 5833
rect 3552 5813 3572 5833
rect 3648 5813 3668 5833
rect 3765 5813 3785 5833
rect 3861 5813 3881 5833
rect 6615 5811 6635 5831
rect 6711 5811 6731 5831
rect 6828 5811 6848 5831
rect 6924 5811 6944 5831
rect 7036 5811 7056 5831
rect 7132 5811 7152 5831
rect 7242 5811 7262 5831
rect 7338 5811 7358 5831
rect 8419 5792 8439 5812
rect 321 5598 341 5618
rect 417 5598 437 5618
rect 534 5598 554 5618
rect 630 5598 650 5618
rect 742 5598 762 5618
rect 838 5598 858 5618
rect 948 5598 968 5618
rect 4150 5632 4170 5652
rect 1044 5598 1064 5618
rect 4246 5632 4266 5652
rect 4356 5632 4376 5652
rect 4452 5632 4472 5652
rect 4564 5632 4584 5652
rect 4660 5632 4680 5652
rect 4777 5632 4797 5652
rect 8515 5792 8535 5812
rect 8625 5792 8645 5812
rect 8721 5792 8741 5812
rect 8833 5792 8853 5812
rect 8929 5792 8949 5812
rect 9046 5792 9066 5812
rect 9142 5792 9162 5812
rect 4873 5632 4893 5652
rect 5602 5577 5622 5597
rect 5698 5577 5718 5597
rect 5815 5577 5835 5597
rect 5911 5577 5931 5597
rect 6023 5577 6043 5597
rect 6119 5577 6139 5597
rect 6229 5577 6249 5597
rect 9431 5611 9451 5631
rect 6325 5577 6345 5597
rect 9527 5611 9547 5631
rect 9637 5611 9657 5631
rect 9733 5611 9753 5631
rect 9845 5611 9865 5631
rect 9941 5611 9961 5631
rect 10058 5611 10078 5631
rect 10154 5611 10174 5631
rect 3088 5393 3108 5413
rect 3184 5393 3204 5413
rect 3294 5393 3314 5413
rect 3390 5393 3410 5413
rect 3502 5393 3522 5413
rect 3598 5393 3618 5413
rect 3715 5393 3735 5413
rect 3811 5393 3831 5413
rect 8369 5372 8389 5392
rect 8465 5372 8485 5392
rect 8575 5372 8595 5392
rect 8671 5372 8691 5392
rect 8783 5372 8803 5392
rect 8879 5372 8899 5392
rect 8996 5372 9016 5392
rect 9092 5372 9112 5392
rect 1389 5271 1409 5291
rect 1485 5271 1505 5291
rect 1602 5271 1622 5291
rect 1698 5271 1718 5291
rect 1810 5271 1830 5291
rect 1906 5271 1926 5291
rect 2016 5271 2036 5291
rect 2112 5271 2132 5291
rect 6670 5250 6690 5270
rect 6766 5250 6786 5270
rect 6883 5250 6903 5270
rect 6979 5250 6999 5270
rect 7091 5250 7111 5270
rect 7187 5250 7207 5270
rect 7297 5250 7317 5270
rect 7393 5250 7413 5270
rect 327 5032 347 5052
rect 423 5032 443 5052
rect 540 5032 560 5052
rect 636 5032 656 5052
rect 748 5032 768 5052
rect 844 5032 864 5052
rect 954 5032 974 5052
rect 4156 5066 4176 5086
rect 1050 5032 1070 5052
rect 4252 5066 4272 5086
rect 4362 5066 4382 5086
rect 4458 5066 4478 5086
rect 4570 5066 4590 5086
rect 4666 5066 4686 5086
rect 4783 5066 4803 5086
rect 4879 5066 4899 5086
rect 5608 5011 5628 5031
rect 1339 4851 1359 4871
rect 1435 4851 1455 4871
rect 1552 4851 1572 4871
rect 1648 4851 1668 4871
rect 1760 4851 1780 4871
rect 1856 4851 1876 4871
rect 1966 4851 1986 4871
rect 5704 5011 5724 5031
rect 5821 5011 5841 5031
rect 5917 5011 5937 5031
rect 6029 5011 6049 5031
rect 6125 5011 6145 5031
rect 6235 5011 6255 5031
rect 9437 5045 9457 5065
rect 6331 5011 6351 5031
rect 9533 5045 9553 5065
rect 9643 5045 9663 5065
rect 9739 5045 9759 5065
rect 9851 5045 9871 5065
rect 9947 5045 9967 5065
rect 10064 5045 10084 5065
rect 10160 5045 10180 5065
rect 2062 4851 2082 4871
rect 3143 4832 3163 4852
rect 3239 4832 3259 4852
rect 3349 4832 3369 4852
rect 3445 4832 3465 4852
rect 3557 4832 3577 4852
rect 3653 4832 3673 4852
rect 3770 4832 3790 4852
rect 3866 4832 3886 4852
rect 6620 4830 6640 4850
rect 6716 4830 6736 4850
rect 6833 4830 6853 4850
rect 6929 4830 6949 4850
rect 7041 4830 7061 4850
rect 7137 4830 7157 4850
rect 7247 4830 7267 4850
rect 7343 4830 7363 4850
rect 8424 4811 8444 4831
rect 326 4617 346 4637
rect 422 4617 442 4637
rect 539 4617 559 4637
rect 635 4617 655 4637
rect 747 4617 767 4637
rect 843 4617 863 4637
rect 953 4617 973 4637
rect 4155 4651 4175 4671
rect 1049 4617 1069 4637
rect 4251 4651 4271 4671
rect 4361 4651 4381 4671
rect 4457 4651 4477 4671
rect 4569 4651 4589 4671
rect 4665 4651 4685 4671
rect 4782 4651 4802 4671
rect 8520 4811 8540 4831
rect 8630 4811 8650 4831
rect 8726 4811 8746 4831
rect 8838 4811 8858 4831
rect 8934 4811 8954 4831
rect 9051 4811 9071 4831
rect 9147 4811 9167 4831
rect 4878 4651 4898 4671
rect 5607 4596 5627 4616
rect 5703 4596 5723 4616
rect 5820 4596 5840 4616
rect 5916 4596 5936 4616
rect 6028 4596 6048 4616
rect 6124 4596 6144 4616
rect 6234 4596 6254 4616
rect 9436 4630 9456 4650
rect 6330 4596 6350 4616
rect 9532 4630 9552 4650
rect 9642 4630 9662 4650
rect 9738 4630 9758 4650
rect 9850 4630 9870 4650
rect 9946 4630 9966 4650
rect 10063 4630 10083 4650
rect 10159 4630 10179 4650
rect 2848 4400 2868 4420
rect 1637 4307 1657 4327
rect 1733 4307 1753 4327
rect 1850 4307 1870 4327
rect 1946 4307 1966 4327
rect 2058 4307 2078 4327
rect 2154 4307 2174 4327
rect 2264 4307 2284 4327
rect 2944 4400 2964 4420
rect 3054 4400 3074 4420
rect 3150 4400 3170 4420
rect 3262 4400 3282 4420
rect 3358 4400 3378 4420
rect 3475 4400 3495 4420
rect 3571 4400 3591 4420
rect 8129 4379 8149 4399
rect 2360 4307 2380 4327
rect 6918 4286 6938 4306
rect 7014 4286 7034 4306
rect 7131 4286 7151 4306
rect 7227 4286 7247 4306
rect 7339 4286 7359 4306
rect 7435 4286 7455 4306
rect 7545 4286 7565 4306
rect 8225 4379 8245 4399
rect 8335 4379 8355 4399
rect 8431 4379 8451 4399
rect 8543 4379 8563 4399
rect 8639 4379 8659 4399
rect 8756 4379 8776 4399
rect 8852 4379 8872 4399
rect 7641 4286 7661 4306
rect 330 4056 350 4076
rect 426 4056 446 4076
rect 543 4056 563 4076
rect 639 4056 659 4076
rect 751 4056 771 4076
rect 847 4056 867 4076
rect 957 4056 977 4076
rect 4159 4090 4179 4110
rect 1053 4056 1073 4076
rect 4255 4090 4275 4110
rect 4365 4090 4385 4110
rect 4461 4090 4481 4110
rect 4573 4090 4593 4110
rect 4669 4090 4689 4110
rect 4786 4090 4806 4110
rect 4882 4090 4902 4110
rect 5611 4035 5631 4055
rect 1342 3875 1362 3895
rect 1438 3875 1458 3895
rect 1555 3875 1575 3895
rect 1651 3875 1671 3895
rect 1763 3875 1783 3895
rect 1859 3875 1879 3895
rect 1969 3875 1989 3895
rect 5707 4035 5727 4055
rect 5824 4035 5844 4055
rect 5920 4035 5940 4055
rect 6032 4035 6052 4055
rect 6128 4035 6148 4055
rect 6238 4035 6258 4055
rect 9440 4069 9460 4089
rect 6334 4035 6354 4055
rect 9536 4069 9556 4089
rect 9646 4069 9666 4089
rect 9742 4069 9762 4089
rect 9854 4069 9874 4089
rect 9950 4069 9970 4089
rect 10067 4069 10087 4089
rect 10163 4069 10183 4089
rect 2065 3875 2085 3895
rect 3146 3856 3166 3876
rect 3242 3856 3262 3876
rect 3352 3856 3372 3876
rect 3448 3856 3468 3876
rect 3560 3856 3580 3876
rect 3656 3856 3676 3876
rect 3773 3856 3793 3876
rect 3869 3856 3889 3876
rect 6623 3854 6643 3874
rect 6719 3854 6739 3874
rect 6836 3854 6856 3874
rect 6932 3854 6952 3874
rect 7044 3854 7064 3874
rect 7140 3854 7160 3874
rect 7250 3854 7270 3874
rect 7346 3854 7366 3874
rect 8427 3835 8447 3855
rect 329 3641 349 3661
rect 425 3641 445 3661
rect 542 3641 562 3661
rect 638 3641 658 3661
rect 750 3641 770 3661
rect 846 3641 866 3661
rect 956 3641 976 3661
rect 4158 3675 4178 3695
rect 1052 3641 1072 3661
rect 4254 3675 4274 3695
rect 4364 3675 4384 3695
rect 4460 3675 4480 3695
rect 4572 3675 4592 3695
rect 4668 3675 4688 3695
rect 4785 3675 4805 3695
rect 8523 3835 8543 3855
rect 8633 3835 8653 3855
rect 8729 3835 8749 3855
rect 8841 3835 8861 3855
rect 8937 3835 8957 3855
rect 9054 3835 9074 3855
rect 9150 3835 9170 3855
rect 4881 3675 4901 3695
rect 5610 3620 5630 3640
rect 5706 3620 5726 3640
rect 5823 3620 5843 3640
rect 5919 3620 5939 3640
rect 6031 3620 6051 3640
rect 6127 3620 6147 3640
rect 6237 3620 6257 3640
rect 9439 3654 9459 3674
rect 6333 3620 6353 3640
rect 9535 3654 9555 3674
rect 9645 3654 9665 3674
rect 9741 3654 9761 3674
rect 9853 3654 9873 3674
rect 9949 3654 9969 3674
rect 10066 3654 10086 3674
rect 10162 3654 10182 3674
rect 3096 3436 3116 3456
rect 3192 3436 3212 3456
rect 3302 3436 3322 3456
rect 3398 3436 3418 3456
rect 3510 3436 3530 3456
rect 3606 3436 3626 3456
rect 3723 3436 3743 3456
rect 3819 3436 3839 3456
rect 8377 3415 8397 3435
rect 8473 3415 8493 3435
rect 8583 3415 8603 3435
rect 8679 3415 8699 3435
rect 8791 3415 8811 3435
rect 8887 3415 8907 3435
rect 9004 3415 9024 3435
rect 9100 3415 9120 3435
rect 1397 3314 1417 3334
rect 1493 3314 1513 3334
rect 1610 3314 1630 3334
rect 1706 3314 1726 3334
rect 1818 3314 1838 3334
rect 1914 3314 1934 3334
rect 2024 3314 2044 3334
rect 2120 3314 2140 3334
rect 6678 3293 6698 3313
rect 6774 3293 6794 3313
rect 6891 3293 6911 3313
rect 6987 3293 7007 3313
rect 7099 3293 7119 3313
rect 7195 3293 7215 3313
rect 7305 3293 7325 3313
rect 7401 3293 7421 3313
rect 335 3075 355 3095
rect 431 3075 451 3095
rect 548 3075 568 3095
rect 644 3075 664 3095
rect 756 3075 776 3095
rect 852 3075 872 3095
rect 962 3075 982 3095
rect 4164 3109 4184 3129
rect 1058 3075 1078 3095
rect 4260 3109 4280 3129
rect 4370 3109 4390 3129
rect 4466 3109 4486 3129
rect 4578 3109 4598 3129
rect 4674 3109 4694 3129
rect 4791 3109 4811 3129
rect 4887 3109 4907 3129
rect 5616 3054 5636 3074
rect 1347 2894 1367 2914
rect 1443 2894 1463 2914
rect 1560 2894 1580 2914
rect 1656 2894 1676 2914
rect 1768 2894 1788 2914
rect 1864 2894 1884 2914
rect 1974 2894 1994 2914
rect 5712 3054 5732 3074
rect 5829 3054 5849 3074
rect 5925 3054 5945 3074
rect 6037 3054 6057 3074
rect 6133 3054 6153 3074
rect 6243 3054 6263 3074
rect 9445 3088 9465 3108
rect 6339 3054 6359 3074
rect 9541 3088 9561 3108
rect 9651 3088 9671 3108
rect 9747 3088 9767 3108
rect 9859 3088 9879 3108
rect 9955 3088 9975 3108
rect 10072 3088 10092 3108
rect 10168 3088 10188 3108
rect 2070 2894 2090 2914
rect 3151 2875 3171 2895
rect 3247 2875 3267 2895
rect 3357 2875 3377 2895
rect 3453 2875 3473 2895
rect 3565 2875 3585 2895
rect 3661 2875 3681 2895
rect 3778 2875 3798 2895
rect 3874 2875 3894 2895
rect 6628 2873 6648 2893
rect 6724 2873 6744 2893
rect 6841 2873 6861 2893
rect 6937 2873 6957 2893
rect 7049 2873 7069 2893
rect 7145 2873 7165 2893
rect 7255 2873 7275 2893
rect 7351 2873 7371 2893
rect 8432 2854 8452 2874
rect 334 2660 354 2680
rect 430 2660 450 2680
rect 547 2660 567 2680
rect 643 2660 663 2680
rect 755 2660 775 2680
rect 851 2660 871 2680
rect 961 2660 981 2680
rect 4163 2694 4183 2714
rect 1057 2660 1077 2680
rect 4259 2694 4279 2714
rect 4369 2694 4389 2714
rect 4465 2694 4485 2714
rect 4577 2694 4597 2714
rect 4673 2694 4693 2714
rect 4790 2694 4810 2714
rect 8528 2854 8548 2874
rect 8638 2854 8658 2874
rect 8734 2854 8754 2874
rect 8846 2854 8866 2874
rect 8942 2854 8962 2874
rect 9059 2854 9079 2874
rect 9155 2854 9175 2874
rect 4886 2694 4906 2714
rect 5615 2639 5635 2659
rect 5711 2639 5731 2659
rect 5828 2639 5848 2659
rect 5924 2639 5944 2659
rect 6036 2639 6056 2659
rect 6132 2639 6152 2659
rect 6242 2639 6262 2659
rect 9444 2673 9464 2693
rect 6338 2639 6358 2659
rect 9540 2673 9560 2693
rect 9650 2673 9670 2693
rect 9746 2673 9766 2693
rect 9858 2673 9878 2693
rect 9954 2673 9974 2693
rect 10071 2673 10091 2693
rect 10167 2673 10187 2693
rect 1562 2382 1582 2402
rect 1658 2382 1678 2402
rect 1775 2382 1795 2402
rect 1871 2382 1891 2402
rect 1983 2382 2003 2402
rect 2079 2382 2099 2402
rect 2189 2382 2209 2402
rect 2285 2382 2305 2402
rect 2943 2408 2963 2428
rect 3039 2408 3059 2428
rect 3149 2408 3169 2428
rect 3245 2408 3265 2428
rect 3357 2408 3377 2428
rect 3453 2408 3473 2428
rect 3570 2408 3590 2428
rect 3666 2408 3686 2428
rect 6843 2361 6863 2381
rect 6939 2361 6959 2381
rect 7056 2361 7076 2381
rect 7152 2361 7172 2381
rect 7264 2361 7284 2381
rect 7360 2361 7380 2381
rect 7470 2361 7490 2381
rect 7566 2361 7586 2381
rect 8224 2387 8244 2407
rect 8320 2387 8340 2407
rect 8430 2387 8450 2407
rect 8526 2387 8546 2407
rect 8638 2387 8658 2407
rect 8734 2387 8754 2407
rect 8851 2387 8871 2407
rect 8947 2387 8967 2407
rect 342 2096 362 2116
rect 438 2096 458 2116
rect 555 2096 575 2116
rect 651 2096 671 2116
rect 763 2096 783 2116
rect 859 2096 879 2116
rect 969 2096 989 2116
rect 4171 2130 4191 2150
rect 1065 2096 1085 2116
rect 4267 2130 4287 2150
rect 4377 2130 4397 2150
rect 4473 2130 4493 2150
rect 4585 2130 4605 2150
rect 4681 2130 4701 2150
rect 4798 2130 4818 2150
rect 4894 2130 4914 2150
rect 5623 2075 5643 2095
rect 1354 1915 1374 1935
rect 1450 1915 1470 1935
rect 1567 1915 1587 1935
rect 1663 1915 1683 1935
rect 1775 1915 1795 1935
rect 1871 1915 1891 1935
rect 1981 1915 2001 1935
rect 5719 2075 5739 2095
rect 5836 2075 5856 2095
rect 5932 2075 5952 2095
rect 6044 2075 6064 2095
rect 6140 2075 6160 2095
rect 6250 2075 6270 2095
rect 9452 2109 9472 2129
rect 6346 2075 6366 2095
rect 9548 2109 9568 2129
rect 9658 2109 9678 2129
rect 9754 2109 9774 2129
rect 9866 2109 9886 2129
rect 9962 2109 9982 2129
rect 10079 2109 10099 2129
rect 10175 2109 10195 2129
rect 2077 1915 2097 1935
rect 3158 1896 3178 1916
rect 3254 1896 3274 1916
rect 3364 1896 3384 1916
rect 3460 1896 3480 1916
rect 3572 1896 3592 1916
rect 3668 1896 3688 1916
rect 3785 1896 3805 1916
rect 3881 1896 3901 1916
rect 6635 1894 6655 1914
rect 6731 1894 6751 1914
rect 6848 1894 6868 1914
rect 6944 1894 6964 1914
rect 7056 1894 7076 1914
rect 7152 1894 7172 1914
rect 7262 1894 7282 1914
rect 7358 1894 7378 1914
rect 8439 1875 8459 1895
rect 341 1681 361 1701
rect 437 1681 457 1701
rect 554 1681 574 1701
rect 650 1681 670 1701
rect 762 1681 782 1701
rect 858 1681 878 1701
rect 968 1681 988 1701
rect 4170 1715 4190 1735
rect 1064 1681 1084 1701
rect 4266 1715 4286 1735
rect 4376 1715 4396 1735
rect 4472 1715 4492 1735
rect 4584 1715 4604 1735
rect 4680 1715 4700 1735
rect 4797 1715 4817 1735
rect 8535 1875 8555 1895
rect 8645 1875 8665 1895
rect 8741 1875 8761 1895
rect 8853 1875 8873 1895
rect 8949 1875 8969 1895
rect 9066 1875 9086 1895
rect 9162 1875 9182 1895
rect 4893 1715 4913 1735
rect 5622 1660 5642 1680
rect 5718 1660 5738 1680
rect 5835 1660 5855 1680
rect 5931 1660 5951 1680
rect 6043 1660 6063 1680
rect 6139 1660 6159 1680
rect 6249 1660 6269 1680
rect 9451 1694 9471 1714
rect 6345 1660 6365 1680
rect 9547 1694 9567 1714
rect 9657 1694 9677 1714
rect 9753 1694 9773 1714
rect 9865 1694 9885 1714
rect 9961 1694 9981 1714
rect 10078 1694 10098 1714
rect 10174 1694 10194 1714
rect 3108 1476 3128 1496
rect 3204 1476 3224 1496
rect 3314 1476 3334 1496
rect 3410 1476 3430 1496
rect 3522 1476 3542 1496
rect 3618 1476 3638 1496
rect 3735 1476 3755 1496
rect 3831 1476 3851 1496
rect 8389 1455 8409 1475
rect 8485 1455 8505 1475
rect 8595 1455 8615 1475
rect 8691 1455 8711 1475
rect 8803 1455 8823 1475
rect 8899 1455 8919 1475
rect 9016 1455 9036 1475
rect 9112 1455 9132 1475
rect 1409 1354 1429 1374
rect 1505 1354 1525 1374
rect 1622 1354 1642 1374
rect 1718 1354 1738 1374
rect 1830 1354 1850 1374
rect 1926 1354 1946 1374
rect 2036 1354 2056 1374
rect 2132 1354 2152 1374
rect 6690 1333 6710 1353
rect 6786 1333 6806 1353
rect 6903 1333 6923 1353
rect 6999 1333 7019 1353
rect 7111 1333 7131 1353
rect 7207 1333 7227 1353
rect 7317 1333 7337 1353
rect 7413 1333 7433 1353
rect 347 1115 367 1135
rect 443 1115 463 1135
rect 560 1115 580 1135
rect 656 1115 676 1135
rect 768 1115 788 1135
rect 864 1115 884 1135
rect 974 1115 994 1135
rect 4176 1149 4196 1169
rect 1070 1115 1090 1135
rect 4272 1149 4292 1169
rect 4382 1149 4402 1169
rect 4478 1149 4498 1169
rect 4590 1149 4610 1169
rect 4686 1149 4706 1169
rect 4803 1149 4823 1169
rect 4899 1149 4919 1169
rect 5628 1094 5648 1114
rect 1359 934 1379 954
rect 1455 934 1475 954
rect 1572 934 1592 954
rect 1668 934 1688 954
rect 1780 934 1800 954
rect 1876 934 1896 954
rect 1986 934 2006 954
rect 5724 1094 5744 1114
rect 5841 1094 5861 1114
rect 5937 1094 5957 1114
rect 6049 1094 6069 1114
rect 6145 1094 6165 1114
rect 6255 1094 6275 1114
rect 9457 1128 9477 1148
rect 6351 1094 6371 1114
rect 9553 1128 9573 1148
rect 9663 1128 9683 1148
rect 9759 1128 9779 1148
rect 9871 1128 9891 1148
rect 9967 1128 9987 1148
rect 10084 1128 10104 1148
rect 10180 1128 10200 1148
rect 2082 934 2102 954
rect 3163 915 3183 935
rect 3259 915 3279 935
rect 3369 915 3389 935
rect 3465 915 3485 935
rect 3577 915 3597 935
rect 3673 915 3693 935
rect 3790 915 3810 935
rect 3886 915 3906 935
rect 6640 913 6660 933
rect 6736 913 6756 933
rect 6853 913 6873 933
rect 6949 913 6969 933
rect 7061 913 7081 933
rect 7157 913 7177 933
rect 7267 913 7287 933
rect 7363 913 7383 933
rect 8444 894 8464 914
rect 346 700 366 720
rect 442 700 462 720
rect 559 700 579 720
rect 655 700 675 720
rect 767 700 787 720
rect 863 700 883 720
rect 973 700 993 720
rect 4175 734 4195 754
rect 1069 700 1089 720
rect 4271 734 4291 754
rect 4381 734 4401 754
rect 4477 734 4497 754
rect 4589 734 4609 754
rect 4685 734 4705 754
rect 4802 734 4822 754
rect 8540 894 8560 914
rect 8650 894 8670 914
rect 8746 894 8766 914
rect 8858 894 8878 914
rect 8954 894 8974 914
rect 9071 894 9091 914
rect 9167 894 9187 914
rect 4898 734 4918 754
rect 5627 679 5647 699
rect 5723 679 5743 699
rect 5840 679 5860 699
rect 5936 679 5956 699
rect 6048 679 6068 699
rect 6144 679 6164 699
rect 6254 679 6274 699
rect 9456 713 9476 733
rect 6350 679 6370 699
rect 9552 713 9572 733
rect 9662 713 9682 733
rect 9758 713 9778 733
rect 9870 713 9890 733
rect 9966 713 9986 733
rect 10083 713 10103 733
rect 10179 713 10199 733
rect 1749 219 1769 239
rect 1845 219 1865 239
rect 1962 219 1982 239
rect 2058 219 2078 239
rect 2170 219 2190 239
rect 2266 219 2286 239
rect 2376 219 2396 239
rect 2472 219 2492 239
rect 7030 198 7050 218
rect 4839 131 4859 151
rect 4935 131 4955 151
rect 5052 131 5072 151
rect 5148 131 5168 151
rect 5260 131 5280 151
rect 5356 131 5376 151
rect 5466 131 5486 151
rect 7126 198 7146 218
rect 7243 198 7263 218
rect 7339 198 7359 218
rect 7451 198 7471 218
rect 7547 198 7567 218
rect 7657 198 7677 218
rect 7753 198 7773 218
rect 5562 131 5582 151
<< poly >>
rect 4171 8188 4221 8204
rect 4379 8188 4429 8204
rect 4587 8188 4637 8204
rect 4800 8188 4850 8204
rect 4171 8121 4221 8146
rect 4171 8095 4177 8121
rect 4203 8095 4221 8121
rect 4171 8069 4221 8095
rect 4379 8117 4429 8146
rect 4379 8093 4393 8117
rect 4417 8093 4429 8117
rect 4379 8069 4429 8093
rect 4587 8122 4637 8146
rect 4587 8098 4602 8122
rect 4626 8098 4637 8122
rect 4587 8069 4637 8098
rect 4800 8117 4850 8146
rect 9452 8167 9502 8183
rect 9660 8167 9710 8183
rect 9868 8167 9918 8183
rect 10081 8167 10131 8183
rect 4800 8097 4817 8117
rect 4837 8097 4850 8117
rect 4800 8069 4850 8097
rect 342 8031 392 8044
rect 555 8031 605 8044
rect 763 8031 813 8044
rect 971 8031 1021 8044
rect 3158 7954 3208 7970
rect 3366 7954 3416 7970
rect 3574 7954 3624 7970
rect 3787 7954 3837 7970
rect 9452 8100 9502 8125
rect 9452 8074 9458 8100
rect 9484 8074 9502 8100
rect 9452 8048 9502 8074
rect 9660 8096 9710 8125
rect 9660 8072 9674 8096
rect 9698 8072 9710 8096
rect 9660 8048 9710 8072
rect 9868 8101 9918 8125
rect 9868 8077 9883 8101
rect 9907 8077 9918 8101
rect 9868 8048 9918 8077
rect 10081 8096 10131 8125
rect 10081 8076 10098 8096
rect 10118 8076 10131 8096
rect 10081 8048 10131 8076
rect 5623 8010 5673 8023
rect 5836 8010 5886 8023
rect 6044 8010 6094 8023
rect 6252 8010 6302 8023
rect 4171 7956 4221 7969
rect 4379 7956 4429 7969
rect 4587 7956 4637 7969
rect 4800 7956 4850 7969
rect 342 7903 392 7931
rect 342 7883 355 7903
rect 375 7883 392 7903
rect 342 7854 392 7883
rect 555 7902 605 7931
rect 555 7878 566 7902
rect 590 7878 605 7902
rect 555 7854 605 7878
rect 763 7907 813 7931
rect 763 7883 775 7907
rect 799 7883 813 7907
rect 763 7854 813 7883
rect 971 7905 1021 7931
rect 971 7879 989 7905
rect 1015 7879 1021 7905
rect 971 7854 1021 7879
rect 3158 7887 3208 7912
rect 1354 7850 1404 7863
rect 1567 7850 1617 7863
rect 1775 7850 1825 7863
rect 1983 7850 2033 7863
rect 3158 7861 3164 7887
rect 3190 7861 3208 7887
rect 342 7796 392 7812
rect 555 7796 605 7812
rect 763 7796 813 7812
rect 971 7796 1021 7812
rect 3158 7835 3208 7861
rect 3366 7883 3416 7912
rect 3366 7859 3380 7883
rect 3404 7859 3416 7883
rect 3366 7835 3416 7859
rect 3574 7888 3624 7912
rect 3574 7864 3589 7888
rect 3613 7864 3624 7888
rect 3574 7835 3624 7864
rect 3787 7883 3837 7912
rect 3787 7863 3804 7883
rect 3824 7863 3837 7883
rect 3787 7835 3837 7863
rect 8439 7933 8489 7949
rect 8647 7933 8697 7949
rect 8855 7933 8905 7949
rect 9068 7933 9118 7949
rect 9452 7935 9502 7948
rect 9660 7935 9710 7948
rect 9868 7935 9918 7948
rect 10081 7935 10131 7948
rect 5623 7882 5673 7910
rect 5623 7862 5636 7882
rect 5656 7862 5673 7882
rect 1354 7722 1404 7750
rect 1354 7702 1367 7722
rect 1387 7702 1404 7722
rect 1354 7673 1404 7702
rect 1567 7721 1617 7750
rect 1567 7697 1578 7721
rect 1602 7697 1617 7721
rect 1567 7673 1617 7697
rect 1775 7726 1825 7750
rect 1775 7702 1787 7726
rect 1811 7702 1825 7726
rect 1775 7673 1825 7702
rect 1983 7724 2033 7750
rect 5623 7833 5673 7862
rect 5836 7881 5886 7910
rect 5836 7857 5847 7881
rect 5871 7857 5886 7881
rect 5836 7833 5886 7857
rect 6044 7886 6094 7910
rect 6044 7862 6056 7886
rect 6080 7862 6094 7886
rect 6044 7833 6094 7862
rect 6252 7884 6302 7910
rect 6252 7858 6270 7884
rect 6296 7858 6302 7884
rect 6252 7833 6302 7858
rect 8439 7866 8489 7891
rect 6635 7829 6685 7842
rect 6848 7829 6898 7842
rect 7056 7829 7106 7842
rect 7264 7829 7314 7842
rect 8439 7840 8445 7866
rect 8471 7840 8489 7866
rect 4170 7773 4220 7789
rect 4378 7773 4428 7789
rect 4586 7773 4636 7789
rect 4799 7773 4849 7789
rect 5623 7775 5673 7791
rect 5836 7775 5886 7791
rect 6044 7775 6094 7791
rect 6252 7775 6302 7791
rect 1983 7698 2001 7724
rect 2027 7698 2033 7724
rect 3158 7722 3208 7735
rect 3366 7722 3416 7735
rect 3574 7722 3624 7735
rect 3787 7722 3837 7735
rect 1983 7673 2033 7698
rect 4170 7706 4220 7731
rect 4170 7680 4176 7706
rect 4202 7680 4220 7706
rect 4170 7654 4220 7680
rect 4378 7702 4428 7731
rect 4378 7678 4392 7702
rect 4416 7678 4428 7702
rect 4378 7654 4428 7678
rect 4586 7707 4636 7731
rect 4586 7683 4601 7707
rect 4625 7683 4636 7707
rect 4586 7654 4636 7683
rect 4799 7702 4849 7731
rect 8439 7814 8489 7840
rect 8647 7862 8697 7891
rect 8647 7838 8661 7862
rect 8685 7838 8697 7862
rect 8647 7814 8697 7838
rect 8855 7867 8905 7891
rect 8855 7843 8870 7867
rect 8894 7843 8905 7867
rect 8855 7814 8905 7843
rect 9068 7862 9118 7891
rect 9068 7842 9085 7862
rect 9105 7842 9118 7862
rect 9068 7814 9118 7842
rect 4799 7682 4816 7702
rect 4836 7682 4849 7702
rect 4799 7654 4849 7682
rect 341 7616 391 7629
rect 554 7616 604 7629
rect 762 7616 812 7629
rect 970 7616 1020 7629
rect 1354 7615 1404 7631
rect 1567 7615 1617 7631
rect 1775 7615 1825 7631
rect 1983 7615 2033 7631
rect 6635 7701 6685 7729
rect 6635 7681 6648 7701
rect 6668 7681 6685 7701
rect 6635 7652 6685 7681
rect 6848 7700 6898 7729
rect 6848 7676 6859 7700
rect 6883 7676 6898 7700
rect 6848 7652 6898 7676
rect 7056 7705 7106 7729
rect 7056 7681 7068 7705
rect 7092 7681 7106 7705
rect 7056 7652 7106 7681
rect 7264 7703 7314 7729
rect 9451 7752 9501 7768
rect 9659 7752 9709 7768
rect 9867 7752 9917 7768
rect 10080 7752 10130 7768
rect 7264 7677 7282 7703
rect 7308 7677 7314 7703
rect 8439 7701 8489 7714
rect 8647 7701 8697 7714
rect 8855 7701 8905 7714
rect 9068 7701 9118 7714
rect 7264 7652 7314 7677
rect 9451 7685 9501 7710
rect 9451 7659 9457 7685
rect 9483 7659 9501 7685
rect 9451 7633 9501 7659
rect 9659 7681 9709 7710
rect 9659 7657 9673 7681
rect 9697 7657 9709 7681
rect 9659 7633 9709 7657
rect 9867 7686 9917 7710
rect 9867 7662 9882 7686
rect 9906 7662 9917 7686
rect 9867 7633 9917 7662
rect 10080 7681 10130 7710
rect 10080 7661 10097 7681
rect 10117 7661 10130 7681
rect 10080 7633 10130 7661
rect 5622 7595 5672 7608
rect 5835 7595 5885 7608
rect 6043 7595 6093 7608
rect 6251 7595 6301 7608
rect 3108 7534 3158 7550
rect 3316 7534 3366 7550
rect 3524 7534 3574 7550
rect 3737 7534 3787 7550
rect 4170 7541 4220 7554
rect 4378 7541 4428 7554
rect 4586 7541 4636 7554
rect 4799 7541 4849 7554
rect 341 7488 391 7516
rect 341 7468 354 7488
rect 374 7468 391 7488
rect 341 7439 391 7468
rect 554 7487 604 7516
rect 554 7463 565 7487
rect 589 7463 604 7487
rect 554 7439 604 7463
rect 762 7492 812 7516
rect 762 7468 774 7492
rect 798 7468 812 7492
rect 762 7439 812 7468
rect 970 7490 1020 7516
rect 970 7464 988 7490
rect 1014 7464 1020 7490
rect 970 7439 1020 7464
rect 3108 7467 3158 7492
rect 3108 7441 3114 7467
rect 3140 7441 3158 7467
rect 3108 7415 3158 7441
rect 3316 7463 3366 7492
rect 3316 7439 3330 7463
rect 3354 7439 3366 7463
rect 3316 7415 3366 7439
rect 3524 7468 3574 7492
rect 3524 7444 3539 7468
rect 3563 7444 3574 7468
rect 3524 7415 3574 7444
rect 3737 7463 3787 7492
rect 3737 7443 3754 7463
rect 3774 7443 3787 7463
rect 3737 7415 3787 7443
rect 6635 7594 6685 7610
rect 6848 7594 6898 7610
rect 7056 7594 7106 7610
rect 7264 7594 7314 7610
rect 8389 7513 8439 7529
rect 8597 7513 8647 7529
rect 8805 7513 8855 7529
rect 9018 7513 9068 7529
rect 9451 7520 9501 7533
rect 9659 7520 9709 7533
rect 9867 7520 9917 7533
rect 10080 7520 10130 7533
rect 5622 7467 5672 7495
rect 341 7381 391 7397
rect 554 7381 604 7397
rect 762 7381 812 7397
rect 970 7381 1020 7397
rect 5622 7447 5635 7467
rect 5655 7447 5672 7467
rect 5622 7418 5672 7447
rect 5835 7466 5885 7495
rect 5835 7442 5846 7466
rect 5870 7442 5885 7466
rect 5835 7418 5885 7442
rect 6043 7471 6093 7495
rect 6043 7447 6055 7471
rect 6079 7447 6093 7471
rect 6043 7418 6093 7447
rect 6251 7469 6301 7495
rect 6251 7443 6269 7469
rect 6295 7443 6301 7469
rect 6251 7418 6301 7443
rect 8389 7446 8439 7471
rect 8389 7420 8395 7446
rect 8421 7420 8439 7446
rect 8389 7394 8439 7420
rect 8597 7442 8647 7471
rect 8597 7418 8611 7442
rect 8635 7418 8647 7442
rect 8597 7394 8647 7418
rect 8805 7447 8855 7471
rect 8805 7423 8820 7447
rect 8844 7423 8855 7447
rect 8805 7394 8855 7423
rect 9018 7442 9068 7471
rect 9018 7422 9035 7442
rect 9055 7422 9068 7442
rect 9018 7394 9068 7422
rect 5622 7360 5672 7376
rect 5835 7360 5885 7376
rect 6043 7360 6093 7376
rect 6251 7360 6301 7376
rect 3108 7302 3158 7315
rect 3316 7302 3366 7315
rect 3524 7302 3574 7315
rect 3737 7302 3787 7315
rect 1409 7289 1459 7302
rect 1622 7289 1672 7302
rect 1830 7289 1880 7302
rect 2038 7289 2088 7302
rect 8389 7281 8439 7294
rect 8597 7281 8647 7294
rect 8805 7281 8855 7294
rect 9018 7281 9068 7294
rect 6690 7268 6740 7281
rect 6903 7268 6953 7281
rect 7111 7268 7161 7281
rect 7319 7268 7369 7281
rect 4176 7207 4226 7223
rect 4384 7207 4434 7223
rect 4592 7207 4642 7223
rect 4805 7207 4855 7223
rect 1409 7161 1459 7189
rect 1409 7141 1422 7161
rect 1442 7141 1459 7161
rect 1409 7112 1459 7141
rect 1622 7160 1672 7189
rect 1622 7136 1633 7160
rect 1657 7136 1672 7160
rect 1622 7112 1672 7136
rect 1830 7165 1880 7189
rect 1830 7141 1842 7165
rect 1866 7141 1880 7165
rect 1830 7112 1880 7141
rect 2038 7163 2088 7189
rect 2038 7137 2056 7163
rect 2082 7137 2088 7163
rect 2038 7112 2088 7137
rect 4176 7140 4226 7165
rect 4176 7114 4182 7140
rect 4208 7114 4226 7140
rect 4176 7088 4226 7114
rect 4384 7136 4434 7165
rect 4384 7112 4398 7136
rect 4422 7112 4434 7136
rect 4384 7088 4434 7112
rect 4592 7141 4642 7165
rect 4592 7117 4607 7141
rect 4631 7117 4642 7141
rect 4592 7088 4642 7117
rect 4805 7136 4855 7165
rect 4805 7116 4822 7136
rect 4842 7116 4855 7136
rect 9457 7186 9507 7202
rect 9665 7186 9715 7202
rect 9873 7186 9923 7202
rect 10086 7186 10136 7202
rect 4805 7088 4855 7116
rect 347 7050 397 7063
rect 560 7050 610 7063
rect 768 7050 818 7063
rect 976 7050 1026 7063
rect 1409 7054 1459 7070
rect 1622 7054 1672 7070
rect 1830 7054 1880 7070
rect 2038 7054 2088 7070
rect 3163 6973 3213 6989
rect 3371 6973 3421 6989
rect 3579 6973 3629 6989
rect 3792 6973 3842 6989
rect 6690 7140 6740 7168
rect 6690 7120 6703 7140
rect 6723 7120 6740 7140
rect 6690 7091 6740 7120
rect 6903 7139 6953 7168
rect 6903 7115 6914 7139
rect 6938 7115 6953 7139
rect 6903 7091 6953 7115
rect 7111 7144 7161 7168
rect 7111 7120 7123 7144
rect 7147 7120 7161 7144
rect 7111 7091 7161 7120
rect 7319 7142 7369 7168
rect 7319 7116 7337 7142
rect 7363 7116 7369 7142
rect 7319 7091 7369 7116
rect 9457 7119 9507 7144
rect 9457 7093 9463 7119
rect 9489 7093 9507 7119
rect 9457 7067 9507 7093
rect 9665 7115 9715 7144
rect 9665 7091 9679 7115
rect 9703 7091 9715 7115
rect 9665 7067 9715 7091
rect 9873 7120 9923 7144
rect 9873 7096 9888 7120
rect 9912 7096 9923 7120
rect 9873 7067 9923 7096
rect 10086 7115 10136 7144
rect 10086 7095 10103 7115
rect 10123 7095 10136 7115
rect 10086 7067 10136 7095
rect 5628 7029 5678 7042
rect 5841 7029 5891 7042
rect 6049 7029 6099 7042
rect 6257 7029 6307 7042
rect 6690 7033 6740 7049
rect 6903 7033 6953 7049
rect 7111 7033 7161 7049
rect 7319 7033 7369 7049
rect 4176 6975 4226 6988
rect 4384 6975 4434 6988
rect 4592 6975 4642 6988
rect 4805 6975 4855 6988
rect 347 6922 397 6950
rect 347 6902 360 6922
rect 380 6902 397 6922
rect 347 6873 397 6902
rect 560 6921 610 6950
rect 560 6897 571 6921
rect 595 6897 610 6921
rect 560 6873 610 6897
rect 768 6926 818 6950
rect 768 6902 780 6926
rect 804 6902 818 6926
rect 768 6873 818 6902
rect 976 6924 1026 6950
rect 976 6898 994 6924
rect 1020 6898 1026 6924
rect 976 6873 1026 6898
rect 3163 6906 3213 6931
rect 1359 6869 1409 6882
rect 1572 6869 1622 6882
rect 1780 6869 1830 6882
rect 1988 6869 2038 6882
rect 3163 6880 3169 6906
rect 3195 6880 3213 6906
rect 347 6815 397 6831
rect 560 6815 610 6831
rect 768 6815 818 6831
rect 976 6815 1026 6831
rect 3163 6854 3213 6880
rect 3371 6902 3421 6931
rect 3371 6878 3385 6902
rect 3409 6878 3421 6902
rect 3371 6854 3421 6878
rect 3579 6907 3629 6931
rect 3579 6883 3594 6907
rect 3618 6883 3629 6907
rect 3579 6854 3629 6883
rect 3792 6902 3842 6931
rect 3792 6882 3809 6902
rect 3829 6882 3842 6902
rect 3792 6854 3842 6882
rect 8444 6952 8494 6968
rect 8652 6952 8702 6968
rect 8860 6952 8910 6968
rect 9073 6952 9123 6968
rect 9457 6954 9507 6967
rect 9665 6954 9715 6967
rect 9873 6954 9923 6967
rect 10086 6954 10136 6967
rect 5628 6901 5678 6929
rect 5628 6881 5641 6901
rect 5661 6881 5678 6901
rect 1359 6741 1409 6769
rect 1359 6721 1372 6741
rect 1392 6721 1409 6741
rect 1359 6692 1409 6721
rect 1572 6740 1622 6769
rect 1572 6716 1583 6740
rect 1607 6716 1622 6740
rect 1572 6692 1622 6716
rect 1780 6745 1830 6769
rect 1780 6721 1792 6745
rect 1816 6721 1830 6745
rect 1780 6692 1830 6721
rect 1988 6743 2038 6769
rect 5628 6852 5678 6881
rect 5841 6900 5891 6929
rect 5841 6876 5852 6900
rect 5876 6876 5891 6900
rect 5841 6852 5891 6876
rect 6049 6905 6099 6929
rect 6049 6881 6061 6905
rect 6085 6881 6099 6905
rect 6049 6852 6099 6881
rect 6257 6903 6307 6929
rect 6257 6877 6275 6903
rect 6301 6877 6307 6903
rect 6257 6852 6307 6877
rect 8444 6885 8494 6910
rect 6640 6848 6690 6861
rect 6853 6848 6903 6861
rect 7061 6848 7111 6861
rect 7269 6848 7319 6861
rect 8444 6859 8450 6885
rect 8476 6859 8494 6885
rect 4175 6792 4225 6808
rect 4383 6792 4433 6808
rect 4591 6792 4641 6808
rect 4804 6792 4854 6808
rect 5628 6794 5678 6810
rect 5841 6794 5891 6810
rect 6049 6794 6099 6810
rect 6257 6794 6307 6810
rect 1988 6717 2006 6743
rect 2032 6717 2038 6743
rect 3163 6741 3213 6754
rect 3371 6741 3421 6754
rect 3579 6741 3629 6754
rect 3792 6741 3842 6754
rect 1988 6692 2038 6717
rect 4175 6725 4225 6750
rect 4175 6699 4181 6725
rect 4207 6699 4225 6725
rect 4175 6673 4225 6699
rect 4383 6721 4433 6750
rect 4383 6697 4397 6721
rect 4421 6697 4433 6721
rect 4383 6673 4433 6697
rect 4591 6726 4641 6750
rect 4591 6702 4606 6726
rect 4630 6702 4641 6726
rect 4591 6673 4641 6702
rect 4804 6721 4854 6750
rect 8444 6833 8494 6859
rect 8652 6881 8702 6910
rect 8652 6857 8666 6881
rect 8690 6857 8702 6881
rect 8652 6833 8702 6857
rect 8860 6886 8910 6910
rect 8860 6862 8875 6886
rect 8899 6862 8910 6886
rect 8860 6833 8910 6862
rect 9073 6881 9123 6910
rect 9073 6861 9090 6881
rect 9110 6861 9123 6881
rect 9073 6833 9123 6861
rect 4804 6701 4821 6721
rect 4841 6701 4854 6721
rect 4804 6673 4854 6701
rect 346 6635 396 6648
rect 559 6635 609 6648
rect 767 6635 817 6648
rect 975 6635 1025 6648
rect 1359 6634 1409 6650
rect 1572 6634 1622 6650
rect 1780 6634 1830 6650
rect 1988 6634 2038 6650
rect 6640 6720 6690 6748
rect 6640 6700 6653 6720
rect 6673 6700 6690 6720
rect 6640 6671 6690 6700
rect 6853 6719 6903 6748
rect 6853 6695 6864 6719
rect 6888 6695 6903 6719
rect 6853 6671 6903 6695
rect 7061 6724 7111 6748
rect 7061 6700 7073 6724
rect 7097 6700 7111 6724
rect 7061 6671 7111 6700
rect 7269 6722 7319 6748
rect 9456 6771 9506 6787
rect 9664 6771 9714 6787
rect 9872 6771 9922 6787
rect 10085 6771 10135 6787
rect 7269 6696 7287 6722
rect 7313 6696 7319 6722
rect 8444 6720 8494 6733
rect 8652 6720 8702 6733
rect 8860 6720 8910 6733
rect 9073 6720 9123 6733
rect 7269 6671 7319 6696
rect 9456 6704 9506 6729
rect 9456 6678 9462 6704
rect 9488 6678 9506 6704
rect 9456 6652 9506 6678
rect 9664 6700 9714 6729
rect 9664 6676 9678 6700
rect 9702 6676 9714 6700
rect 9664 6652 9714 6676
rect 9872 6705 9922 6729
rect 9872 6681 9887 6705
rect 9911 6681 9922 6705
rect 9872 6652 9922 6681
rect 10085 6700 10135 6729
rect 10085 6680 10102 6700
rect 10122 6680 10135 6700
rect 10085 6652 10135 6680
rect 5627 6614 5677 6627
rect 5840 6614 5890 6627
rect 6048 6614 6098 6627
rect 6256 6614 6306 6627
rect 4175 6560 4225 6573
rect 4383 6560 4433 6573
rect 4591 6560 4641 6573
rect 4804 6560 4854 6573
rect 346 6507 396 6535
rect 346 6487 359 6507
rect 379 6487 396 6507
rect 346 6458 396 6487
rect 559 6506 609 6535
rect 559 6482 570 6506
rect 594 6482 609 6506
rect 559 6458 609 6482
rect 767 6511 817 6535
rect 767 6487 779 6511
rect 803 6487 817 6511
rect 767 6458 817 6487
rect 975 6509 1025 6535
rect 975 6483 993 6509
rect 1019 6483 1025 6509
rect 2955 6506 3005 6522
rect 3163 6506 3213 6522
rect 3371 6506 3421 6522
rect 3584 6506 3634 6522
rect 975 6458 1025 6483
rect 6640 6613 6690 6629
rect 6853 6613 6903 6629
rect 7061 6613 7111 6629
rect 7269 6613 7319 6629
rect 9456 6539 9506 6552
rect 9664 6539 9714 6552
rect 9872 6539 9922 6552
rect 10085 6539 10135 6552
rect 2955 6439 3005 6464
rect 346 6400 396 6416
rect 559 6400 609 6416
rect 767 6400 817 6416
rect 975 6400 1025 6416
rect 2955 6413 2961 6439
rect 2987 6413 3005 6439
rect 2955 6387 3005 6413
rect 3163 6435 3213 6464
rect 3163 6411 3177 6435
rect 3201 6411 3213 6435
rect 3163 6387 3213 6411
rect 3371 6440 3421 6464
rect 3371 6416 3386 6440
rect 3410 6416 3421 6440
rect 3371 6387 3421 6416
rect 3584 6435 3634 6464
rect 5627 6486 5677 6514
rect 3584 6415 3601 6435
rect 3621 6415 3634 6435
rect 5627 6466 5640 6486
rect 5660 6466 5677 6486
rect 3584 6387 3634 6415
rect 5627 6437 5677 6466
rect 5840 6485 5890 6514
rect 5840 6461 5851 6485
rect 5875 6461 5890 6485
rect 5840 6437 5890 6461
rect 6048 6490 6098 6514
rect 6048 6466 6060 6490
rect 6084 6466 6098 6490
rect 6048 6437 6098 6466
rect 6256 6488 6306 6514
rect 6256 6462 6274 6488
rect 6300 6462 6306 6488
rect 8236 6485 8286 6501
rect 8444 6485 8494 6501
rect 8652 6485 8702 6501
rect 8865 6485 8915 6501
rect 6256 6437 6306 6462
rect 1574 6357 1624 6370
rect 1787 6357 1837 6370
rect 1995 6357 2045 6370
rect 2203 6357 2253 6370
rect 8236 6418 8286 6443
rect 5627 6379 5677 6395
rect 5840 6379 5890 6395
rect 6048 6379 6098 6395
rect 6256 6379 6306 6395
rect 8236 6392 8242 6418
rect 8268 6392 8286 6418
rect 8236 6366 8286 6392
rect 8444 6414 8494 6443
rect 8444 6390 8458 6414
rect 8482 6390 8494 6414
rect 8444 6366 8494 6390
rect 8652 6419 8702 6443
rect 8652 6395 8667 6419
rect 8691 6395 8702 6419
rect 8652 6366 8702 6395
rect 8865 6414 8915 6443
rect 8865 6394 8882 6414
rect 8902 6394 8915 6414
rect 8865 6366 8915 6394
rect 6855 6336 6905 6349
rect 7068 6336 7118 6349
rect 7276 6336 7326 6349
rect 7484 6336 7534 6349
rect 2955 6274 3005 6287
rect 3163 6274 3213 6287
rect 3371 6274 3421 6287
rect 3584 6274 3634 6287
rect 1574 6229 1624 6257
rect 1574 6209 1587 6229
rect 1607 6209 1624 6229
rect 1574 6180 1624 6209
rect 1787 6228 1837 6257
rect 1787 6204 1798 6228
rect 1822 6204 1837 6228
rect 1787 6180 1837 6204
rect 1995 6233 2045 6257
rect 1995 6209 2007 6233
rect 2031 6209 2045 6233
rect 1995 6180 2045 6209
rect 2203 6231 2253 6257
rect 2203 6205 2221 6231
rect 2247 6205 2253 6231
rect 4183 6228 4233 6244
rect 4391 6228 4441 6244
rect 4599 6228 4649 6244
rect 4812 6228 4862 6244
rect 2203 6180 2253 6205
rect 8236 6253 8286 6266
rect 8444 6253 8494 6266
rect 8652 6253 8702 6266
rect 8865 6253 8915 6266
rect 4183 6161 4233 6186
rect 1574 6122 1624 6138
rect 1787 6122 1837 6138
rect 1995 6122 2045 6138
rect 2203 6122 2253 6138
rect 4183 6135 4189 6161
rect 4215 6135 4233 6161
rect 4183 6109 4233 6135
rect 4391 6157 4441 6186
rect 4391 6133 4405 6157
rect 4429 6133 4441 6157
rect 4391 6109 4441 6133
rect 4599 6162 4649 6186
rect 4599 6138 4614 6162
rect 4638 6138 4649 6162
rect 4599 6109 4649 6138
rect 4812 6157 4862 6186
rect 6855 6208 6905 6236
rect 4812 6137 4829 6157
rect 4849 6137 4862 6157
rect 6855 6188 6868 6208
rect 6888 6188 6905 6208
rect 4812 6109 4862 6137
rect 6855 6159 6905 6188
rect 7068 6207 7118 6236
rect 7068 6183 7079 6207
rect 7103 6183 7118 6207
rect 7068 6159 7118 6183
rect 7276 6212 7326 6236
rect 7276 6188 7288 6212
rect 7312 6188 7326 6212
rect 7276 6159 7326 6188
rect 7484 6210 7534 6236
rect 7484 6184 7502 6210
rect 7528 6184 7534 6210
rect 9464 6207 9514 6223
rect 9672 6207 9722 6223
rect 9880 6207 9930 6223
rect 10093 6207 10143 6223
rect 7484 6159 7534 6184
rect 354 6071 404 6084
rect 567 6071 617 6084
rect 775 6071 825 6084
rect 983 6071 1033 6084
rect 3170 5994 3220 6010
rect 3378 5994 3428 6010
rect 3586 5994 3636 6010
rect 3799 5994 3849 6010
rect 9464 6140 9514 6165
rect 6855 6101 6905 6117
rect 7068 6101 7118 6117
rect 7276 6101 7326 6117
rect 7484 6101 7534 6117
rect 9464 6114 9470 6140
rect 9496 6114 9514 6140
rect 9464 6088 9514 6114
rect 9672 6136 9722 6165
rect 9672 6112 9686 6136
rect 9710 6112 9722 6136
rect 9672 6088 9722 6112
rect 9880 6141 9930 6165
rect 9880 6117 9895 6141
rect 9919 6117 9930 6141
rect 9880 6088 9930 6117
rect 10093 6136 10143 6165
rect 10093 6116 10110 6136
rect 10130 6116 10143 6136
rect 10093 6088 10143 6116
rect 5635 6050 5685 6063
rect 5848 6050 5898 6063
rect 6056 6050 6106 6063
rect 6264 6050 6314 6063
rect 4183 5996 4233 6009
rect 4391 5996 4441 6009
rect 4599 5996 4649 6009
rect 4812 5996 4862 6009
rect 354 5943 404 5971
rect 354 5923 367 5943
rect 387 5923 404 5943
rect 354 5894 404 5923
rect 567 5942 617 5971
rect 567 5918 578 5942
rect 602 5918 617 5942
rect 567 5894 617 5918
rect 775 5947 825 5971
rect 775 5923 787 5947
rect 811 5923 825 5947
rect 775 5894 825 5923
rect 983 5945 1033 5971
rect 983 5919 1001 5945
rect 1027 5919 1033 5945
rect 983 5894 1033 5919
rect 3170 5927 3220 5952
rect 1366 5890 1416 5903
rect 1579 5890 1629 5903
rect 1787 5890 1837 5903
rect 1995 5890 2045 5903
rect 3170 5901 3176 5927
rect 3202 5901 3220 5927
rect 354 5836 404 5852
rect 567 5836 617 5852
rect 775 5836 825 5852
rect 983 5836 1033 5852
rect 3170 5875 3220 5901
rect 3378 5923 3428 5952
rect 3378 5899 3392 5923
rect 3416 5899 3428 5923
rect 3378 5875 3428 5899
rect 3586 5928 3636 5952
rect 3586 5904 3601 5928
rect 3625 5904 3636 5928
rect 3586 5875 3636 5904
rect 3799 5923 3849 5952
rect 3799 5903 3816 5923
rect 3836 5903 3849 5923
rect 3799 5875 3849 5903
rect 8451 5973 8501 5989
rect 8659 5973 8709 5989
rect 8867 5973 8917 5989
rect 9080 5973 9130 5989
rect 9464 5975 9514 5988
rect 9672 5975 9722 5988
rect 9880 5975 9930 5988
rect 10093 5975 10143 5988
rect 5635 5922 5685 5950
rect 5635 5902 5648 5922
rect 5668 5902 5685 5922
rect 1366 5762 1416 5790
rect 1366 5742 1379 5762
rect 1399 5742 1416 5762
rect 1366 5713 1416 5742
rect 1579 5761 1629 5790
rect 1579 5737 1590 5761
rect 1614 5737 1629 5761
rect 1579 5713 1629 5737
rect 1787 5766 1837 5790
rect 1787 5742 1799 5766
rect 1823 5742 1837 5766
rect 1787 5713 1837 5742
rect 1995 5764 2045 5790
rect 5635 5873 5685 5902
rect 5848 5921 5898 5950
rect 5848 5897 5859 5921
rect 5883 5897 5898 5921
rect 5848 5873 5898 5897
rect 6056 5926 6106 5950
rect 6056 5902 6068 5926
rect 6092 5902 6106 5926
rect 6056 5873 6106 5902
rect 6264 5924 6314 5950
rect 6264 5898 6282 5924
rect 6308 5898 6314 5924
rect 6264 5873 6314 5898
rect 8451 5906 8501 5931
rect 6647 5869 6697 5882
rect 6860 5869 6910 5882
rect 7068 5869 7118 5882
rect 7276 5869 7326 5882
rect 8451 5880 8457 5906
rect 8483 5880 8501 5906
rect 4182 5813 4232 5829
rect 4390 5813 4440 5829
rect 4598 5813 4648 5829
rect 4811 5813 4861 5829
rect 5635 5815 5685 5831
rect 5848 5815 5898 5831
rect 6056 5815 6106 5831
rect 6264 5815 6314 5831
rect 1995 5738 2013 5764
rect 2039 5738 2045 5764
rect 3170 5762 3220 5775
rect 3378 5762 3428 5775
rect 3586 5762 3636 5775
rect 3799 5762 3849 5775
rect 1995 5713 2045 5738
rect 4182 5746 4232 5771
rect 4182 5720 4188 5746
rect 4214 5720 4232 5746
rect 4182 5694 4232 5720
rect 4390 5742 4440 5771
rect 4390 5718 4404 5742
rect 4428 5718 4440 5742
rect 4390 5694 4440 5718
rect 4598 5747 4648 5771
rect 4598 5723 4613 5747
rect 4637 5723 4648 5747
rect 4598 5694 4648 5723
rect 4811 5742 4861 5771
rect 8451 5854 8501 5880
rect 8659 5902 8709 5931
rect 8659 5878 8673 5902
rect 8697 5878 8709 5902
rect 8659 5854 8709 5878
rect 8867 5907 8917 5931
rect 8867 5883 8882 5907
rect 8906 5883 8917 5907
rect 8867 5854 8917 5883
rect 9080 5902 9130 5931
rect 9080 5882 9097 5902
rect 9117 5882 9130 5902
rect 9080 5854 9130 5882
rect 4811 5722 4828 5742
rect 4848 5722 4861 5742
rect 4811 5694 4861 5722
rect 353 5656 403 5669
rect 566 5656 616 5669
rect 774 5656 824 5669
rect 982 5656 1032 5669
rect 1366 5655 1416 5671
rect 1579 5655 1629 5671
rect 1787 5655 1837 5671
rect 1995 5655 2045 5671
rect 6647 5741 6697 5769
rect 6647 5721 6660 5741
rect 6680 5721 6697 5741
rect 6647 5692 6697 5721
rect 6860 5740 6910 5769
rect 6860 5716 6871 5740
rect 6895 5716 6910 5740
rect 6860 5692 6910 5716
rect 7068 5745 7118 5769
rect 7068 5721 7080 5745
rect 7104 5721 7118 5745
rect 7068 5692 7118 5721
rect 7276 5743 7326 5769
rect 9463 5792 9513 5808
rect 9671 5792 9721 5808
rect 9879 5792 9929 5808
rect 10092 5792 10142 5808
rect 7276 5717 7294 5743
rect 7320 5717 7326 5743
rect 8451 5741 8501 5754
rect 8659 5741 8709 5754
rect 8867 5741 8917 5754
rect 9080 5741 9130 5754
rect 7276 5692 7326 5717
rect 9463 5725 9513 5750
rect 9463 5699 9469 5725
rect 9495 5699 9513 5725
rect 9463 5673 9513 5699
rect 9671 5721 9721 5750
rect 9671 5697 9685 5721
rect 9709 5697 9721 5721
rect 9671 5673 9721 5697
rect 9879 5726 9929 5750
rect 9879 5702 9894 5726
rect 9918 5702 9929 5726
rect 9879 5673 9929 5702
rect 10092 5721 10142 5750
rect 10092 5701 10109 5721
rect 10129 5701 10142 5721
rect 10092 5673 10142 5701
rect 5634 5635 5684 5648
rect 5847 5635 5897 5648
rect 6055 5635 6105 5648
rect 6263 5635 6313 5648
rect 3120 5574 3170 5590
rect 3328 5574 3378 5590
rect 3536 5574 3586 5590
rect 3749 5574 3799 5590
rect 4182 5581 4232 5594
rect 4390 5581 4440 5594
rect 4598 5581 4648 5594
rect 4811 5581 4861 5594
rect 353 5528 403 5556
rect 353 5508 366 5528
rect 386 5508 403 5528
rect 353 5479 403 5508
rect 566 5527 616 5556
rect 566 5503 577 5527
rect 601 5503 616 5527
rect 566 5479 616 5503
rect 774 5532 824 5556
rect 774 5508 786 5532
rect 810 5508 824 5532
rect 774 5479 824 5508
rect 982 5530 1032 5556
rect 982 5504 1000 5530
rect 1026 5504 1032 5530
rect 982 5479 1032 5504
rect 3120 5507 3170 5532
rect 3120 5481 3126 5507
rect 3152 5481 3170 5507
rect 3120 5455 3170 5481
rect 3328 5503 3378 5532
rect 3328 5479 3342 5503
rect 3366 5479 3378 5503
rect 3328 5455 3378 5479
rect 3536 5508 3586 5532
rect 3536 5484 3551 5508
rect 3575 5484 3586 5508
rect 3536 5455 3586 5484
rect 3749 5503 3799 5532
rect 3749 5483 3766 5503
rect 3786 5483 3799 5503
rect 3749 5455 3799 5483
rect 6647 5634 6697 5650
rect 6860 5634 6910 5650
rect 7068 5634 7118 5650
rect 7276 5634 7326 5650
rect 8401 5553 8451 5569
rect 8609 5553 8659 5569
rect 8817 5553 8867 5569
rect 9030 5553 9080 5569
rect 9463 5560 9513 5573
rect 9671 5560 9721 5573
rect 9879 5560 9929 5573
rect 10092 5560 10142 5573
rect 5634 5507 5684 5535
rect 353 5421 403 5437
rect 566 5421 616 5437
rect 774 5421 824 5437
rect 982 5421 1032 5437
rect 5634 5487 5647 5507
rect 5667 5487 5684 5507
rect 5634 5458 5684 5487
rect 5847 5506 5897 5535
rect 5847 5482 5858 5506
rect 5882 5482 5897 5506
rect 5847 5458 5897 5482
rect 6055 5511 6105 5535
rect 6055 5487 6067 5511
rect 6091 5487 6105 5511
rect 6055 5458 6105 5487
rect 6263 5509 6313 5535
rect 6263 5483 6281 5509
rect 6307 5483 6313 5509
rect 6263 5458 6313 5483
rect 8401 5486 8451 5511
rect 8401 5460 8407 5486
rect 8433 5460 8451 5486
rect 8401 5434 8451 5460
rect 8609 5482 8659 5511
rect 8609 5458 8623 5482
rect 8647 5458 8659 5482
rect 8609 5434 8659 5458
rect 8817 5487 8867 5511
rect 8817 5463 8832 5487
rect 8856 5463 8867 5487
rect 8817 5434 8867 5463
rect 9030 5482 9080 5511
rect 9030 5462 9047 5482
rect 9067 5462 9080 5482
rect 9030 5434 9080 5462
rect 5634 5400 5684 5416
rect 5847 5400 5897 5416
rect 6055 5400 6105 5416
rect 6263 5400 6313 5416
rect 3120 5342 3170 5355
rect 3328 5342 3378 5355
rect 3536 5342 3586 5355
rect 3749 5342 3799 5355
rect 1421 5329 1471 5342
rect 1634 5329 1684 5342
rect 1842 5329 1892 5342
rect 2050 5329 2100 5342
rect 8401 5321 8451 5334
rect 8609 5321 8659 5334
rect 8817 5321 8867 5334
rect 9030 5321 9080 5334
rect 6702 5308 6752 5321
rect 6915 5308 6965 5321
rect 7123 5308 7173 5321
rect 7331 5308 7381 5321
rect 4188 5247 4238 5263
rect 4396 5247 4446 5263
rect 4604 5247 4654 5263
rect 4817 5247 4867 5263
rect 1421 5201 1471 5229
rect 1421 5181 1434 5201
rect 1454 5181 1471 5201
rect 1421 5152 1471 5181
rect 1634 5200 1684 5229
rect 1634 5176 1645 5200
rect 1669 5176 1684 5200
rect 1634 5152 1684 5176
rect 1842 5205 1892 5229
rect 1842 5181 1854 5205
rect 1878 5181 1892 5205
rect 1842 5152 1892 5181
rect 2050 5203 2100 5229
rect 2050 5177 2068 5203
rect 2094 5177 2100 5203
rect 2050 5152 2100 5177
rect 4188 5180 4238 5205
rect 4188 5154 4194 5180
rect 4220 5154 4238 5180
rect 4188 5128 4238 5154
rect 4396 5176 4446 5205
rect 4396 5152 4410 5176
rect 4434 5152 4446 5176
rect 4396 5128 4446 5152
rect 4604 5181 4654 5205
rect 4604 5157 4619 5181
rect 4643 5157 4654 5181
rect 4604 5128 4654 5157
rect 4817 5176 4867 5205
rect 4817 5156 4834 5176
rect 4854 5156 4867 5176
rect 9469 5226 9519 5242
rect 9677 5226 9727 5242
rect 9885 5226 9935 5242
rect 10098 5226 10148 5242
rect 4817 5128 4867 5156
rect 359 5090 409 5103
rect 572 5090 622 5103
rect 780 5090 830 5103
rect 988 5090 1038 5103
rect 1421 5094 1471 5110
rect 1634 5094 1684 5110
rect 1842 5094 1892 5110
rect 2050 5094 2100 5110
rect 3175 5013 3225 5029
rect 3383 5013 3433 5029
rect 3591 5013 3641 5029
rect 3804 5013 3854 5029
rect 6702 5180 6752 5208
rect 6702 5160 6715 5180
rect 6735 5160 6752 5180
rect 6702 5131 6752 5160
rect 6915 5179 6965 5208
rect 6915 5155 6926 5179
rect 6950 5155 6965 5179
rect 6915 5131 6965 5155
rect 7123 5184 7173 5208
rect 7123 5160 7135 5184
rect 7159 5160 7173 5184
rect 7123 5131 7173 5160
rect 7331 5182 7381 5208
rect 7331 5156 7349 5182
rect 7375 5156 7381 5182
rect 7331 5131 7381 5156
rect 9469 5159 9519 5184
rect 9469 5133 9475 5159
rect 9501 5133 9519 5159
rect 9469 5107 9519 5133
rect 9677 5155 9727 5184
rect 9677 5131 9691 5155
rect 9715 5131 9727 5155
rect 9677 5107 9727 5131
rect 9885 5160 9935 5184
rect 9885 5136 9900 5160
rect 9924 5136 9935 5160
rect 9885 5107 9935 5136
rect 10098 5155 10148 5184
rect 10098 5135 10115 5155
rect 10135 5135 10148 5155
rect 10098 5107 10148 5135
rect 5640 5069 5690 5082
rect 5853 5069 5903 5082
rect 6061 5069 6111 5082
rect 6269 5069 6319 5082
rect 6702 5073 6752 5089
rect 6915 5073 6965 5089
rect 7123 5073 7173 5089
rect 7331 5073 7381 5089
rect 4188 5015 4238 5028
rect 4396 5015 4446 5028
rect 4604 5015 4654 5028
rect 4817 5015 4867 5028
rect 359 4962 409 4990
rect 359 4942 372 4962
rect 392 4942 409 4962
rect 359 4913 409 4942
rect 572 4961 622 4990
rect 572 4937 583 4961
rect 607 4937 622 4961
rect 572 4913 622 4937
rect 780 4966 830 4990
rect 780 4942 792 4966
rect 816 4942 830 4966
rect 780 4913 830 4942
rect 988 4964 1038 4990
rect 988 4938 1006 4964
rect 1032 4938 1038 4964
rect 988 4913 1038 4938
rect 3175 4946 3225 4971
rect 1371 4909 1421 4922
rect 1584 4909 1634 4922
rect 1792 4909 1842 4922
rect 2000 4909 2050 4922
rect 3175 4920 3181 4946
rect 3207 4920 3225 4946
rect 359 4855 409 4871
rect 572 4855 622 4871
rect 780 4855 830 4871
rect 988 4855 1038 4871
rect 3175 4894 3225 4920
rect 3383 4942 3433 4971
rect 3383 4918 3397 4942
rect 3421 4918 3433 4942
rect 3383 4894 3433 4918
rect 3591 4947 3641 4971
rect 3591 4923 3606 4947
rect 3630 4923 3641 4947
rect 3591 4894 3641 4923
rect 3804 4942 3854 4971
rect 3804 4922 3821 4942
rect 3841 4922 3854 4942
rect 3804 4894 3854 4922
rect 8456 4992 8506 5008
rect 8664 4992 8714 5008
rect 8872 4992 8922 5008
rect 9085 4992 9135 5008
rect 9469 4994 9519 5007
rect 9677 4994 9727 5007
rect 9885 4994 9935 5007
rect 10098 4994 10148 5007
rect 5640 4941 5690 4969
rect 5640 4921 5653 4941
rect 5673 4921 5690 4941
rect 1371 4781 1421 4809
rect 1371 4761 1384 4781
rect 1404 4761 1421 4781
rect 1371 4732 1421 4761
rect 1584 4780 1634 4809
rect 1584 4756 1595 4780
rect 1619 4756 1634 4780
rect 1584 4732 1634 4756
rect 1792 4785 1842 4809
rect 1792 4761 1804 4785
rect 1828 4761 1842 4785
rect 1792 4732 1842 4761
rect 2000 4783 2050 4809
rect 5640 4892 5690 4921
rect 5853 4940 5903 4969
rect 5853 4916 5864 4940
rect 5888 4916 5903 4940
rect 5853 4892 5903 4916
rect 6061 4945 6111 4969
rect 6061 4921 6073 4945
rect 6097 4921 6111 4945
rect 6061 4892 6111 4921
rect 6269 4943 6319 4969
rect 6269 4917 6287 4943
rect 6313 4917 6319 4943
rect 6269 4892 6319 4917
rect 8456 4925 8506 4950
rect 6652 4888 6702 4901
rect 6865 4888 6915 4901
rect 7073 4888 7123 4901
rect 7281 4888 7331 4901
rect 8456 4899 8462 4925
rect 8488 4899 8506 4925
rect 4187 4832 4237 4848
rect 4395 4832 4445 4848
rect 4603 4832 4653 4848
rect 4816 4832 4866 4848
rect 5640 4834 5690 4850
rect 5853 4834 5903 4850
rect 6061 4834 6111 4850
rect 6269 4834 6319 4850
rect 2000 4757 2018 4783
rect 2044 4757 2050 4783
rect 3175 4781 3225 4794
rect 3383 4781 3433 4794
rect 3591 4781 3641 4794
rect 3804 4781 3854 4794
rect 2000 4732 2050 4757
rect 4187 4765 4237 4790
rect 4187 4739 4193 4765
rect 4219 4739 4237 4765
rect 4187 4713 4237 4739
rect 4395 4761 4445 4790
rect 4395 4737 4409 4761
rect 4433 4737 4445 4761
rect 4395 4713 4445 4737
rect 4603 4766 4653 4790
rect 4603 4742 4618 4766
rect 4642 4742 4653 4766
rect 4603 4713 4653 4742
rect 4816 4761 4866 4790
rect 8456 4873 8506 4899
rect 8664 4921 8714 4950
rect 8664 4897 8678 4921
rect 8702 4897 8714 4921
rect 8664 4873 8714 4897
rect 8872 4926 8922 4950
rect 8872 4902 8887 4926
rect 8911 4902 8922 4926
rect 8872 4873 8922 4902
rect 9085 4921 9135 4950
rect 9085 4901 9102 4921
rect 9122 4901 9135 4921
rect 9085 4873 9135 4901
rect 4816 4741 4833 4761
rect 4853 4741 4866 4761
rect 4816 4713 4866 4741
rect 358 4675 408 4688
rect 571 4675 621 4688
rect 779 4675 829 4688
rect 987 4675 1037 4688
rect 1371 4674 1421 4690
rect 1584 4674 1634 4690
rect 1792 4674 1842 4690
rect 2000 4674 2050 4690
rect 6652 4760 6702 4788
rect 6652 4740 6665 4760
rect 6685 4740 6702 4760
rect 6652 4711 6702 4740
rect 6865 4759 6915 4788
rect 6865 4735 6876 4759
rect 6900 4735 6915 4759
rect 6865 4711 6915 4735
rect 7073 4764 7123 4788
rect 7073 4740 7085 4764
rect 7109 4740 7123 4764
rect 7073 4711 7123 4740
rect 7281 4762 7331 4788
rect 9468 4811 9518 4827
rect 9676 4811 9726 4827
rect 9884 4811 9934 4827
rect 10097 4811 10147 4827
rect 7281 4736 7299 4762
rect 7325 4736 7331 4762
rect 8456 4760 8506 4773
rect 8664 4760 8714 4773
rect 8872 4760 8922 4773
rect 9085 4760 9135 4773
rect 7281 4711 7331 4736
rect 9468 4744 9518 4769
rect 9468 4718 9474 4744
rect 9500 4718 9518 4744
rect 9468 4692 9518 4718
rect 9676 4740 9726 4769
rect 9676 4716 9690 4740
rect 9714 4716 9726 4740
rect 9676 4692 9726 4716
rect 9884 4745 9934 4769
rect 9884 4721 9899 4745
rect 9923 4721 9934 4745
rect 9884 4692 9934 4721
rect 10097 4740 10147 4769
rect 10097 4720 10114 4740
rect 10134 4720 10147 4740
rect 10097 4692 10147 4720
rect 5639 4654 5689 4667
rect 5852 4654 5902 4667
rect 6060 4654 6110 4667
rect 6268 4654 6318 4667
rect 4187 4600 4237 4613
rect 4395 4600 4445 4613
rect 4603 4600 4653 4613
rect 4816 4600 4866 4613
rect 2880 4581 2930 4597
rect 3088 4581 3138 4597
rect 3296 4581 3346 4597
rect 3509 4581 3559 4597
rect 358 4547 408 4575
rect 358 4527 371 4547
rect 391 4527 408 4547
rect 358 4498 408 4527
rect 571 4546 621 4575
rect 571 4522 582 4546
rect 606 4522 621 4546
rect 571 4498 621 4522
rect 779 4551 829 4575
rect 779 4527 791 4551
rect 815 4527 829 4551
rect 779 4498 829 4527
rect 987 4549 1037 4575
rect 987 4523 1005 4549
rect 1031 4523 1037 4549
rect 6652 4653 6702 4669
rect 6865 4653 6915 4669
rect 7073 4653 7123 4669
rect 7281 4653 7331 4669
rect 9468 4579 9518 4592
rect 9676 4579 9726 4592
rect 9884 4579 9934 4592
rect 10097 4579 10147 4592
rect 8161 4560 8211 4576
rect 8369 4560 8419 4576
rect 8577 4560 8627 4576
rect 8790 4560 8840 4576
rect 987 4498 1037 4523
rect 2880 4514 2930 4539
rect 2880 4488 2886 4514
rect 2912 4488 2930 4514
rect 2880 4462 2930 4488
rect 3088 4510 3138 4539
rect 3088 4486 3102 4510
rect 3126 4486 3138 4510
rect 3088 4462 3138 4486
rect 3296 4515 3346 4539
rect 3296 4491 3311 4515
rect 3335 4491 3346 4515
rect 3296 4462 3346 4491
rect 3509 4510 3559 4539
rect 3509 4490 3526 4510
rect 3546 4490 3559 4510
rect 5639 4526 5689 4554
rect 3509 4462 3559 4490
rect 358 4440 408 4456
rect 571 4440 621 4456
rect 779 4440 829 4456
rect 987 4440 1037 4456
rect 1669 4365 1719 4378
rect 1882 4365 1932 4378
rect 2090 4365 2140 4378
rect 2298 4365 2348 4378
rect 5639 4506 5652 4526
rect 5672 4506 5689 4526
rect 5639 4477 5689 4506
rect 5852 4525 5902 4554
rect 5852 4501 5863 4525
rect 5887 4501 5902 4525
rect 5852 4477 5902 4501
rect 6060 4530 6110 4554
rect 6060 4506 6072 4530
rect 6096 4506 6110 4530
rect 6060 4477 6110 4506
rect 6268 4528 6318 4554
rect 6268 4502 6286 4528
rect 6312 4502 6318 4528
rect 6268 4477 6318 4502
rect 8161 4493 8211 4518
rect 8161 4467 8167 4493
rect 8193 4467 8211 4493
rect 8161 4441 8211 4467
rect 8369 4489 8419 4518
rect 8369 4465 8383 4489
rect 8407 4465 8419 4489
rect 8369 4441 8419 4465
rect 8577 4494 8627 4518
rect 8577 4470 8592 4494
rect 8616 4470 8627 4494
rect 8577 4441 8627 4470
rect 8790 4489 8840 4518
rect 8790 4469 8807 4489
rect 8827 4469 8840 4489
rect 8790 4441 8840 4469
rect 5639 4419 5689 4435
rect 5852 4419 5902 4435
rect 6060 4419 6110 4435
rect 6268 4419 6318 4435
rect 2880 4349 2930 4362
rect 3088 4349 3138 4362
rect 3296 4349 3346 4362
rect 3509 4349 3559 4362
rect 6950 4344 7000 4357
rect 7163 4344 7213 4357
rect 7371 4344 7421 4357
rect 7579 4344 7629 4357
rect 4191 4271 4241 4287
rect 4399 4271 4449 4287
rect 4607 4271 4657 4287
rect 4820 4271 4870 4287
rect 1669 4237 1719 4265
rect 1669 4217 1682 4237
rect 1702 4217 1719 4237
rect 1669 4188 1719 4217
rect 1882 4236 1932 4265
rect 1882 4212 1893 4236
rect 1917 4212 1932 4236
rect 1882 4188 1932 4212
rect 2090 4241 2140 4265
rect 2090 4217 2102 4241
rect 2126 4217 2140 4241
rect 2090 4188 2140 4217
rect 2298 4239 2348 4265
rect 2298 4213 2316 4239
rect 2342 4213 2348 4239
rect 2298 4188 2348 4213
rect 4191 4204 4241 4229
rect 4191 4178 4197 4204
rect 4223 4178 4241 4204
rect 4191 4152 4241 4178
rect 4399 4200 4449 4229
rect 4399 4176 4413 4200
rect 4437 4176 4449 4200
rect 4399 4152 4449 4176
rect 4607 4205 4657 4229
rect 4607 4181 4622 4205
rect 4646 4181 4657 4205
rect 4607 4152 4657 4181
rect 4820 4200 4870 4229
rect 4820 4180 4837 4200
rect 4857 4180 4870 4200
rect 8161 4328 8211 4341
rect 8369 4328 8419 4341
rect 8577 4328 8627 4341
rect 8790 4328 8840 4341
rect 9472 4250 9522 4266
rect 9680 4250 9730 4266
rect 9888 4250 9938 4266
rect 10101 4250 10151 4266
rect 6950 4216 7000 4244
rect 4820 4152 4870 4180
rect 6950 4196 6963 4216
rect 6983 4196 7000 4216
rect 6950 4167 7000 4196
rect 7163 4215 7213 4244
rect 7163 4191 7174 4215
rect 7198 4191 7213 4215
rect 7163 4167 7213 4191
rect 7371 4220 7421 4244
rect 7371 4196 7383 4220
rect 7407 4196 7421 4220
rect 7371 4167 7421 4196
rect 7579 4218 7629 4244
rect 7579 4192 7597 4218
rect 7623 4192 7629 4218
rect 7579 4167 7629 4192
rect 9472 4183 9522 4208
rect 1669 4130 1719 4146
rect 1882 4130 1932 4146
rect 2090 4130 2140 4146
rect 2298 4130 2348 4146
rect 362 4114 412 4127
rect 575 4114 625 4127
rect 783 4114 833 4127
rect 991 4114 1041 4127
rect 3178 4037 3228 4053
rect 3386 4037 3436 4053
rect 3594 4037 3644 4053
rect 3807 4037 3857 4053
rect 9472 4157 9478 4183
rect 9504 4157 9522 4183
rect 9472 4131 9522 4157
rect 9680 4179 9730 4208
rect 9680 4155 9694 4179
rect 9718 4155 9730 4179
rect 9680 4131 9730 4155
rect 9888 4184 9938 4208
rect 9888 4160 9903 4184
rect 9927 4160 9938 4184
rect 9888 4131 9938 4160
rect 10101 4179 10151 4208
rect 10101 4159 10118 4179
rect 10138 4159 10151 4179
rect 10101 4131 10151 4159
rect 6950 4109 7000 4125
rect 7163 4109 7213 4125
rect 7371 4109 7421 4125
rect 7579 4109 7629 4125
rect 5643 4093 5693 4106
rect 5856 4093 5906 4106
rect 6064 4093 6114 4106
rect 6272 4093 6322 4106
rect 4191 4039 4241 4052
rect 4399 4039 4449 4052
rect 4607 4039 4657 4052
rect 4820 4039 4870 4052
rect 362 3986 412 4014
rect 362 3966 375 3986
rect 395 3966 412 3986
rect 362 3937 412 3966
rect 575 3985 625 4014
rect 575 3961 586 3985
rect 610 3961 625 3985
rect 575 3937 625 3961
rect 783 3990 833 4014
rect 783 3966 795 3990
rect 819 3966 833 3990
rect 783 3937 833 3966
rect 991 3988 1041 4014
rect 991 3962 1009 3988
rect 1035 3962 1041 3988
rect 991 3937 1041 3962
rect 3178 3970 3228 3995
rect 1374 3933 1424 3946
rect 1587 3933 1637 3946
rect 1795 3933 1845 3946
rect 2003 3933 2053 3946
rect 3178 3944 3184 3970
rect 3210 3944 3228 3970
rect 362 3879 412 3895
rect 575 3879 625 3895
rect 783 3879 833 3895
rect 991 3879 1041 3895
rect 3178 3918 3228 3944
rect 3386 3966 3436 3995
rect 3386 3942 3400 3966
rect 3424 3942 3436 3966
rect 3386 3918 3436 3942
rect 3594 3971 3644 3995
rect 3594 3947 3609 3971
rect 3633 3947 3644 3971
rect 3594 3918 3644 3947
rect 3807 3966 3857 3995
rect 3807 3946 3824 3966
rect 3844 3946 3857 3966
rect 3807 3918 3857 3946
rect 8459 4016 8509 4032
rect 8667 4016 8717 4032
rect 8875 4016 8925 4032
rect 9088 4016 9138 4032
rect 9472 4018 9522 4031
rect 9680 4018 9730 4031
rect 9888 4018 9938 4031
rect 10101 4018 10151 4031
rect 5643 3965 5693 3993
rect 5643 3945 5656 3965
rect 5676 3945 5693 3965
rect 1374 3805 1424 3833
rect 1374 3785 1387 3805
rect 1407 3785 1424 3805
rect 1374 3756 1424 3785
rect 1587 3804 1637 3833
rect 1587 3780 1598 3804
rect 1622 3780 1637 3804
rect 1587 3756 1637 3780
rect 1795 3809 1845 3833
rect 1795 3785 1807 3809
rect 1831 3785 1845 3809
rect 1795 3756 1845 3785
rect 2003 3807 2053 3833
rect 5643 3916 5693 3945
rect 5856 3964 5906 3993
rect 5856 3940 5867 3964
rect 5891 3940 5906 3964
rect 5856 3916 5906 3940
rect 6064 3969 6114 3993
rect 6064 3945 6076 3969
rect 6100 3945 6114 3969
rect 6064 3916 6114 3945
rect 6272 3967 6322 3993
rect 6272 3941 6290 3967
rect 6316 3941 6322 3967
rect 6272 3916 6322 3941
rect 8459 3949 8509 3974
rect 6655 3912 6705 3925
rect 6868 3912 6918 3925
rect 7076 3912 7126 3925
rect 7284 3912 7334 3925
rect 8459 3923 8465 3949
rect 8491 3923 8509 3949
rect 4190 3856 4240 3872
rect 4398 3856 4448 3872
rect 4606 3856 4656 3872
rect 4819 3856 4869 3872
rect 5643 3858 5693 3874
rect 5856 3858 5906 3874
rect 6064 3858 6114 3874
rect 6272 3858 6322 3874
rect 2003 3781 2021 3807
rect 2047 3781 2053 3807
rect 3178 3805 3228 3818
rect 3386 3805 3436 3818
rect 3594 3805 3644 3818
rect 3807 3805 3857 3818
rect 2003 3756 2053 3781
rect 4190 3789 4240 3814
rect 4190 3763 4196 3789
rect 4222 3763 4240 3789
rect 4190 3737 4240 3763
rect 4398 3785 4448 3814
rect 4398 3761 4412 3785
rect 4436 3761 4448 3785
rect 4398 3737 4448 3761
rect 4606 3790 4656 3814
rect 4606 3766 4621 3790
rect 4645 3766 4656 3790
rect 4606 3737 4656 3766
rect 4819 3785 4869 3814
rect 8459 3897 8509 3923
rect 8667 3945 8717 3974
rect 8667 3921 8681 3945
rect 8705 3921 8717 3945
rect 8667 3897 8717 3921
rect 8875 3950 8925 3974
rect 8875 3926 8890 3950
rect 8914 3926 8925 3950
rect 8875 3897 8925 3926
rect 9088 3945 9138 3974
rect 9088 3925 9105 3945
rect 9125 3925 9138 3945
rect 9088 3897 9138 3925
rect 4819 3765 4836 3785
rect 4856 3765 4869 3785
rect 4819 3737 4869 3765
rect 361 3699 411 3712
rect 574 3699 624 3712
rect 782 3699 832 3712
rect 990 3699 1040 3712
rect 1374 3698 1424 3714
rect 1587 3698 1637 3714
rect 1795 3698 1845 3714
rect 2003 3698 2053 3714
rect 6655 3784 6705 3812
rect 6655 3764 6668 3784
rect 6688 3764 6705 3784
rect 6655 3735 6705 3764
rect 6868 3783 6918 3812
rect 6868 3759 6879 3783
rect 6903 3759 6918 3783
rect 6868 3735 6918 3759
rect 7076 3788 7126 3812
rect 7076 3764 7088 3788
rect 7112 3764 7126 3788
rect 7076 3735 7126 3764
rect 7284 3786 7334 3812
rect 9471 3835 9521 3851
rect 9679 3835 9729 3851
rect 9887 3835 9937 3851
rect 10100 3835 10150 3851
rect 7284 3760 7302 3786
rect 7328 3760 7334 3786
rect 8459 3784 8509 3797
rect 8667 3784 8717 3797
rect 8875 3784 8925 3797
rect 9088 3784 9138 3797
rect 7284 3735 7334 3760
rect 9471 3768 9521 3793
rect 9471 3742 9477 3768
rect 9503 3742 9521 3768
rect 9471 3716 9521 3742
rect 9679 3764 9729 3793
rect 9679 3740 9693 3764
rect 9717 3740 9729 3764
rect 9679 3716 9729 3740
rect 9887 3769 9937 3793
rect 9887 3745 9902 3769
rect 9926 3745 9937 3769
rect 9887 3716 9937 3745
rect 10100 3764 10150 3793
rect 10100 3744 10117 3764
rect 10137 3744 10150 3764
rect 10100 3716 10150 3744
rect 5642 3678 5692 3691
rect 5855 3678 5905 3691
rect 6063 3678 6113 3691
rect 6271 3678 6321 3691
rect 3128 3617 3178 3633
rect 3336 3617 3386 3633
rect 3544 3617 3594 3633
rect 3757 3617 3807 3633
rect 4190 3624 4240 3637
rect 4398 3624 4448 3637
rect 4606 3624 4656 3637
rect 4819 3624 4869 3637
rect 361 3571 411 3599
rect 361 3551 374 3571
rect 394 3551 411 3571
rect 361 3522 411 3551
rect 574 3570 624 3599
rect 574 3546 585 3570
rect 609 3546 624 3570
rect 574 3522 624 3546
rect 782 3575 832 3599
rect 782 3551 794 3575
rect 818 3551 832 3575
rect 782 3522 832 3551
rect 990 3573 1040 3599
rect 990 3547 1008 3573
rect 1034 3547 1040 3573
rect 990 3522 1040 3547
rect 3128 3550 3178 3575
rect 3128 3524 3134 3550
rect 3160 3524 3178 3550
rect 3128 3498 3178 3524
rect 3336 3546 3386 3575
rect 3336 3522 3350 3546
rect 3374 3522 3386 3546
rect 3336 3498 3386 3522
rect 3544 3551 3594 3575
rect 3544 3527 3559 3551
rect 3583 3527 3594 3551
rect 3544 3498 3594 3527
rect 3757 3546 3807 3575
rect 3757 3526 3774 3546
rect 3794 3526 3807 3546
rect 3757 3498 3807 3526
rect 6655 3677 6705 3693
rect 6868 3677 6918 3693
rect 7076 3677 7126 3693
rect 7284 3677 7334 3693
rect 8409 3596 8459 3612
rect 8617 3596 8667 3612
rect 8825 3596 8875 3612
rect 9038 3596 9088 3612
rect 9471 3603 9521 3616
rect 9679 3603 9729 3616
rect 9887 3603 9937 3616
rect 10100 3603 10150 3616
rect 5642 3550 5692 3578
rect 361 3464 411 3480
rect 574 3464 624 3480
rect 782 3464 832 3480
rect 990 3464 1040 3480
rect 5642 3530 5655 3550
rect 5675 3530 5692 3550
rect 5642 3501 5692 3530
rect 5855 3549 5905 3578
rect 5855 3525 5866 3549
rect 5890 3525 5905 3549
rect 5855 3501 5905 3525
rect 6063 3554 6113 3578
rect 6063 3530 6075 3554
rect 6099 3530 6113 3554
rect 6063 3501 6113 3530
rect 6271 3552 6321 3578
rect 6271 3526 6289 3552
rect 6315 3526 6321 3552
rect 6271 3501 6321 3526
rect 8409 3529 8459 3554
rect 8409 3503 8415 3529
rect 8441 3503 8459 3529
rect 8409 3477 8459 3503
rect 8617 3525 8667 3554
rect 8617 3501 8631 3525
rect 8655 3501 8667 3525
rect 8617 3477 8667 3501
rect 8825 3530 8875 3554
rect 8825 3506 8840 3530
rect 8864 3506 8875 3530
rect 8825 3477 8875 3506
rect 9038 3525 9088 3554
rect 9038 3505 9055 3525
rect 9075 3505 9088 3525
rect 9038 3477 9088 3505
rect 5642 3443 5692 3459
rect 5855 3443 5905 3459
rect 6063 3443 6113 3459
rect 6271 3443 6321 3459
rect 3128 3385 3178 3398
rect 3336 3385 3386 3398
rect 3544 3385 3594 3398
rect 3757 3385 3807 3398
rect 1429 3372 1479 3385
rect 1642 3372 1692 3385
rect 1850 3372 1900 3385
rect 2058 3372 2108 3385
rect 8409 3364 8459 3377
rect 8617 3364 8667 3377
rect 8825 3364 8875 3377
rect 9038 3364 9088 3377
rect 6710 3351 6760 3364
rect 6923 3351 6973 3364
rect 7131 3351 7181 3364
rect 7339 3351 7389 3364
rect 4196 3290 4246 3306
rect 4404 3290 4454 3306
rect 4612 3290 4662 3306
rect 4825 3290 4875 3306
rect 1429 3244 1479 3272
rect 1429 3224 1442 3244
rect 1462 3224 1479 3244
rect 1429 3195 1479 3224
rect 1642 3243 1692 3272
rect 1642 3219 1653 3243
rect 1677 3219 1692 3243
rect 1642 3195 1692 3219
rect 1850 3248 1900 3272
rect 1850 3224 1862 3248
rect 1886 3224 1900 3248
rect 1850 3195 1900 3224
rect 2058 3246 2108 3272
rect 2058 3220 2076 3246
rect 2102 3220 2108 3246
rect 2058 3195 2108 3220
rect 4196 3223 4246 3248
rect 4196 3197 4202 3223
rect 4228 3197 4246 3223
rect 4196 3171 4246 3197
rect 4404 3219 4454 3248
rect 4404 3195 4418 3219
rect 4442 3195 4454 3219
rect 4404 3171 4454 3195
rect 4612 3224 4662 3248
rect 4612 3200 4627 3224
rect 4651 3200 4662 3224
rect 4612 3171 4662 3200
rect 4825 3219 4875 3248
rect 4825 3199 4842 3219
rect 4862 3199 4875 3219
rect 9477 3269 9527 3285
rect 9685 3269 9735 3285
rect 9893 3269 9943 3285
rect 10106 3269 10156 3285
rect 4825 3171 4875 3199
rect 367 3133 417 3146
rect 580 3133 630 3146
rect 788 3133 838 3146
rect 996 3133 1046 3146
rect 1429 3137 1479 3153
rect 1642 3137 1692 3153
rect 1850 3137 1900 3153
rect 2058 3137 2108 3153
rect 3183 3056 3233 3072
rect 3391 3056 3441 3072
rect 3599 3056 3649 3072
rect 3812 3056 3862 3072
rect 6710 3223 6760 3251
rect 6710 3203 6723 3223
rect 6743 3203 6760 3223
rect 6710 3174 6760 3203
rect 6923 3222 6973 3251
rect 6923 3198 6934 3222
rect 6958 3198 6973 3222
rect 6923 3174 6973 3198
rect 7131 3227 7181 3251
rect 7131 3203 7143 3227
rect 7167 3203 7181 3227
rect 7131 3174 7181 3203
rect 7339 3225 7389 3251
rect 7339 3199 7357 3225
rect 7383 3199 7389 3225
rect 7339 3174 7389 3199
rect 9477 3202 9527 3227
rect 9477 3176 9483 3202
rect 9509 3176 9527 3202
rect 9477 3150 9527 3176
rect 9685 3198 9735 3227
rect 9685 3174 9699 3198
rect 9723 3174 9735 3198
rect 9685 3150 9735 3174
rect 9893 3203 9943 3227
rect 9893 3179 9908 3203
rect 9932 3179 9943 3203
rect 9893 3150 9943 3179
rect 10106 3198 10156 3227
rect 10106 3178 10123 3198
rect 10143 3178 10156 3198
rect 10106 3150 10156 3178
rect 5648 3112 5698 3125
rect 5861 3112 5911 3125
rect 6069 3112 6119 3125
rect 6277 3112 6327 3125
rect 6710 3116 6760 3132
rect 6923 3116 6973 3132
rect 7131 3116 7181 3132
rect 7339 3116 7389 3132
rect 4196 3058 4246 3071
rect 4404 3058 4454 3071
rect 4612 3058 4662 3071
rect 4825 3058 4875 3071
rect 367 3005 417 3033
rect 367 2985 380 3005
rect 400 2985 417 3005
rect 367 2956 417 2985
rect 580 3004 630 3033
rect 580 2980 591 3004
rect 615 2980 630 3004
rect 580 2956 630 2980
rect 788 3009 838 3033
rect 788 2985 800 3009
rect 824 2985 838 3009
rect 788 2956 838 2985
rect 996 3007 1046 3033
rect 996 2981 1014 3007
rect 1040 2981 1046 3007
rect 996 2956 1046 2981
rect 3183 2989 3233 3014
rect 1379 2952 1429 2965
rect 1592 2952 1642 2965
rect 1800 2952 1850 2965
rect 2008 2952 2058 2965
rect 3183 2963 3189 2989
rect 3215 2963 3233 2989
rect 367 2898 417 2914
rect 580 2898 630 2914
rect 788 2898 838 2914
rect 996 2898 1046 2914
rect 3183 2937 3233 2963
rect 3391 2985 3441 3014
rect 3391 2961 3405 2985
rect 3429 2961 3441 2985
rect 3391 2937 3441 2961
rect 3599 2990 3649 3014
rect 3599 2966 3614 2990
rect 3638 2966 3649 2990
rect 3599 2937 3649 2966
rect 3812 2985 3862 3014
rect 3812 2965 3829 2985
rect 3849 2965 3862 2985
rect 3812 2937 3862 2965
rect 8464 3035 8514 3051
rect 8672 3035 8722 3051
rect 8880 3035 8930 3051
rect 9093 3035 9143 3051
rect 9477 3037 9527 3050
rect 9685 3037 9735 3050
rect 9893 3037 9943 3050
rect 10106 3037 10156 3050
rect 5648 2984 5698 3012
rect 5648 2964 5661 2984
rect 5681 2964 5698 2984
rect 1379 2824 1429 2852
rect 1379 2804 1392 2824
rect 1412 2804 1429 2824
rect 1379 2775 1429 2804
rect 1592 2823 1642 2852
rect 1592 2799 1603 2823
rect 1627 2799 1642 2823
rect 1592 2775 1642 2799
rect 1800 2828 1850 2852
rect 1800 2804 1812 2828
rect 1836 2804 1850 2828
rect 1800 2775 1850 2804
rect 2008 2826 2058 2852
rect 5648 2935 5698 2964
rect 5861 2983 5911 3012
rect 5861 2959 5872 2983
rect 5896 2959 5911 2983
rect 5861 2935 5911 2959
rect 6069 2988 6119 3012
rect 6069 2964 6081 2988
rect 6105 2964 6119 2988
rect 6069 2935 6119 2964
rect 6277 2986 6327 3012
rect 6277 2960 6295 2986
rect 6321 2960 6327 2986
rect 6277 2935 6327 2960
rect 8464 2968 8514 2993
rect 6660 2931 6710 2944
rect 6873 2931 6923 2944
rect 7081 2931 7131 2944
rect 7289 2931 7339 2944
rect 8464 2942 8470 2968
rect 8496 2942 8514 2968
rect 4195 2875 4245 2891
rect 4403 2875 4453 2891
rect 4611 2875 4661 2891
rect 4824 2875 4874 2891
rect 5648 2877 5698 2893
rect 5861 2877 5911 2893
rect 6069 2877 6119 2893
rect 6277 2877 6327 2893
rect 2008 2800 2026 2826
rect 2052 2800 2058 2826
rect 3183 2824 3233 2837
rect 3391 2824 3441 2837
rect 3599 2824 3649 2837
rect 3812 2824 3862 2837
rect 2008 2775 2058 2800
rect 4195 2808 4245 2833
rect 4195 2782 4201 2808
rect 4227 2782 4245 2808
rect 4195 2756 4245 2782
rect 4403 2804 4453 2833
rect 4403 2780 4417 2804
rect 4441 2780 4453 2804
rect 4403 2756 4453 2780
rect 4611 2809 4661 2833
rect 4611 2785 4626 2809
rect 4650 2785 4661 2809
rect 4611 2756 4661 2785
rect 4824 2804 4874 2833
rect 8464 2916 8514 2942
rect 8672 2964 8722 2993
rect 8672 2940 8686 2964
rect 8710 2940 8722 2964
rect 8672 2916 8722 2940
rect 8880 2969 8930 2993
rect 8880 2945 8895 2969
rect 8919 2945 8930 2969
rect 8880 2916 8930 2945
rect 9093 2964 9143 2993
rect 9093 2944 9110 2964
rect 9130 2944 9143 2964
rect 9093 2916 9143 2944
rect 4824 2784 4841 2804
rect 4861 2784 4874 2804
rect 4824 2756 4874 2784
rect 366 2718 416 2731
rect 579 2718 629 2731
rect 787 2718 837 2731
rect 995 2718 1045 2731
rect 1379 2717 1429 2733
rect 1592 2717 1642 2733
rect 1800 2717 1850 2733
rect 2008 2717 2058 2733
rect 6660 2803 6710 2831
rect 6660 2783 6673 2803
rect 6693 2783 6710 2803
rect 6660 2754 6710 2783
rect 6873 2802 6923 2831
rect 6873 2778 6884 2802
rect 6908 2778 6923 2802
rect 6873 2754 6923 2778
rect 7081 2807 7131 2831
rect 7081 2783 7093 2807
rect 7117 2783 7131 2807
rect 7081 2754 7131 2783
rect 7289 2805 7339 2831
rect 9476 2854 9526 2870
rect 9684 2854 9734 2870
rect 9892 2854 9942 2870
rect 10105 2854 10155 2870
rect 7289 2779 7307 2805
rect 7333 2779 7339 2805
rect 8464 2803 8514 2816
rect 8672 2803 8722 2816
rect 8880 2803 8930 2816
rect 9093 2803 9143 2816
rect 7289 2754 7339 2779
rect 9476 2787 9526 2812
rect 9476 2761 9482 2787
rect 9508 2761 9526 2787
rect 9476 2735 9526 2761
rect 9684 2783 9734 2812
rect 9684 2759 9698 2783
rect 9722 2759 9734 2783
rect 9684 2735 9734 2759
rect 9892 2788 9942 2812
rect 9892 2764 9907 2788
rect 9931 2764 9942 2788
rect 9892 2735 9942 2764
rect 10105 2783 10155 2812
rect 10105 2763 10122 2783
rect 10142 2763 10155 2783
rect 10105 2735 10155 2763
rect 5647 2697 5697 2710
rect 5860 2697 5910 2710
rect 6068 2697 6118 2710
rect 6276 2697 6326 2710
rect 4195 2643 4245 2656
rect 4403 2643 4453 2656
rect 4611 2643 4661 2656
rect 4824 2643 4874 2656
rect 366 2590 416 2618
rect 366 2570 379 2590
rect 399 2570 416 2590
rect 366 2541 416 2570
rect 579 2589 629 2618
rect 579 2565 590 2589
rect 614 2565 629 2589
rect 579 2541 629 2565
rect 787 2594 837 2618
rect 787 2570 799 2594
rect 823 2570 837 2594
rect 787 2541 837 2570
rect 995 2592 1045 2618
rect 995 2566 1013 2592
rect 1039 2566 1045 2592
rect 2975 2589 3025 2605
rect 3183 2589 3233 2605
rect 3391 2589 3441 2605
rect 3604 2589 3654 2605
rect 995 2541 1045 2566
rect 6660 2696 6710 2712
rect 6873 2696 6923 2712
rect 7081 2696 7131 2712
rect 7289 2696 7339 2712
rect 9476 2622 9526 2635
rect 9684 2622 9734 2635
rect 9892 2622 9942 2635
rect 10105 2622 10155 2635
rect 2975 2522 3025 2547
rect 366 2483 416 2499
rect 579 2483 629 2499
rect 787 2483 837 2499
rect 995 2483 1045 2499
rect 2975 2496 2981 2522
rect 3007 2496 3025 2522
rect 2975 2470 3025 2496
rect 3183 2518 3233 2547
rect 3183 2494 3197 2518
rect 3221 2494 3233 2518
rect 3183 2470 3233 2494
rect 3391 2523 3441 2547
rect 3391 2499 3406 2523
rect 3430 2499 3441 2523
rect 3391 2470 3441 2499
rect 3604 2518 3654 2547
rect 5647 2569 5697 2597
rect 3604 2498 3621 2518
rect 3641 2498 3654 2518
rect 5647 2549 5660 2569
rect 5680 2549 5697 2569
rect 3604 2470 3654 2498
rect 5647 2520 5697 2549
rect 5860 2568 5910 2597
rect 5860 2544 5871 2568
rect 5895 2544 5910 2568
rect 5860 2520 5910 2544
rect 6068 2573 6118 2597
rect 6068 2549 6080 2573
rect 6104 2549 6118 2573
rect 6068 2520 6118 2549
rect 6276 2571 6326 2597
rect 6276 2545 6294 2571
rect 6320 2545 6326 2571
rect 8256 2568 8306 2584
rect 8464 2568 8514 2584
rect 8672 2568 8722 2584
rect 8885 2568 8935 2584
rect 6276 2520 6326 2545
rect 1594 2440 1644 2453
rect 1807 2440 1857 2453
rect 2015 2440 2065 2453
rect 2223 2440 2273 2453
rect 8256 2501 8306 2526
rect 5647 2462 5697 2478
rect 5860 2462 5910 2478
rect 6068 2462 6118 2478
rect 6276 2462 6326 2478
rect 8256 2475 8262 2501
rect 8288 2475 8306 2501
rect 8256 2449 8306 2475
rect 8464 2497 8514 2526
rect 8464 2473 8478 2497
rect 8502 2473 8514 2497
rect 8464 2449 8514 2473
rect 8672 2502 8722 2526
rect 8672 2478 8687 2502
rect 8711 2478 8722 2502
rect 8672 2449 8722 2478
rect 8885 2497 8935 2526
rect 8885 2477 8902 2497
rect 8922 2477 8935 2497
rect 8885 2449 8935 2477
rect 6875 2419 6925 2432
rect 7088 2419 7138 2432
rect 7296 2419 7346 2432
rect 7504 2419 7554 2432
rect 2975 2357 3025 2370
rect 3183 2357 3233 2370
rect 3391 2357 3441 2370
rect 3604 2357 3654 2370
rect 1594 2312 1644 2340
rect 1594 2292 1607 2312
rect 1627 2292 1644 2312
rect 1594 2263 1644 2292
rect 1807 2311 1857 2340
rect 1807 2287 1818 2311
rect 1842 2287 1857 2311
rect 1807 2263 1857 2287
rect 2015 2316 2065 2340
rect 2015 2292 2027 2316
rect 2051 2292 2065 2316
rect 2015 2263 2065 2292
rect 2223 2314 2273 2340
rect 2223 2288 2241 2314
rect 2267 2288 2273 2314
rect 4203 2311 4253 2327
rect 4411 2311 4461 2327
rect 4619 2311 4669 2327
rect 4832 2311 4882 2327
rect 2223 2263 2273 2288
rect 8256 2336 8306 2349
rect 8464 2336 8514 2349
rect 8672 2336 8722 2349
rect 8885 2336 8935 2349
rect 4203 2244 4253 2269
rect 1594 2205 1644 2221
rect 1807 2205 1857 2221
rect 2015 2205 2065 2221
rect 2223 2205 2273 2221
rect 4203 2218 4209 2244
rect 4235 2218 4253 2244
rect 4203 2192 4253 2218
rect 4411 2240 4461 2269
rect 4411 2216 4425 2240
rect 4449 2216 4461 2240
rect 4411 2192 4461 2216
rect 4619 2245 4669 2269
rect 4619 2221 4634 2245
rect 4658 2221 4669 2245
rect 4619 2192 4669 2221
rect 4832 2240 4882 2269
rect 6875 2291 6925 2319
rect 4832 2220 4849 2240
rect 4869 2220 4882 2240
rect 6875 2271 6888 2291
rect 6908 2271 6925 2291
rect 4832 2192 4882 2220
rect 6875 2242 6925 2271
rect 7088 2290 7138 2319
rect 7088 2266 7099 2290
rect 7123 2266 7138 2290
rect 7088 2242 7138 2266
rect 7296 2295 7346 2319
rect 7296 2271 7308 2295
rect 7332 2271 7346 2295
rect 7296 2242 7346 2271
rect 7504 2293 7554 2319
rect 7504 2267 7522 2293
rect 7548 2267 7554 2293
rect 9484 2290 9534 2306
rect 9692 2290 9742 2306
rect 9900 2290 9950 2306
rect 10113 2290 10163 2306
rect 7504 2242 7554 2267
rect 374 2154 424 2167
rect 587 2154 637 2167
rect 795 2154 845 2167
rect 1003 2154 1053 2167
rect 3190 2077 3240 2093
rect 3398 2077 3448 2093
rect 3606 2077 3656 2093
rect 3819 2077 3869 2093
rect 9484 2223 9534 2248
rect 6875 2184 6925 2200
rect 7088 2184 7138 2200
rect 7296 2184 7346 2200
rect 7504 2184 7554 2200
rect 9484 2197 9490 2223
rect 9516 2197 9534 2223
rect 9484 2171 9534 2197
rect 9692 2219 9742 2248
rect 9692 2195 9706 2219
rect 9730 2195 9742 2219
rect 9692 2171 9742 2195
rect 9900 2224 9950 2248
rect 9900 2200 9915 2224
rect 9939 2200 9950 2224
rect 9900 2171 9950 2200
rect 10113 2219 10163 2248
rect 10113 2199 10130 2219
rect 10150 2199 10163 2219
rect 10113 2171 10163 2199
rect 5655 2133 5705 2146
rect 5868 2133 5918 2146
rect 6076 2133 6126 2146
rect 6284 2133 6334 2146
rect 4203 2079 4253 2092
rect 4411 2079 4461 2092
rect 4619 2079 4669 2092
rect 4832 2079 4882 2092
rect 374 2026 424 2054
rect 374 2006 387 2026
rect 407 2006 424 2026
rect 374 1977 424 2006
rect 587 2025 637 2054
rect 587 2001 598 2025
rect 622 2001 637 2025
rect 587 1977 637 2001
rect 795 2030 845 2054
rect 795 2006 807 2030
rect 831 2006 845 2030
rect 795 1977 845 2006
rect 1003 2028 1053 2054
rect 1003 2002 1021 2028
rect 1047 2002 1053 2028
rect 1003 1977 1053 2002
rect 3190 2010 3240 2035
rect 1386 1973 1436 1986
rect 1599 1973 1649 1986
rect 1807 1973 1857 1986
rect 2015 1973 2065 1986
rect 3190 1984 3196 2010
rect 3222 1984 3240 2010
rect 374 1919 424 1935
rect 587 1919 637 1935
rect 795 1919 845 1935
rect 1003 1919 1053 1935
rect 3190 1958 3240 1984
rect 3398 2006 3448 2035
rect 3398 1982 3412 2006
rect 3436 1982 3448 2006
rect 3398 1958 3448 1982
rect 3606 2011 3656 2035
rect 3606 1987 3621 2011
rect 3645 1987 3656 2011
rect 3606 1958 3656 1987
rect 3819 2006 3869 2035
rect 3819 1986 3836 2006
rect 3856 1986 3869 2006
rect 3819 1958 3869 1986
rect 8471 2056 8521 2072
rect 8679 2056 8729 2072
rect 8887 2056 8937 2072
rect 9100 2056 9150 2072
rect 9484 2058 9534 2071
rect 9692 2058 9742 2071
rect 9900 2058 9950 2071
rect 10113 2058 10163 2071
rect 5655 2005 5705 2033
rect 5655 1985 5668 2005
rect 5688 1985 5705 2005
rect 1386 1845 1436 1873
rect 1386 1825 1399 1845
rect 1419 1825 1436 1845
rect 1386 1796 1436 1825
rect 1599 1844 1649 1873
rect 1599 1820 1610 1844
rect 1634 1820 1649 1844
rect 1599 1796 1649 1820
rect 1807 1849 1857 1873
rect 1807 1825 1819 1849
rect 1843 1825 1857 1849
rect 1807 1796 1857 1825
rect 2015 1847 2065 1873
rect 5655 1956 5705 1985
rect 5868 2004 5918 2033
rect 5868 1980 5879 2004
rect 5903 1980 5918 2004
rect 5868 1956 5918 1980
rect 6076 2009 6126 2033
rect 6076 1985 6088 2009
rect 6112 1985 6126 2009
rect 6076 1956 6126 1985
rect 6284 2007 6334 2033
rect 6284 1981 6302 2007
rect 6328 1981 6334 2007
rect 6284 1956 6334 1981
rect 8471 1989 8521 2014
rect 6667 1952 6717 1965
rect 6880 1952 6930 1965
rect 7088 1952 7138 1965
rect 7296 1952 7346 1965
rect 8471 1963 8477 1989
rect 8503 1963 8521 1989
rect 4202 1896 4252 1912
rect 4410 1896 4460 1912
rect 4618 1896 4668 1912
rect 4831 1896 4881 1912
rect 5655 1898 5705 1914
rect 5868 1898 5918 1914
rect 6076 1898 6126 1914
rect 6284 1898 6334 1914
rect 2015 1821 2033 1847
rect 2059 1821 2065 1847
rect 3190 1845 3240 1858
rect 3398 1845 3448 1858
rect 3606 1845 3656 1858
rect 3819 1845 3869 1858
rect 2015 1796 2065 1821
rect 4202 1829 4252 1854
rect 4202 1803 4208 1829
rect 4234 1803 4252 1829
rect 4202 1777 4252 1803
rect 4410 1825 4460 1854
rect 4410 1801 4424 1825
rect 4448 1801 4460 1825
rect 4410 1777 4460 1801
rect 4618 1830 4668 1854
rect 4618 1806 4633 1830
rect 4657 1806 4668 1830
rect 4618 1777 4668 1806
rect 4831 1825 4881 1854
rect 8471 1937 8521 1963
rect 8679 1985 8729 2014
rect 8679 1961 8693 1985
rect 8717 1961 8729 1985
rect 8679 1937 8729 1961
rect 8887 1990 8937 2014
rect 8887 1966 8902 1990
rect 8926 1966 8937 1990
rect 8887 1937 8937 1966
rect 9100 1985 9150 2014
rect 9100 1965 9117 1985
rect 9137 1965 9150 1985
rect 9100 1937 9150 1965
rect 4831 1805 4848 1825
rect 4868 1805 4881 1825
rect 4831 1777 4881 1805
rect 373 1739 423 1752
rect 586 1739 636 1752
rect 794 1739 844 1752
rect 1002 1739 1052 1752
rect 1386 1738 1436 1754
rect 1599 1738 1649 1754
rect 1807 1738 1857 1754
rect 2015 1738 2065 1754
rect 6667 1824 6717 1852
rect 6667 1804 6680 1824
rect 6700 1804 6717 1824
rect 6667 1775 6717 1804
rect 6880 1823 6930 1852
rect 6880 1799 6891 1823
rect 6915 1799 6930 1823
rect 6880 1775 6930 1799
rect 7088 1828 7138 1852
rect 7088 1804 7100 1828
rect 7124 1804 7138 1828
rect 7088 1775 7138 1804
rect 7296 1826 7346 1852
rect 9483 1875 9533 1891
rect 9691 1875 9741 1891
rect 9899 1875 9949 1891
rect 10112 1875 10162 1891
rect 7296 1800 7314 1826
rect 7340 1800 7346 1826
rect 8471 1824 8521 1837
rect 8679 1824 8729 1837
rect 8887 1824 8937 1837
rect 9100 1824 9150 1837
rect 7296 1775 7346 1800
rect 9483 1808 9533 1833
rect 9483 1782 9489 1808
rect 9515 1782 9533 1808
rect 9483 1756 9533 1782
rect 9691 1804 9741 1833
rect 9691 1780 9705 1804
rect 9729 1780 9741 1804
rect 9691 1756 9741 1780
rect 9899 1809 9949 1833
rect 9899 1785 9914 1809
rect 9938 1785 9949 1809
rect 9899 1756 9949 1785
rect 10112 1804 10162 1833
rect 10112 1784 10129 1804
rect 10149 1784 10162 1804
rect 10112 1756 10162 1784
rect 5654 1718 5704 1731
rect 5867 1718 5917 1731
rect 6075 1718 6125 1731
rect 6283 1718 6333 1731
rect 3140 1657 3190 1673
rect 3348 1657 3398 1673
rect 3556 1657 3606 1673
rect 3769 1657 3819 1673
rect 4202 1664 4252 1677
rect 4410 1664 4460 1677
rect 4618 1664 4668 1677
rect 4831 1664 4881 1677
rect 373 1611 423 1639
rect 373 1591 386 1611
rect 406 1591 423 1611
rect 373 1562 423 1591
rect 586 1610 636 1639
rect 586 1586 597 1610
rect 621 1586 636 1610
rect 586 1562 636 1586
rect 794 1615 844 1639
rect 794 1591 806 1615
rect 830 1591 844 1615
rect 794 1562 844 1591
rect 1002 1613 1052 1639
rect 1002 1587 1020 1613
rect 1046 1587 1052 1613
rect 1002 1562 1052 1587
rect 3140 1590 3190 1615
rect 3140 1564 3146 1590
rect 3172 1564 3190 1590
rect 3140 1538 3190 1564
rect 3348 1586 3398 1615
rect 3348 1562 3362 1586
rect 3386 1562 3398 1586
rect 3348 1538 3398 1562
rect 3556 1591 3606 1615
rect 3556 1567 3571 1591
rect 3595 1567 3606 1591
rect 3556 1538 3606 1567
rect 3769 1586 3819 1615
rect 3769 1566 3786 1586
rect 3806 1566 3819 1586
rect 3769 1538 3819 1566
rect 6667 1717 6717 1733
rect 6880 1717 6930 1733
rect 7088 1717 7138 1733
rect 7296 1717 7346 1733
rect 8421 1636 8471 1652
rect 8629 1636 8679 1652
rect 8837 1636 8887 1652
rect 9050 1636 9100 1652
rect 9483 1643 9533 1656
rect 9691 1643 9741 1656
rect 9899 1643 9949 1656
rect 10112 1643 10162 1656
rect 5654 1590 5704 1618
rect 373 1504 423 1520
rect 586 1504 636 1520
rect 794 1504 844 1520
rect 1002 1504 1052 1520
rect 5654 1570 5667 1590
rect 5687 1570 5704 1590
rect 5654 1541 5704 1570
rect 5867 1589 5917 1618
rect 5867 1565 5878 1589
rect 5902 1565 5917 1589
rect 5867 1541 5917 1565
rect 6075 1594 6125 1618
rect 6075 1570 6087 1594
rect 6111 1570 6125 1594
rect 6075 1541 6125 1570
rect 6283 1592 6333 1618
rect 6283 1566 6301 1592
rect 6327 1566 6333 1592
rect 6283 1541 6333 1566
rect 8421 1569 8471 1594
rect 8421 1543 8427 1569
rect 8453 1543 8471 1569
rect 8421 1517 8471 1543
rect 8629 1565 8679 1594
rect 8629 1541 8643 1565
rect 8667 1541 8679 1565
rect 8629 1517 8679 1541
rect 8837 1570 8887 1594
rect 8837 1546 8852 1570
rect 8876 1546 8887 1570
rect 8837 1517 8887 1546
rect 9050 1565 9100 1594
rect 9050 1545 9067 1565
rect 9087 1545 9100 1565
rect 9050 1517 9100 1545
rect 5654 1483 5704 1499
rect 5867 1483 5917 1499
rect 6075 1483 6125 1499
rect 6283 1483 6333 1499
rect 3140 1425 3190 1438
rect 3348 1425 3398 1438
rect 3556 1425 3606 1438
rect 3769 1425 3819 1438
rect 1441 1412 1491 1425
rect 1654 1412 1704 1425
rect 1862 1412 1912 1425
rect 2070 1412 2120 1425
rect 8421 1404 8471 1417
rect 8629 1404 8679 1417
rect 8837 1404 8887 1417
rect 9050 1404 9100 1417
rect 6722 1391 6772 1404
rect 6935 1391 6985 1404
rect 7143 1391 7193 1404
rect 7351 1391 7401 1404
rect 4208 1330 4258 1346
rect 4416 1330 4466 1346
rect 4624 1330 4674 1346
rect 4837 1330 4887 1346
rect 1441 1284 1491 1312
rect 1441 1264 1454 1284
rect 1474 1264 1491 1284
rect 1441 1235 1491 1264
rect 1654 1283 1704 1312
rect 1654 1259 1665 1283
rect 1689 1259 1704 1283
rect 1654 1235 1704 1259
rect 1862 1288 1912 1312
rect 1862 1264 1874 1288
rect 1898 1264 1912 1288
rect 1862 1235 1912 1264
rect 2070 1286 2120 1312
rect 2070 1260 2088 1286
rect 2114 1260 2120 1286
rect 2070 1235 2120 1260
rect 4208 1263 4258 1288
rect 4208 1237 4214 1263
rect 4240 1237 4258 1263
rect 4208 1211 4258 1237
rect 4416 1259 4466 1288
rect 4416 1235 4430 1259
rect 4454 1235 4466 1259
rect 4416 1211 4466 1235
rect 4624 1264 4674 1288
rect 4624 1240 4639 1264
rect 4663 1240 4674 1264
rect 4624 1211 4674 1240
rect 4837 1259 4887 1288
rect 4837 1239 4854 1259
rect 4874 1239 4887 1259
rect 9489 1309 9539 1325
rect 9697 1309 9747 1325
rect 9905 1309 9955 1325
rect 10118 1309 10168 1325
rect 4837 1211 4887 1239
rect 379 1173 429 1186
rect 592 1173 642 1186
rect 800 1173 850 1186
rect 1008 1173 1058 1186
rect 1441 1177 1491 1193
rect 1654 1177 1704 1193
rect 1862 1177 1912 1193
rect 2070 1177 2120 1193
rect 3195 1096 3245 1112
rect 3403 1096 3453 1112
rect 3611 1096 3661 1112
rect 3824 1096 3874 1112
rect 6722 1263 6772 1291
rect 6722 1243 6735 1263
rect 6755 1243 6772 1263
rect 6722 1214 6772 1243
rect 6935 1262 6985 1291
rect 6935 1238 6946 1262
rect 6970 1238 6985 1262
rect 6935 1214 6985 1238
rect 7143 1267 7193 1291
rect 7143 1243 7155 1267
rect 7179 1243 7193 1267
rect 7143 1214 7193 1243
rect 7351 1265 7401 1291
rect 7351 1239 7369 1265
rect 7395 1239 7401 1265
rect 7351 1214 7401 1239
rect 9489 1242 9539 1267
rect 9489 1216 9495 1242
rect 9521 1216 9539 1242
rect 9489 1190 9539 1216
rect 9697 1238 9747 1267
rect 9697 1214 9711 1238
rect 9735 1214 9747 1238
rect 9697 1190 9747 1214
rect 9905 1243 9955 1267
rect 9905 1219 9920 1243
rect 9944 1219 9955 1243
rect 9905 1190 9955 1219
rect 10118 1238 10168 1267
rect 10118 1218 10135 1238
rect 10155 1218 10168 1238
rect 10118 1190 10168 1218
rect 5660 1152 5710 1165
rect 5873 1152 5923 1165
rect 6081 1152 6131 1165
rect 6289 1152 6339 1165
rect 6722 1156 6772 1172
rect 6935 1156 6985 1172
rect 7143 1156 7193 1172
rect 7351 1156 7401 1172
rect 4208 1098 4258 1111
rect 4416 1098 4466 1111
rect 4624 1098 4674 1111
rect 4837 1098 4887 1111
rect 379 1045 429 1073
rect 379 1025 392 1045
rect 412 1025 429 1045
rect 379 996 429 1025
rect 592 1044 642 1073
rect 592 1020 603 1044
rect 627 1020 642 1044
rect 592 996 642 1020
rect 800 1049 850 1073
rect 800 1025 812 1049
rect 836 1025 850 1049
rect 800 996 850 1025
rect 1008 1047 1058 1073
rect 1008 1021 1026 1047
rect 1052 1021 1058 1047
rect 1008 996 1058 1021
rect 3195 1029 3245 1054
rect 1391 992 1441 1005
rect 1604 992 1654 1005
rect 1812 992 1862 1005
rect 2020 992 2070 1005
rect 3195 1003 3201 1029
rect 3227 1003 3245 1029
rect 379 938 429 954
rect 592 938 642 954
rect 800 938 850 954
rect 1008 938 1058 954
rect 3195 977 3245 1003
rect 3403 1025 3453 1054
rect 3403 1001 3417 1025
rect 3441 1001 3453 1025
rect 3403 977 3453 1001
rect 3611 1030 3661 1054
rect 3611 1006 3626 1030
rect 3650 1006 3661 1030
rect 3611 977 3661 1006
rect 3824 1025 3874 1054
rect 3824 1005 3841 1025
rect 3861 1005 3874 1025
rect 3824 977 3874 1005
rect 8476 1075 8526 1091
rect 8684 1075 8734 1091
rect 8892 1075 8942 1091
rect 9105 1075 9155 1091
rect 9489 1077 9539 1090
rect 9697 1077 9747 1090
rect 9905 1077 9955 1090
rect 10118 1077 10168 1090
rect 5660 1024 5710 1052
rect 5660 1004 5673 1024
rect 5693 1004 5710 1024
rect 1391 864 1441 892
rect 1391 844 1404 864
rect 1424 844 1441 864
rect 1391 815 1441 844
rect 1604 863 1654 892
rect 1604 839 1615 863
rect 1639 839 1654 863
rect 1604 815 1654 839
rect 1812 868 1862 892
rect 1812 844 1824 868
rect 1848 844 1862 868
rect 1812 815 1862 844
rect 2020 866 2070 892
rect 5660 975 5710 1004
rect 5873 1023 5923 1052
rect 5873 999 5884 1023
rect 5908 999 5923 1023
rect 5873 975 5923 999
rect 6081 1028 6131 1052
rect 6081 1004 6093 1028
rect 6117 1004 6131 1028
rect 6081 975 6131 1004
rect 6289 1026 6339 1052
rect 6289 1000 6307 1026
rect 6333 1000 6339 1026
rect 6289 975 6339 1000
rect 8476 1008 8526 1033
rect 6672 971 6722 984
rect 6885 971 6935 984
rect 7093 971 7143 984
rect 7301 971 7351 984
rect 8476 982 8482 1008
rect 8508 982 8526 1008
rect 4207 915 4257 931
rect 4415 915 4465 931
rect 4623 915 4673 931
rect 4836 915 4886 931
rect 5660 917 5710 933
rect 5873 917 5923 933
rect 6081 917 6131 933
rect 6289 917 6339 933
rect 2020 840 2038 866
rect 2064 840 2070 866
rect 3195 864 3245 877
rect 3403 864 3453 877
rect 3611 864 3661 877
rect 3824 864 3874 877
rect 2020 815 2070 840
rect 4207 848 4257 873
rect 4207 822 4213 848
rect 4239 822 4257 848
rect 4207 796 4257 822
rect 4415 844 4465 873
rect 4415 820 4429 844
rect 4453 820 4465 844
rect 4415 796 4465 820
rect 4623 849 4673 873
rect 4623 825 4638 849
rect 4662 825 4673 849
rect 4623 796 4673 825
rect 4836 844 4886 873
rect 8476 956 8526 982
rect 8684 1004 8734 1033
rect 8684 980 8698 1004
rect 8722 980 8734 1004
rect 8684 956 8734 980
rect 8892 1009 8942 1033
rect 8892 985 8907 1009
rect 8931 985 8942 1009
rect 8892 956 8942 985
rect 9105 1004 9155 1033
rect 9105 984 9122 1004
rect 9142 984 9155 1004
rect 9105 956 9155 984
rect 4836 824 4853 844
rect 4873 824 4886 844
rect 4836 796 4886 824
rect 378 758 428 771
rect 591 758 641 771
rect 799 758 849 771
rect 1007 758 1057 771
rect 1391 757 1441 773
rect 1604 757 1654 773
rect 1812 757 1862 773
rect 2020 757 2070 773
rect 6672 843 6722 871
rect 6672 823 6685 843
rect 6705 823 6722 843
rect 6672 794 6722 823
rect 6885 842 6935 871
rect 6885 818 6896 842
rect 6920 818 6935 842
rect 6885 794 6935 818
rect 7093 847 7143 871
rect 7093 823 7105 847
rect 7129 823 7143 847
rect 7093 794 7143 823
rect 7301 845 7351 871
rect 9488 894 9538 910
rect 9696 894 9746 910
rect 9904 894 9954 910
rect 10117 894 10167 910
rect 7301 819 7319 845
rect 7345 819 7351 845
rect 8476 843 8526 856
rect 8684 843 8734 856
rect 8892 843 8942 856
rect 9105 843 9155 856
rect 7301 794 7351 819
rect 9488 827 9538 852
rect 9488 801 9494 827
rect 9520 801 9538 827
rect 9488 775 9538 801
rect 9696 823 9746 852
rect 9696 799 9710 823
rect 9734 799 9746 823
rect 9696 775 9746 799
rect 9904 828 9954 852
rect 9904 804 9919 828
rect 9943 804 9954 828
rect 9904 775 9954 804
rect 10117 823 10167 852
rect 10117 803 10134 823
rect 10154 803 10167 823
rect 10117 775 10167 803
rect 5659 737 5709 750
rect 5872 737 5922 750
rect 6080 737 6130 750
rect 6288 737 6338 750
rect 4207 683 4257 696
rect 4415 683 4465 696
rect 4623 683 4673 696
rect 4836 683 4886 696
rect 378 630 428 658
rect 378 610 391 630
rect 411 610 428 630
rect 378 581 428 610
rect 591 629 641 658
rect 591 605 602 629
rect 626 605 641 629
rect 591 581 641 605
rect 799 634 849 658
rect 799 610 811 634
rect 835 610 849 634
rect 799 581 849 610
rect 1007 632 1057 658
rect 1007 606 1025 632
rect 1051 606 1057 632
rect 1007 581 1057 606
rect 6672 736 6722 752
rect 6885 736 6935 752
rect 7093 736 7143 752
rect 7301 736 7351 752
rect 9488 662 9538 675
rect 9696 662 9746 675
rect 9904 662 9954 675
rect 10117 662 10167 675
rect 5659 609 5709 637
rect 5659 589 5672 609
rect 5692 589 5709 609
rect 378 523 428 539
rect 591 523 641 539
rect 799 523 849 539
rect 1007 523 1057 539
rect 5659 560 5709 589
rect 5872 608 5922 637
rect 5872 584 5883 608
rect 5907 584 5922 608
rect 5872 560 5922 584
rect 6080 613 6130 637
rect 6080 589 6092 613
rect 6116 589 6130 613
rect 6080 560 6130 589
rect 6288 611 6338 637
rect 6288 585 6306 611
rect 6332 585 6338 611
rect 6288 560 6338 585
rect 5659 502 5709 518
rect 5872 502 5922 518
rect 6080 502 6130 518
rect 6288 502 6338 518
rect 1781 277 1831 290
rect 1994 277 2044 290
rect 2202 277 2252 290
rect 2410 277 2460 290
rect 7062 256 7112 269
rect 7275 256 7325 269
rect 7483 256 7533 269
rect 7691 256 7741 269
rect 4871 189 4921 202
rect 5084 189 5134 202
rect 5292 189 5342 202
rect 5500 189 5550 202
rect 1781 149 1831 177
rect 1781 129 1794 149
rect 1814 129 1831 149
rect 1781 100 1831 129
rect 1994 148 2044 177
rect 1994 124 2005 148
rect 2029 124 2044 148
rect 1994 100 2044 124
rect 2202 153 2252 177
rect 2202 129 2214 153
rect 2238 129 2252 153
rect 2202 100 2252 129
rect 2410 151 2460 177
rect 2410 125 2428 151
rect 2454 125 2460 151
rect 2410 100 2460 125
rect 7062 128 7112 156
rect 7062 108 7075 128
rect 7095 108 7112 128
rect 4871 61 4921 89
rect 1781 42 1831 58
rect 1994 42 2044 58
rect 2202 42 2252 58
rect 2410 42 2460 58
rect 4871 41 4884 61
rect 4904 41 4921 61
rect 4871 12 4921 41
rect 5084 60 5134 89
rect 5084 36 5095 60
rect 5119 36 5134 60
rect 5084 12 5134 36
rect 5292 65 5342 89
rect 5292 41 5304 65
rect 5328 41 5342 65
rect 5292 12 5342 41
rect 5500 63 5550 89
rect 7062 79 7112 108
rect 7275 127 7325 156
rect 7275 103 7286 127
rect 7310 103 7325 127
rect 7275 79 7325 103
rect 7483 132 7533 156
rect 7483 108 7495 132
rect 7519 108 7533 132
rect 7483 79 7533 108
rect 7691 130 7741 156
rect 7691 104 7709 130
rect 7735 104 7741 130
rect 7691 79 7741 104
rect 5500 37 5518 63
rect 5544 37 5550 63
rect 5500 12 5550 37
rect 7062 21 7112 37
rect 7275 21 7325 37
rect 7483 21 7533 37
rect 7691 21 7741 37
rect 4871 -46 4921 -30
rect 5084 -46 5134 -30
rect 5292 -46 5342 -30
rect 5500 -46 5550 -30
<< polycont >>
rect 4177 8095 4203 8121
rect 4393 8093 4417 8117
rect 4602 8098 4626 8122
rect 4817 8097 4837 8117
rect 9458 8074 9484 8100
rect 9674 8072 9698 8096
rect 9883 8077 9907 8101
rect 10098 8076 10118 8096
rect 355 7883 375 7903
rect 566 7878 590 7902
rect 775 7883 799 7907
rect 989 7879 1015 7905
rect 3164 7861 3190 7887
rect 3380 7859 3404 7883
rect 3589 7864 3613 7888
rect 3804 7863 3824 7883
rect 5636 7862 5656 7882
rect 1367 7702 1387 7722
rect 1578 7697 1602 7721
rect 1787 7702 1811 7726
rect 5847 7857 5871 7881
rect 6056 7862 6080 7886
rect 6270 7858 6296 7884
rect 8445 7840 8471 7866
rect 2001 7698 2027 7724
rect 4176 7680 4202 7706
rect 4392 7678 4416 7702
rect 4601 7683 4625 7707
rect 8661 7838 8685 7862
rect 8870 7843 8894 7867
rect 9085 7842 9105 7862
rect 4816 7682 4836 7702
rect 6648 7681 6668 7701
rect 6859 7676 6883 7700
rect 7068 7681 7092 7705
rect 7282 7677 7308 7703
rect 9457 7659 9483 7685
rect 9673 7657 9697 7681
rect 9882 7662 9906 7686
rect 10097 7661 10117 7681
rect 354 7468 374 7488
rect 565 7463 589 7487
rect 774 7468 798 7492
rect 988 7464 1014 7490
rect 3114 7441 3140 7467
rect 3330 7439 3354 7463
rect 3539 7444 3563 7468
rect 3754 7443 3774 7463
rect 5635 7447 5655 7467
rect 5846 7442 5870 7466
rect 6055 7447 6079 7471
rect 6269 7443 6295 7469
rect 8395 7420 8421 7446
rect 8611 7418 8635 7442
rect 8820 7423 8844 7447
rect 9035 7422 9055 7442
rect 1422 7141 1442 7161
rect 1633 7136 1657 7160
rect 1842 7141 1866 7165
rect 2056 7137 2082 7163
rect 4182 7114 4208 7140
rect 4398 7112 4422 7136
rect 4607 7117 4631 7141
rect 4822 7116 4842 7136
rect 6703 7120 6723 7140
rect 6914 7115 6938 7139
rect 7123 7120 7147 7144
rect 7337 7116 7363 7142
rect 9463 7093 9489 7119
rect 9679 7091 9703 7115
rect 9888 7096 9912 7120
rect 10103 7095 10123 7115
rect 360 6902 380 6922
rect 571 6897 595 6921
rect 780 6902 804 6926
rect 994 6898 1020 6924
rect 3169 6880 3195 6906
rect 3385 6878 3409 6902
rect 3594 6883 3618 6907
rect 3809 6882 3829 6902
rect 5641 6881 5661 6901
rect 1372 6721 1392 6741
rect 1583 6716 1607 6740
rect 1792 6721 1816 6745
rect 5852 6876 5876 6900
rect 6061 6881 6085 6905
rect 6275 6877 6301 6903
rect 8450 6859 8476 6885
rect 2006 6717 2032 6743
rect 4181 6699 4207 6725
rect 4397 6697 4421 6721
rect 4606 6702 4630 6726
rect 8666 6857 8690 6881
rect 8875 6862 8899 6886
rect 9090 6861 9110 6881
rect 4821 6701 4841 6721
rect 6653 6700 6673 6720
rect 6864 6695 6888 6719
rect 7073 6700 7097 6724
rect 7287 6696 7313 6722
rect 9462 6678 9488 6704
rect 9678 6676 9702 6700
rect 9887 6681 9911 6705
rect 10102 6680 10122 6700
rect 359 6487 379 6507
rect 570 6482 594 6506
rect 779 6487 803 6511
rect 993 6483 1019 6509
rect 2961 6413 2987 6439
rect 3177 6411 3201 6435
rect 3386 6416 3410 6440
rect 3601 6415 3621 6435
rect 5640 6466 5660 6486
rect 5851 6461 5875 6485
rect 6060 6466 6084 6490
rect 6274 6462 6300 6488
rect 8242 6392 8268 6418
rect 8458 6390 8482 6414
rect 8667 6395 8691 6419
rect 8882 6394 8902 6414
rect 1587 6209 1607 6229
rect 1798 6204 1822 6228
rect 2007 6209 2031 6233
rect 2221 6205 2247 6231
rect 4189 6135 4215 6161
rect 4405 6133 4429 6157
rect 4614 6138 4638 6162
rect 4829 6137 4849 6157
rect 6868 6188 6888 6208
rect 7079 6183 7103 6207
rect 7288 6188 7312 6212
rect 7502 6184 7528 6210
rect 9470 6114 9496 6140
rect 9686 6112 9710 6136
rect 9895 6117 9919 6141
rect 10110 6116 10130 6136
rect 367 5923 387 5943
rect 578 5918 602 5942
rect 787 5923 811 5947
rect 1001 5919 1027 5945
rect 3176 5901 3202 5927
rect 3392 5899 3416 5923
rect 3601 5904 3625 5928
rect 3816 5903 3836 5923
rect 5648 5902 5668 5922
rect 1379 5742 1399 5762
rect 1590 5737 1614 5761
rect 1799 5742 1823 5766
rect 5859 5897 5883 5921
rect 6068 5902 6092 5926
rect 6282 5898 6308 5924
rect 8457 5880 8483 5906
rect 2013 5738 2039 5764
rect 4188 5720 4214 5746
rect 4404 5718 4428 5742
rect 4613 5723 4637 5747
rect 8673 5878 8697 5902
rect 8882 5883 8906 5907
rect 9097 5882 9117 5902
rect 4828 5722 4848 5742
rect 6660 5721 6680 5741
rect 6871 5716 6895 5740
rect 7080 5721 7104 5745
rect 7294 5717 7320 5743
rect 9469 5699 9495 5725
rect 9685 5697 9709 5721
rect 9894 5702 9918 5726
rect 10109 5701 10129 5721
rect 366 5508 386 5528
rect 577 5503 601 5527
rect 786 5508 810 5532
rect 1000 5504 1026 5530
rect 3126 5481 3152 5507
rect 3342 5479 3366 5503
rect 3551 5484 3575 5508
rect 3766 5483 3786 5503
rect 5647 5487 5667 5507
rect 5858 5482 5882 5506
rect 6067 5487 6091 5511
rect 6281 5483 6307 5509
rect 8407 5460 8433 5486
rect 8623 5458 8647 5482
rect 8832 5463 8856 5487
rect 9047 5462 9067 5482
rect 1434 5181 1454 5201
rect 1645 5176 1669 5200
rect 1854 5181 1878 5205
rect 2068 5177 2094 5203
rect 4194 5154 4220 5180
rect 4410 5152 4434 5176
rect 4619 5157 4643 5181
rect 4834 5156 4854 5176
rect 6715 5160 6735 5180
rect 6926 5155 6950 5179
rect 7135 5160 7159 5184
rect 7349 5156 7375 5182
rect 9475 5133 9501 5159
rect 9691 5131 9715 5155
rect 9900 5136 9924 5160
rect 10115 5135 10135 5155
rect 372 4942 392 4962
rect 583 4937 607 4961
rect 792 4942 816 4966
rect 1006 4938 1032 4964
rect 3181 4920 3207 4946
rect 3397 4918 3421 4942
rect 3606 4923 3630 4947
rect 3821 4922 3841 4942
rect 5653 4921 5673 4941
rect 1384 4761 1404 4781
rect 1595 4756 1619 4780
rect 1804 4761 1828 4785
rect 5864 4916 5888 4940
rect 6073 4921 6097 4945
rect 6287 4917 6313 4943
rect 8462 4899 8488 4925
rect 2018 4757 2044 4783
rect 4193 4739 4219 4765
rect 4409 4737 4433 4761
rect 4618 4742 4642 4766
rect 8678 4897 8702 4921
rect 8887 4902 8911 4926
rect 9102 4901 9122 4921
rect 4833 4741 4853 4761
rect 6665 4740 6685 4760
rect 6876 4735 6900 4759
rect 7085 4740 7109 4764
rect 7299 4736 7325 4762
rect 9474 4718 9500 4744
rect 9690 4716 9714 4740
rect 9899 4721 9923 4745
rect 10114 4720 10134 4740
rect 371 4527 391 4547
rect 582 4522 606 4546
rect 791 4527 815 4551
rect 1005 4523 1031 4549
rect 2886 4488 2912 4514
rect 3102 4486 3126 4510
rect 3311 4491 3335 4515
rect 3526 4490 3546 4510
rect 5652 4506 5672 4526
rect 5863 4501 5887 4525
rect 6072 4506 6096 4530
rect 6286 4502 6312 4528
rect 8167 4467 8193 4493
rect 8383 4465 8407 4489
rect 8592 4470 8616 4494
rect 8807 4469 8827 4489
rect 1682 4217 1702 4237
rect 1893 4212 1917 4236
rect 2102 4217 2126 4241
rect 2316 4213 2342 4239
rect 4197 4178 4223 4204
rect 4413 4176 4437 4200
rect 4622 4181 4646 4205
rect 4837 4180 4857 4200
rect 6963 4196 6983 4216
rect 7174 4191 7198 4215
rect 7383 4196 7407 4220
rect 7597 4192 7623 4218
rect 9478 4157 9504 4183
rect 9694 4155 9718 4179
rect 9903 4160 9927 4184
rect 10118 4159 10138 4179
rect 375 3966 395 3986
rect 586 3961 610 3985
rect 795 3966 819 3990
rect 1009 3962 1035 3988
rect 3184 3944 3210 3970
rect 3400 3942 3424 3966
rect 3609 3947 3633 3971
rect 3824 3946 3844 3966
rect 5656 3945 5676 3965
rect 1387 3785 1407 3805
rect 1598 3780 1622 3804
rect 1807 3785 1831 3809
rect 5867 3940 5891 3964
rect 6076 3945 6100 3969
rect 6290 3941 6316 3967
rect 8465 3923 8491 3949
rect 2021 3781 2047 3807
rect 4196 3763 4222 3789
rect 4412 3761 4436 3785
rect 4621 3766 4645 3790
rect 8681 3921 8705 3945
rect 8890 3926 8914 3950
rect 9105 3925 9125 3945
rect 4836 3765 4856 3785
rect 6668 3764 6688 3784
rect 6879 3759 6903 3783
rect 7088 3764 7112 3788
rect 7302 3760 7328 3786
rect 9477 3742 9503 3768
rect 9693 3740 9717 3764
rect 9902 3745 9926 3769
rect 10117 3744 10137 3764
rect 374 3551 394 3571
rect 585 3546 609 3570
rect 794 3551 818 3575
rect 1008 3547 1034 3573
rect 3134 3524 3160 3550
rect 3350 3522 3374 3546
rect 3559 3527 3583 3551
rect 3774 3526 3794 3546
rect 5655 3530 5675 3550
rect 5866 3525 5890 3549
rect 6075 3530 6099 3554
rect 6289 3526 6315 3552
rect 8415 3503 8441 3529
rect 8631 3501 8655 3525
rect 8840 3506 8864 3530
rect 9055 3505 9075 3525
rect 1442 3224 1462 3244
rect 1653 3219 1677 3243
rect 1862 3224 1886 3248
rect 2076 3220 2102 3246
rect 4202 3197 4228 3223
rect 4418 3195 4442 3219
rect 4627 3200 4651 3224
rect 4842 3199 4862 3219
rect 6723 3203 6743 3223
rect 6934 3198 6958 3222
rect 7143 3203 7167 3227
rect 7357 3199 7383 3225
rect 9483 3176 9509 3202
rect 9699 3174 9723 3198
rect 9908 3179 9932 3203
rect 10123 3178 10143 3198
rect 380 2985 400 3005
rect 591 2980 615 3004
rect 800 2985 824 3009
rect 1014 2981 1040 3007
rect 3189 2963 3215 2989
rect 3405 2961 3429 2985
rect 3614 2966 3638 2990
rect 3829 2965 3849 2985
rect 5661 2964 5681 2984
rect 1392 2804 1412 2824
rect 1603 2799 1627 2823
rect 1812 2804 1836 2828
rect 5872 2959 5896 2983
rect 6081 2964 6105 2988
rect 6295 2960 6321 2986
rect 8470 2942 8496 2968
rect 2026 2800 2052 2826
rect 4201 2782 4227 2808
rect 4417 2780 4441 2804
rect 4626 2785 4650 2809
rect 8686 2940 8710 2964
rect 8895 2945 8919 2969
rect 9110 2944 9130 2964
rect 4841 2784 4861 2804
rect 6673 2783 6693 2803
rect 6884 2778 6908 2802
rect 7093 2783 7117 2807
rect 7307 2779 7333 2805
rect 9482 2761 9508 2787
rect 9698 2759 9722 2783
rect 9907 2764 9931 2788
rect 10122 2763 10142 2783
rect 379 2570 399 2590
rect 590 2565 614 2589
rect 799 2570 823 2594
rect 1013 2566 1039 2592
rect 2981 2496 3007 2522
rect 3197 2494 3221 2518
rect 3406 2499 3430 2523
rect 3621 2498 3641 2518
rect 5660 2549 5680 2569
rect 5871 2544 5895 2568
rect 6080 2549 6104 2573
rect 6294 2545 6320 2571
rect 8262 2475 8288 2501
rect 8478 2473 8502 2497
rect 8687 2478 8711 2502
rect 8902 2477 8922 2497
rect 1607 2292 1627 2312
rect 1818 2287 1842 2311
rect 2027 2292 2051 2316
rect 2241 2288 2267 2314
rect 4209 2218 4235 2244
rect 4425 2216 4449 2240
rect 4634 2221 4658 2245
rect 4849 2220 4869 2240
rect 6888 2271 6908 2291
rect 7099 2266 7123 2290
rect 7308 2271 7332 2295
rect 7522 2267 7548 2293
rect 9490 2197 9516 2223
rect 9706 2195 9730 2219
rect 9915 2200 9939 2224
rect 10130 2199 10150 2219
rect 387 2006 407 2026
rect 598 2001 622 2025
rect 807 2006 831 2030
rect 1021 2002 1047 2028
rect 3196 1984 3222 2010
rect 3412 1982 3436 2006
rect 3621 1987 3645 2011
rect 3836 1986 3856 2006
rect 5668 1985 5688 2005
rect 1399 1825 1419 1845
rect 1610 1820 1634 1844
rect 1819 1825 1843 1849
rect 5879 1980 5903 2004
rect 6088 1985 6112 2009
rect 6302 1981 6328 2007
rect 8477 1963 8503 1989
rect 2033 1821 2059 1847
rect 4208 1803 4234 1829
rect 4424 1801 4448 1825
rect 4633 1806 4657 1830
rect 8693 1961 8717 1985
rect 8902 1966 8926 1990
rect 9117 1965 9137 1985
rect 4848 1805 4868 1825
rect 6680 1804 6700 1824
rect 6891 1799 6915 1823
rect 7100 1804 7124 1828
rect 7314 1800 7340 1826
rect 9489 1782 9515 1808
rect 9705 1780 9729 1804
rect 9914 1785 9938 1809
rect 10129 1784 10149 1804
rect 386 1591 406 1611
rect 597 1586 621 1610
rect 806 1591 830 1615
rect 1020 1587 1046 1613
rect 3146 1564 3172 1590
rect 3362 1562 3386 1586
rect 3571 1567 3595 1591
rect 3786 1566 3806 1586
rect 5667 1570 5687 1590
rect 5878 1565 5902 1589
rect 6087 1570 6111 1594
rect 6301 1566 6327 1592
rect 8427 1543 8453 1569
rect 8643 1541 8667 1565
rect 8852 1546 8876 1570
rect 9067 1545 9087 1565
rect 1454 1264 1474 1284
rect 1665 1259 1689 1283
rect 1874 1264 1898 1288
rect 2088 1260 2114 1286
rect 4214 1237 4240 1263
rect 4430 1235 4454 1259
rect 4639 1240 4663 1264
rect 4854 1239 4874 1259
rect 6735 1243 6755 1263
rect 6946 1238 6970 1262
rect 7155 1243 7179 1267
rect 7369 1239 7395 1265
rect 9495 1216 9521 1242
rect 9711 1214 9735 1238
rect 9920 1219 9944 1243
rect 10135 1218 10155 1238
rect 392 1025 412 1045
rect 603 1020 627 1044
rect 812 1025 836 1049
rect 1026 1021 1052 1047
rect 3201 1003 3227 1029
rect 3417 1001 3441 1025
rect 3626 1006 3650 1030
rect 3841 1005 3861 1025
rect 5673 1004 5693 1024
rect 1404 844 1424 864
rect 1615 839 1639 863
rect 1824 844 1848 868
rect 5884 999 5908 1023
rect 6093 1004 6117 1028
rect 6307 1000 6333 1026
rect 8482 982 8508 1008
rect 2038 840 2064 866
rect 4213 822 4239 848
rect 4429 820 4453 844
rect 4638 825 4662 849
rect 8698 980 8722 1004
rect 8907 985 8931 1009
rect 9122 984 9142 1004
rect 4853 824 4873 844
rect 6685 823 6705 843
rect 6896 818 6920 842
rect 7105 823 7129 847
rect 7319 819 7345 845
rect 9494 801 9520 827
rect 9710 799 9734 823
rect 9919 804 9943 828
rect 10134 803 10154 823
rect 391 610 411 630
rect 602 605 626 629
rect 811 610 835 634
rect 1025 606 1051 632
rect 5672 589 5692 609
rect 5883 584 5907 608
rect 6092 589 6116 613
rect 6306 585 6332 611
rect 1794 129 1814 149
rect 2005 124 2029 148
rect 2214 129 2238 153
rect 2428 125 2454 151
rect 7075 108 7095 128
rect 4884 41 4904 61
rect 5095 36 5119 60
rect 5304 41 5328 65
rect 7286 103 7310 127
rect 7495 108 7519 132
rect 7709 104 7735 130
rect 5518 37 5544 63
<< ndiffres >>
rect 97 8226 154 8245
rect 97 8223 118 8226
rect 3 8208 118 8223
rect 136 8208 154 8226
rect 3 8185 154 8208
rect 5378 8205 5435 8224
rect 5378 8202 5399 8205
rect 3 8149 45 8185
rect 2 8148 102 8149
rect 2 8127 158 8148
rect 5028 8177 5089 8193
rect 5284 8187 5399 8202
rect 5417 8187 5435 8205
rect 5028 8173 5184 8177
rect 5028 8155 5048 8173
rect 5066 8155 5184 8173
rect 2 8109 120 8127
rect 138 8109 158 8127
rect 2 8105 158 8109
rect 97 8089 158 8105
rect 5028 8134 5184 8155
rect 5084 8133 5184 8134
rect 5284 8164 5435 8187
rect 5141 8097 5183 8133
rect 5284 8128 5326 8164
rect 5032 8074 5183 8097
rect 5283 8127 5383 8128
rect 5283 8106 5439 8127
rect 10309 8156 10370 8172
rect 10309 8152 10465 8156
rect 10309 8134 10329 8152
rect 10347 8134 10465 8152
rect 5283 8088 5401 8106
rect 5419 8088 5439 8106
rect 5283 8084 5439 8088
rect 95 8012 152 8031
rect 95 8009 116 8012
rect 1 7994 116 8009
rect 134 7994 152 8012
rect 1 7971 152 7994
rect 1 7935 43 7971
rect 0 7934 100 7935
rect 0 7913 156 7934
rect 5032 8056 5050 8074
rect 5068 8059 5183 8074
rect 5378 8068 5439 8084
rect 5068 8056 5089 8059
rect 5032 8037 5089 8056
rect 10309 8113 10465 8134
rect 10365 8112 10465 8113
rect 10422 8076 10464 8112
rect 10313 8053 10464 8076
rect 5035 7976 5096 7992
rect 5376 7991 5433 8010
rect 5376 7988 5397 7991
rect 5035 7972 5191 7976
rect 5035 7954 5055 7972
rect 5073 7954 5191 7972
rect 0 7895 118 7913
rect 136 7895 156 7913
rect 0 7891 156 7895
rect 95 7875 156 7891
rect 5035 7933 5191 7954
rect 5091 7932 5191 7933
rect 5282 7973 5397 7988
rect 5415 7973 5433 7991
rect 5282 7950 5433 7973
rect 5148 7896 5190 7932
rect 5282 7914 5324 7950
rect 5039 7873 5190 7896
rect 5039 7855 5057 7873
rect 5075 7858 5190 7873
rect 5281 7913 5381 7914
rect 5281 7892 5437 7913
rect 10313 8035 10331 8053
rect 10349 8038 10464 8053
rect 10349 8035 10370 8038
rect 10313 8016 10370 8035
rect 10316 7955 10377 7971
rect 10316 7951 10472 7955
rect 10316 7933 10336 7951
rect 10354 7933 10472 7951
rect 5281 7874 5399 7892
rect 5417 7874 5437 7892
rect 5281 7870 5437 7874
rect 5075 7855 5096 7858
rect 5039 7836 5096 7855
rect 5376 7854 5437 7870
rect 95 7730 152 7749
rect 95 7727 116 7730
rect 1 7712 116 7727
rect 134 7712 152 7730
rect 1 7689 152 7712
rect 1 7653 43 7689
rect 10316 7912 10472 7933
rect 10372 7911 10472 7912
rect 0 7652 100 7653
rect 0 7631 156 7652
rect 10429 7875 10471 7911
rect 10320 7852 10471 7875
rect 10320 7834 10338 7852
rect 10356 7837 10471 7852
rect 10356 7834 10377 7837
rect 10320 7815 10377 7834
rect 5035 7694 5096 7710
rect 5376 7709 5433 7728
rect 5376 7706 5397 7709
rect 5035 7690 5191 7694
rect 5035 7672 5055 7690
rect 5073 7672 5191 7690
rect 0 7613 118 7631
rect 136 7613 156 7631
rect 0 7609 156 7613
rect 95 7593 156 7609
rect 102 7529 159 7548
rect 102 7526 123 7529
rect 8 7511 123 7526
rect 141 7511 159 7529
rect 5035 7651 5191 7672
rect 5091 7650 5191 7651
rect 5282 7691 5397 7706
rect 5415 7691 5433 7709
rect 5282 7668 5433 7691
rect 5148 7614 5190 7650
rect 5282 7632 5324 7668
rect 5039 7591 5190 7614
rect 5039 7573 5057 7591
rect 5075 7576 5190 7591
rect 5281 7631 5381 7632
rect 5281 7610 5437 7631
rect 10316 7673 10377 7689
rect 10316 7669 10472 7673
rect 10316 7651 10336 7669
rect 10354 7651 10472 7669
rect 5281 7592 5399 7610
rect 5417 7592 5437 7610
rect 5281 7588 5437 7592
rect 5075 7573 5096 7576
rect 5039 7554 5096 7573
rect 5376 7572 5437 7588
rect 8 7488 159 7511
rect 8 7452 50 7488
rect 7 7451 107 7452
rect 7 7430 163 7451
rect 5383 7508 5440 7527
rect 5383 7505 5404 7508
rect 7 7412 125 7430
rect 143 7412 163 7430
rect 7 7408 163 7412
rect 102 7392 163 7408
rect 5033 7480 5094 7496
rect 5289 7490 5404 7505
rect 5422 7490 5440 7508
rect 10316 7630 10472 7651
rect 10372 7629 10472 7630
rect 10429 7593 10471 7629
rect 10320 7570 10471 7593
rect 10320 7552 10338 7570
rect 10356 7555 10471 7570
rect 10356 7552 10377 7555
rect 10320 7533 10377 7552
rect 5033 7476 5189 7480
rect 5033 7458 5053 7476
rect 5071 7458 5189 7476
rect 5033 7437 5189 7458
rect 5089 7436 5189 7437
rect 5289 7467 5440 7490
rect 5146 7400 5188 7436
rect 5289 7431 5331 7467
rect 5037 7377 5188 7400
rect 5288 7430 5388 7431
rect 5288 7409 5444 7430
rect 5288 7391 5406 7409
rect 5424 7391 5444 7409
rect 5288 7387 5444 7391
rect 5037 7359 5055 7377
rect 5073 7362 5188 7377
rect 5383 7371 5444 7387
rect 10314 7459 10375 7475
rect 10314 7455 10470 7459
rect 10314 7437 10334 7455
rect 10352 7437 10470 7455
rect 10314 7416 10470 7437
rect 10370 7415 10470 7416
rect 5073 7359 5094 7362
rect 5037 7340 5094 7359
rect 10427 7379 10469 7415
rect 10318 7356 10469 7379
rect 10318 7338 10336 7356
rect 10354 7341 10469 7356
rect 10354 7338 10375 7341
rect 10318 7319 10375 7338
rect 102 7245 159 7264
rect 102 7242 123 7245
rect 8 7227 123 7242
rect 141 7227 159 7245
rect 8 7204 159 7227
rect 8 7168 50 7204
rect 5383 7224 5440 7243
rect 5383 7221 5404 7224
rect 7 7167 107 7168
rect 7 7146 163 7167
rect 7 7128 125 7146
rect 143 7128 163 7146
rect 7 7124 163 7128
rect 102 7108 163 7124
rect 5033 7196 5094 7212
rect 5289 7206 5404 7221
rect 5422 7206 5440 7224
rect 5033 7192 5189 7196
rect 5033 7174 5053 7192
rect 5071 7174 5189 7192
rect 5033 7153 5189 7174
rect 5089 7152 5189 7153
rect 5289 7183 5440 7206
rect 5146 7116 5188 7152
rect 5289 7147 5331 7183
rect 5037 7093 5188 7116
rect 5288 7146 5388 7147
rect 5288 7125 5444 7146
rect 5288 7107 5406 7125
rect 5424 7107 5444 7125
rect 5288 7103 5444 7107
rect 100 7031 157 7050
rect 100 7028 121 7031
rect 6 7013 121 7028
rect 139 7013 157 7031
rect 6 6990 157 7013
rect 6 6954 48 6990
rect 5 6953 105 6954
rect 5 6932 161 6953
rect 5037 7075 5055 7093
rect 5073 7078 5188 7093
rect 5383 7087 5444 7103
rect 10314 7175 10375 7191
rect 10314 7171 10470 7175
rect 10314 7153 10334 7171
rect 10352 7153 10470 7171
rect 5073 7075 5094 7078
rect 5037 7056 5094 7075
rect 10314 7132 10470 7153
rect 10370 7131 10470 7132
rect 10427 7095 10469 7131
rect 10318 7072 10469 7095
rect 5040 6995 5101 7011
rect 5381 7010 5438 7029
rect 5381 7007 5402 7010
rect 5040 6991 5196 6995
rect 5040 6973 5060 6991
rect 5078 6973 5196 6991
rect 5 6914 123 6932
rect 141 6914 161 6932
rect 5 6910 161 6914
rect 100 6894 161 6910
rect 5040 6952 5196 6973
rect 5096 6951 5196 6952
rect 5287 6992 5402 7007
rect 5420 6992 5438 7010
rect 5287 6969 5438 6992
rect 5153 6915 5195 6951
rect 5287 6933 5329 6969
rect 5044 6892 5195 6915
rect 5044 6874 5062 6892
rect 5080 6877 5195 6892
rect 5286 6932 5386 6933
rect 5286 6911 5442 6932
rect 10318 7054 10336 7072
rect 10354 7057 10469 7072
rect 10354 7054 10375 7057
rect 10318 7035 10375 7054
rect 10321 6974 10382 6990
rect 10321 6970 10477 6974
rect 10321 6952 10341 6970
rect 10359 6952 10477 6970
rect 5286 6893 5404 6911
rect 5422 6893 5442 6911
rect 5286 6889 5442 6893
rect 5080 6874 5101 6877
rect 5044 6855 5101 6874
rect 5381 6873 5442 6889
rect 100 6749 157 6768
rect 100 6746 121 6749
rect 6 6731 121 6746
rect 139 6731 157 6749
rect 6 6708 157 6731
rect 6 6672 48 6708
rect 10321 6931 10477 6952
rect 10377 6930 10477 6931
rect 5 6671 105 6672
rect 5 6650 161 6671
rect 10434 6894 10476 6930
rect 10325 6871 10476 6894
rect 10325 6853 10343 6871
rect 10361 6856 10476 6871
rect 10361 6853 10382 6856
rect 10325 6834 10382 6853
rect 5040 6713 5101 6729
rect 5381 6728 5438 6747
rect 5381 6725 5402 6728
rect 5040 6709 5196 6713
rect 5040 6691 5060 6709
rect 5078 6691 5196 6709
rect 5 6632 123 6650
rect 141 6632 161 6650
rect 5 6628 161 6632
rect 100 6612 161 6628
rect 107 6548 164 6567
rect 107 6545 128 6548
rect 13 6530 128 6545
rect 146 6530 164 6548
rect 5040 6670 5196 6691
rect 5096 6669 5196 6670
rect 5287 6710 5402 6725
rect 5420 6710 5438 6728
rect 5287 6687 5438 6710
rect 5153 6633 5195 6669
rect 5287 6651 5329 6687
rect 5044 6610 5195 6633
rect 5044 6592 5062 6610
rect 5080 6595 5195 6610
rect 5286 6650 5386 6651
rect 5286 6629 5442 6650
rect 10321 6692 10382 6708
rect 10321 6688 10477 6692
rect 10321 6670 10341 6688
rect 10359 6670 10477 6688
rect 5286 6611 5404 6629
rect 5422 6611 5442 6629
rect 5286 6607 5442 6611
rect 5080 6592 5101 6595
rect 5044 6573 5101 6592
rect 5381 6591 5442 6607
rect 13 6507 164 6530
rect 13 6471 55 6507
rect 12 6470 112 6471
rect 12 6449 168 6470
rect 5388 6527 5445 6546
rect 5388 6524 5409 6527
rect 5038 6499 5099 6515
rect 5294 6509 5409 6524
rect 5427 6509 5445 6527
rect 10321 6649 10477 6670
rect 10377 6648 10477 6649
rect 10434 6612 10476 6648
rect 10325 6589 10476 6612
rect 10325 6571 10343 6589
rect 10361 6574 10476 6589
rect 10361 6571 10382 6574
rect 10325 6552 10382 6571
rect 5038 6495 5194 6499
rect 5038 6477 5058 6495
rect 5076 6477 5194 6495
rect 12 6431 130 6449
rect 148 6431 168 6449
rect 12 6427 168 6431
rect 107 6411 168 6427
rect 5038 6456 5194 6477
rect 5094 6455 5194 6456
rect 5294 6486 5445 6509
rect 5151 6419 5193 6455
rect 5294 6450 5336 6486
rect 5042 6396 5193 6419
rect 5293 6449 5393 6450
rect 5293 6428 5449 6449
rect 10319 6478 10380 6494
rect 10319 6474 10475 6478
rect 10319 6456 10339 6474
rect 10357 6456 10475 6474
rect 5293 6410 5411 6428
rect 5429 6410 5449 6428
rect 5293 6406 5449 6410
rect 109 6266 166 6285
rect 109 6263 130 6266
rect 15 6248 130 6263
rect 148 6248 166 6266
rect 5042 6378 5060 6396
rect 5078 6381 5193 6396
rect 5388 6390 5449 6406
rect 5078 6378 5099 6381
rect 5042 6359 5099 6378
rect 10319 6435 10475 6456
rect 10375 6434 10475 6435
rect 10432 6398 10474 6434
rect 10323 6375 10474 6398
rect 15 6225 166 6248
rect 15 6189 57 6225
rect 14 6188 114 6189
rect 14 6167 170 6188
rect 5390 6245 5447 6264
rect 5390 6242 5411 6245
rect 5040 6217 5101 6233
rect 5296 6227 5411 6242
rect 5429 6227 5447 6245
rect 10323 6357 10341 6375
rect 10359 6360 10474 6375
rect 10359 6357 10380 6360
rect 10323 6338 10380 6357
rect 5040 6213 5196 6217
rect 5040 6195 5060 6213
rect 5078 6195 5196 6213
rect 14 6149 132 6167
rect 150 6149 170 6167
rect 14 6145 170 6149
rect 109 6129 170 6145
rect 5040 6174 5196 6195
rect 5096 6173 5196 6174
rect 5296 6204 5447 6227
rect 5153 6137 5195 6173
rect 5296 6168 5338 6204
rect 5044 6114 5195 6137
rect 5295 6167 5395 6168
rect 5295 6146 5451 6167
rect 10321 6196 10382 6212
rect 10321 6192 10477 6196
rect 10321 6174 10341 6192
rect 10359 6174 10477 6192
rect 5295 6128 5413 6146
rect 5431 6128 5451 6146
rect 5295 6124 5451 6128
rect 107 6052 164 6071
rect 107 6049 128 6052
rect 13 6034 128 6049
rect 146 6034 164 6052
rect 13 6011 164 6034
rect 13 5975 55 6011
rect 12 5974 112 5975
rect 12 5953 168 5974
rect 5044 6096 5062 6114
rect 5080 6099 5195 6114
rect 5390 6108 5451 6124
rect 5080 6096 5101 6099
rect 5044 6077 5101 6096
rect 10321 6153 10477 6174
rect 10377 6152 10477 6153
rect 10434 6116 10476 6152
rect 10325 6093 10476 6116
rect 5047 6016 5108 6032
rect 5388 6031 5445 6050
rect 5388 6028 5409 6031
rect 5047 6012 5203 6016
rect 5047 5994 5067 6012
rect 5085 5994 5203 6012
rect 12 5935 130 5953
rect 148 5935 168 5953
rect 12 5931 168 5935
rect 107 5915 168 5931
rect 5047 5973 5203 5994
rect 5103 5972 5203 5973
rect 5294 6013 5409 6028
rect 5427 6013 5445 6031
rect 5294 5990 5445 6013
rect 5160 5936 5202 5972
rect 5294 5954 5336 5990
rect 5051 5913 5202 5936
rect 5051 5895 5069 5913
rect 5087 5898 5202 5913
rect 5293 5953 5393 5954
rect 5293 5932 5449 5953
rect 10325 6075 10343 6093
rect 10361 6078 10476 6093
rect 10361 6075 10382 6078
rect 10325 6056 10382 6075
rect 10328 5995 10389 6011
rect 10328 5991 10484 5995
rect 10328 5973 10348 5991
rect 10366 5973 10484 5991
rect 5293 5914 5411 5932
rect 5429 5914 5449 5932
rect 5293 5910 5449 5914
rect 5087 5895 5108 5898
rect 5051 5876 5108 5895
rect 5388 5894 5449 5910
rect 107 5770 164 5789
rect 107 5767 128 5770
rect 13 5752 128 5767
rect 146 5752 164 5770
rect 13 5729 164 5752
rect 13 5693 55 5729
rect 10328 5952 10484 5973
rect 10384 5951 10484 5952
rect 12 5692 112 5693
rect 12 5671 168 5692
rect 10441 5915 10483 5951
rect 10332 5892 10483 5915
rect 10332 5874 10350 5892
rect 10368 5877 10483 5892
rect 10368 5874 10389 5877
rect 10332 5855 10389 5874
rect 5047 5734 5108 5750
rect 5388 5749 5445 5768
rect 5388 5746 5409 5749
rect 5047 5730 5203 5734
rect 5047 5712 5067 5730
rect 5085 5712 5203 5730
rect 12 5653 130 5671
rect 148 5653 168 5671
rect 12 5649 168 5653
rect 107 5633 168 5649
rect 114 5569 171 5588
rect 114 5566 135 5569
rect 20 5551 135 5566
rect 153 5551 171 5569
rect 5047 5691 5203 5712
rect 5103 5690 5203 5691
rect 5294 5731 5409 5746
rect 5427 5731 5445 5749
rect 5294 5708 5445 5731
rect 5160 5654 5202 5690
rect 5294 5672 5336 5708
rect 5051 5631 5202 5654
rect 5051 5613 5069 5631
rect 5087 5616 5202 5631
rect 5293 5671 5393 5672
rect 5293 5650 5449 5671
rect 10328 5713 10389 5729
rect 10328 5709 10484 5713
rect 10328 5691 10348 5709
rect 10366 5691 10484 5709
rect 5293 5632 5411 5650
rect 5429 5632 5449 5650
rect 5293 5628 5449 5632
rect 5087 5613 5108 5616
rect 5051 5594 5108 5613
rect 5388 5612 5449 5628
rect 20 5528 171 5551
rect 20 5492 62 5528
rect 19 5491 119 5492
rect 19 5470 175 5491
rect 5395 5548 5452 5567
rect 5395 5545 5416 5548
rect 19 5452 137 5470
rect 155 5452 175 5470
rect 19 5448 175 5452
rect 114 5432 175 5448
rect 5045 5520 5106 5536
rect 5301 5530 5416 5545
rect 5434 5530 5452 5548
rect 10328 5670 10484 5691
rect 10384 5669 10484 5670
rect 10441 5633 10483 5669
rect 10332 5610 10483 5633
rect 10332 5592 10350 5610
rect 10368 5595 10483 5610
rect 10368 5592 10389 5595
rect 10332 5573 10389 5592
rect 5045 5516 5201 5520
rect 5045 5498 5065 5516
rect 5083 5498 5201 5516
rect 5045 5477 5201 5498
rect 5101 5476 5201 5477
rect 5301 5507 5452 5530
rect 5158 5440 5200 5476
rect 5301 5471 5343 5507
rect 5049 5417 5200 5440
rect 5300 5470 5400 5471
rect 5300 5449 5456 5470
rect 5300 5431 5418 5449
rect 5436 5431 5456 5449
rect 5300 5427 5456 5431
rect 5049 5399 5067 5417
rect 5085 5402 5200 5417
rect 5395 5411 5456 5427
rect 10326 5499 10387 5515
rect 10326 5495 10482 5499
rect 10326 5477 10346 5495
rect 10364 5477 10482 5495
rect 10326 5456 10482 5477
rect 10382 5455 10482 5456
rect 5085 5399 5106 5402
rect 5049 5380 5106 5399
rect 10439 5419 10481 5455
rect 10330 5396 10481 5419
rect 10330 5378 10348 5396
rect 10366 5381 10481 5396
rect 10366 5378 10387 5381
rect 10330 5359 10387 5378
rect 114 5285 171 5304
rect 114 5282 135 5285
rect 20 5267 135 5282
rect 153 5267 171 5285
rect 20 5244 171 5267
rect 20 5208 62 5244
rect 5395 5264 5452 5283
rect 5395 5261 5416 5264
rect 19 5207 119 5208
rect 19 5186 175 5207
rect 19 5168 137 5186
rect 155 5168 175 5186
rect 19 5164 175 5168
rect 114 5148 175 5164
rect 5045 5236 5106 5252
rect 5301 5246 5416 5261
rect 5434 5246 5452 5264
rect 5045 5232 5201 5236
rect 5045 5214 5065 5232
rect 5083 5214 5201 5232
rect 5045 5193 5201 5214
rect 5101 5192 5201 5193
rect 5301 5223 5452 5246
rect 5158 5156 5200 5192
rect 5301 5187 5343 5223
rect 5049 5133 5200 5156
rect 5300 5186 5400 5187
rect 5300 5165 5456 5186
rect 5300 5147 5418 5165
rect 5436 5147 5456 5165
rect 5300 5143 5456 5147
rect 112 5071 169 5090
rect 112 5068 133 5071
rect 18 5053 133 5068
rect 151 5053 169 5071
rect 18 5030 169 5053
rect 18 4994 60 5030
rect 17 4993 117 4994
rect 17 4972 173 4993
rect 5049 5115 5067 5133
rect 5085 5118 5200 5133
rect 5395 5127 5456 5143
rect 10326 5215 10387 5231
rect 10326 5211 10482 5215
rect 10326 5193 10346 5211
rect 10364 5193 10482 5211
rect 5085 5115 5106 5118
rect 5049 5096 5106 5115
rect 10326 5172 10482 5193
rect 10382 5171 10482 5172
rect 10439 5135 10481 5171
rect 10330 5112 10481 5135
rect 5052 5035 5113 5051
rect 5393 5050 5450 5069
rect 5393 5047 5414 5050
rect 5052 5031 5208 5035
rect 5052 5013 5072 5031
rect 5090 5013 5208 5031
rect 17 4954 135 4972
rect 153 4954 173 4972
rect 17 4950 173 4954
rect 112 4934 173 4950
rect 5052 4992 5208 5013
rect 5108 4991 5208 4992
rect 5299 5032 5414 5047
rect 5432 5032 5450 5050
rect 5299 5009 5450 5032
rect 5165 4955 5207 4991
rect 5299 4973 5341 5009
rect 5056 4932 5207 4955
rect 5056 4914 5074 4932
rect 5092 4917 5207 4932
rect 5298 4972 5398 4973
rect 5298 4951 5454 4972
rect 10330 5094 10348 5112
rect 10366 5097 10481 5112
rect 10366 5094 10387 5097
rect 10330 5075 10387 5094
rect 10333 5014 10394 5030
rect 10333 5010 10489 5014
rect 10333 4992 10353 5010
rect 10371 4992 10489 5010
rect 5298 4933 5416 4951
rect 5434 4933 5454 4951
rect 5298 4929 5454 4933
rect 5092 4914 5113 4917
rect 5056 4895 5113 4914
rect 5393 4913 5454 4929
rect 112 4789 169 4808
rect 112 4786 133 4789
rect 18 4771 133 4786
rect 151 4771 169 4789
rect 18 4748 169 4771
rect 18 4712 60 4748
rect 10333 4971 10489 4992
rect 10389 4970 10489 4971
rect 17 4711 117 4712
rect 17 4690 173 4711
rect 10446 4934 10488 4970
rect 10337 4911 10488 4934
rect 10337 4893 10355 4911
rect 10373 4896 10488 4911
rect 10373 4893 10394 4896
rect 10337 4874 10394 4893
rect 5052 4753 5113 4769
rect 5393 4768 5450 4787
rect 5393 4765 5414 4768
rect 5052 4749 5208 4753
rect 5052 4731 5072 4749
rect 5090 4731 5208 4749
rect 17 4672 135 4690
rect 153 4672 173 4690
rect 17 4668 173 4672
rect 112 4652 173 4668
rect 119 4588 176 4607
rect 119 4585 140 4588
rect 25 4570 140 4585
rect 158 4570 176 4588
rect 5052 4710 5208 4731
rect 5108 4709 5208 4710
rect 5299 4750 5414 4765
rect 5432 4750 5450 4768
rect 5299 4727 5450 4750
rect 5165 4673 5207 4709
rect 5299 4691 5341 4727
rect 5056 4650 5207 4673
rect 5056 4632 5074 4650
rect 5092 4635 5207 4650
rect 5298 4690 5398 4691
rect 5298 4669 5454 4690
rect 10333 4732 10394 4748
rect 10333 4728 10489 4732
rect 10333 4710 10353 4728
rect 10371 4710 10489 4728
rect 5298 4651 5416 4669
rect 5434 4651 5454 4669
rect 5298 4647 5454 4651
rect 5092 4632 5113 4635
rect 5056 4613 5113 4632
rect 5393 4631 5454 4647
rect 25 4547 176 4570
rect 25 4511 67 4547
rect 24 4510 124 4511
rect 24 4489 180 4510
rect 5400 4567 5457 4586
rect 5400 4564 5421 4567
rect 5050 4539 5111 4555
rect 5306 4549 5421 4564
rect 5439 4549 5457 4567
rect 10333 4689 10489 4710
rect 10389 4688 10489 4689
rect 10446 4652 10488 4688
rect 10337 4629 10488 4652
rect 10337 4611 10355 4629
rect 10373 4614 10488 4629
rect 10373 4611 10394 4614
rect 10337 4592 10394 4611
rect 24 4471 142 4489
rect 160 4471 180 4489
rect 24 4467 180 4471
rect 119 4451 180 4467
rect 5050 4535 5206 4539
rect 5050 4517 5070 4535
rect 5088 4517 5206 4535
rect 5050 4496 5206 4517
rect 5106 4495 5206 4496
rect 5306 4526 5457 4549
rect 117 4309 174 4328
rect 117 4306 138 4309
rect 23 4291 138 4306
rect 156 4291 174 4309
rect 23 4268 174 4291
rect 23 4232 65 4268
rect 5163 4459 5205 4495
rect 5306 4490 5348 4526
rect 5054 4436 5205 4459
rect 5305 4489 5405 4490
rect 5305 4468 5461 4489
rect 10331 4518 10392 4534
rect 5305 4450 5423 4468
rect 5441 4450 5461 4468
rect 5305 4446 5461 4450
rect 5054 4418 5072 4436
rect 5090 4421 5205 4436
rect 5400 4430 5461 4446
rect 10331 4514 10487 4518
rect 10331 4496 10351 4514
rect 10369 4496 10487 4514
rect 10331 4475 10487 4496
rect 10387 4474 10487 4475
rect 5090 4418 5111 4421
rect 5054 4399 5111 4418
rect 5398 4288 5455 4307
rect 5398 4285 5419 4288
rect 22 4231 122 4232
rect 22 4210 178 4231
rect 22 4192 140 4210
rect 158 4192 178 4210
rect 22 4188 178 4192
rect 5048 4260 5109 4276
rect 5304 4270 5419 4285
rect 5437 4270 5455 4288
rect 5048 4256 5204 4260
rect 5048 4238 5068 4256
rect 5086 4238 5204 4256
rect 117 4172 178 4188
rect 5048 4217 5204 4238
rect 5104 4216 5204 4217
rect 5304 4247 5455 4270
rect 5161 4180 5203 4216
rect 5304 4211 5346 4247
rect 10444 4438 10486 4474
rect 10335 4415 10486 4438
rect 10335 4397 10353 4415
rect 10371 4400 10486 4415
rect 10371 4397 10392 4400
rect 10335 4378 10392 4397
rect 5052 4157 5203 4180
rect 5303 4210 5403 4211
rect 5303 4189 5459 4210
rect 5303 4171 5421 4189
rect 5439 4171 5459 4189
rect 5303 4167 5459 4171
rect 10329 4239 10390 4255
rect 10329 4235 10485 4239
rect 10329 4217 10349 4235
rect 10367 4217 10485 4235
rect 115 4095 172 4114
rect 115 4092 136 4095
rect 21 4077 136 4092
rect 154 4077 172 4095
rect 21 4054 172 4077
rect 21 4018 63 4054
rect 20 4017 120 4018
rect 20 3996 176 4017
rect 5052 4139 5070 4157
rect 5088 4142 5203 4157
rect 5398 4151 5459 4167
rect 5088 4139 5109 4142
rect 5052 4120 5109 4139
rect 10329 4196 10485 4217
rect 10385 4195 10485 4196
rect 10442 4159 10484 4195
rect 10333 4136 10484 4159
rect 5055 4059 5116 4075
rect 5396 4074 5453 4093
rect 5396 4071 5417 4074
rect 5055 4055 5211 4059
rect 5055 4037 5075 4055
rect 5093 4037 5211 4055
rect 20 3978 138 3996
rect 156 3978 176 3996
rect 20 3974 176 3978
rect 115 3958 176 3974
rect 5055 4016 5211 4037
rect 5111 4015 5211 4016
rect 5302 4056 5417 4071
rect 5435 4056 5453 4074
rect 5302 4033 5453 4056
rect 5168 3979 5210 4015
rect 5302 3997 5344 4033
rect 5059 3956 5210 3979
rect 5059 3938 5077 3956
rect 5095 3941 5210 3956
rect 5301 3996 5401 3997
rect 5301 3975 5457 3996
rect 10333 4118 10351 4136
rect 10369 4121 10484 4136
rect 10369 4118 10390 4121
rect 10333 4099 10390 4118
rect 10336 4038 10397 4054
rect 10336 4034 10492 4038
rect 10336 4016 10356 4034
rect 10374 4016 10492 4034
rect 5301 3957 5419 3975
rect 5437 3957 5457 3975
rect 5301 3953 5457 3957
rect 5095 3938 5116 3941
rect 5059 3919 5116 3938
rect 5396 3937 5457 3953
rect 115 3813 172 3832
rect 115 3810 136 3813
rect 21 3795 136 3810
rect 154 3795 172 3813
rect 21 3772 172 3795
rect 21 3736 63 3772
rect 10336 3995 10492 4016
rect 10392 3994 10492 3995
rect 20 3735 120 3736
rect 20 3714 176 3735
rect 10449 3958 10491 3994
rect 10340 3935 10491 3958
rect 10340 3917 10358 3935
rect 10376 3920 10491 3935
rect 10376 3917 10397 3920
rect 10340 3898 10397 3917
rect 5055 3777 5116 3793
rect 5396 3792 5453 3811
rect 5396 3789 5417 3792
rect 5055 3773 5211 3777
rect 5055 3755 5075 3773
rect 5093 3755 5211 3773
rect 20 3696 138 3714
rect 156 3696 176 3714
rect 20 3692 176 3696
rect 115 3676 176 3692
rect 122 3612 179 3631
rect 122 3609 143 3612
rect 28 3594 143 3609
rect 161 3594 179 3612
rect 5055 3734 5211 3755
rect 5111 3733 5211 3734
rect 5302 3774 5417 3789
rect 5435 3774 5453 3792
rect 5302 3751 5453 3774
rect 5168 3697 5210 3733
rect 5302 3715 5344 3751
rect 5059 3674 5210 3697
rect 5059 3656 5077 3674
rect 5095 3659 5210 3674
rect 5301 3714 5401 3715
rect 5301 3693 5457 3714
rect 10336 3756 10397 3772
rect 10336 3752 10492 3756
rect 10336 3734 10356 3752
rect 10374 3734 10492 3752
rect 5301 3675 5419 3693
rect 5437 3675 5457 3693
rect 5301 3671 5457 3675
rect 5095 3656 5116 3659
rect 5059 3637 5116 3656
rect 5396 3655 5457 3671
rect 28 3571 179 3594
rect 28 3535 70 3571
rect 27 3534 127 3535
rect 27 3513 183 3534
rect 5403 3591 5460 3610
rect 5403 3588 5424 3591
rect 27 3495 145 3513
rect 163 3495 183 3513
rect 27 3491 183 3495
rect 122 3475 183 3491
rect 5053 3563 5114 3579
rect 5309 3573 5424 3588
rect 5442 3573 5460 3591
rect 10336 3713 10492 3734
rect 10392 3712 10492 3713
rect 10449 3676 10491 3712
rect 10340 3653 10491 3676
rect 10340 3635 10358 3653
rect 10376 3638 10491 3653
rect 10376 3635 10397 3638
rect 10340 3616 10397 3635
rect 5053 3559 5209 3563
rect 5053 3541 5073 3559
rect 5091 3541 5209 3559
rect 5053 3520 5209 3541
rect 5109 3519 5209 3520
rect 5309 3550 5460 3573
rect 5166 3483 5208 3519
rect 5309 3514 5351 3550
rect 5057 3460 5208 3483
rect 5308 3513 5408 3514
rect 5308 3492 5464 3513
rect 5308 3474 5426 3492
rect 5444 3474 5464 3492
rect 5308 3470 5464 3474
rect 5057 3442 5075 3460
rect 5093 3445 5208 3460
rect 5403 3454 5464 3470
rect 10334 3542 10395 3558
rect 10334 3538 10490 3542
rect 10334 3520 10354 3538
rect 10372 3520 10490 3538
rect 10334 3499 10490 3520
rect 10390 3498 10490 3499
rect 5093 3442 5114 3445
rect 5057 3423 5114 3442
rect 10447 3462 10489 3498
rect 10338 3439 10489 3462
rect 10338 3421 10356 3439
rect 10374 3424 10489 3439
rect 10374 3421 10395 3424
rect 10338 3402 10395 3421
rect 122 3328 179 3347
rect 122 3325 143 3328
rect 28 3310 143 3325
rect 161 3310 179 3328
rect 28 3287 179 3310
rect 28 3251 70 3287
rect 5403 3307 5460 3326
rect 5403 3304 5424 3307
rect 27 3250 127 3251
rect 27 3229 183 3250
rect 27 3211 145 3229
rect 163 3211 183 3229
rect 27 3207 183 3211
rect 122 3191 183 3207
rect 5053 3279 5114 3295
rect 5309 3289 5424 3304
rect 5442 3289 5460 3307
rect 5053 3275 5209 3279
rect 5053 3257 5073 3275
rect 5091 3257 5209 3275
rect 5053 3236 5209 3257
rect 5109 3235 5209 3236
rect 5309 3266 5460 3289
rect 5166 3199 5208 3235
rect 5309 3230 5351 3266
rect 5057 3176 5208 3199
rect 5308 3229 5408 3230
rect 5308 3208 5464 3229
rect 5308 3190 5426 3208
rect 5444 3190 5464 3208
rect 5308 3186 5464 3190
rect 120 3114 177 3133
rect 120 3111 141 3114
rect 26 3096 141 3111
rect 159 3096 177 3114
rect 26 3073 177 3096
rect 26 3037 68 3073
rect 25 3036 125 3037
rect 25 3015 181 3036
rect 5057 3158 5075 3176
rect 5093 3161 5208 3176
rect 5403 3170 5464 3186
rect 10334 3258 10395 3274
rect 10334 3254 10490 3258
rect 10334 3236 10354 3254
rect 10372 3236 10490 3254
rect 5093 3158 5114 3161
rect 5057 3139 5114 3158
rect 10334 3215 10490 3236
rect 10390 3214 10490 3215
rect 10447 3178 10489 3214
rect 10338 3155 10489 3178
rect 5060 3078 5121 3094
rect 5401 3093 5458 3112
rect 5401 3090 5422 3093
rect 5060 3074 5216 3078
rect 5060 3056 5080 3074
rect 5098 3056 5216 3074
rect 25 2997 143 3015
rect 161 2997 181 3015
rect 25 2993 181 2997
rect 120 2977 181 2993
rect 5060 3035 5216 3056
rect 5116 3034 5216 3035
rect 5307 3075 5422 3090
rect 5440 3075 5458 3093
rect 5307 3052 5458 3075
rect 5173 2998 5215 3034
rect 5307 3016 5349 3052
rect 5064 2975 5215 2998
rect 5064 2957 5082 2975
rect 5100 2960 5215 2975
rect 5306 3015 5406 3016
rect 5306 2994 5462 3015
rect 10338 3137 10356 3155
rect 10374 3140 10489 3155
rect 10374 3137 10395 3140
rect 10338 3118 10395 3137
rect 10341 3057 10402 3073
rect 10341 3053 10497 3057
rect 10341 3035 10361 3053
rect 10379 3035 10497 3053
rect 5306 2976 5424 2994
rect 5442 2976 5462 2994
rect 5306 2972 5462 2976
rect 5100 2957 5121 2960
rect 5064 2938 5121 2957
rect 5401 2956 5462 2972
rect 120 2832 177 2851
rect 120 2829 141 2832
rect 26 2814 141 2829
rect 159 2814 177 2832
rect 26 2791 177 2814
rect 26 2755 68 2791
rect 10341 3014 10497 3035
rect 10397 3013 10497 3014
rect 25 2754 125 2755
rect 25 2733 181 2754
rect 10454 2977 10496 3013
rect 10345 2954 10496 2977
rect 10345 2936 10363 2954
rect 10381 2939 10496 2954
rect 10381 2936 10402 2939
rect 10345 2917 10402 2936
rect 5060 2796 5121 2812
rect 5401 2811 5458 2830
rect 5401 2808 5422 2811
rect 5060 2792 5216 2796
rect 5060 2774 5080 2792
rect 5098 2774 5216 2792
rect 25 2715 143 2733
rect 161 2715 181 2733
rect 25 2711 181 2715
rect 120 2695 181 2711
rect 127 2631 184 2650
rect 127 2628 148 2631
rect 33 2613 148 2628
rect 166 2613 184 2631
rect 5060 2753 5216 2774
rect 5116 2752 5216 2753
rect 5307 2793 5422 2808
rect 5440 2793 5458 2811
rect 5307 2770 5458 2793
rect 5173 2716 5215 2752
rect 5307 2734 5349 2770
rect 5064 2693 5215 2716
rect 5064 2675 5082 2693
rect 5100 2678 5215 2693
rect 5306 2733 5406 2734
rect 5306 2712 5462 2733
rect 10341 2775 10402 2791
rect 10341 2771 10497 2775
rect 10341 2753 10361 2771
rect 10379 2753 10497 2771
rect 5306 2694 5424 2712
rect 5442 2694 5462 2712
rect 5306 2690 5462 2694
rect 5100 2675 5121 2678
rect 5064 2656 5121 2675
rect 5401 2674 5462 2690
rect 33 2590 184 2613
rect 33 2554 75 2590
rect 32 2553 132 2554
rect 32 2532 188 2553
rect 5408 2610 5465 2629
rect 5408 2607 5429 2610
rect 5058 2582 5119 2598
rect 5314 2592 5429 2607
rect 5447 2592 5465 2610
rect 10341 2732 10497 2753
rect 10397 2731 10497 2732
rect 10454 2695 10496 2731
rect 10345 2672 10496 2695
rect 10345 2654 10363 2672
rect 10381 2657 10496 2672
rect 10381 2654 10402 2657
rect 10345 2635 10402 2654
rect 5058 2578 5214 2582
rect 5058 2560 5078 2578
rect 5096 2560 5214 2578
rect 32 2514 150 2532
rect 168 2514 188 2532
rect 32 2510 188 2514
rect 127 2494 188 2510
rect 5058 2539 5214 2560
rect 5114 2538 5214 2539
rect 5314 2569 5465 2592
rect 5171 2502 5213 2538
rect 5314 2533 5356 2569
rect 5062 2479 5213 2502
rect 5313 2532 5413 2533
rect 5313 2511 5469 2532
rect 10339 2561 10400 2577
rect 10339 2557 10495 2561
rect 10339 2539 10359 2557
rect 10377 2539 10495 2557
rect 5313 2493 5431 2511
rect 5449 2493 5469 2511
rect 5313 2489 5469 2493
rect 129 2349 186 2368
rect 129 2346 150 2349
rect 35 2331 150 2346
rect 168 2331 186 2349
rect 5062 2461 5080 2479
rect 5098 2464 5213 2479
rect 5408 2473 5469 2489
rect 5098 2461 5119 2464
rect 5062 2442 5119 2461
rect 10339 2518 10495 2539
rect 10395 2517 10495 2518
rect 10452 2481 10494 2517
rect 10343 2458 10494 2481
rect 35 2308 186 2331
rect 35 2272 77 2308
rect 34 2271 134 2272
rect 34 2250 190 2271
rect 5410 2328 5467 2347
rect 5410 2325 5431 2328
rect 5060 2300 5121 2316
rect 5316 2310 5431 2325
rect 5449 2310 5467 2328
rect 10343 2440 10361 2458
rect 10379 2443 10494 2458
rect 10379 2440 10400 2443
rect 10343 2421 10400 2440
rect 5060 2296 5216 2300
rect 5060 2278 5080 2296
rect 5098 2278 5216 2296
rect 34 2232 152 2250
rect 170 2232 190 2250
rect 34 2228 190 2232
rect 129 2212 190 2228
rect 5060 2257 5216 2278
rect 5116 2256 5216 2257
rect 5316 2287 5467 2310
rect 5173 2220 5215 2256
rect 5316 2251 5358 2287
rect 5064 2197 5215 2220
rect 5315 2250 5415 2251
rect 5315 2229 5471 2250
rect 10341 2279 10402 2295
rect 10341 2275 10497 2279
rect 10341 2257 10361 2275
rect 10379 2257 10497 2275
rect 5315 2211 5433 2229
rect 5451 2211 5471 2229
rect 5315 2207 5471 2211
rect 127 2135 184 2154
rect 127 2132 148 2135
rect 33 2117 148 2132
rect 166 2117 184 2135
rect 33 2094 184 2117
rect 33 2058 75 2094
rect 32 2057 132 2058
rect 32 2036 188 2057
rect 5064 2179 5082 2197
rect 5100 2182 5215 2197
rect 5410 2191 5471 2207
rect 5100 2179 5121 2182
rect 5064 2160 5121 2179
rect 10341 2236 10497 2257
rect 10397 2235 10497 2236
rect 10454 2199 10496 2235
rect 10345 2176 10496 2199
rect 5067 2099 5128 2115
rect 5408 2114 5465 2133
rect 5408 2111 5429 2114
rect 5067 2095 5223 2099
rect 5067 2077 5087 2095
rect 5105 2077 5223 2095
rect 32 2018 150 2036
rect 168 2018 188 2036
rect 32 2014 188 2018
rect 127 1998 188 2014
rect 5067 2056 5223 2077
rect 5123 2055 5223 2056
rect 5314 2096 5429 2111
rect 5447 2096 5465 2114
rect 5314 2073 5465 2096
rect 5180 2019 5222 2055
rect 5314 2037 5356 2073
rect 5071 1996 5222 2019
rect 5071 1978 5089 1996
rect 5107 1981 5222 1996
rect 5313 2036 5413 2037
rect 5313 2015 5469 2036
rect 10345 2158 10363 2176
rect 10381 2161 10496 2176
rect 10381 2158 10402 2161
rect 10345 2139 10402 2158
rect 10348 2078 10409 2094
rect 10348 2074 10504 2078
rect 10348 2056 10368 2074
rect 10386 2056 10504 2074
rect 5313 1997 5431 2015
rect 5449 1997 5469 2015
rect 5313 1993 5469 1997
rect 5107 1978 5128 1981
rect 5071 1959 5128 1978
rect 5408 1977 5469 1993
rect 127 1853 184 1872
rect 127 1850 148 1853
rect 33 1835 148 1850
rect 166 1835 184 1853
rect 33 1812 184 1835
rect 33 1776 75 1812
rect 10348 2035 10504 2056
rect 10404 2034 10504 2035
rect 32 1775 132 1776
rect 32 1754 188 1775
rect 10461 1998 10503 2034
rect 10352 1975 10503 1998
rect 10352 1957 10370 1975
rect 10388 1960 10503 1975
rect 10388 1957 10409 1960
rect 10352 1938 10409 1957
rect 5067 1817 5128 1833
rect 5408 1832 5465 1851
rect 5408 1829 5429 1832
rect 5067 1813 5223 1817
rect 5067 1795 5087 1813
rect 5105 1795 5223 1813
rect 32 1736 150 1754
rect 168 1736 188 1754
rect 32 1732 188 1736
rect 127 1716 188 1732
rect 134 1652 191 1671
rect 134 1649 155 1652
rect 40 1634 155 1649
rect 173 1634 191 1652
rect 5067 1774 5223 1795
rect 5123 1773 5223 1774
rect 5314 1814 5429 1829
rect 5447 1814 5465 1832
rect 5314 1791 5465 1814
rect 5180 1737 5222 1773
rect 5314 1755 5356 1791
rect 5071 1714 5222 1737
rect 5071 1696 5089 1714
rect 5107 1699 5222 1714
rect 5313 1754 5413 1755
rect 5313 1733 5469 1754
rect 10348 1796 10409 1812
rect 10348 1792 10504 1796
rect 10348 1774 10368 1792
rect 10386 1774 10504 1792
rect 5313 1715 5431 1733
rect 5449 1715 5469 1733
rect 5313 1711 5469 1715
rect 5107 1696 5128 1699
rect 5071 1677 5128 1696
rect 5408 1695 5469 1711
rect 40 1611 191 1634
rect 40 1575 82 1611
rect 39 1574 139 1575
rect 39 1553 195 1574
rect 5415 1631 5472 1650
rect 5415 1628 5436 1631
rect 39 1535 157 1553
rect 175 1535 195 1553
rect 39 1531 195 1535
rect 134 1515 195 1531
rect 5065 1603 5126 1619
rect 5321 1613 5436 1628
rect 5454 1613 5472 1631
rect 10348 1753 10504 1774
rect 10404 1752 10504 1753
rect 10461 1716 10503 1752
rect 10352 1693 10503 1716
rect 10352 1675 10370 1693
rect 10388 1678 10503 1693
rect 10388 1675 10409 1678
rect 10352 1656 10409 1675
rect 5065 1599 5221 1603
rect 5065 1581 5085 1599
rect 5103 1581 5221 1599
rect 5065 1560 5221 1581
rect 5121 1559 5221 1560
rect 5321 1590 5472 1613
rect 5178 1523 5220 1559
rect 5321 1554 5363 1590
rect 5069 1500 5220 1523
rect 5320 1553 5420 1554
rect 5320 1532 5476 1553
rect 5320 1514 5438 1532
rect 5456 1514 5476 1532
rect 5320 1510 5476 1514
rect 5069 1482 5087 1500
rect 5105 1485 5220 1500
rect 5415 1494 5476 1510
rect 10346 1582 10407 1598
rect 10346 1578 10502 1582
rect 10346 1560 10366 1578
rect 10384 1560 10502 1578
rect 10346 1539 10502 1560
rect 10402 1538 10502 1539
rect 5105 1482 5126 1485
rect 5069 1463 5126 1482
rect 10459 1502 10501 1538
rect 10350 1479 10501 1502
rect 10350 1461 10368 1479
rect 10386 1464 10501 1479
rect 10386 1461 10407 1464
rect 10350 1442 10407 1461
rect 134 1368 191 1387
rect 134 1365 155 1368
rect 40 1350 155 1365
rect 173 1350 191 1368
rect 40 1327 191 1350
rect 40 1291 82 1327
rect 5415 1347 5472 1366
rect 5415 1344 5436 1347
rect 39 1290 139 1291
rect 39 1269 195 1290
rect 39 1251 157 1269
rect 175 1251 195 1269
rect 39 1247 195 1251
rect 134 1231 195 1247
rect 5065 1319 5126 1335
rect 5321 1329 5436 1344
rect 5454 1329 5472 1347
rect 5065 1315 5221 1319
rect 5065 1297 5085 1315
rect 5103 1297 5221 1315
rect 5065 1276 5221 1297
rect 5121 1275 5221 1276
rect 5321 1306 5472 1329
rect 5178 1239 5220 1275
rect 5321 1270 5363 1306
rect 5069 1216 5220 1239
rect 5320 1269 5420 1270
rect 5320 1248 5476 1269
rect 5320 1230 5438 1248
rect 5456 1230 5476 1248
rect 5320 1226 5476 1230
rect 132 1154 189 1173
rect 132 1151 153 1154
rect 38 1136 153 1151
rect 171 1136 189 1154
rect 38 1113 189 1136
rect 38 1077 80 1113
rect 37 1076 137 1077
rect 37 1055 193 1076
rect 5069 1198 5087 1216
rect 5105 1201 5220 1216
rect 5415 1210 5476 1226
rect 10346 1298 10407 1314
rect 10346 1294 10502 1298
rect 10346 1276 10366 1294
rect 10384 1276 10502 1294
rect 5105 1198 5126 1201
rect 5069 1179 5126 1198
rect 10346 1255 10502 1276
rect 10402 1254 10502 1255
rect 10459 1218 10501 1254
rect 10350 1195 10501 1218
rect 5072 1118 5133 1134
rect 5413 1133 5470 1152
rect 5413 1130 5434 1133
rect 5072 1114 5228 1118
rect 5072 1096 5092 1114
rect 5110 1096 5228 1114
rect 37 1037 155 1055
rect 173 1037 193 1055
rect 37 1033 193 1037
rect 132 1017 193 1033
rect 5072 1075 5228 1096
rect 5128 1074 5228 1075
rect 5319 1115 5434 1130
rect 5452 1115 5470 1133
rect 5319 1092 5470 1115
rect 5185 1038 5227 1074
rect 5319 1056 5361 1092
rect 5076 1015 5227 1038
rect 5076 997 5094 1015
rect 5112 1000 5227 1015
rect 5318 1055 5418 1056
rect 5318 1034 5474 1055
rect 10350 1177 10368 1195
rect 10386 1180 10501 1195
rect 10386 1177 10407 1180
rect 10350 1158 10407 1177
rect 10353 1097 10414 1113
rect 10353 1093 10509 1097
rect 10353 1075 10373 1093
rect 10391 1075 10509 1093
rect 5318 1016 5436 1034
rect 5454 1016 5474 1034
rect 5318 1012 5474 1016
rect 5112 997 5133 1000
rect 5076 978 5133 997
rect 5413 996 5474 1012
rect 132 872 189 891
rect 132 869 153 872
rect 38 854 153 869
rect 171 854 189 872
rect 38 831 189 854
rect 38 795 80 831
rect 10353 1054 10509 1075
rect 10409 1053 10509 1054
rect 37 794 137 795
rect 37 773 193 794
rect 10466 1017 10508 1053
rect 10357 994 10508 1017
rect 10357 976 10375 994
rect 10393 979 10508 994
rect 10393 976 10414 979
rect 10357 957 10414 976
rect 5072 836 5133 852
rect 5413 851 5470 870
rect 5413 848 5434 851
rect 5072 832 5228 836
rect 5072 814 5092 832
rect 5110 814 5228 832
rect 37 755 155 773
rect 173 755 193 773
rect 37 751 193 755
rect 132 735 193 751
rect 139 671 196 690
rect 139 668 160 671
rect 45 653 160 668
rect 178 653 196 671
rect 5072 793 5228 814
rect 5128 792 5228 793
rect 5319 833 5434 848
rect 5452 833 5470 851
rect 5319 810 5470 833
rect 5185 756 5227 792
rect 5319 774 5361 810
rect 5076 733 5227 756
rect 5076 715 5094 733
rect 5112 718 5227 733
rect 5318 773 5418 774
rect 5318 752 5474 773
rect 10353 815 10414 831
rect 10353 811 10509 815
rect 10353 793 10373 811
rect 10391 793 10509 811
rect 5318 734 5436 752
rect 5454 734 5474 752
rect 5318 730 5474 734
rect 5112 715 5133 718
rect 5076 696 5133 715
rect 5413 714 5474 730
rect 45 630 196 653
rect 45 594 87 630
rect 44 593 144 594
rect 44 572 200 593
rect 5420 650 5477 669
rect 5420 647 5441 650
rect 5070 622 5131 638
rect 5326 632 5441 647
rect 5459 632 5477 650
rect 10353 772 10509 793
rect 10409 771 10509 772
rect 10466 735 10508 771
rect 10357 712 10508 735
rect 10357 694 10375 712
rect 10393 697 10508 712
rect 10393 694 10414 697
rect 10357 675 10414 694
rect 5070 618 5226 622
rect 5070 600 5090 618
rect 5108 600 5226 618
rect 44 554 162 572
rect 180 554 200 572
rect 44 550 200 554
rect 139 534 200 550
rect 5070 579 5226 600
rect 5126 578 5226 579
rect 5326 609 5477 632
rect 5183 542 5225 578
rect 5326 573 5368 609
rect 5074 519 5225 542
rect 5325 572 5425 573
rect 5325 551 5481 572
rect 10351 601 10412 617
rect 10351 597 10507 601
rect 10351 579 10371 597
rect 10389 579 10507 597
rect 5325 533 5443 551
rect 5461 533 5481 551
rect 5325 529 5481 533
rect 5074 501 5092 519
rect 5110 504 5225 519
rect 5420 513 5481 529
rect 10351 558 10507 579
rect 10407 557 10507 558
rect 10464 521 10506 557
rect 5110 501 5131 504
rect 5074 482 5131 501
rect 10355 498 10506 521
rect 10355 480 10373 498
rect 10391 483 10506 498
rect 10391 480 10412 483
rect 10355 461 10412 480
<< locali >>
rect 110 8235 145 8283
rect 5038 8277 5434 8283
rect 4449 8259 5434 8277
rect 108 8226 145 8235
rect 108 8208 118 8226
rect 136 8208 145 8226
rect 108 8198 145 8208
rect 4031 8242 4199 8243
rect 4450 8242 4474 8259
rect 5038 8251 5434 8259
rect 10319 8256 10357 8262
rect 4031 8216 4475 8242
rect 4031 8214 4199 8216
rect 111 8134 148 8136
rect 111 8133 759 8134
rect 110 8127 759 8133
rect 110 8109 120 8127
rect 138 8113 759 8127
rect 138 8109 148 8113
rect 589 8112 759 8113
rect 110 8099 148 8109
rect 110 8021 145 8099
rect 722 8089 759 8112
rect 106 8012 145 8021
rect 106 7994 116 8012
rect 134 7994 145 8012
rect 106 7988 145 7994
rect 301 8064 551 8088
rect 301 7993 338 8064
rect 453 8003 484 8004
rect 106 7984 143 7988
rect 301 7973 310 7993
rect 330 7973 338 7993
rect 301 7963 338 7973
rect 397 7993 484 8003
rect 397 7973 406 7993
rect 426 7973 484 7993
rect 397 7964 484 7973
rect 397 7963 434 7964
rect 109 7913 146 7922
rect 107 7895 118 7913
rect 136 7895 146 7913
rect 453 7911 484 7964
rect 514 7993 551 8064
rect 722 8069 1115 8089
rect 1135 8069 1138 8089
rect 722 8064 1138 8069
rect 722 8063 1063 8064
rect 666 8003 697 8004
rect 514 7973 523 7993
rect 543 7973 551 7993
rect 514 7963 551 7973
rect 610 7996 697 8003
rect 610 7993 671 7996
rect 610 7973 619 7993
rect 639 7976 671 7993
rect 692 7976 697 7996
rect 639 7973 697 7976
rect 610 7966 697 7973
rect 722 7993 759 8063
rect 1025 8062 1062 8063
rect 4031 8036 4058 8214
rect 4098 8176 4162 8188
rect 4438 8184 4475 8216
rect 4646 8215 4895 8237
rect 4646 8184 4683 8215
rect 4859 8213 4895 8215
rect 5038 8218 5076 8251
rect 4859 8184 4896 8213
rect 4098 8175 4133 8176
rect 4075 8170 4133 8175
rect 4075 8150 4078 8170
rect 4098 8156 4133 8170
rect 4153 8156 4162 8176
rect 4098 8148 4162 8156
rect 4124 8147 4162 8148
rect 4125 8146 4162 8147
rect 4228 8180 4264 8181
rect 4336 8180 4372 8181
rect 4228 8174 4372 8180
rect 4228 8172 4294 8174
rect 4228 8152 4236 8172
rect 4256 8153 4294 8172
rect 4316 8172 4372 8174
rect 4316 8153 4344 8172
rect 4256 8152 4344 8153
rect 4364 8152 4372 8172
rect 4228 8146 4372 8152
rect 4438 8176 4476 8184
rect 4544 8180 4580 8181
rect 4438 8156 4447 8176
rect 4467 8156 4476 8176
rect 4438 8147 4476 8156
rect 4495 8173 4580 8180
rect 4495 8153 4502 8173
rect 4523 8172 4580 8173
rect 4523 8153 4552 8172
rect 4495 8152 4552 8153
rect 4572 8152 4580 8172
rect 4438 8146 4475 8147
rect 4495 8146 4580 8152
rect 4646 8176 4684 8184
rect 4757 8180 4793 8181
rect 4646 8156 4655 8176
rect 4675 8156 4684 8176
rect 4646 8147 4684 8156
rect 4708 8172 4793 8180
rect 4708 8152 4765 8172
rect 4785 8152 4793 8172
rect 4646 8146 4683 8147
rect 4708 8146 4793 8152
rect 4859 8176 4897 8184
rect 4859 8156 4868 8176
rect 4888 8156 4897 8176
rect 4859 8147 4897 8156
rect 5038 8183 5074 8218
rect 5391 8214 5426 8251
rect 9730 8238 10357 8256
rect 5389 8205 5426 8214
rect 5389 8187 5399 8205
rect 5417 8187 5426 8205
rect 5038 8173 5075 8183
rect 5389 8177 5426 8187
rect 9312 8221 9480 8222
rect 9731 8221 9755 8238
rect 9312 8195 9756 8221
rect 9312 8193 9480 8195
rect 5038 8155 5048 8173
rect 5066 8155 5075 8173
rect 4859 8146 4896 8147
rect 5038 8146 5075 8155
rect 4282 8125 4318 8146
rect 4708 8125 4739 8146
rect 4115 8121 4215 8125
rect 4115 8117 4177 8121
rect 4115 8091 4122 8117
rect 4148 8095 4177 8117
rect 4203 8095 4215 8121
rect 4148 8091 4215 8095
rect 4115 8088 4215 8091
rect 4283 8088 4318 8125
rect 4380 8122 4739 8125
rect 4380 8117 4602 8122
rect 4380 8093 4393 8117
rect 4417 8098 4602 8117
rect 4626 8098 4739 8122
rect 4417 8093 4739 8098
rect 4380 8089 4739 8093
rect 4806 8117 4955 8125
rect 4806 8097 4817 8117
rect 4837 8097 4955 8117
rect 5392 8113 5429 8115
rect 5392 8112 6040 8113
rect 4806 8090 4955 8097
rect 5391 8106 6040 8112
rect 4806 8089 4847 8090
rect 4130 8036 4167 8037
rect 4226 8036 4263 8037
rect 4282 8036 4318 8088
rect 4337 8036 4374 8037
rect 4030 8027 4168 8036
rect 2966 8009 2997 8012
rect 874 8003 910 8004
rect 722 7973 731 7993
rect 751 7973 759 7993
rect 610 7964 666 7966
rect 610 7963 647 7964
rect 722 7963 759 7973
rect 818 7993 966 8003
rect 1066 8000 1162 8002
rect 818 7973 827 7993
rect 847 7973 937 7993
rect 957 7973 966 7993
rect 818 7964 966 7973
rect 1024 7993 1162 8000
rect 1024 7973 1033 7993
rect 1053 7973 1162 7993
rect 1024 7964 1162 7973
rect 2966 7983 2973 8009
rect 2992 7983 2997 8009
rect 818 7963 855 7964
rect 874 7912 910 7964
rect 929 7963 966 7964
rect 1025 7963 1062 7964
rect 345 7910 386 7911
rect 107 7746 146 7895
rect 237 7903 386 7910
rect 237 7883 355 7903
rect 375 7883 386 7903
rect 237 7875 386 7883
rect 453 7907 812 7911
rect 453 7902 775 7907
rect 453 7878 566 7902
rect 590 7883 775 7902
rect 799 7883 812 7907
rect 590 7878 812 7883
rect 453 7875 812 7878
rect 874 7875 909 7912
rect 977 7909 1077 7912
rect 977 7905 1044 7909
rect 977 7879 989 7905
rect 1015 7883 1044 7905
rect 1070 7883 1077 7909
rect 1015 7879 1077 7883
rect 977 7875 1077 7879
rect 453 7854 484 7875
rect 874 7854 910 7875
rect 296 7853 333 7854
rect 295 7844 333 7853
rect 295 7824 304 7844
rect 324 7824 333 7844
rect 295 7816 333 7824
rect 399 7848 484 7854
rect 509 7853 546 7854
rect 399 7828 407 7848
rect 427 7828 484 7848
rect 399 7820 484 7828
rect 508 7844 546 7853
rect 508 7824 517 7844
rect 537 7824 546 7844
rect 399 7819 435 7820
rect 508 7816 546 7824
rect 612 7848 697 7854
rect 717 7853 754 7854
rect 612 7828 620 7848
rect 640 7847 697 7848
rect 640 7828 669 7847
rect 612 7827 669 7828
rect 690 7827 697 7847
rect 612 7820 697 7827
rect 716 7844 754 7853
rect 716 7824 725 7844
rect 745 7824 754 7844
rect 612 7819 648 7820
rect 716 7816 754 7824
rect 820 7849 964 7854
rect 820 7848 885 7849
rect 820 7828 828 7848
rect 848 7828 885 7848
rect 907 7848 964 7849
rect 907 7828 936 7848
rect 956 7828 964 7848
rect 820 7820 964 7828
rect 820 7819 856 7820
rect 928 7819 964 7820
rect 1030 7853 1067 7854
rect 1030 7852 1068 7853
rect 1030 7844 1094 7852
rect 1030 7824 1039 7844
rect 1059 7830 1094 7844
rect 1114 7830 1117 7850
rect 1059 7825 1117 7830
rect 1059 7824 1094 7825
rect 296 7787 333 7816
rect 297 7785 333 7787
rect 509 7785 546 7816
rect 297 7763 546 7785
rect 717 7784 754 7816
rect 1030 7812 1094 7824
rect 1134 7786 1161 7964
rect 993 7784 1161 7786
rect 717 7758 1161 7784
rect 1313 7883 1563 7907
rect 1313 7812 1350 7883
rect 1465 7822 1496 7823
rect 1313 7792 1322 7812
rect 1342 7792 1350 7812
rect 1313 7782 1350 7792
rect 1409 7812 1496 7822
rect 1409 7792 1418 7812
rect 1438 7792 1496 7812
rect 1409 7783 1496 7792
rect 1409 7782 1446 7783
rect 717 7748 739 7758
rect 993 7757 1161 7758
rect 677 7746 739 7748
rect 107 7739 739 7746
rect 106 7730 739 7739
rect 1465 7730 1496 7783
rect 1526 7812 1563 7883
rect 1734 7888 2127 7908
rect 2147 7888 2150 7908
rect 1734 7883 2150 7888
rect 1734 7882 2075 7883
rect 1678 7822 1709 7823
rect 1526 7792 1535 7812
rect 1555 7792 1563 7812
rect 1526 7782 1563 7792
rect 1622 7815 1709 7822
rect 1622 7812 1683 7815
rect 1622 7792 1631 7812
rect 1651 7795 1683 7812
rect 1704 7795 1709 7815
rect 1651 7792 1709 7795
rect 1622 7785 1709 7792
rect 1734 7812 1771 7882
rect 2037 7881 2074 7882
rect 1886 7822 1922 7823
rect 1734 7792 1743 7812
rect 1763 7792 1771 7812
rect 1622 7783 1678 7785
rect 1622 7782 1659 7783
rect 1734 7782 1771 7792
rect 1830 7812 1978 7822
rect 2078 7819 2174 7821
rect 1830 7792 1839 7812
rect 1859 7792 1949 7812
rect 1969 7792 1978 7812
rect 1830 7783 1978 7792
rect 2036 7812 2174 7819
rect 2036 7792 2045 7812
rect 2065 7792 2174 7812
rect 2036 7783 2174 7792
rect 1830 7782 1867 7783
rect 1886 7731 1922 7783
rect 1941 7782 1978 7783
rect 2037 7782 2074 7783
rect 106 7712 116 7730
rect 134 7729 739 7730
rect 1357 7729 1398 7730
rect 134 7724 155 7729
rect 134 7712 146 7724
rect 1249 7722 1398 7729
rect 106 7704 146 7712
rect 189 7711 215 7712
rect 106 7702 143 7704
rect 189 7693 743 7711
rect 1249 7702 1367 7722
rect 1387 7702 1398 7722
rect 1249 7694 1398 7702
rect 1465 7726 1824 7730
rect 1465 7721 1787 7726
rect 1465 7697 1578 7721
rect 1602 7702 1787 7721
rect 1811 7702 1824 7726
rect 1602 7697 1824 7702
rect 1465 7694 1824 7697
rect 1886 7694 1921 7731
rect 1989 7728 2089 7731
rect 1989 7724 2056 7728
rect 1989 7698 2001 7724
rect 2027 7702 2056 7724
rect 2082 7702 2089 7728
rect 2027 7698 2089 7702
rect 1989 7694 2089 7698
rect 109 7634 146 7640
rect 189 7634 215 7693
rect 722 7674 743 7693
rect 109 7631 215 7634
rect 109 7613 118 7631
rect 136 7617 215 7631
rect 300 7649 550 7673
rect 136 7615 212 7617
rect 136 7613 146 7615
rect 109 7603 146 7613
rect 114 7538 145 7603
rect 300 7578 337 7649
rect 452 7588 483 7589
rect 300 7558 309 7578
rect 329 7558 337 7578
rect 300 7548 337 7558
rect 396 7578 483 7588
rect 396 7558 405 7578
rect 425 7558 483 7578
rect 396 7549 483 7558
rect 396 7548 433 7549
rect 113 7529 150 7538
rect 113 7511 123 7529
rect 141 7511 150 7529
rect 113 7501 150 7511
rect 452 7496 483 7549
rect 513 7578 550 7649
rect 721 7654 1114 7674
rect 1134 7654 1137 7674
rect 1465 7673 1496 7694
rect 1886 7673 1922 7694
rect 1308 7672 1345 7673
rect 721 7649 1137 7654
rect 1307 7663 1345 7672
rect 721 7648 1062 7649
rect 665 7588 696 7589
rect 513 7558 522 7578
rect 542 7558 550 7578
rect 513 7548 550 7558
rect 609 7581 696 7588
rect 609 7578 670 7581
rect 609 7558 618 7578
rect 638 7561 670 7578
rect 691 7561 696 7581
rect 638 7558 696 7561
rect 609 7551 696 7558
rect 721 7578 758 7648
rect 1024 7647 1061 7648
rect 1307 7643 1316 7663
rect 1336 7643 1345 7663
rect 1307 7635 1345 7643
rect 1411 7667 1496 7673
rect 1521 7672 1558 7673
rect 1411 7647 1419 7667
rect 1439 7647 1496 7667
rect 1411 7639 1496 7647
rect 1520 7663 1558 7672
rect 1520 7643 1529 7663
rect 1549 7643 1558 7663
rect 1411 7638 1447 7639
rect 1520 7635 1558 7643
rect 1624 7667 1709 7673
rect 1729 7672 1766 7673
rect 1624 7647 1632 7667
rect 1652 7666 1709 7667
rect 1652 7647 1681 7666
rect 1624 7646 1681 7647
rect 1702 7646 1709 7666
rect 1624 7639 1709 7646
rect 1728 7663 1766 7672
rect 1728 7643 1737 7663
rect 1757 7643 1766 7663
rect 1624 7638 1660 7639
rect 1728 7635 1766 7643
rect 1832 7667 1976 7673
rect 1832 7647 1840 7667
rect 1860 7647 1892 7667
rect 1916 7647 1948 7667
rect 1968 7647 1976 7667
rect 1832 7639 1976 7647
rect 1832 7638 1868 7639
rect 1940 7638 1976 7639
rect 2042 7672 2079 7673
rect 2042 7671 2080 7672
rect 2042 7663 2106 7671
rect 2042 7643 2051 7663
rect 2071 7649 2106 7663
rect 2126 7649 2129 7669
rect 2071 7644 2129 7649
rect 2071 7643 2106 7644
rect 1308 7606 1345 7635
rect 1309 7604 1345 7606
rect 1521 7604 1558 7635
rect 873 7588 909 7589
rect 721 7558 730 7578
rect 750 7558 758 7578
rect 609 7549 665 7551
rect 609 7548 646 7549
rect 721 7548 758 7558
rect 817 7578 965 7588
rect 1065 7585 1161 7587
rect 817 7558 826 7578
rect 846 7558 936 7578
rect 956 7558 965 7578
rect 817 7549 965 7558
rect 1023 7578 1161 7585
rect 1309 7582 1558 7604
rect 1729 7603 1766 7635
rect 2042 7631 2106 7643
rect 2146 7605 2173 7783
rect 2005 7603 2173 7605
rect 1729 7599 2173 7603
rect 1023 7558 1032 7578
rect 1052 7558 1161 7578
rect 1729 7580 1778 7599
rect 1798 7580 2173 7599
rect 1729 7577 2173 7580
rect 2005 7576 2173 7577
rect 2873 7590 2902 7592
rect 2873 7585 2905 7590
rect 2873 7567 2880 7585
rect 2900 7567 2905 7585
rect 2966 7589 2997 7983
rect 3018 8008 3186 8009
rect 3018 8005 3462 8008
rect 3018 7986 3393 8005
rect 3413 7986 3462 8005
rect 4030 8007 4139 8027
rect 4159 8007 4168 8027
rect 3018 7982 3462 7986
rect 3018 7980 3186 7982
rect 3018 7802 3045 7980
rect 3085 7942 3149 7954
rect 3425 7950 3462 7982
rect 3633 7981 3882 8003
rect 4030 8000 4168 8007
rect 4226 8027 4374 8036
rect 4226 8007 4235 8027
rect 4255 8007 4345 8027
rect 4365 8007 4374 8027
rect 4030 7998 4126 8000
rect 4226 7997 4374 8007
rect 4433 8027 4470 8037
rect 4545 8036 4582 8037
rect 4526 8034 4582 8036
rect 4433 8007 4441 8027
rect 4461 8007 4470 8027
rect 4282 7996 4318 7997
rect 3633 7950 3670 7981
rect 3846 7979 3882 7981
rect 3846 7950 3883 7979
rect 3085 7941 3120 7942
rect 3062 7936 3120 7941
rect 3062 7916 3065 7936
rect 3085 7922 3120 7936
rect 3140 7922 3149 7942
rect 3085 7914 3149 7922
rect 3111 7913 3149 7914
rect 3112 7912 3149 7913
rect 3215 7946 3251 7947
rect 3323 7946 3359 7947
rect 3215 7938 3359 7946
rect 3215 7918 3223 7938
rect 3243 7937 3331 7938
rect 3243 7918 3276 7937
rect 3215 7917 3276 7918
rect 3300 7918 3331 7937
rect 3351 7918 3359 7938
rect 3300 7917 3359 7918
rect 3215 7912 3359 7917
rect 3425 7942 3463 7950
rect 3531 7946 3567 7947
rect 3425 7922 3434 7942
rect 3454 7922 3463 7942
rect 3425 7913 3463 7922
rect 3482 7939 3567 7946
rect 3482 7919 3489 7939
rect 3510 7938 3567 7939
rect 3510 7919 3539 7938
rect 3482 7918 3539 7919
rect 3559 7918 3567 7938
rect 3425 7912 3462 7913
rect 3482 7912 3567 7918
rect 3633 7942 3671 7950
rect 3744 7946 3780 7947
rect 3633 7922 3642 7942
rect 3662 7922 3671 7942
rect 3633 7913 3671 7922
rect 3695 7938 3780 7946
rect 3695 7918 3752 7938
rect 3772 7918 3780 7938
rect 3633 7912 3670 7913
rect 3695 7912 3780 7918
rect 3846 7942 3884 7950
rect 3846 7922 3855 7942
rect 3875 7922 3884 7942
rect 4130 7937 4167 7938
rect 4433 7937 4470 8007
rect 4495 8027 4582 8034
rect 4495 8024 4553 8027
rect 4495 8004 4500 8024
rect 4521 8007 4553 8024
rect 4573 8007 4582 8027
rect 4521 8004 4582 8007
rect 4495 7997 4582 8004
rect 4641 8027 4678 8037
rect 4641 8007 4649 8027
rect 4669 8007 4678 8027
rect 4495 7996 4526 7997
rect 4129 7936 4470 7937
rect 3846 7913 3884 7922
rect 4054 7931 4470 7936
rect 3846 7912 3883 7913
rect 3269 7891 3305 7912
rect 3695 7891 3726 7912
rect 4054 7911 4057 7931
rect 4077 7911 4470 7931
rect 4641 7936 4678 8007
rect 4708 8036 4739 8089
rect 5391 8088 5401 8106
rect 5419 8092 6040 8106
rect 5419 8088 5429 8092
rect 5870 8091 6040 8092
rect 5041 8074 5078 8084
rect 5041 8056 5050 8074
rect 5068 8056 5078 8074
rect 5041 8047 5078 8056
rect 5391 8078 5429 8088
rect 4758 8036 4795 8037
rect 4708 8027 4795 8036
rect 4708 8007 4766 8027
rect 4786 8007 4795 8027
rect 4708 7997 4795 8007
rect 4854 8027 4891 8037
rect 4854 8007 4862 8027
rect 4882 8007 4891 8027
rect 4708 7996 4739 7997
rect 4854 7936 4891 8007
rect 5046 7982 5077 8047
rect 5391 8000 5426 8078
rect 6003 8068 6040 8091
rect 5387 7991 5426 8000
rect 5045 7972 5082 7982
rect 5045 7970 5055 7972
rect 4979 7968 5055 7970
rect 4641 7912 4891 7936
rect 4976 7954 5055 7968
rect 5073 7954 5082 7972
rect 5387 7973 5397 7991
rect 5415 7973 5426 7991
rect 5387 7967 5426 7973
rect 5582 8043 5832 8067
rect 5582 7972 5619 8043
rect 5734 7982 5765 7983
rect 5387 7963 5424 7967
rect 4976 7951 5082 7954
rect 4448 7892 4469 7911
rect 4976 7892 5002 7951
rect 5045 7945 5082 7951
rect 5582 7952 5591 7972
rect 5611 7952 5619 7972
rect 5582 7942 5619 7952
rect 5678 7972 5765 7982
rect 5678 7952 5687 7972
rect 5707 7952 5765 7972
rect 5678 7943 5765 7952
rect 5678 7942 5715 7943
rect 5390 7892 5427 7901
rect 3102 7887 3202 7891
rect 3102 7883 3164 7887
rect 3102 7857 3109 7883
rect 3135 7861 3164 7883
rect 3190 7861 3202 7887
rect 3135 7857 3202 7861
rect 3102 7854 3202 7857
rect 3270 7854 3305 7891
rect 3367 7888 3726 7891
rect 3367 7883 3589 7888
rect 3367 7859 3380 7883
rect 3404 7864 3589 7883
rect 3613 7864 3726 7888
rect 3404 7859 3726 7864
rect 3367 7855 3726 7859
rect 3793 7883 3942 7891
rect 3793 7863 3804 7883
rect 3824 7863 3942 7883
rect 4448 7874 5002 7892
rect 5048 7881 5085 7883
rect 4976 7873 5002 7874
rect 5045 7873 5085 7881
rect 3793 7856 3942 7863
rect 5045 7861 5057 7873
rect 5036 7856 5057 7861
rect 3793 7855 3834 7856
rect 4452 7855 5057 7856
rect 5075 7855 5085 7873
rect 3117 7802 3154 7803
rect 3213 7802 3250 7803
rect 3269 7802 3305 7854
rect 3324 7802 3361 7803
rect 3017 7793 3155 7802
rect 3017 7773 3126 7793
rect 3146 7773 3155 7793
rect 3017 7766 3155 7773
rect 3213 7793 3361 7802
rect 3213 7773 3222 7793
rect 3242 7773 3332 7793
rect 3352 7773 3361 7793
rect 3017 7764 3113 7766
rect 3213 7763 3361 7773
rect 3420 7793 3457 7803
rect 3532 7802 3569 7803
rect 3513 7800 3569 7802
rect 3420 7773 3428 7793
rect 3448 7773 3457 7793
rect 3269 7762 3305 7763
rect 3117 7703 3154 7704
rect 3420 7703 3457 7773
rect 3482 7793 3569 7800
rect 3482 7790 3540 7793
rect 3482 7770 3487 7790
rect 3508 7773 3540 7790
rect 3560 7773 3569 7793
rect 3508 7770 3569 7773
rect 3482 7763 3569 7770
rect 3628 7793 3665 7803
rect 3628 7773 3636 7793
rect 3656 7773 3665 7793
rect 3482 7762 3513 7763
rect 3116 7702 3457 7703
rect 3041 7697 3457 7702
rect 3041 7677 3044 7697
rect 3064 7677 3457 7697
rect 3628 7702 3665 7773
rect 3695 7802 3726 7855
rect 4452 7846 5085 7855
rect 5388 7874 5399 7892
rect 5417 7874 5427 7892
rect 5734 7890 5765 7943
rect 5795 7972 5832 8043
rect 6003 8048 6396 8068
rect 6416 8048 6419 8068
rect 6003 8043 6419 8048
rect 6003 8042 6344 8043
rect 5947 7982 5978 7983
rect 5795 7952 5804 7972
rect 5824 7952 5832 7972
rect 5795 7942 5832 7952
rect 5891 7975 5978 7982
rect 5891 7972 5952 7975
rect 5891 7952 5900 7972
rect 5920 7955 5952 7972
rect 5973 7955 5978 7975
rect 5920 7952 5978 7955
rect 5891 7945 5978 7952
rect 6003 7972 6040 8042
rect 6306 8041 6343 8042
rect 9312 8015 9339 8193
rect 9379 8155 9443 8167
rect 9719 8163 9756 8195
rect 9927 8194 10176 8216
rect 9927 8163 9964 8194
rect 10140 8192 10176 8194
rect 10319 8197 10357 8238
rect 10140 8163 10177 8192
rect 9379 8154 9414 8155
rect 9356 8149 9414 8154
rect 9356 8129 9359 8149
rect 9379 8135 9414 8149
rect 9434 8135 9443 8155
rect 9379 8127 9443 8135
rect 9405 8126 9443 8127
rect 9406 8125 9443 8126
rect 9509 8159 9545 8160
rect 9617 8159 9653 8160
rect 9509 8153 9653 8159
rect 9509 8151 9575 8153
rect 9509 8131 9517 8151
rect 9537 8132 9575 8151
rect 9597 8151 9653 8153
rect 9597 8132 9625 8151
rect 9537 8131 9625 8132
rect 9645 8131 9653 8151
rect 9509 8125 9653 8131
rect 9719 8155 9757 8163
rect 9825 8159 9861 8160
rect 9719 8135 9728 8155
rect 9748 8135 9757 8155
rect 9719 8126 9757 8135
rect 9776 8152 9861 8159
rect 9776 8132 9783 8152
rect 9804 8151 9861 8152
rect 9804 8132 9833 8151
rect 9776 8131 9833 8132
rect 9853 8131 9861 8151
rect 9719 8125 9756 8126
rect 9776 8125 9861 8131
rect 9927 8155 9965 8163
rect 10038 8159 10074 8160
rect 9927 8135 9936 8155
rect 9956 8135 9965 8155
rect 9927 8126 9965 8135
rect 9989 8151 10074 8159
rect 9989 8131 10046 8151
rect 10066 8131 10074 8151
rect 9927 8125 9964 8126
rect 9989 8125 10074 8131
rect 10140 8155 10178 8163
rect 10140 8135 10149 8155
rect 10169 8135 10178 8155
rect 10140 8126 10178 8135
rect 10319 8162 10355 8197
rect 10319 8152 10356 8162
rect 10319 8134 10329 8152
rect 10347 8134 10356 8152
rect 10140 8125 10177 8126
rect 10319 8125 10356 8134
rect 9563 8104 9599 8125
rect 9989 8104 10020 8125
rect 9396 8100 9496 8104
rect 9396 8096 9458 8100
rect 9396 8070 9403 8096
rect 9429 8074 9458 8096
rect 9484 8074 9496 8100
rect 9429 8070 9496 8074
rect 9396 8067 9496 8070
rect 9564 8067 9599 8104
rect 9661 8101 10020 8104
rect 9661 8096 9883 8101
rect 9661 8072 9674 8096
rect 9698 8077 9883 8096
rect 9907 8077 10020 8101
rect 9698 8072 10020 8077
rect 9661 8068 10020 8072
rect 10087 8096 10236 8104
rect 10087 8076 10098 8096
rect 10118 8076 10236 8096
rect 10087 8069 10236 8076
rect 10087 8068 10128 8069
rect 9411 8015 9448 8016
rect 9507 8015 9544 8016
rect 9563 8015 9599 8067
rect 9618 8015 9655 8016
rect 9311 8006 9449 8015
rect 8247 7988 8278 7991
rect 6155 7982 6191 7983
rect 6003 7952 6012 7972
rect 6032 7952 6040 7972
rect 5891 7943 5947 7945
rect 5891 7942 5928 7943
rect 6003 7942 6040 7952
rect 6099 7972 6247 7982
rect 6347 7979 6443 7981
rect 6099 7952 6108 7972
rect 6128 7952 6218 7972
rect 6238 7952 6247 7972
rect 6099 7943 6247 7952
rect 6305 7972 6443 7979
rect 6305 7952 6314 7972
rect 6334 7952 6443 7972
rect 6305 7943 6443 7952
rect 8247 7962 8254 7988
rect 8273 7962 8278 7988
rect 6099 7942 6136 7943
rect 6155 7891 6191 7943
rect 6210 7942 6247 7943
rect 6306 7942 6343 7943
rect 5626 7889 5667 7890
rect 4452 7839 5084 7846
rect 4452 7837 4514 7839
rect 4030 7827 4198 7828
rect 4452 7827 4474 7837
rect 3745 7802 3782 7803
rect 3695 7793 3782 7802
rect 3695 7773 3753 7793
rect 3773 7773 3782 7793
rect 3695 7763 3782 7773
rect 3841 7793 3878 7803
rect 3841 7773 3849 7793
rect 3869 7773 3878 7793
rect 3695 7762 3726 7763
rect 3841 7702 3878 7773
rect 3628 7678 3878 7702
rect 4030 7801 4474 7827
rect 4030 7799 4198 7801
rect 4030 7621 4057 7799
rect 4097 7761 4161 7773
rect 4437 7769 4474 7801
rect 4645 7800 4894 7822
rect 4645 7769 4682 7800
rect 4858 7798 4894 7800
rect 4858 7769 4895 7798
rect 4097 7760 4132 7761
rect 4074 7755 4132 7760
rect 4074 7735 4077 7755
rect 4097 7741 4132 7755
rect 4152 7741 4161 7761
rect 4097 7733 4161 7741
rect 4123 7732 4161 7733
rect 4124 7731 4161 7732
rect 4227 7765 4263 7766
rect 4335 7765 4371 7766
rect 4227 7757 4371 7765
rect 4227 7737 4235 7757
rect 4255 7737 4284 7757
rect 4227 7736 4284 7737
rect 4306 7737 4343 7757
rect 4363 7737 4371 7757
rect 4306 7736 4371 7737
rect 4227 7731 4371 7736
rect 4437 7761 4475 7769
rect 4543 7765 4579 7766
rect 4437 7741 4446 7761
rect 4466 7741 4475 7761
rect 4437 7732 4475 7741
rect 4494 7758 4579 7765
rect 4494 7738 4501 7758
rect 4522 7757 4579 7758
rect 4522 7738 4551 7757
rect 4494 7737 4551 7738
rect 4571 7737 4579 7757
rect 4437 7731 4474 7732
rect 4494 7731 4579 7737
rect 4645 7761 4683 7769
rect 4756 7765 4792 7766
rect 4645 7741 4654 7761
rect 4674 7741 4683 7761
rect 4645 7732 4683 7741
rect 4707 7757 4792 7765
rect 4707 7737 4764 7757
rect 4784 7737 4792 7757
rect 4645 7731 4682 7732
rect 4707 7731 4792 7737
rect 4858 7761 4896 7769
rect 4858 7741 4867 7761
rect 4887 7741 4896 7761
rect 4858 7732 4896 7741
rect 4858 7731 4895 7732
rect 4281 7710 4317 7731
rect 4707 7710 4738 7731
rect 4114 7706 4214 7710
rect 4114 7702 4176 7706
rect 4114 7676 4121 7702
rect 4147 7680 4176 7702
rect 4202 7680 4214 7706
rect 4147 7676 4214 7680
rect 4114 7673 4214 7676
rect 4282 7673 4317 7710
rect 4379 7707 4738 7710
rect 4379 7702 4601 7707
rect 4379 7678 4392 7702
rect 4416 7683 4601 7702
rect 4625 7683 4738 7707
rect 4416 7678 4738 7683
rect 4379 7674 4738 7678
rect 4805 7702 4954 7710
rect 4805 7682 4816 7702
rect 4836 7682 4954 7702
rect 4805 7675 4954 7682
rect 5045 7690 5084 7839
rect 5388 7725 5427 7874
rect 5518 7882 5667 7889
rect 5518 7862 5636 7882
rect 5656 7862 5667 7882
rect 5518 7854 5667 7862
rect 5734 7886 6093 7890
rect 5734 7881 6056 7886
rect 5734 7857 5847 7881
rect 5871 7862 6056 7881
rect 6080 7862 6093 7886
rect 5871 7857 6093 7862
rect 5734 7854 6093 7857
rect 6155 7854 6190 7891
rect 6258 7888 6358 7891
rect 6258 7884 6325 7888
rect 6258 7858 6270 7884
rect 6296 7862 6325 7884
rect 6351 7862 6358 7888
rect 6296 7858 6358 7862
rect 6258 7854 6358 7858
rect 5734 7833 5765 7854
rect 6155 7833 6191 7854
rect 5577 7832 5614 7833
rect 5576 7823 5614 7832
rect 5576 7803 5585 7823
rect 5605 7803 5614 7823
rect 5576 7795 5614 7803
rect 5680 7827 5765 7833
rect 5790 7832 5827 7833
rect 5680 7807 5688 7827
rect 5708 7807 5765 7827
rect 5680 7799 5765 7807
rect 5789 7823 5827 7832
rect 5789 7803 5798 7823
rect 5818 7803 5827 7823
rect 5680 7798 5716 7799
rect 5789 7795 5827 7803
rect 5893 7827 5978 7833
rect 5998 7832 6035 7833
rect 5893 7807 5901 7827
rect 5921 7826 5978 7827
rect 5921 7807 5950 7826
rect 5893 7806 5950 7807
rect 5971 7806 5978 7826
rect 5893 7799 5978 7806
rect 5997 7823 6035 7832
rect 5997 7803 6006 7823
rect 6026 7803 6035 7823
rect 5893 7798 5929 7799
rect 5997 7795 6035 7803
rect 6101 7828 6245 7833
rect 6101 7827 6166 7828
rect 6101 7807 6109 7827
rect 6129 7807 6166 7827
rect 6188 7827 6245 7828
rect 6188 7807 6217 7827
rect 6237 7807 6245 7827
rect 6101 7799 6245 7807
rect 6101 7798 6137 7799
rect 6209 7798 6245 7799
rect 6311 7832 6348 7833
rect 6311 7831 6349 7832
rect 6311 7823 6375 7831
rect 6311 7803 6320 7823
rect 6340 7809 6375 7823
rect 6395 7809 6398 7829
rect 6340 7804 6398 7809
rect 6340 7803 6375 7804
rect 5577 7766 5614 7795
rect 5578 7764 5614 7766
rect 5790 7764 5827 7795
rect 5578 7742 5827 7764
rect 5998 7763 6035 7795
rect 6311 7791 6375 7803
rect 6415 7765 6442 7943
rect 6274 7763 6442 7765
rect 5998 7737 6442 7763
rect 6594 7862 6844 7886
rect 6594 7791 6631 7862
rect 6746 7801 6777 7802
rect 6594 7771 6603 7791
rect 6623 7771 6631 7791
rect 6594 7761 6631 7771
rect 6690 7791 6777 7801
rect 6690 7771 6699 7791
rect 6719 7771 6777 7791
rect 6690 7762 6777 7771
rect 6690 7761 6727 7762
rect 5998 7727 6020 7737
rect 6274 7736 6442 7737
rect 5958 7725 6020 7727
rect 5388 7718 6020 7725
rect 4805 7674 4846 7675
rect 4129 7621 4166 7622
rect 4225 7621 4262 7622
rect 4281 7621 4317 7673
rect 4336 7621 4373 7622
rect 4029 7612 4167 7621
rect 4029 7592 4138 7612
rect 4158 7592 4167 7612
rect 2966 7588 3136 7589
rect 2966 7573 3412 7588
rect 4029 7585 4167 7592
rect 4225 7612 4373 7621
rect 4225 7592 4234 7612
rect 4254 7592 4344 7612
rect 4364 7592 4373 7612
rect 4029 7583 4125 7585
rect 2873 7562 2905 7567
rect 1023 7549 1161 7558
rect 817 7548 854 7549
rect 873 7497 909 7549
rect 928 7548 965 7549
rect 1024 7548 1061 7549
rect 344 7495 385 7496
rect 236 7488 385 7495
rect 236 7468 354 7488
rect 374 7468 385 7488
rect 236 7460 385 7468
rect 452 7492 811 7496
rect 452 7487 774 7492
rect 452 7463 565 7487
rect 589 7468 774 7487
rect 798 7468 811 7492
rect 589 7463 811 7468
rect 452 7460 811 7463
rect 873 7460 908 7497
rect 976 7494 1076 7497
rect 976 7490 1043 7494
rect 976 7464 988 7490
rect 1014 7468 1043 7490
rect 1069 7468 1076 7494
rect 1014 7464 1076 7468
rect 976 7460 1076 7464
rect 452 7439 483 7460
rect 873 7439 909 7460
rect 116 7430 153 7439
rect 295 7438 332 7439
rect 116 7412 125 7430
rect 143 7412 153 7430
rect 116 7402 153 7412
rect 117 7367 153 7402
rect 294 7429 332 7438
rect 294 7409 303 7429
rect 323 7409 332 7429
rect 294 7401 332 7409
rect 398 7433 483 7439
rect 508 7438 545 7439
rect 398 7413 406 7433
rect 426 7413 483 7433
rect 398 7405 483 7413
rect 507 7429 545 7438
rect 507 7409 516 7429
rect 536 7409 545 7429
rect 398 7404 434 7405
rect 507 7401 545 7409
rect 611 7433 696 7439
rect 716 7438 753 7439
rect 611 7413 619 7433
rect 639 7432 696 7433
rect 639 7413 668 7432
rect 611 7412 668 7413
rect 689 7412 696 7432
rect 611 7405 696 7412
rect 715 7429 753 7438
rect 715 7409 724 7429
rect 744 7409 753 7429
rect 611 7404 647 7405
rect 715 7401 753 7409
rect 819 7433 963 7439
rect 819 7413 827 7433
rect 847 7432 935 7433
rect 847 7413 875 7432
rect 819 7411 875 7413
rect 897 7413 935 7432
rect 955 7413 963 7433
rect 897 7411 963 7413
rect 819 7405 963 7411
rect 819 7404 855 7405
rect 927 7404 963 7405
rect 1029 7438 1066 7439
rect 1029 7437 1067 7438
rect 1029 7429 1093 7437
rect 1029 7409 1038 7429
rect 1058 7415 1093 7429
rect 1113 7415 1116 7435
rect 1058 7410 1116 7415
rect 1058 7409 1093 7410
rect 295 7372 332 7401
rect 115 7326 153 7367
rect 296 7370 332 7372
rect 508 7370 545 7401
rect 296 7348 545 7370
rect 716 7369 753 7401
rect 1029 7397 1093 7409
rect 1133 7371 1160 7549
rect 992 7369 1160 7371
rect 716 7343 1160 7369
rect 717 7326 741 7343
rect 992 7342 1160 7343
rect 115 7308 742 7326
rect 1368 7322 1618 7346
rect 115 7302 153 7308
rect 115 7278 152 7302
rect 115 7254 150 7278
rect 113 7245 150 7254
rect 113 7227 123 7245
rect 141 7227 150 7245
rect 113 7217 150 7227
rect 1368 7251 1405 7322
rect 1520 7261 1551 7262
rect 1368 7231 1377 7251
rect 1397 7231 1405 7251
rect 1368 7221 1405 7231
rect 1464 7251 1551 7261
rect 1464 7231 1473 7251
rect 1493 7231 1551 7251
rect 1464 7222 1551 7231
rect 1464 7221 1501 7222
rect 1520 7169 1551 7222
rect 1581 7251 1618 7322
rect 1789 7327 2182 7347
rect 2202 7327 2205 7347
rect 1789 7322 2205 7327
rect 1789 7321 2130 7322
rect 1733 7261 1764 7262
rect 1581 7231 1590 7251
rect 1610 7231 1618 7251
rect 1581 7221 1618 7231
rect 1677 7254 1764 7261
rect 1677 7251 1738 7254
rect 1677 7231 1686 7251
rect 1706 7234 1738 7251
rect 1759 7234 1764 7254
rect 1706 7231 1764 7234
rect 1677 7224 1764 7231
rect 1789 7251 1826 7321
rect 2092 7320 2129 7321
rect 1941 7261 1977 7262
rect 1789 7231 1798 7251
rect 1818 7231 1826 7251
rect 1677 7222 1733 7224
rect 1677 7221 1714 7222
rect 1789 7221 1826 7231
rect 1885 7251 2033 7261
rect 2133 7258 2229 7260
rect 1885 7231 1894 7251
rect 1914 7231 2004 7251
rect 2024 7231 2033 7251
rect 1885 7222 2033 7231
rect 2091 7251 2229 7258
rect 2091 7231 2100 7251
rect 2120 7231 2229 7251
rect 2091 7222 2229 7231
rect 1885 7221 1922 7222
rect 1941 7170 1977 7222
rect 1996 7221 2033 7222
rect 2092 7221 2129 7222
rect 1412 7168 1453 7169
rect 1304 7161 1453 7168
rect 116 7153 153 7155
rect 116 7152 764 7153
rect 115 7146 764 7152
rect 115 7128 125 7146
rect 143 7132 764 7146
rect 1304 7141 1422 7161
rect 1442 7141 1453 7161
rect 1304 7133 1453 7141
rect 1520 7165 1879 7169
rect 1520 7160 1842 7165
rect 1520 7136 1633 7160
rect 1657 7141 1842 7160
rect 1866 7141 1879 7165
rect 1657 7136 1879 7141
rect 1520 7133 1879 7136
rect 1941 7133 1976 7170
rect 2044 7167 2144 7170
rect 2044 7163 2111 7167
rect 2044 7137 2056 7163
rect 2082 7141 2111 7163
rect 2137 7141 2144 7167
rect 2082 7137 2144 7141
rect 2044 7133 2144 7137
rect 143 7128 153 7132
rect 594 7131 764 7132
rect 115 7118 153 7128
rect 115 7040 150 7118
rect 727 7108 764 7131
rect 1520 7112 1551 7133
rect 1941 7112 1977 7133
rect 1363 7111 1400 7112
rect 111 7031 150 7040
rect 111 7013 121 7031
rect 139 7013 150 7031
rect 111 7007 150 7013
rect 306 7083 556 7107
rect 306 7012 343 7083
rect 458 7022 489 7023
rect 111 7003 148 7007
rect 306 6992 315 7012
rect 335 6992 343 7012
rect 306 6982 343 6992
rect 402 7012 489 7022
rect 402 6992 411 7012
rect 431 6992 489 7012
rect 402 6983 489 6992
rect 402 6982 439 6983
rect 114 6932 151 6941
rect 112 6914 123 6932
rect 141 6914 151 6932
rect 458 6930 489 6983
rect 519 7012 556 7083
rect 727 7088 1120 7108
rect 1140 7088 1143 7108
rect 727 7083 1143 7088
rect 1362 7102 1400 7111
rect 727 7082 1068 7083
rect 1362 7082 1371 7102
rect 1391 7082 1400 7102
rect 671 7022 702 7023
rect 519 6992 528 7012
rect 548 6992 556 7012
rect 519 6982 556 6992
rect 615 7015 702 7022
rect 615 7012 676 7015
rect 615 6992 624 7012
rect 644 6995 676 7012
rect 697 6995 702 7015
rect 644 6992 702 6995
rect 615 6985 702 6992
rect 727 7012 764 7082
rect 1030 7081 1067 7082
rect 1362 7074 1400 7082
rect 1466 7106 1551 7112
rect 1576 7111 1613 7112
rect 1466 7086 1474 7106
rect 1494 7086 1551 7106
rect 1466 7078 1551 7086
rect 1575 7102 1613 7111
rect 1575 7082 1584 7102
rect 1604 7082 1613 7102
rect 1466 7077 1502 7078
rect 1575 7074 1613 7082
rect 1679 7106 1764 7112
rect 1784 7111 1821 7112
rect 1679 7086 1687 7106
rect 1707 7105 1764 7106
rect 1707 7086 1736 7105
rect 1679 7085 1736 7086
rect 1757 7085 1764 7105
rect 1679 7078 1764 7085
rect 1783 7102 1821 7111
rect 1783 7082 1792 7102
rect 1812 7082 1821 7102
rect 1679 7077 1715 7078
rect 1783 7074 1821 7082
rect 1887 7106 2031 7112
rect 1887 7086 1895 7106
rect 1915 7104 2003 7106
rect 1915 7087 1951 7104
rect 1975 7087 2003 7104
rect 1915 7086 2003 7087
rect 2023 7086 2031 7106
rect 1887 7078 2031 7086
rect 1887 7077 1923 7078
rect 1995 7077 2031 7078
rect 2097 7111 2134 7112
rect 2097 7110 2135 7111
rect 2097 7102 2161 7110
rect 2097 7082 2106 7102
rect 2126 7088 2161 7102
rect 2181 7088 2184 7108
rect 2126 7083 2184 7088
rect 2126 7082 2161 7083
rect 1363 7045 1400 7074
rect 1364 7043 1400 7045
rect 1576 7043 1613 7074
rect 879 7022 915 7023
rect 727 6992 736 7012
rect 756 6992 764 7012
rect 615 6983 671 6985
rect 615 6982 652 6983
rect 727 6982 764 6992
rect 823 7012 971 7022
rect 1364 7021 1613 7043
rect 1784 7042 1821 7074
rect 2097 7070 2161 7082
rect 2201 7044 2228 7222
rect 2060 7042 2228 7044
rect 1784 7031 2228 7042
rect 1071 7019 1167 7021
rect 823 6992 832 7012
rect 852 6992 942 7012
rect 962 6992 971 7012
rect 823 6983 971 6992
rect 1029 7012 1167 7019
rect 1784 7016 2230 7031
rect 2060 7015 2230 7016
rect 1029 6992 1038 7012
rect 1058 6992 1167 7012
rect 1029 6983 1167 6992
rect 823 6982 860 6983
rect 879 6931 915 6983
rect 934 6982 971 6983
rect 1030 6982 1067 6983
rect 350 6929 391 6930
rect 112 6765 151 6914
rect 242 6922 391 6929
rect 242 6902 360 6922
rect 380 6902 391 6922
rect 242 6894 391 6902
rect 458 6926 817 6930
rect 458 6921 780 6926
rect 458 6897 571 6921
rect 595 6902 780 6921
rect 804 6902 817 6926
rect 595 6897 817 6902
rect 458 6894 817 6897
rect 879 6894 914 6931
rect 982 6928 1082 6931
rect 982 6924 1049 6928
rect 982 6898 994 6924
rect 1020 6902 1049 6924
rect 1075 6902 1082 6928
rect 1020 6898 1082 6902
rect 982 6894 1082 6898
rect 458 6873 489 6894
rect 879 6873 915 6894
rect 301 6872 338 6873
rect 300 6863 338 6872
rect 300 6843 309 6863
rect 329 6843 338 6863
rect 300 6835 338 6843
rect 404 6867 489 6873
rect 514 6872 551 6873
rect 404 6847 412 6867
rect 432 6847 489 6867
rect 404 6839 489 6847
rect 513 6863 551 6872
rect 513 6843 522 6863
rect 542 6843 551 6863
rect 404 6838 440 6839
rect 513 6835 551 6843
rect 617 6867 702 6873
rect 722 6872 759 6873
rect 617 6847 625 6867
rect 645 6866 702 6867
rect 645 6847 674 6866
rect 617 6846 674 6847
rect 695 6846 702 6866
rect 617 6839 702 6846
rect 721 6863 759 6872
rect 721 6843 730 6863
rect 750 6843 759 6863
rect 617 6838 653 6839
rect 721 6835 759 6843
rect 825 6868 969 6873
rect 825 6867 890 6868
rect 825 6847 833 6867
rect 853 6847 890 6867
rect 912 6867 969 6868
rect 912 6847 941 6867
rect 961 6847 969 6867
rect 825 6839 969 6847
rect 825 6838 861 6839
rect 933 6838 969 6839
rect 1035 6872 1072 6873
rect 1035 6871 1073 6872
rect 1035 6863 1099 6871
rect 1035 6843 1044 6863
rect 1064 6849 1099 6863
rect 1119 6849 1122 6869
rect 1064 6844 1122 6849
rect 1064 6843 1099 6844
rect 301 6806 338 6835
rect 302 6804 338 6806
rect 514 6804 551 6835
rect 302 6782 551 6804
rect 722 6803 759 6835
rect 1035 6831 1099 6843
rect 1139 6805 1166 6983
rect 998 6803 1166 6805
rect 722 6777 1166 6803
rect 1318 6902 1568 6926
rect 1318 6831 1355 6902
rect 1470 6841 1501 6842
rect 1318 6811 1327 6831
rect 1347 6811 1355 6831
rect 1318 6801 1355 6811
rect 1414 6831 1501 6841
rect 1414 6811 1423 6831
rect 1443 6811 1501 6831
rect 1414 6802 1501 6811
rect 1414 6801 1451 6802
rect 722 6767 744 6777
rect 998 6776 1166 6777
rect 682 6765 744 6767
rect 112 6758 744 6765
rect 111 6749 744 6758
rect 1470 6749 1501 6802
rect 1531 6831 1568 6902
rect 1739 6907 2132 6927
rect 2152 6907 2155 6927
rect 1739 6902 2155 6907
rect 1739 6901 2080 6902
rect 1683 6841 1714 6842
rect 1531 6811 1540 6831
rect 1560 6811 1568 6831
rect 1531 6801 1568 6811
rect 1627 6834 1714 6841
rect 1627 6831 1688 6834
rect 1627 6811 1636 6831
rect 1656 6814 1688 6831
rect 1709 6814 1714 6834
rect 1656 6811 1714 6814
rect 1627 6804 1714 6811
rect 1739 6831 1776 6901
rect 2042 6900 2079 6901
rect 1891 6841 1927 6842
rect 1739 6811 1748 6831
rect 1768 6811 1776 6831
rect 1627 6802 1683 6804
rect 1627 6801 1664 6802
rect 1739 6801 1776 6811
rect 1835 6831 1983 6841
rect 2083 6838 2179 6840
rect 1835 6811 1844 6831
rect 1864 6811 1954 6831
rect 1974 6811 1983 6831
rect 1835 6802 1983 6811
rect 2041 6831 2179 6838
rect 2041 6811 2050 6831
rect 2070 6811 2179 6831
rect 2041 6802 2179 6811
rect 1835 6801 1872 6802
rect 1891 6750 1927 6802
rect 1946 6801 1983 6802
rect 2042 6801 2079 6802
rect 111 6731 121 6749
rect 139 6748 744 6749
rect 1362 6748 1403 6749
rect 139 6743 160 6748
rect 139 6731 151 6743
rect 1254 6741 1403 6748
rect 111 6723 151 6731
rect 194 6730 220 6731
rect 111 6721 148 6723
rect 194 6712 748 6730
rect 1254 6721 1372 6741
rect 1392 6721 1403 6741
rect 1254 6713 1403 6721
rect 1470 6745 1829 6749
rect 1470 6740 1792 6745
rect 1470 6716 1583 6740
rect 1607 6721 1792 6740
rect 1816 6721 1829 6745
rect 1607 6716 1829 6721
rect 1470 6713 1829 6716
rect 1891 6713 1926 6750
rect 1994 6747 2094 6750
rect 1994 6743 2061 6747
rect 1994 6717 2006 6743
rect 2032 6721 2061 6743
rect 2087 6721 2094 6747
rect 2032 6717 2094 6721
rect 1994 6713 2094 6717
rect 114 6653 151 6659
rect 194 6653 220 6712
rect 727 6693 748 6712
rect 114 6650 220 6653
rect 114 6632 123 6650
rect 141 6636 220 6650
rect 305 6668 555 6692
rect 141 6634 217 6636
rect 141 6632 151 6634
rect 114 6622 151 6632
rect 119 6557 150 6622
rect 305 6597 342 6668
rect 457 6607 488 6608
rect 305 6577 314 6597
rect 334 6577 342 6597
rect 305 6567 342 6577
rect 401 6597 488 6607
rect 401 6577 410 6597
rect 430 6577 488 6597
rect 401 6568 488 6577
rect 401 6567 438 6568
rect 118 6548 155 6557
rect 118 6530 128 6548
rect 146 6530 155 6548
rect 118 6520 155 6530
rect 457 6515 488 6568
rect 518 6597 555 6668
rect 726 6673 1119 6693
rect 1139 6673 1142 6693
rect 1470 6692 1501 6713
rect 1891 6692 1927 6713
rect 1313 6691 1350 6692
rect 726 6668 1142 6673
rect 1312 6682 1350 6691
rect 726 6667 1067 6668
rect 670 6607 701 6608
rect 518 6577 527 6597
rect 547 6577 555 6597
rect 518 6567 555 6577
rect 614 6600 701 6607
rect 614 6597 675 6600
rect 614 6577 623 6597
rect 643 6580 675 6597
rect 696 6580 701 6600
rect 643 6577 701 6580
rect 614 6570 701 6577
rect 726 6597 763 6667
rect 1029 6666 1066 6667
rect 1312 6662 1321 6682
rect 1341 6662 1350 6682
rect 1312 6654 1350 6662
rect 1416 6686 1501 6692
rect 1526 6691 1563 6692
rect 1416 6666 1424 6686
rect 1444 6666 1501 6686
rect 1416 6658 1501 6666
rect 1525 6682 1563 6691
rect 1525 6662 1534 6682
rect 1554 6662 1563 6682
rect 1416 6657 1452 6658
rect 1525 6654 1563 6662
rect 1629 6686 1714 6692
rect 1734 6691 1771 6692
rect 1629 6666 1637 6686
rect 1657 6685 1714 6686
rect 1657 6666 1686 6685
rect 1629 6665 1686 6666
rect 1707 6665 1714 6685
rect 1629 6658 1714 6665
rect 1733 6682 1771 6691
rect 1733 6662 1742 6682
rect 1762 6662 1771 6682
rect 1629 6657 1665 6658
rect 1733 6654 1771 6662
rect 1837 6687 1981 6692
rect 1837 6686 1896 6687
rect 1837 6666 1845 6686
rect 1865 6667 1896 6686
rect 1920 6686 1981 6687
rect 1920 6667 1953 6686
rect 1865 6666 1953 6667
rect 1973 6666 1981 6686
rect 1837 6658 1981 6666
rect 1837 6657 1873 6658
rect 1945 6657 1981 6658
rect 2047 6691 2084 6692
rect 2047 6690 2085 6691
rect 2047 6682 2111 6690
rect 2047 6662 2056 6682
rect 2076 6668 2111 6682
rect 2131 6668 2134 6688
rect 2076 6663 2134 6668
rect 2076 6662 2111 6663
rect 1313 6625 1350 6654
rect 1314 6623 1350 6625
rect 1526 6623 1563 6654
rect 878 6607 914 6608
rect 726 6577 735 6597
rect 755 6577 763 6597
rect 614 6568 670 6570
rect 614 6567 651 6568
rect 726 6567 763 6577
rect 822 6597 970 6607
rect 1070 6604 1166 6606
rect 822 6577 831 6597
rect 851 6577 941 6597
rect 961 6577 970 6597
rect 822 6568 970 6577
rect 1028 6597 1166 6604
rect 1314 6601 1563 6623
rect 1734 6622 1771 6654
rect 2047 6650 2111 6662
rect 2151 6624 2178 6802
rect 2010 6622 2178 6624
rect 1734 6618 2178 6622
rect 1028 6577 1037 6597
rect 1057 6577 1166 6597
rect 1734 6599 1783 6618
rect 1803 6599 2178 6618
rect 1734 6596 2178 6599
rect 2010 6595 2178 6596
rect 2199 6621 2230 7015
rect 2199 6595 2204 6621
rect 2223 6595 2230 6621
rect 2199 6592 2230 6595
rect 1028 6568 1166 6577
rect 822 6567 859 6568
rect 878 6516 914 6568
rect 933 6567 970 6568
rect 1029 6567 1066 6568
rect 349 6514 390 6515
rect 241 6507 390 6514
rect 241 6487 359 6507
rect 379 6487 390 6507
rect 241 6479 390 6487
rect 457 6511 816 6515
rect 457 6506 779 6511
rect 457 6482 570 6506
rect 594 6487 779 6506
rect 803 6487 816 6511
rect 594 6482 816 6487
rect 457 6479 816 6482
rect 878 6479 913 6516
rect 981 6513 1081 6516
rect 981 6509 1048 6513
rect 981 6483 993 6509
rect 1019 6487 1048 6509
rect 1074 6487 1081 6513
rect 1019 6483 1081 6487
rect 981 6479 1081 6483
rect 457 6458 488 6479
rect 878 6458 914 6479
rect 121 6449 158 6458
rect 300 6457 337 6458
rect 121 6431 130 6449
rect 148 6431 158 6449
rect 121 6421 158 6431
rect 122 6386 158 6421
rect 299 6448 337 6457
rect 299 6428 308 6448
rect 328 6428 337 6448
rect 299 6420 337 6428
rect 403 6452 488 6458
rect 513 6457 550 6458
rect 403 6432 411 6452
rect 431 6432 488 6452
rect 403 6424 488 6432
rect 512 6448 550 6457
rect 512 6428 521 6448
rect 541 6428 550 6448
rect 403 6423 439 6424
rect 512 6420 550 6428
rect 616 6452 701 6458
rect 721 6457 758 6458
rect 616 6432 624 6452
rect 644 6451 701 6452
rect 644 6432 673 6451
rect 616 6431 673 6432
rect 694 6431 701 6451
rect 616 6424 701 6431
rect 720 6448 758 6457
rect 720 6428 729 6448
rect 749 6428 758 6448
rect 616 6423 652 6424
rect 720 6420 758 6428
rect 824 6452 968 6458
rect 824 6432 832 6452
rect 852 6451 940 6452
rect 852 6432 880 6451
rect 824 6430 880 6432
rect 902 6432 940 6451
rect 960 6432 968 6452
rect 902 6430 968 6432
rect 824 6424 968 6430
rect 824 6423 860 6424
rect 932 6423 968 6424
rect 1034 6457 1071 6458
rect 1034 6456 1072 6457
rect 1034 6448 1098 6456
rect 1034 6428 1043 6448
rect 1063 6434 1098 6448
rect 1118 6434 1121 6454
rect 1063 6429 1121 6434
rect 1063 6428 1098 6429
rect 300 6391 337 6420
rect 120 6345 158 6386
rect 301 6389 337 6391
rect 513 6389 550 6420
rect 301 6367 550 6389
rect 721 6388 758 6420
rect 1034 6416 1098 6428
rect 1138 6390 1165 6568
rect 2749 6557 2786 6568
rect 2875 6561 2905 7562
rect 2968 7562 3412 7573
rect 2968 7560 3136 7562
rect 2968 7382 2995 7560
rect 3035 7522 3099 7534
rect 3375 7530 3412 7562
rect 3583 7561 3832 7583
rect 4225 7582 4373 7592
rect 4432 7612 4469 7622
rect 4544 7621 4581 7622
rect 4525 7619 4581 7621
rect 4432 7592 4440 7612
rect 4460 7592 4469 7612
rect 4281 7581 4317 7582
rect 3583 7530 3620 7561
rect 3796 7559 3832 7561
rect 3796 7530 3833 7559
rect 3035 7521 3070 7522
rect 3012 7516 3070 7521
rect 3012 7496 3015 7516
rect 3035 7502 3070 7516
rect 3090 7502 3099 7522
rect 3035 7494 3099 7502
rect 3061 7493 3099 7494
rect 3062 7492 3099 7493
rect 3165 7526 3201 7527
rect 3273 7526 3309 7527
rect 3165 7518 3309 7526
rect 3165 7498 3173 7518
rect 3193 7499 3225 7518
rect 3248 7499 3281 7518
rect 3193 7498 3281 7499
rect 3301 7498 3309 7518
rect 3165 7492 3309 7498
rect 3375 7522 3413 7530
rect 3481 7526 3517 7527
rect 3375 7502 3384 7522
rect 3404 7502 3413 7522
rect 3375 7493 3413 7502
rect 3432 7519 3517 7526
rect 3432 7499 3439 7519
rect 3460 7518 3517 7519
rect 3460 7499 3489 7518
rect 3432 7498 3489 7499
rect 3509 7498 3517 7518
rect 3375 7492 3412 7493
rect 3432 7492 3517 7498
rect 3583 7522 3621 7530
rect 3694 7526 3730 7527
rect 3583 7502 3592 7522
rect 3612 7502 3621 7522
rect 3583 7493 3621 7502
rect 3645 7518 3730 7526
rect 3645 7498 3702 7518
rect 3722 7498 3730 7518
rect 3583 7492 3620 7493
rect 3645 7492 3730 7498
rect 3796 7522 3834 7530
rect 4129 7522 4166 7523
rect 4432 7522 4469 7592
rect 4494 7612 4581 7619
rect 4494 7609 4552 7612
rect 4494 7589 4499 7609
rect 4520 7592 4552 7609
rect 4572 7592 4581 7612
rect 4520 7589 4581 7592
rect 4494 7582 4581 7589
rect 4640 7612 4677 7622
rect 4640 7592 4648 7612
rect 4668 7592 4677 7612
rect 4494 7581 4525 7582
rect 3796 7502 3805 7522
rect 3825 7502 3834 7522
rect 4128 7521 4469 7522
rect 3796 7493 3834 7502
rect 4053 7516 4469 7521
rect 4053 7496 4056 7516
rect 4076 7496 4469 7516
rect 4640 7521 4677 7592
rect 4707 7621 4738 7674
rect 5045 7672 5055 7690
rect 5073 7672 5084 7690
rect 5387 7709 6020 7718
rect 6746 7709 6777 7762
rect 6807 7791 6844 7862
rect 7015 7867 7408 7887
rect 7428 7867 7431 7887
rect 7015 7862 7431 7867
rect 7015 7861 7356 7862
rect 6959 7801 6990 7802
rect 6807 7771 6816 7791
rect 6836 7771 6844 7791
rect 6807 7761 6844 7771
rect 6903 7794 6990 7801
rect 6903 7791 6964 7794
rect 6903 7771 6912 7791
rect 6932 7774 6964 7791
rect 6985 7774 6990 7794
rect 6932 7771 6990 7774
rect 6903 7764 6990 7771
rect 7015 7791 7052 7861
rect 7318 7860 7355 7861
rect 7167 7801 7203 7802
rect 7015 7771 7024 7791
rect 7044 7771 7052 7791
rect 6903 7762 6959 7764
rect 6903 7761 6940 7762
rect 7015 7761 7052 7771
rect 7111 7791 7259 7801
rect 7359 7798 7455 7800
rect 7111 7771 7120 7791
rect 7140 7771 7230 7791
rect 7250 7771 7259 7791
rect 7111 7762 7259 7771
rect 7317 7791 7455 7798
rect 7317 7771 7326 7791
rect 7346 7771 7455 7791
rect 7317 7762 7455 7771
rect 7111 7761 7148 7762
rect 7167 7710 7203 7762
rect 7222 7761 7259 7762
rect 7318 7761 7355 7762
rect 5387 7691 5397 7709
rect 5415 7708 6020 7709
rect 6638 7708 6679 7709
rect 5415 7703 5436 7708
rect 5415 7691 5427 7703
rect 6530 7701 6679 7708
rect 5387 7683 5427 7691
rect 5470 7690 5496 7691
rect 5387 7681 5424 7683
rect 5470 7672 6024 7690
rect 6530 7681 6648 7701
rect 6668 7681 6679 7701
rect 6530 7673 6679 7681
rect 6746 7705 7105 7709
rect 6746 7700 7068 7705
rect 6746 7676 6859 7700
rect 6883 7681 7068 7700
rect 7092 7681 7105 7705
rect 6883 7676 7105 7681
rect 6746 7673 7105 7676
rect 7167 7673 7202 7710
rect 7270 7707 7370 7710
rect 7270 7703 7337 7707
rect 7270 7677 7282 7703
rect 7308 7681 7337 7703
rect 7363 7681 7370 7707
rect 7308 7677 7370 7681
rect 7270 7673 7370 7677
rect 5045 7663 5082 7672
rect 4757 7621 4794 7622
rect 4707 7612 4794 7621
rect 4707 7592 4765 7612
rect 4785 7592 4794 7612
rect 4707 7582 4794 7592
rect 4853 7612 4890 7622
rect 4853 7592 4861 7612
rect 4881 7592 4890 7612
rect 5390 7613 5427 7619
rect 5470 7613 5496 7672
rect 6003 7653 6024 7672
rect 5390 7610 5496 7613
rect 5048 7597 5085 7601
rect 4707 7581 4738 7582
rect 4853 7521 4890 7592
rect 4640 7497 4890 7521
rect 5046 7591 5085 7597
rect 5046 7573 5057 7591
rect 5075 7573 5085 7591
rect 5390 7592 5399 7610
rect 5417 7596 5496 7610
rect 5581 7628 5831 7652
rect 5417 7594 5493 7596
rect 5417 7592 5427 7594
rect 5390 7582 5427 7592
rect 5046 7564 5085 7573
rect 3796 7492 3833 7493
rect 3219 7471 3255 7492
rect 3645 7471 3676 7492
rect 4432 7473 4469 7496
rect 5046 7486 5081 7564
rect 5395 7517 5426 7582
rect 5581 7557 5618 7628
rect 5733 7567 5764 7568
rect 5581 7537 5590 7557
rect 5610 7537 5618 7557
rect 5581 7527 5618 7537
rect 5677 7557 5764 7567
rect 5677 7537 5686 7557
rect 5706 7537 5764 7557
rect 5677 7528 5764 7537
rect 5677 7527 5714 7528
rect 5043 7476 5081 7486
rect 5394 7508 5431 7517
rect 5394 7490 5404 7508
rect 5422 7490 5431 7508
rect 5394 7480 5431 7490
rect 4432 7472 4602 7473
rect 5043 7472 5053 7476
rect 3052 7467 3152 7471
rect 3052 7463 3114 7467
rect 3052 7437 3059 7463
rect 3085 7441 3114 7463
rect 3140 7441 3152 7467
rect 3085 7437 3152 7441
rect 3052 7434 3152 7437
rect 3220 7434 3255 7471
rect 3317 7468 3676 7471
rect 3317 7463 3539 7468
rect 3317 7439 3330 7463
rect 3354 7444 3539 7463
rect 3563 7444 3676 7468
rect 3354 7439 3676 7444
rect 3317 7435 3676 7439
rect 3743 7463 3892 7471
rect 3743 7443 3754 7463
rect 3774 7443 3892 7463
rect 4432 7458 5053 7472
rect 5071 7458 5081 7476
rect 5733 7475 5764 7528
rect 5794 7557 5831 7628
rect 6002 7633 6395 7653
rect 6415 7633 6418 7653
rect 6746 7652 6777 7673
rect 7167 7652 7203 7673
rect 6589 7651 6626 7652
rect 6002 7628 6418 7633
rect 6588 7642 6626 7651
rect 6002 7627 6343 7628
rect 5946 7567 5977 7568
rect 5794 7537 5803 7557
rect 5823 7537 5831 7557
rect 5794 7527 5831 7537
rect 5890 7560 5977 7567
rect 5890 7557 5951 7560
rect 5890 7537 5899 7557
rect 5919 7540 5951 7557
rect 5972 7540 5977 7560
rect 5919 7537 5977 7540
rect 5890 7530 5977 7537
rect 6002 7557 6039 7627
rect 6305 7626 6342 7627
rect 6588 7622 6597 7642
rect 6617 7622 6626 7642
rect 6588 7614 6626 7622
rect 6692 7646 6777 7652
rect 6802 7651 6839 7652
rect 6692 7626 6700 7646
rect 6720 7626 6777 7646
rect 6692 7618 6777 7626
rect 6801 7642 6839 7651
rect 6801 7622 6810 7642
rect 6830 7622 6839 7642
rect 6692 7617 6728 7618
rect 6801 7614 6839 7622
rect 6905 7646 6990 7652
rect 7010 7651 7047 7652
rect 6905 7626 6913 7646
rect 6933 7645 6990 7646
rect 6933 7626 6962 7645
rect 6905 7625 6962 7626
rect 6983 7625 6990 7645
rect 6905 7618 6990 7625
rect 7009 7642 7047 7651
rect 7009 7622 7018 7642
rect 7038 7622 7047 7642
rect 6905 7617 6941 7618
rect 7009 7614 7047 7622
rect 7113 7646 7257 7652
rect 7113 7626 7121 7646
rect 7141 7626 7173 7646
rect 7197 7626 7229 7646
rect 7249 7626 7257 7646
rect 7113 7618 7257 7626
rect 7113 7617 7149 7618
rect 7221 7617 7257 7618
rect 7323 7651 7360 7652
rect 7323 7650 7361 7651
rect 7323 7642 7387 7650
rect 7323 7622 7332 7642
rect 7352 7628 7387 7642
rect 7407 7628 7410 7648
rect 7352 7623 7410 7628
rect 7352 7622 7387 7623
rect 6589 7585 6626 7614
rect 6590 7583 6626 7585
rect 6802 7583 6839 7614
rect 6154 7567 6190 7568
rect 6002 7537 6011 7557
rect 6031 7537 6039 7557
rect 5890 7528 5946 7530
rect 5890 7527 5927 7528
rect 6002 7527 6039 7537
rect 6098 7557 6246 7567
rect 6346 7564 6442 7566
rect 6098 7537 6107 7557
rect 6127 7537 6217 7557
rect 6237 7537 6246 7557
rect 6098 7528 6246 7537
rect 6304 7557 6442 7564
rect 6590 7561 6839 7583
rect 7010 7582 7047 7614
rect 7323 7610 7387 7622
rect 7427 7584 7454 7762
rect 7286 7582 7454 7584
rect 7010 7578 7454 7582
rect 6304 7537 6313 7557
rect 6333 7537 6442 7557
rect 7010 7559 7059 7578
rect 7079 7559 7454 7578
rect 7010 7556 7454 7559
rect 7286 7555 7454 7556
rect 8154 7569 8183 7571
rect 8154 7564 8186 7569
rect 8154 7546 8161 7564
rect 8181 7546 8186 7564
rect 8247 7568 8278 7962
rect 8299 7987 8467 7988
rect 8299 7984 8743 7987
rect 8299 7965 8674 7984
rect 8694 7965 8743 7984
rect 9311 7986 9420 8006
rect 9440 7986 9449 8006
rect 8299 7961 8743 7965
rect 8299 7959 8467 7961
rect 8299 7781 8326 7959
rect 8366 7921 8430 7933
rect 8706 7929 8743 7961
rect 8914 7960 9163 7982
rect 9311 7979 9449 7986
rect 9507 8006 9655 8015
rect 9507 7986 9516 8006
rect 9536 7986 9626 8006
rect 9646 7986 9655 8006
rect 9311 7977 9407 7979
rect 9507 7976 9655 7986
rect 9714 8006 9751 8016
rect 9826 8015 9863 8016
rect 9807 8013 9863 8015
rect 9714 7986 9722 8006
rect 9742 7986 9751 8006
rect 9563 7975 9599 7976
rect 8914 7929 8951 7960
rect 9127 7958 9163 7960
rect 9127 7929 9164 7958
rect 8366 7920 8401 7921
rect 8343 7915 8401 7920
rect 8343 7895 8346 7915
rect 8366 7901 8401 7915
rect 8421 7901 8430 7921
rect 8366 7893 8430 7901
rect 8392 7892 8430 7893
rect 8393 7891 8430 7892
rect 8496 7925 8532 7926
rect 8604 7925 8640 7926
rect 8496 7917 8640 7925
rect 8496 7897 8504 7917
rect 8524 7916 8612 7917
rect 8524 7897 8557 7916
rect 8496 7896 8557 7897
rect 8581 7897 8612 7916
rect 8632 7897 8640 7917
rect 8581 7896 8640 7897
rect 8496 7891 8640 7896
rect 8706 7921 8744 7929
rect 8812 7925 8848 7926
rect 8706 7901 8715 7921
rect 8735 7901 8744 7921
rect 8706 7892 8744 7901
rect 8763 7918 8848 7925
rect 8763 7898 8770 7918
rect 8791 7917 8848 7918
rect 8791 7898 8820 7917
rect 8763 7897 8820 7898
rect 8840 7897 8848 7917
rect 8706 7891 8743 7892
rect 8763 7891 8848 7897
rect 8914 7921 8952 7929
rect 9025 7925 9061 7926
rect 8914 7901 8923 7921
rect 8943 7901 8952 7921
rect 8914 7892 8952 7901
rect 8976 7917 9061 7925
rect 8976 7897 9033 7917
rect 9053 7897 9061 7917
rect 8914 7891 8951 7892
rect 8976 7891 9061 7897
rect 9127 7921 9165 7929
rect 9127 7901 9136 7921
rect 9156 7901 9165 7921
rect 9411 7916 9448 7917
rect 9714 7916 9751 7986
rect 9776 8006 9863 8013
rect 9776 8003 9834 8006
rect 9776 7983 9781 8003
rect 9802 7986 9834 8003
rect 9854 7986 9863 8006
rect 9802 7983 9863 7986
rect 9776 7976 9863 7983
rect 9922 8006 9959 8016
rect 9922 7986 9930 8006
rect 9950 7986 9959 8006
rect 9776 7975 9807 7976
rect 9410 7915 9751 7916
rect 9127 7892 9165 7901
rect 9335 7910 9751 7915
rect 9127 7891 9164 7892
rect 8550 7870 8586 7891
rect 8976 7870 9007 7891
rect 9335 7890 9338 7910
rect 9358 7890 9751 7910
rect 9922 7915 9959 7986
rect 9989 8015 10020 8068
rect 10322 8053 10359 8063
rect 10322 8035 10331 8053
rect 10349 8035 10359 8053
rect 10322 8026 10359 8035
rect 10039 8015 10076 8016
rect 9989 8006 10076 8015
rect 9989 7986 10047 8006
rect 10067 7986 10076 8006
rect 9989 7976 10076 7986
rect 10135 8006 10172 8016
rect 10135 7986 10143 8006
rect 10163 7986 10172 8006
rect 9989 7975 10020 7976
rect 10135 7915 10172 7986
rect 10327 7961 10358 8026
rect 10326 7951 10363 7961
rect 10326 7949 10336 7951
rect 10260 7947 10336 7949
rect 9922 7891 10172 7915
rect 10257 7933 10336 7947
rect 10354 7933 10363 7951
rect 10257 7930 10363 7933
rect 9729 7871 9750 7890
rect 10257 7871 10283 7930
rect 10326 7924 10363 7930
rect 8383 7866 8483 7870
rect 8383 7862 8445 7866
rect 8383 7836 8390 7862
rect 8416 7840 8445 7862
rect 8471 7840 8483 7866
rect 8416 7836 8483 7840
rect 8383 7833 8483 7836
rect 8551 7833 8586 7870
rect 8648 7867 9007 7870
rect 8648 7862 8870 7867
rect 8648 7838 8661 7862
rect 8685 7843 8870 7862
rect 8894 7843 9007 7867
rect 8685 7838 9007 7843
rect 8648 7834 9007 7838
rect 9074 7862 9223 7870
rect 9074 7842 9085 7862
rect 9105 7842 9223 7862
rect 9729 7853 10283 7871
rect 10329 7860 10366 7862
rect 10257 7852 10283 7853
rect 10326 7852 10366 7860
rect 9074 7835 9223 7842
rect 10326 7840 10338 7852
rect 10317 7835 10338 7840
rect 9074 7834 9115 7835
rect 9733 7834 10338 7835
rect 10356 7834 10366 7852
rect 8398 7781 8435 7782
rect 8494 7781 8531 7782
rect 8550 7781 8586 7833
rect 8605 7781 8642 7782
rect 8298 7772 8436 7781
rect 8298 7752 8407 7772
rect 8427 7752 8436 7772
rect 8298 7745 8436 7752
rect 8494 7772 8642 7781
rect 8494 7752 8503 7772
rect 8523 7752 8613 7772
rect 8633 7752 8642 7772
rect 8298 7743 8394 7745
rect 8494 7742 8642 7752
rect 8701 7772 8738 7782
rect 8813 7781 8850 7782
rect 8794 7779 8850 7781
rect 8701 7752 8709 7772
rect 8729 7752 8738 7772
rect 8550 7741 8586 7742
rect 8398 7682 8435 7683
rect 8701 7682 8738 7752
rect 8763 7772 8850 7779
rect 8763 7769 8821 7772
rect 8763 7749 8768 7769
rect 8789 7752 8821 7769
rect 8841 7752 8850 7772
rect 8789 7749 8850 7752
rect 8763 7742 8850 7749
rect 8909 7772 8946 7782
rect 8909 7752 8917 7772
rect 8937 7752 8946 7772
rect 8763 7741 8794 7742
rect 8397 7681 8738 7682
rect 8322 7676 8738 7681
rect 8322 7656 8325 7676
rect 8345 7656 8738 7676
rect 8909 7681 8946 7752
rect 8976 7781 9007 7834
rect 9733 7825 10366 7834
rect 9733 7818 10365 7825
rect 9733 7816 9795 7818
rect 9311 7806 9479 7807
rect 9733 7806 9755 7816
rect 9026 7781 9063 7782
rect 8976 7772 9063 7781
rect 8976 7752 9034 7772
rect 9054 7752 9063 7772
rect 8976 7742 9063 7752
rect 9122 7772 9159 7782
rect 9122 7752 9130 7772
rect 9150 7752 9159 7772
rect 8976 7741 9007 7742
rect 9122 7681 9159 7752
rect 8909 7657 9159 7681
rect 9311 7780 9755 7806
rect 9311 7778 9479 7780
rect 9311 7600 9338 7778
rect 9378 7740 9442 7752
rect 9718 7748 9755 7780
rect 9926 7779 10175 7801
rect 9926 7748 9963 7779
rect 10139 7777 10175 7779
rect 10139 7748 10176 7777
rect 9378 7739 9413 7740
rect 9355 7734 9413 7739
rect 9355 7714 9358 7734
rect 9378 7720 9413 7734
rect 9433 7720 9442 7740
rect 9378 7712 9442 7720
rect 9404 7711 9442 7712
rect 9405 7710 9442 7711
rect 9508 7744 9544 7745
rect 9616 7744 9652 7745
rect 9508 7736 9652 7744
rect 9508 7716 9516 7736
rect 9536 7716 9565 7736
rect 9508 7715 9565 7716
rect 9587 7716 9624 7736
rect 9644 7716 9652 7736
rect 9587 7715 9652 7716
rect 9508 7710 9652 7715
rect 9718 7740 9756 7748
rect 9824 7744 9860 7745
rect 9718 7720 9727 7740
rect 9747 7720 9756 7740
rect 9718 7711 9756 7720
rect 9775 7737 9860 7744
rect 9775 7717 9782 7737
rect 9803 7736 9860 7737
rect 9803 7717 9832 7736
rect 9775 7716 9832 7717
rect 9852 7716 9860 7736
rect 9718 7710 9755 7711
rect 9775 7710 9860 7716
rect 9926 7740 9964 7748
rect 10037 7744 10073 7745
rect 9926 7720 9935 7740
rect 9955 7720 9964 7740
rect 9926 7711 9964 7720
rect 9988 7736 10073 7744
rect 9988 7716 10045 7736
rect 10065 7716 10073 7736
rect 9926 7710 9963 7711
rect 9988 7710 10073 7716
rect 10139 7740 10177 7748
rect 10139 7720 10148 7740
rect 10168 7720 10177 7740
rect 10139 7711 10177 7720
rect 10139 7710 10176 7711
rect 9562 7689 9598 7710
rect 9988 7689 10019 7710
rect 9395 7685 9495 7689
rect 9395 7681 9457 7685
rect 9395 7655 9402 7681
rect 9428 7659 9457 7681
rect 9483 7659 9495 7685
rect 9428 7655 9495 7659
rect 9395 7652 9495 7655
rect 9563 7652 9598 7689
rect 9660 7686 10019 7689
rect 9660 7681 9882 7686
rect 9660 7657 9673 7681
rect 9697 7662 9882 7681
rect 9906 7662 10019 7686
rect 9697 7657 10019 7662
rect 9660 7653 10019 7657
rect 10086 7681 10235 7689
rect 10086 7661 10097 7681
rect 10117 7661 10235 7681
rect 10086 7654 10235 7661
rect 10326 7669 10365 7818
rect 10086 7653 10127 7654
rect 9410 7600 9447 7601
rect 9506 7600 9543 7601
rect 9562 7600 9598 7652
rect 9617 7600 9654 7601
rect 9310 7591 9448 7600
rect 9310 7571 9419 7591
rect 9439 7571 9448 7591
rect 8247 7567 8417 7568
rect 8247 7552 8693 7567
rect 9310 7564 9448 7571
rect 9506 7591 9654 7600
rect 9506 7571 9515 7591
rect 9535 7571 9625 7591
rect 9645 7571 9654 7591
rect 9310 7562 9406 7564
rect 8154 7541 8186 7546
rect 6304 7528 6442 7537
rect 6098 7527 6135 7528
rect 6154 7476 6190 7528
rect 6209 7527 6246 7528
rect 6305 7527 6342 7528
rect 5625 7474 5666 7475
rect 4432 7452 5081 7458
rect 5517 7467 5666 7474
rect 4432 7451 5080 7452
rect 5043 7449 5080 7451
rect 3743 7436 3892 7443
rect 5517 7447 5635 7467
rect 5655 7447 5666 7467
rect 5517 7439 5666 7447
rect 5733 7471 6092 7475
rect 5733 7466 6055 7471
rect 5733 7442 5846 7466
rect 5870 7447 6055 7466
rect 6079 7447 6092 7471
rect 5870 7442 6092 7447
rect 5733 7439 6092 7442
rect 6154 7439 6189 7476
rect 6257 7473 6357 7476
rect 6257 7469 6324 7473
rect 6257 7443 6269 7469
rect 6295 7447 6324 7469
rect 6350 7447 6357 7473
rect 6295 7443 6357 7447
rect 6257 7439 6357 7443
rect 3743 7435 3784 7436
rect 3067 7382 3104 7383
rect 3163 7382 3200 7383
rect 3219 7382 3255 7434
rect 3274 7382 3311 7383
rect 2967 7373 3105 7382
rect 2967 7353 3076 7373
rect 3096 7353 3105 7373
rect 2967 7346 3105 7353
rect 3163 7373 3311 7382
rect 3163 7353 3172 7373
rect 3192 7353 3282 7373
rect 3302 7353 3311 7373
rect 2967 7344 3063 7346
rect 3163 7343 3311 7353
rect 3370 7373 3407 7383
rect 3482 7382 3519 7383
rect 3463 7380 3519 7382
rect 3370 7353 3378 7373
rect 3398 7353 3407 7373
rect 3219 7342 3255 7343
rect 3067 7283 3104 7284
rect 3370 7283 3407 7353
rect 3432 7373 3519 7380
rect 3432 7370 3490 7373
rect 3432 7350 3437 7370
rect 3458 7353 3490 7370
rect 3510 7353 3519 7373
rect 3458 7350 3519 7353
rect 3432 7343 3519 7350
rect 3578 7373 3615 7383
rect 3578 7353 3586 7373
rect 3606 7353 3615 7373
rect 3432 7342 3463 7343
rect 3066 7282 3407 7283
rect 2991 7277 3407 7282
rect 2991 7257 2994 7277
rect 3014 7257 3407 7277
rect 3578 7282 3615 7353
rect 3645 7382 3676 7435
rect 5733 7418 5764 7439
rect 6154 7418 6190 7439
rect 5397 7409 5434 7418
rect 5576 7417 5613 7418
rect 5397 7391 5406 7409
rect 5424 7391 5434 7409
rect 3695 7382 3732 7383
rect 3645 7373 3732 7382
rect 3645 7353 3703 7373
rect 3723 7353 3732 7373
rect 3645 7343 3732 7353
rect 3791 7373 3828 7383
rect 3791 7353 3799 7373
rect 3819 7353 3828 7373
rect 3645 7342 3676 7343
rect 3791 7282 3828 7353
rect 5046 7377 5083 7387
rect 5397 7381 5434 7391
rect 5046 7359 5055 7377
rect 5073 7359 5083 7377
rect 5046 7350 5083 7359
rect 5046 7326 5081 7350
rect 5398 7346 5434 7381
rect 5575 7408 5613 7417
rect 5575 7388 5584 7408
rect 5604 7388 5613 7408
rect 5575 7380 5613 7388
rect 5679 7412 5764 7418
rect 5789 7417 5826 7418
rect 5679 7392 5687 7412
rect 5707 7392 5764 7412
rect 5679 7384 5764 7392
rect 5788 7408 5826 7417
rect 5788 7388 5797 7408
rect 5817 7388 5826 7408
rect 5679 7383 5715 7384
rect 5788 7380 5826 7388
rect 5892 7412 5977 7418
rect 5997 7417 6034 7418
rect 5892 7392 5900 7412
rect 5920 7411 5977 7412
rect 5920 7392 5949 7411
rect 5892 7391 5949 7392
rect 5970 7391 5977 7411
rect 5892 7384 5977 7391
rect 5996 7408 6034 7417
rect 5996 7388 6005 7408
rect 6025 7388 6034 7408
rect 5892 7383 5928 7384
rect 5996 7380 6034 7388
rect 6100 7412 6244 7418
rect 6100 7392 6108 7412
rect 6128 7411 6216 7412
rect 6128 7392 6156 7411
rect 6100 7390 6156 7392
rect 6178 7392 6216 7411
rect 6236 7392 6244 7412
rect 6178 7390 6244 7392
rect 6100 7384 6244 7390
rect 6100 7383 6136 7384
rect 6208 7383 6244 7384
rect 6310 7417 6347 7418
rect 6310 7416 6348 7417
rect 6310 7408 6374 7416
rect 6310 7388 6319 7408
rect 6339 7394 6374 7408
rect 6394 7394 6397 7414
rect 6339 7389 6397 7394
rect 6339 7388 6374 7389
rect 5576 7351 5613 7380
rect 5044 7302 5081 7326
rect 5043 7296 5081 7302
rect 3578 7258 3828 7282
rect 4454 7278 5081 7296
rect 4036 7261 4204 7262
rect 4455 7261 4479 7278
rect 4036 7235 4480 7261
rect 4036 7233 4204 7235
rect 4036 7055 4063 7233
rect 4103 7195 4167 7207
rect 4443 7203 4480 7235
rect 4651 7234 4900 7256
rect 4651 7203 4688 7234
rect 4864 7232 4900 7234
rect 5043 7237 5081 7278
rect 5396 7305 5434 7346
rect 5577 7349 5613 7351
rect 5789 7349 5826 7380
rect 5577 7327 5826 7349
rect 5997 7348 6034 7380
rect 6310 7376 6374 7388
rect 6414 7350 6441 7528
rect 6273 7348 6441 7350
rect 5997 7322 6441 7348
rect 5998 7305 6022 7322
rect 6273 7321 6441 7322
rect 5396 7287 6023 7305
rect 6649 7301 6899 7325
rect 5396 7281 5434 7287
rect 5396 7257 5433 7281
rect 4864 7203 4901 7232
rect 4103 7194 4138 7195
rect 4080 7189 4138 7194
rect 4080 7169 4083 7189
rect 4103 7175 4138 7189
rect 4158 7175 4167 7195
rect 4103 7167 4167 7175
rect 4129 7166 4167 7167
rect 4130 7165 4167 7166
rect 4233 7199 4269 7200
rect 4341 7199 4377 7200
rect 4233 7193 4377 7199
rect 4233 7191 4299 7193
rect 4233 7171 4241 7191
rect 4261 7172 4299 7191
rect 4321 7191 4377 7193
rect 4321 7172 4349 7191
rect 4261 7171 4349 7172
rect 4369 7171 4377 7191
rect 4233 7165 4377 7171
rect 4443 7195 4481 7203
rect 4549 7199 4585 7200
rect 4443 7175 4452 7195
rect 4472 7175 4481 7195
rect 4443 7166 4481 7175
rect 4500 7192 4585 7199
rect 4500 7172 4507 7192
rect 4528 7191 4585 7192
rect 4528 7172 4557 7191
rect 4500 7171 4557 7172
rect 4577 7171 4585 7191
rect 4443 7165 4480 7166
rect 4500 7165 4585 7171
rect 4651 7195 4689 7203
rect 4762 7199 4798 7200
rect 4651 7175 4660 7195
rect 4680 7175 4689 7195
rect 4651 7166 4689 7175
rect 4713 7191 4798 7199
rect 4713 7171 4770 7191
rect 4790 7171 4798 7191
rect 4651 7165 4688 7166
rect 4713 7165 4798 7171
rect 4864 7195 4902 7203
rect 4864 7175 4873 7195
rect 4893 7175 4902 7195
rect 4864 7166 4902 7175
rect 5043 7202 5079 7237
rect 5396 7233 5431 7257
rect 5394 7224 5431 7233
rect 5394 7206 5404 7224
rect 5422 7206 5431 7224
rect 5043 7192 5080 7202
rect 5394 7196 5431 7206
rect 6649 7230 6686 7301
rect 6801 7240 6832 7241
rect 6649 7210 6658 7230
rect 6678 7210 6686 7230
rect 6649 7200 6686 7210
rect 6745 7230 6832 7240
rect 6745 7210 6754 7230
rect 6774 7210 6832 7230
rect 6745 7201 6832 7210
rect 6745 7200 6782 7201
rect 5043 7174 5053 7192
rect 5071 7174 5080 7192
rect 4864 7165 4901 7166
rect 5043 7165 5080 7174
rect 4287 7144 4323 7165
rect 4713 7144 4744 7165
rect 6801 7148 6832 7201
rect 6862 7230 6899 7301
rect 7070 7306 7463 7326
rect 7483 7306 7486 7326
rect 7070 7301 7486 7306
rect 7070 7300 7411 7301
rect 7014 7240 7045 7241
rect 6862 7210 6871 7230
rect 6891 7210 6899 7230
rect 6862 7200 6899 7210
rect 6958 7233 7045 7240
rect 6958 7230 7019 7233
rect 6958 7210 6967 7230
rect 6987 7213 7019 7230
rect 7040 7213 7045 7233
rect 6987 7210 7045 7213
rect 6958 7203 7045 7210
rect 7070 7230 7107 7300
rect 7373 7299 7410 7300
rect 7222 7240 7258 7241
rect 7070 7210 7079 7230
rect 7099 7210 7107 7230
rect 6958 7201 7014 7203
rect 6958 7200 6995 7201
rect 7070 7200 7107 7210
rect 7166 7230 7314 7240
rect 7414 7237 7510 7239
rect 7166 7210 7175 7230
rect 7195 7210 7285 7230
rect 7305 7210 7314 7230
rect 7166 7201 7314 7210
rect 7372 7230 7510 7237
rect 7372 7210 7381 7230
rect 7401 7210 7510 7230
rect 7372 7201 7510 7210
rect 7166 7200 7203 7201
rect 7222 7149 7258 7201
rect 7277 7200 7314 7201
rect 7373 7200 7410 7201
rect 6693 7147 6734 7148
rect 4120 7140 4220 7144
rect 4120 7136 4182 7140
rect 4120 7110 4127 7136
rect 4153 7114 4182 7136
rect 4208 7114 4220 7140
rect 4153 7110 4220 7114
rect 4120 7107 4220 7110
rect 4288 7107 4323 7144
rect 4385 7141 4744 7144
rect 4385 7136 4607 7141
rect 4385 7112 4398 7136
rect 4422 7117 4607 7136
rect 4631 7117 4744 7141
rect 4422 7112 4744 7117
rect 4385 7108 4744 7112
rect 4811 7136 4960 7144
rect 4811 7116 4822 7136
rect 4842 7116 4960 7136
rect 6585 7140 6734 7147
rect 5397 7132 5434 7134
rect 5397 7131 6045 7132
rect 4811 7109 4960 7116
rect 5396 7125 6045 7131
rect 4811 7108 4852 7109
rect 4135 7055 4172 7056
rect 4231 7055 4268 7056
rect 4287 7055 4323 7107
rect 4342 7055 4379 7056
rect 4035 7046 4173 7055
rect 3023 7027 3191 7028
rect 3023 7024 3467 7027
rect 3023 7005 3398 7024
rect 3418 7005 3467 7024
rect 4035 7026 4144 7046
rect 4164 7026 4173 7046
rect 3023 7001 3467 7005
rect 3023 6999 3191 7001
rect 3023 6821 3050 6999
rect 3090 6961 3154 6973
rect 3430 6969 3467 7001
rect 3638 7000 3887 7022
rect 4035 7019 4173 7026
rect 4231 7046 4379 7055
rect 4231 7026 4240 7046
rect 4260 7026 4350 7046
rect 4370 7026 4379 7046
rect 4035 7017 4131 7019
rect 4231 7016 4379 7026
rect 4438 7046 4475 7056
rect 4550 7055 4587 7056
rect 4531 7053 4587 7055
rect 4438 7026 4446 7046
rect 4466 7026 4475 7046
rect 4287 7015 4323 7016
rect 3638 6969 3675 7000
rect 3851 6998 3887 7000
rect 3851 6969 3888 6998
rect 3090 6960 3125 6961
rect 3067 6955 3125 6960
rect 3067 6935 3070 6955
rect 3090 6941 3125 6955
rect 3145 6941 3154 6961
rect 3090 6933 3154 6941
rect 3116 6932 3154 6933
rect 3117 6931 3154 6932
rect 3220 6965 3256 6966
rect 3328 6965 3364 6966
rect 3220 6957 3364 6965
rect 3220 6937 3228 6957
rect 3248 6937 3280 6957
rect 3304 6937 3336 6957
rect 3356 6937 3364 6957
rect 3220 6931 3364 6937
rect 3430 6961 3468 6969
rect 3536 6965 3572 6966
rect 3430 6941 3439 6961
rect 3459 6941 3468 6961
rect 3430 6932 3468 6941
rect 3487 6958 3572 6965
rect 3487 6938 3494 6958
rect 3515 6957 3572 6958
rect 3515 6938 3544 6957
rect 3487 6937 3544 6938
rect 3564 6937 3572 6957
rect 3430 6931 3467 6932
rect 3487 6931 3572 6937
rect 3638 6961 3676 6969
rect 3749 6965 3785 6966
rect 3638 6941 3647 6961
rect 3667 6941 3676 6961
rect 3638 6932 3676 6941
rect 3700 6957 3785 6965
rect 3700 6937 3757 6957
rect 3777 6937 3785 6957
rect 3638 6931 3675 6932
rect 3700 6931 3785 6937
rect 3851 6961 3889 6969
rect 3851 6941 3860 6961
rect 3880 6941 3889 6961
rect 4135 6956 4172 6957
rect 4438 6956 4475 7026
rect 4500 7046 4587 7053
rect 4500 7043 4558 7046
rect 4500 7023 4505 7043
rect 4526 7026 4558 7043
rect 4578 7026 4587 7046
rect 4526 7023 4587 7026
rect 4500 7016 4587 7023
rect 4646 7046 4683 7056
rect 4646 7026 4654 7046
rect 4674 7026 4683 7046
rect 4500 7015 4531 7016
rect 4134 6955 4475 6956
rect 3851 6932 3889 6941
rect 4059 6950 4475 6955
rect 3851 6931 3888 6932
rect 3274 6910 3310 6931
rect 3700 6910 3731 6931
rect 4059 6930 4062 6950
rect 4082 6930 4475 6950
rect 4646 6955 4683 7026
rect 4713 7055 4744 7108
rect 5396 7107 5406 7125
rect 5424 7111 6045 7125
rect 6585 7120 6703 7140
rect 6723 7120 6734 7140
rect 6585 7112 6734 7120
rect 6801 7144 7160 7148
rect 6801 7139 7123 7144
rect 6801 7115 6914 7139
rect 6938 7120 7123 7139
rect 7147 7120 7160 7144
rect 6938 7115 7160 7120
rect 6801 7112 7160 7115
rect 7222 7112 7257 7149
rect 7325 7146 7425 7149
rect 7325 7142 7392 7146
rect 7325 7116 7337 7142
rect 7363 7120 7392 7142
rect 7418 7120 7425 7146
rect 7363 7116 7425 7120
rect 7325 7112 7425 7116
rect 5424 7107 5434 7111
rect 5875 7110 6045 7111
rect 5046 7093 5083 7103
rect 5046 7075 5055 7093
rect 5073 7075 5083 7093
rect 5046 7066 5083 7075
rect 5396 7097 5434 7107
rect 4763 7055 4800 7056
rect 4713 7046 4800 7055
rect 4713 7026 4771 7046
rect 4791 7026 4800 7046
rect 4713 7016 4800 7026
rect 4859 7046 4896 7056
rect 4859 7026 4867 7046
rect 4887 7026 4896 7046
rect 4713 7015 4744 7016
rect 4859 6955 4896 7026
rect 5051 7001 5082 7066
rect 5396 7019 5431 7097
rect 6008 7087 6045 7110
rect 6801 7091 6832 7112
rect 7222 7091 7258 7112
rect 6644 7090 6681 7091
rect 5392 7010 5431 7019
rect 5050 6991 5087 7001
rect 5050 6989 5060 6991
rect 4984 6987 5060 6989
rect 4646 6931 4896 6955
rect 4981 6973 5060 6987
rect 5078 6973 5087 6991
rect 5392 6992 5402 7010
rect 5420 6992 5431 7010
rect 5392 6986 5431 6992
rect 5587 7062 5837 7086
rect 5587 6991 5624 7062
rect 5739 7001 5770 7002
rect 5392 6982 5429 6986
rect 4981 6970 5087 6973
rect 4453 6911 4474 6930
rect 4981 6911 5007 6970
rect 5050 6964 5087 6970
rect 5587 6971 5596 6991
rect 5616 6971 5624 6991
rect 5587 6961 5624 6971
rect 5683 6991 5770 7001
rect 5683 6971 5692 6991
rect 5712 6971 5770 6991
rect 5683 6962 5770 6971
rect 5683 6961 5720 6962
rect 5395 6911 5432 6920
rect 3107 6906 3207 6910
rect 3107 6902 3169 6906
rect 3107 6876 3114 6902
rect 3140 6880 3169 6902
rect 3195 6880 3207 6906
rect 3140 6876 3207 6880
rect 3107 6873 3207 6876
rect 3275 6873 3310 6910
rect 3372 6907 3731 6910
rect 3372 6902 3594 6907
rect 3372 6878 3385 6902
rect 3409 6883 3594 6902
rect 3618 6883 3731 6907
rect 3409 6878 3731 6883
rect 3372 6874 3731 6878
rect 3798 6902 3947 6910
rect 3798 6882 3809 6902
rect 3829 6882 3947 6902
rect 4453 6893 5007 6911
rect 5053 6900 5090 6902
rect 4981 6892 5007 6893
rect 5050 6892 5090 6900
rect 3798 6875 3947 6882
rect 5050 6880 5062 6892
rect 5041 6875 5062 6880
rect 3798 6874 3839 6875
rect 4457 6874 5062 6875
rect 5080 6874 5090 6892
rect 3122 6821 3159 6822
rect 3218 6821 3255 6822
rect 3274 6821 3310 6873
rect 3329 6821 3366 6822
rect 3022 6812 3160 6821
rect 3022 6792 3131 6812
rect 3151 6792 3160 6812
rect 3022 6785 3160 6792
rect 3218 6812 3366 6821
rect 3218 6792 3227 6812
rect 3247 6792 3337 6812
rect 3357 6792 3366 6812
rect 3022 6783 3118 6785
rect 3218 6782 3366 6792
rect 3425 6812 3462 6822
rect 3537 6821 3574 6822
rect 3518 6819 3574 6821
rect 3425 6792 3433 6812
rect 3453 6792 3462 6812
rect 3274 6781 3310 6782
rect 3122 6722 3159 6723
rect 3425 6722 3462 6792
rect 3487 6812 3574 6819
rect 3487 6809 3545 6812
rect 3487 6789 3492 6809
rect 3513 6792 3545 6809
rect 3565 6792 3574 6812
rect 3513 6789 3574 6792
rect 3487 6782 3574 6789
rect 3633 6812 3670 6822
rect 3633 6792 3641 6812
rect 3661 6792 3670 6812
rect 3487 6781 3518 6782
rect 3121 6721 3462 6722
rect 3046 6716 3462 6721
rect 3046 6696 3049 6716
rect 3069 6696 3462 6716
rect 3633 6721 3670 6792
rect 3700 6821 3731 6874
rect 4457 6865 5090 6874
rect 5393 6893 5404 6911
rect 5422 6893 5432 6911
rect 5739 6909 5770 6962
rect 5800 6991 5837 7062
rect 6008 7067 6401 7087
rect 6421 7067 6424 7087
rect 6008 7062 6424 7067
rect 6643 7081 6681 7090
rect 6008 7061 6349 7062
rect 6643 7061 6652 7081
rect 6672 7061 6681 7081
rect 5952 7001 5983 7002
rect 5800 6971 5809 6991
rect 5829 6971 5837 6991
rect 5800 6961 5837 6971
rect 5896 6994 5983 7001
rect 5896 6991 5957 6994
rect 5896 6971 5905 6991
rect 5925 6974 5957 6991
rect 5978 6974 5983 6994
rect 5925 6971 5983 6974
rect 5896 6964 5983 6971
rect 6008 6991 6045 7061
rect 6311 7060 6348 7061
rect 6643 7053 6681 7061
rect 6747 7085 6832 7091
rect 6857 7090 6894 7091
rect 6747 7065 6755 7085
rect 6775 7065 6832 7085
rect 6747 7057 6832 7065
rect 6856 7081 6894 7090
rect 6856 7061 6865 7081
rect 6885 7061 6894 7081
rect 6747 7056 6783 7057
rect 6856 7053 6894 7061
rect 6960 7085 7045 7091
rect 7065 7090 7102 7091
rect 6960 7065 6968 7085
rect 6988 7084 7045 7085
rect 6988 7065 7017 7084
rect 6960 7064 7017 7065
rect 7038 7064 7045 7084
rect 6960 7057 7045 7064
rect 7064 7081 7102 7090
rect 7064 7061 7073 7081
rect 7093 7061 7102 7081
rect 6960 7056 6996 7057
rect 7064 7053 7102 7061
rect 7168 7085 7312 7091
rect 7168 7065 7176 7085
rect 7196 7083 7284 7085
rect 7196 7066 7232 7083
rect 7256 7066 7284 7083
rect 7196 7065 7284 7066
rect 7304 7065 7312 7085
rect 7168 7057 7312 7065
rect 7168 7056 7204 7057
rect 7276 7056 7312 7057
rect 7378 7090 7415 7091
rect 7378 7089 7416 7090
rect 7378 7081 7442 7089
rect 7378 7061 7387 7081
rect 7407 7067 7442 7081
rect 7462 7067 7465 7087
rect 7407 7062 7465 7067
rect 7407 7061 7442 7062
rect 6644 7024 6681 7053
rect 6645 7022 6681 7024
rect 6857 7022 6894 7053
rect 6160 7001 6196 7002
rect 6008 6971 6017 6991
rect 6037 6971 6045 6991
rect 5896 6962 5952 6964
rect 5896 6961 5933 6962
rect 6008 6961 6045 6971
rect 6104 6991 6252 7001
rect 6645 7000 6894 7022
rect 7065 7021 7102 7053
rect 7378 7049 7442 7061
rect 7482 7023 7509 7201
rect 7341 7021 7509 7023
rect 7065 7010 7509 7021
rect 6352 6998 6448 7000
rect 6104 6971 6113 6991
rect 6133 6971 6223 6991
rect 6243 6971 6252 6991
rect 6104 6962 6252 6971
rect 6310 6991 6448 6998
rect 7065 6995 7511 7010
rect 7341 6994 7511 6995
rect 6310 6971 6319 6991
rect 6339 6971 6448 6991
rect 6310 6962 6448 6971
rect 6104 6961 6141 6962
rect 6160 6910 6196 6962
rect 6215 6961 6252 6962
rect 6311 6961 6348 6962
rect 5631 6908 5672 6909
rect 4457 6858 5089 6865
rect 4457 6856 4519 6858
rect 4035 6846 4203 6847
rect 4457 6846 4479 6856
rect 3750 6821 3787 6822
rect 3700 6812 3787 6821
rect 3700 6792 3758 6812
rect 3778 6792 3787 6812
rect 3700 6782 3787 6792
rect 3846 6812 3883 6822
rect 3846 6792 3854 6812
rect 3874 6792 3883 6812
rect 3700 6781 3731 6782
rect 3846 6721 3883 6792
rect 3633 6697 3883 6721
rect 4035 6820 4479 6846
rect 4035 6818 4203 6820
rect 4035 6640 4062 6818
rect 4102 6780 4166 6792
rect 4442 6788 4479 6820
rect 4650 6819 4899 6841
rect 4650 6788 4687 6819
rect 4863 6817 4899 6819
rect 4863 6788 4900 6817
rect 4102 6779 4137 6780
rect 4079 6774 4137 6779
rect 4079 6754 4082 6774
rect 4102 6760 4137 6774
rect 4157 6760 4166 6780
rect 4102 6752 4166 6760
rect 4128 6751 4166 6752
rect 4129 6750 4166 6751
rect 4232 6784 4268 6785
rect 4340 6784 4376 6785
rect 4232 6776 4376 6784
rect 4232 6756 4240 6776
rect 4260 6756 4289 6776
rect 4232 6755 4289 6756
rect 4311 6756 4348 6776
rect 4368 6756 4376 6776
rect 4311 6755 4376 6756
rect 4232 6750 4376 6755
rect 4442 6780 4480 6788
rect 4548 6784 4584 6785
rect 4442 6760 4451 6780
rect 4471 6760 4480 6780
rect 4442 6751 4480 6760
rect 4499 6777 4584 6784
rect 4499 6757 4506 6777
rect 4527 6776 4584 6777
rect 4527 6757 4556 6776
rect 4499 6756 4556 6757
rect 4576 6756 4584 6776
rect 4442 6750 4479 6751
rect 4499 6750 4584 6756
rect 4650 6780 4688 6788
rect 4761 6784 4797 6785
rect 4650 6760 4659 6780
rect 4679 6760 4688 6780
rect 4650 6751 4688 6760
rect 4712 6776 4797 6784
rect 4712 6756 4769 6776
rect 4789 6756 4797 6776
rect 4650 6750 4687 6751
rect 4712 6750 4797 6756
rect 4863 6780 4901 6788
rect 4863 6760 4872 6780
rect 4892 6760 4901 6780
rect 4863 6751 4901 6760
rect 4863 6750 4900 6751
rect 4286 6729 4322 6750
rect 4712 6729 4743 6750
rect 4119 6725 4219 6729
rect 4119 6721 4181 6725
rect 4119 6695 4126 6721
rect 4152 6699 4181 6721
rect 4207 6699 4219 6725
rect 4152 6695 4219 6699
rect 4119 6692 4219 6695
rect 4287 6692 4322 6729
rect 4384 6726 4743 6729
rect 4384 6721 4606 6726
rect 4384 6697 4397 6721
rect 4421 6702 4606 6721
rect 4630 6702 4743 6726
rect 4421 6697 4743 6702
rect 4384 6693 4743 6697
rect 4810 6721 4959 6729
rect 4810 6701 4821 6721
rect 4841 6701 4959 6721
rect 4810 6694 4959 6701
rect 5050 6709 5089 6858
rect 5393 6744 5432 6893
rect 5523 6901 5672 6908
rect 5523 6881 5641 6901
rect 5661 6881 5672 6901
rect 5523 6873 5672 6881
rect 5739 6905 6098 6909
rect 5739 6900 6061 6905
rect 5739 6876 5852 6900
rect 5876 6881 6061 6900
rect 6085 6881 6098 6905
rect 5876 6876 6098 6881
rect 5739 6873 6098 6876
rect 6160 6873 6195 6910
rect 6263 6907 6363 6910
rect 6263 6903 6330 6907
rect 6263 6877 6275 6903
rect 6301 6881 6330 6903
rect 6356 6881 6363 6907
rect 6301 6877 6363 6881
rect 6263 6873 6363 6877
rect 5739 6852 5770 6873
rect 6160 6852 6196 6873
rect 5582 6851 5619 6852
rect 5581 6842 5619 6851
rect 5581 6822 5590 6842
rect 5610 6822 5619 6842
rect 5581 6814 5619 6822
rect 5685 6846 5770 6852
rect 5795 6851 5832 6852
rect 5685 6826 5693 6846
rect 5713 6826 5770 6846
rect 5685 6818 5770 6826
rect 5794 6842 5832 6851
rect 5794 6822 5803 6842
rect 5823 6822 5832 6842
rect 5685 6817 5721 6818
rect 5794 6814 5832 6822
rect 5898 6846 5983 6852
rect 6003 6851 6040 6852
rect 5898 6826 5906 6846
rect 5926 6845 5983 6846
rect 5926 6826 5955 6845
rect 5898 6825 5955 6826
rect 5976 6825 5983 6845
rect 5898 6818 5983 6825
rect 6002 6842 6040 6851
rect 6002 6822 6011 6842
rect 6031 6822 6040 6842
rect 5898 6817 5934 6818
rect 6002 6814 6040 6822
rect 6106 6847 6250 6852
rect 6106 6846 6171 6847
rect 6106 6826 6114 6846
rect 6134 6826 6171 6846
rect 6193 6846 6250 6847
rect 6193 6826 6222 6846
rect 6242 6826 6250 6846
rect 6106 6818 6250 6826
rect 6106 6817 6142 6818
rect 6214 6817 6250 6818
rect 6316 6851 6353 6852
rect 6316 6850 6354 6851
rect 6316 6842 6380 6850
rect 6316 6822 6325 6842
rect 6345 6828 6380 6842
rect 6400 6828 6403 6848
rect 6345 6823 6403 6828
rect 6345 6822 6380 6823
rect 5582 6785 5619 6814
rect 5583 6783 5619 6785
rect 5795 6783 5832 6814
rect 5583 6761 5832 6783
rect 6003 6782 6040 6814
rect 6316 6810 6380 6822
rect 6420 6784 6447 6962
rect 6279 6782 6447 6784
rect 6003 6756 6447 6782
rect 6599 6881 6849 6905
rect 6599 6810 6636 6881
rect 6751 6820 6782 6821
rect 6599 6790 6608 6810
rect 6628 6790 6636 6810
rect 6599 6780 6636 6790
rect 6695 6810 6782 6820
rect 6695 6790 6704 6810
rect 6724 6790 6782 6810
rect 6695 6781 6782 6790
rect 6695 6780 6732 6781
rect 6003 6746 6025 6756
rect 6279 6755 6447 6756
rect 5963 6744 6025 6746
rect 5393 6737 6025 6744
rect 4810 6693 4851 6694
rect 4134 6640 4171 6641
rect 4230 6640 4267 6641
rect 4286 6640 4322 6692
rect 4341 6640 4378 6641
rect 4034 6631 4172 6640
rect 4034 6611 4143 6631
rect 4163 6611 4172 6631
rect 4034 6604 4172 6611
rect 4230 6631 4378 6640
rect 4230 6611 4239 6631
rect 4259 6611 4349 6631
rect 4369 6611 4378 6631
rect 4034 6602 4130 6604
rect 4230 6601 4378 6611
rect 4437 6631 4474 6641
rect 4549 6640 4586 6641
rect 4530 6638 4586 6640
rect 4437 6611 4445 6631
rect 4465 6611 4474 6631
rect 4286 6600 4322 6601
rect 2749 6538 2757 6557
rect 2780 6538 2786 6557
rect 2749 6527 2786 6538
rect 2815 6560 2983 6561
rect 2815 6534 3259 6560
rect 2815 6532 2983 6534
rect 2752 6467 2785 6527
rect 997 6388 1165 6390
rect 721 6362 1165 6388
rect 722 6345 746 6362
rect 997 6361 1165 6362
rect 1533 6390 1783 6414
rect 120 6327 747 6345
rect 120 6321 158 6327
rect 122 6275 157 6321
rect 1533 6319 1570 6390
rect 1685 6329 1716 6330
rect 1533 6299 1542 6319
rect 1562 6299 1570 6319
rect 1533 6289 1570 6299
rect 1629 6319 1716 6329
rect 1629 6299 1638 6319
rect 1658 6299 1716 6319
rect 1629 6290 1716 6299
rect 1629 6289 1666 6290
rect 120 6266 157 6275
rect 120 6248 130 6266
rect 148 6248 157 6266
rect 120 6238 157 6248
rect 1685 6237 1716 6290
rect 1746 6319 1783 6390
rect 1954 6395 2347 6415
rect 2367 6395 2370 6415
rect 1954 6390 2370 6395
rect 1954 6389 2295 6390
rect 1898 6329 1929 6330
rect 1746 6299 1755 6319
rect 1775 6299 1783 6319
rect 1746 6289 1783 6299
rect 1842 6322 1929 6329
rect 1842 6319 1903 6322
rect 1842 6299 1851 6319
rect 1871 6302 1903 6319
rect 1924 6302 1929 6322
rect 1871 6299 1929 6302
rect 1842 6292 1929 6299
rect 1954 6319 1991 6389
rect 2257 6388 2294 6389
rect 2106 6329 2142 6330
rect 1954 6299 1963 6319
rect 1983 6299 1991 6319
rect 1842 6290 1898 6292
rect 1842 6289 1879 6290
rect 1954 6289 1991 6299
rect 2050 6319 2198 6329
rect 2298 6326 2394 6328
rect 2050 6299 2059 6319
rect 2079 6299 2169 6319
rect 2189 6299 2198 6319
rect 2050 6290 2198 6299
rect 2256 6319 2394 6326
rect 2256 6299 2265 6319
rect 2285 6299 2394 6319
rect 2256 6290 2394 6299
rect 2050 6289 2087 6290
rect 2106 6238 2142 6290
rect 2161 6289 2198 6290
rect 2257 6289 2294 6290
rect 1577 6236 1618 6237
rect 1469 6229 1618 6236
rect 1469 6209 1587 6229
rect 1607 6209 1618 6229
rect 1469 6201 1618 6209
rect 1685 6233 2044 6237
rect 1685 6228 2007 6233
rect 1685 6204 1798 6228
rect 1822 6209 2007 6228
rect 2031 6209 2044 6233
rect 1822 6204 2044 6209
rect 1685 6201 2044 6204
rect 2106 6201 2141 6238
rect 2209 6235 2309 6238
rect 2209 6231 2276 6235
rect 2209 6205 2221 6231
rect 2247 6209 2276 6231
rect 2302 6209 2309 6235
rect 2247 6205 2309 6209
rect 2209 6201 2309 6205
rect 1685 6180 1716 6201
rect 2106 6180 2142 6201
rect 1528 6179 1565 6180
rect 123 6174 160 6176
rect 123 6173 771 6174
rect 122 6167 771 6173
rect 122 6149 132 6167
rect 150 6153 771 6167
rect 150 6149 160 6153
rect 601 6152 771 6153
rect 122 6139 160 6149
rect 122 6061 157 6139
rect 734 6129 771 6152
rect 1527 6170 1565 6179
rect 1527 6150 1536 6170
rect 1556 6150 1565 6170
rect 1527 6142 1565 6150
rect 1631 6174 1716 6180
rect 1741 6179 1778 6180
rect 1631 6154 1639 6174
rect 1659 6154 1716 6174
rect 1631 6146 1716 6154
rect 1740 6170 1778 6179
rect 1740 6150 1749 6170
rect 1769 6150 1778 6170
rect 1631 6145 1667 6146
rect 1740 6142 1778 6150
rect 1844 6174 1929 6180
rect 1949 6179 1986 6180
rect 1844 6154 1852 6174
rect 1872 6173 1929 6174
rect 1872 6154 1901 6173
rect 1844 6153 1901 6154
rect 1922 6153 1929 6173
rect 1844 6146 1929 6153
rect 1948 6170 1986 6179
rect 1948 6150 1957 6170
rect 1977 6150 1986 6170
rect 1844 6145 1880 6146
rect 1948 6142 1986 6150
rect 2052 6178 2196 6180
rect 2052 6174 2110 6178
rect 2052 6154 2060 6174
rect 2080 6154 2110 6174
rect 2052 6152 2110 6154
rect 2135 6174 2196 6178
rect 2135 6154 2168 6174
rect 2188 6154 2196 6174
rect 2135 6152 2196 6154
rect 2052 6146 2196 6152
rect 2052 6145 2088 6146
rect 2160 6145 2196 6146
rect 2262 6179 2299 6180
rect 2262 6178 2300 6179
rect 2262 6170 2326 6178
rect 2262 6150 2271 6170
rect 2291 6156 2326 6170
rect 2346 6156 2349 6176
rect 2291 6151 2349 6156
rect 2291 6150 2326 6151
rect 118 6052 157 6061
rect 118 6034 128 6052
rect 146 6034 157 6052
rect 118 6028 157 6034
rect 313 6104 563 6128
rect 313 6033 350 6104
rect 465 6043 496 6044
rect 118 6024 155 6028
rect 313 6013 322 6033
rect 342 6013 350 6033
rect 313 6003 350 6013
rect 409 6033 496 6043
rect 409 6013 418 6033
rect 438 6013 496 6033
rect 409 6004 496 6013
rect 409 6003 446 6004
rect 121 5953 158 5962
rect 119 5935 130 5953
rect 148 5935 158 5953
rect 465 5951 496 6004
rect 526 6033 563 6104
rect 734 6109 1127 6129
rect 1147 6109 1150 6129
rect 1528 6113 1565 6142
rect 734 6104 1150 6109
rect 1529 6111 1565 6113
rect 1741 6111 1778 6142
rect 734 6103 1075 6104
rect 678 6043 709 6044
rect 526 6013 535 6033
rect 555 6013 563 6033
rect 526 6003 563 6013
rect 622 6036 709 6043
rect 622 6033 683 6036
rect 622 6013 631 6033
rect 651 6016 683 6033
rect 704 6016 709 6036
rect 651 6013 709 6016
rect 622 6006 709 6013
rect 734 6033 771 6103
rect 1037 6102 1074 6103
rect 1529 6089 1778 6111
rect 1949 6110 1986 6142
rect 2262 6138 2326 6150
rect 2366 6112 2393 6290
rect 2225 6110 2393 6112
rect 1949 6084 2393 6110
rect 2225 6083 2393 6084
rect 886 6043 922 6044
rect 734 6013 743 6033
rect 763 6013 771 6033
rect 622 6004 678 6006
rect 622 6003 659 6004
rect 734 6003 771 6013
rect 830 6033 978 6043
rect 1078 6040 1174 6042
rect 830 6013 839 6033
rect 859 6013 949 6033
rect 969 6013 978 6033
rect 830 6004 978 6013
rect 1036 6033 1174 6040
rect 1036 6013 1045 6033
rect 1065 6013 1174 6033
rect 1036 6004 1174 6013
rect 830 6003 867 6004
rect 886 5952 922 6004
rect 941 6003 978 6004
rect 1037 6003 1074 6004
rect 357 5950 398 5951
rect 119 5786 158 5935
rect 249 5943 398 5950
rect 249 5923 367 5943
rect 387 5923 398 5943
rect 249 5915 398 5923
rect 465 5947 824 5951
rect 465 5942 787 5947
rect 465 5918 578 5942
rect 602 5923 787 5942
rect 811 5923 824 5947
rect 602 5918 824 5923
rect 465 5915 824 5918
rect 886 5915 921 5952
rect 989 5949 1089 5952
rect 989 5945 1056 5949
rect 989 5919 1001 5945
rect 1027 5923 1056 5945
rect 1082 5923 1089 5949
rect 1027 5919 1089 5923
rect 989 5915 1089 5919
rect 465 5894 496 5915
rect 886 5894 922 5915
rect 308 5893 345 5894
rect 307 5884 345 5893
rect 307 5864 316 5884
rect 336 5864 345 5884
rect 307 5856 345 5864
rect 411 5888 496 5894
rect 521 5893 558 5894
rect 411 5868 419 5888
rect 439 5868 496 5888
rect 411 5860 496 5868
rect 520 5884 558 5893
rect 520 5864 529 5884
rect 549 5864 558 5884
rect 411 5859 447 5860
rect 520 5856 558 5864
rect 624 5888 709 5894
rect 729 5893 766 5894
rect 624 5868 632 5888
rect 652 5887 709 5888
rect 652 5868 681 5887
rect 624 5867 681 5868
rect 702 5867 709 5887
rect 624 5860 709 5867
rect 728 5884 766 5893
rect 728 5864 737 5884
rect 757 5864 766 5884
rect 624 5859 660 5860
rect 728 5856 766 5864
rect 832 5889 976 5894
rect 832 5888 897 5889
rect 832 5868 840 5888
rect 860 5868 897 5888
rect 919 5888 976 5889
rect 919 5868 948 5888
rect 968 5868 976 5888
rect 832 5860 976 5868
rect 832 5859 868 5860
rect 940 5859 976 5860
rect 1042 5893 1079 5894
rect 1042 5892 1080 5893
rect 1042 5884 1106 5892
rect 1042 5864 1051 5884
rect 1071 5870 1106 5884
rect 1126 5870 1129 5890
rect 1071 5865 1129 5870
rect 1071 5864 1106 5865
rect 308 5827 345 5856
rect 309 5825 345 5827
rect 521 5825 558 5856
rect 309 5803 558 5825
rect 729 5824 766 5856
rect 1042 5852 1106 5864
rect 1146 5826 1173 6004
rect 1005 5824 1173 5826
rect 729 5798 1173 5824
rect 1325 5923 1575 5947
rect 1325 5852 1362 5923
rect 1477 5862 1508 5863
rect 1325 5832 1334 5852
rect 1354 5832 1362 5852
rect 1325 5822 1362 5832
rect 1421 5852 1508 5862
rect 1421 5832 1430 5852
rect 1450 5832 1508 5852
rect 1421 5823 1508 5832
rect 1421 5822 1458 5823
rect 729 5788 751 5798
rect 1005 5797 1173 5798
rect 689 5786 751 5788
rect 119 5779 751 5786
rect 118 5770 751 5779
rect 1477 5770 1508 5823
rect 1538 5852 1575 5923
rect 1746 5928 2139 5948
rect 2159 5928 2162 5948
rect 1746 5923 2162 5928
rect 1746 5922 2087 5923
rect 1690 5862 1721 5863
rect 1538 5832 1547 5852
rect 1567 5832 1575 5852
rect 1538 5822 1575 5832
rect 1634 5855 1721 5862
rect 1634 5852 1695 5855
rect 1634 5832 1643 5852
rect 1663 5835 1695 5852
rect 1716 5835 1721 5855
rect 1663 5832 1721 5835
rect 1634 5825 1721 5832
rect 1746 5852 1783 5922
rect 2049 5921 2086 5922
rect 1898 5862 1934 5863
rect 1746 5832 1755 5852
rect 1775 5832 1783 5852
rect 1634 5823 1690 5825
rect 1634 5822 1671 5823
rect 1746 5822 1783 5832
rect 1842 5852 1990 5862
rect 2090 5859 2186 5861
rect 1842 5832 1851 5852
rect 1871 5832 1961 5852
rect 1981 5832 1990 5852
rect 1842 5823 1990 5832
rect 2048 5852 2186 5859
rect 2048 5832 2057 5852
rect 2077 5832 2186 5852
rect 2048 5823 2186 5832
rect 1842 5822 1879 5823
rect 1898 5771 1934 5823
rect 1953 5822 1990 5823
rect 2049 5822 2086 5823
rect 118 5752 128 5770
rect 146 5769 751 5770
rect 1369 5769 1410 5770
rect 146 5764 167 5769
rect 146 5752 158 5764
rect 1261 5762 1410 5769
rect 118 5744 158 5752
rect 201 5751 227 5752
rect 118 5742 155 5744
rect 201 5733 755 5751
rect 1261 5742 1379 5762
rect 1399 5742 1410 5762
rect 1261 5734 1410 5742
rect 1477 5766 1836 5770
rect 1477 5761 1799 5766
rect 1477 5737 1590 5761
rect 1614 5742 1799 5761
rect 1823 5742 1836 5766
rect 1614 5737 1836 5742
rect 1477 5734 1836 5737
rect 1898 5734 1933 5771
rect 2001 5768 2101 5771
rect 2001 5764 2068 5768
rect 2001 5738 2013 5764
rect 2039 5742 2068 5764
rect 2094 5742 2101 5768
rect 2039 5738 2101 5742
rect 2001 5734 2101 5738
rect 121 5674 158 5680
rect 201 5674 227 5733
rect 734 5714 755 5733
rect 121 5671 227 5674
rect 121 5653 130 5671
rect 148 5657 227 5671
rect 312 5689 562 5713
rect 148 5655 224 5657
rect 148 5653 158 5655
rect 121 5643 158 5653
rect 126 5578 157 5643
rect 312 5618 349 5689
rect 464 5628 495 5629
rect 312 5598 321 5618
rect 341 5598 349 5618
rect 312 5588 349 5598
rect 408 5618 495 5628
rect 408 5598 417 5618
rect 437 5598 495 5618
rect 408 5589 495 5598
rect 408 5588 445 5589
rect 125 5569 162 5578
rect 125 5551 135 5569
rect 153 5551 162 5569
rect 125 5541 162 5551
rect 464 5536 495 5589
rect 525 5618 562 5689
rect 733 5694 1126 5714
rect 1146 5694 1149 5714
rect 1477 5713 1508 5734
rect 1898 5713 1934 5734
rect 1320 5712 1357 5713
rect 733 5689 1149 5694
rect 1319 5703 1357 5712
rect 733 5688 1074 5689
rect 677 5628 708 5629
rect 525 5598 534 5618
rect 554 5598 562 5618
rect 525 5588 562 5598
rect 621 5621 708 5628
rect 621 5618 682 5621
rect 621 5598 630 5618
rect 650 5601 682 5618
rect 703 5601 708 5621
rect 650 5598 708 5601
rect 621 5591 708 5598
rect 733 5618 770 5688
rect 1036 5687 1073 5688
rect 1319 5683 1328 5703
rect 1348 5683 1357 5703
rect 1319 5675 1357 5683
rect 1423 5707 1508 5713
rect 1533 5712 1570 5713
rect 1423 5687 1431 5707
rect 1451 5687 1508 5707
rect 1423 5679 1508 5687
rect 1532 5703 1570 5712
rect 1532 5683 1541 5703
rect 1561 5683 1570 5703
rect 1423 5678 1459 5679
rect 1532 5675 1570 5683
rect 1636 5707 1721 5713
rect 1741 5712 1778 5713
rect 1636 5687 1644 5707
rect 1664 5706 1721 5707
rect 1664 5687 1693 5706
rect 1636 5686 1693 5687
rect 1714 5686 1721 5706
rect 1636 5679 1721 5686
rect 1740 5703 1778 5712
rect 1740 5683 1749 5703
rect 1769 5683 1778 5703
rect 1636 5678 1672 5679
rect 1740 5675 1778 5683
rect 1844 5707 1988 5713
rect 1844 5687 1852 5707
rect 1872 5687 1904 5707
rect 1928 5687 1960 5707
rect 1980 5687 1988 5707
rect 1844 5679 1988 5687
rect 1844 5678 1880 5679
rect 1952 5678 1988 5679
rect 2054 5712 2091 5713
rect 2054 5711 2092 5712
rect 2054 5703 2118 5711
rect 2054 5683 2063 5703
rect 2083 5689 2118 5703
rect 2138 5689 2141 5709
rect 2083 5684 2141 5689
rect 2083 5683 2118 5684
rect 1320 5646 1357 5675
rect 1321 5644 1357 5646
rect 1533 5644 1570 5675
rect 885 5628 921 5629
rect 733 5598 742 5618
rect 762 5598 770 5618
rect 621 5589 677 5591
rect 621 5588 658 5589
rect 733 5588 770 5598
rect 829 5618 977 5628
rect 1077 5625 1173 5627
rect 829 5598 838 5618
rect 858 5598 948 5618
rect 968 5598 977 5618
rect 829 5589 977 5598
rect 1035 5618 1173 5625
rect 1321 5622 1570 5644
rect 1741 5643 1778 5675
rect 2054 5671 2118 5683
rect 2158 5645 2185 5823
rect 2017 5643 2185 5645
rect 1741 5639 2185 5643
rect 1035 5598 1044 5618
rect 1064 5598 1173 5618
rect 1741 5620 1790 5639
rect 1810 5620 2185 5639
rect 1741 5617 2185 5620
rect 2017 5616 2185 5617
rect 1035 5589 1173 5598
rect 829 5588 866 5589
rect 885 5537 921 5589
rect 940 5588 977 5589
rect 1036 5588 1073 5589
rect 356 5535 397 5536
rect 248 5528 397 5535
rect 248 5508 366 5528
rect 386 5508 397 5528
rect 248 5500 397 5508
rect 464 5532 823 5536
rect 464 5527 786 5532
rect 464 5503 577 5527
rect 601 5508 786 5527
rect 810 5508 823 5532
rect 601 5503 823 5508
rect 464 5500 823 5503
rect 885 5500 920 5537
rect 988 5534 1088 5537
rect 988 5530 1055 5534
rect 988 5504 1000 5530
rect 1026 5508 1055 5530
rect 1081 5508 1088 5534
rect 1026 5504 1088 5508
rect 988 5500 1088 5504
rect 464 5479 495 5500
rect 885 5479 921 5500
rect 128 5470 165 5479
rect 307 5478 344 5479
rect 128 5452 137 5470
rect 155 5452 165 5470
rect 128 5442 165 5452
rect 129 5407 165 5442
rect 306 5469 344 5478
rect 306 5449 315 5469
rect 335 5449 344 5469
rect 306 5441 344 5449
rect 410 5473 495 5479
rect 520 5478 557 5479
rect 410 5453 418 5473
rect 438 5453 495 5473
rect 410 5445 495 5453
rect 519 5469 557 5478
rect 519 5449 528 5469
rect 548 5449 557 5469
rect 410 5444 446 5445
rect 519 5441 557 5449
rect 623 5473 708 5479
rect 728 5478 765 5479
rect 623 5453 631 5473
rect 651 5472 708 5473
rect 651 5453 680 5472
rect 623 5452 680 5453
rect 701 5452 708 5472
rect 623 5445 708 5452
rect 727 5469 765 5478
rect 727 5449 736 5469
rect 756 5449 765 5469
rect 623 5444 659 5445
rect 727 5441 765 5449
rect 831 5473 975 5479
rect 831 5453 839 5473
rect 859 5472 947 5473
rect 859 5453 887 5472
rect 831 5451 887 5453
rect 909 5453 947 5472
rect 967 5453 975 5473
rect 909 5451 975 5453
rect 831 5445 975 5451
rect 831 5444 867 5445
rect 939 5444 975 5445
rect 1041 5478 1078 5479
rect 1041 5477 1079 5478
rect 1041 5469 1105 5477
rect 1041 5449 1050 5469
rect 1070 5455 1105 5469
rect 1125 5455 1128 5475
rect 1070 5450 1128 5455
rect 1070 5449 1105 5450
rect 307 5412 344 5441
rect 127 5366 165 5407
rect 308 5410 344 5412
rect 520 5410 557 5441
rect 308 5388 557 5410
rect 728 5409 765 5441
rect 1041 5437 1105 5449
rect 1145 5411 1172 5589
rect 1004 5409 1172 5411
rect 728 5383 1172 5409
rect 729 5366 753 5383
rect 1004 5382 1172 5383
rect 127 5348 754 5366
rect 1380 5362 1630 5386
rect 127 5342 165 5348
rect 127 5318 164 5342
rect 127 5294 162 5318
rect 125 5285 162 5294
rect 125 5267 135 5285
rect 153 5267 162 5285
rect 125 5257 162 5267
rect 1380 5291 1417 5362
rect 1532 5301 1563 5302
rect 1380 5271 1389 5291
rect 1409 5271 1417 5291
rect 1380 5261 1417 5271
rect 1476 5291 1563 5301
rect 1476 5271 1485 5291
rect 1505 5271 1563 5291
rect 1476 5262 1563 5271
rect 1476 5261 1513 5262
rect 1532 5209 1563 5262
rect 1593 5291 1630 5362
rect 1801 5367 2194 5387
rect 2214 5367 2217 5387
rect 1801 5362 2217 5367
rect 1801 5361 2142 5362
rect 1745 5301 1776 5302
rect 1593 5271 1602 5291
rect 1622 5271 1630 5291
rect 1593 5261 1630 5271
rect 1689 5294 1776 5301
rect 1689 5291 1750 5294
rect 1689 5271 1698 5291
rect 1718 5274 1750 5291
rect 1771 5274 1776 5294
rect 1718 5271 1776 5274
rect 1689 5264 1776 5271
rect 1801 5291 1838 5361
rect 2104 5360 2141 5361
rect 1953 5301 1989 5302
rect 1801 5271 1810 5291
rect 1830 5271 1838 5291
rect 1689 5262 1745 5264
rect 1689 5261 1726 5262
rect 1801 5261 1838 5271
rect 1897 5291 2045 5301
rect 2145 5298 2241 5300
rect 1897 5271 1906 5291
rect 1926 5271 2016 5291
rect 2036 5271 2045 5291
rect 1897 5262 2045 5271
rect 2103 5291 2241 5298
rect 2103 5271 2112 5291
rect 2132 5271 2241 5291
rect 2103 5262 2241 5271
rect 1897 5261 1934 5262
rect 1953 5210 1989 5262
rect 2008 5261 2045 5262
rect 2104 5261 2141 5262
rect 1424 5208 1465 5209
rect 1316 5201 1465 5208
rect 128 5193 165 5195
rect 128 5192 776 5193
rect 127 5186 776 5192
rect 127 5168 137 5186
rect 155 5172 776 5186
rect 1316 5181 1434 5201
rect 1454 5181 1465 5201
rect 1316 5173 1465 5181
rect 1532 5205 1891 5209
rect 1532 5200 1854 5205
rect 1532 5176 1645 5200
rect 1669 5181 1854 5200
rect 1878 5181 1891 5205
rect 1669 5176 1891 5181
rect 1532 5173 1891 5176
rect 1953 5173 1988 5210
rect 2056 5207 2156 5210
rect 2056 5203 2123 5207
rect 2056 5177 2068 5203
rect 2094 5181 2123 5203
rect 2149 5181 2156 5207
rect 2094 5177 2156 5181
rect 2056 5173 2156 5177
rect 155 5168 165 5172
rect 606 5171 776 5172
rect 127 5158 165 5168
rect 127 5080 162 5158
rect 739 5148 776 5171
rect 1532 5152 1563 5173
rect 1953 5152 1989 5173
rect 1375 5151 1412 5152
rect 123 5071 162 5080
rect 123 5053 133 5071
rect 151 5053 162 5071
rect 123 5047 162 5053
rect 318 5123 568 5147
rect 318 5052 355 5123
rect 470 5062 501 5063
rect 123 5043 160 5047
rect 318 5032 327 5052
rect 347 5032 355 5052
rect 318 5022 355 5032
rect 414 5052 501 5062
rect 414 5032 423 5052
rect 443 5032 501 5052
rect 414 5023 501 5032
rect 414 5022 451 5023
rect 126 4972 163 4981
rect 124 4954 135 4972
rect 153 4954 163 4972
rect 470 4970 501 5023
rect 531 5052 568 5123
rect 739 5128 1132 5148
rect 1152 5128 1155 5148
rect 739 5123 1155 5128
rect 1374 5142 1412 5151
rect 739 5122 1080 5123
rect 1374 5122 1383 5142
rect 1403 5122 1412 5142
rect 683 5062 714 5063
rect 531 5032 540 5052
rect 560 5032 568 5052
rect 531 5022 568 5032
rect 627 5055 714 5062
rect 627 5052 688 5055
rect 627 5032 636 5052
rect 656 5035 688 5052
rect 709 5035 714 5055
rect 656 5032 714 5035
rect 627 5025 714 5032
rect 739 5052 776 5122
rect 1042 5121 1079 5122
rect 1374 5114 1412 5122
rect 1478 5146 1563 5152
rect 1588 5151 1625 5152
rect 1478 5126 1486 5146
rect 1506 5126 1563 5146
rect 1478 5118 1563 5126
rect 1587 5142 1625 5151
rect 1587 5122 1596 5142
rect 1616 5122 1625 5142
rect 1478 5117 1514 5118
rect 1587 5114 1625 5122
rect 1691 5146 1776 5152
rect 1796 5151 1833 5152
rect 1691 5126 1699 5146
rect 1719 5145 1776 5146
rect 1719 5126 1748 5145
rect 1691 5125 1748 5126
rect 1769 5125 1776 5145
rect 1691 5118 1776 5125
rect 1795 5142 1833 5151
rect 1795 5122 1804 5142
rect 1824 5122 1833 5142
rect 1691 5117 1727 5118
rect 1795 5114 1833 5122
rect 1899 5146 2043 5152
rect 1899 5126 1907 5146
rect 1927 5145 2015 5146
rect 1927 5126 1960 5145
rect 1983 5126 2015 5145
rect 2035 5126 2043 5146
rect 1899 5118 2043 5126
rect 1899 5117 1935 5118
rect 2007 5117 2043 5118
rect 2109 5151 2146 5152
rect 2109 5150 2147 5151
rect 2109 5142 2173 5150
rect 2109 5122 2118 5142
rect 2138 5128 2173 5142
rect 2193 5128 2196 5148
rect 2138 5123 2196 5128
rect 2138 5122 2173 5123
rect 1375 5085 1412 5114
rect 1376 5083 1412 5085
rect 1588 5083 1625 5114
rect 891 5062 927 5063
rect 739 5032 748 5052
rect 768 5032 776 5052
rect 627 5023 683 5025
rect 627 5022 664 5023
rect 739 5022 776 5032
rect 835 5052 983 5062
rect 1376 5061 1625 5083
rect 1796 5082 1833 5114
rect 2109 5110 2173 5122
rect 2213 5084 2240 5262
rect 2072 5082 2240 5084
rect 1796 5071 2240 5082
rect 2303 5082 2333 6083
rect 2303 5077 2335 5082
rect 1083 5059 1179 5061
rect 835 5032 844 5052
rect 864 5032 954 5052
rect 974 5032 983 5052
rect 835 5023 983 5032
rect 1041 5052 1179 5059
rect 1796 5056 2242 5071
rect 2072 5055 2242 5056
rect 1041 5032 1050 5052
rect 1070 5032 1179 5052
rect 1041 5023 1179 5032
rect 835 5022 872 5023
rect 891 4971 927 5023
rect 946 5022 983 5023
rect 1042 5022 1079 5023
rect 362 4969 403 4970
rect 124 4805 163 4954
rect 254 4962 403 4969
rect 254 4942 372 4962
rect 392 4942 403 4962
rect 254 4934 403 4942
rect 470 4966 829 4970
rect 470 4961 792 4966
rect 470 4937 583 4961
rect 607 4942 792 4961
rect 816 4942 829 4966
rect 607 4937 829 4942
rect 470 4934 829 4937
rect 891 4934 926 4971
rect 994 4968 1094 4971
rect 994 4964 1061 4968
rect 994 4938 1006 4964
rect 1032 4942 1061 4964
rect 1087 4942 1094 4968
rect 1032 4938 1094 4942
rect 994 4934 1094 4938
rect 470 4913 501 4934
rect 891 4913 927 4934
rect 313 4912 350 4913
rect 312 4903 350 4912
rect 312 4883 321 4903
rect 341 4883 350 4903
rect 312 4875 350 4883
rect 416 4907 501 4913
rect 526 4912 563 4913
rect 416 4887 424 4907
rect 444 4887 501 4907
rect 416 4879 501 4887
rect 525 4903 563 4912
rect 525 4883 534 4903
rect 554 4883 563 4903
rect 416 4878 452 4879
rect 525 4875 563 4883
rect 629 4907 714 4913
rect 734 4912 771 4913
rect 629 4887 637 4907
rect 657 4906 714 4907
rect 657 4887 686 4906
rect 629 4886 686 4887
rect 707 4886 714 4906
rect 629 4879 714 4886
rect 733 4903 771 4912
rect 733 4883 742 4903
rect 762 4883 771 4903
rect 629 4878 665 4879
rect 733 4875 771 4883
rect 837 4908 981 4913
rect 837 4907 902 4908
rect 837 4887 845 4907
rect 865 4887 902 4907
rect 924 4907 981 4908
rect 924 4887 953 4907
rect 973 4887 981 4907
rect 837 4879 981 4887
rect 837 4878 873 4879
rect 945 4878 981 4879
rect 1047 4912 1084 4913
rect 1047 4911 1085 4912
rect 1047 4903 1111 4911
rect 1047 4883 1056 4903
rect 1076 4889 1111 4903
rect 1131 4889 1134 4909
rect 1076 4884 1134 4889
rect 1076 4883 1111 4884
rect 313 4846 350 4875
rect 314 4844 350 4846
rect 526 4844 563 4875
rect 314 4822 563 4844
rect 734 4843 771 4875
rect 1047 4871 1111 4883
rect 1151 4845 1178 5023
rect 1010 4843 1178 4845
rect 734 4817 1178 4843
rect 1330 4942 1580 4966
rect 1330 4871 1367 4942
rect 1482 4881 1513 4882
rect 1330 4851 1339 4871
rect 1359 4851 1367 4871
rect 1330 4841 1367 4851
rect 1426 4871 1513 4881
rect 1426 4851 1435 4871
rect 1455 4851 1513 4871
rect 1426 4842 1513 4851
rect 1426 4841 1463 4842
rect 734 4807 756 4817
rect 1010 4816 1178 4817
rect 694 4805 756 4807
rect 124 4798 756 4805
rect 123 4789 756 4798
rect 1482 4789 1513 4842
rect 1543 4871 1580 4942
rect 1751 4947 2144 4967
rect 2164 4947 2167 4967
rect 1751 4942 2167 4947
rect 1751 4941 2092 4942
rect 1695 4881 1726 4882
rect 1543 4851 1552 4871
rect 1572 4851 1580 4871
rect 1543 4841 1580 4851
rect 1639 4874 1726 4881
rect 1639 4871 1700 4874
rect 1639 4851 1648 4871
rect 1668 4854 1700 4871
rect 1721 4854 1726 4874
rect 1668 4851 1726 4854
rect 1639 4844 1726 4851
rect 1751 4871 1788 4941
rect 2054 4940 2091 4941
rect 1903 4881 1939 4882
rect 1751 4851 1760 4871
rect 1780 4851 1788 4871
rect 1639 4842 1695 4844
rect 1639 4841 1676 4842
rect 1751 4841 1788 4851
rect 1847 4871 1995 4881
rect 2095 4878 2191 4880
rect 1847 4851 1856 4871
rect 1876 4851 1966 4871
rect 1986 4851 1995 4871
rect 1847 4842 1995 4851
rect 2053 4871 2191 4878
rect 2053 4851 2062 4871
rect 2082 4851 2191 4871
rect 2053 4842 2191 4851
rect 1847 4841 1884 4842
rect 1903 4790 1939 4842
rect 1958 4841 1995 4842
rect 2054 4841 2091 4842
rect 123 4771 133 4789
rect 151 4788 756 4789
rect 1374 4788 1415 4789
rect 151 4783 172 4788
rect 151 4771 163 4783
rect 1266 4781 1415 4788
rect 123 4763 163 4771
rect 206 4770 232 4771
rect 123 4761 160 4763
rect 206 4752 760 4770
rect 1266 4761 1384 4781
rect 1404 4761 1415 4781
rect 1266 4753 1415 4761
rect 1482 4785 1841 4789
rect 1482 4780 1804 4785
rect 1482 4756 1595 4780
rect 1619 4761 1804 4780
rect 1828 4761 1841 4785
rect 1619 4756 1841 4761
rect 1482 4753 1841 4756
rect 1903 4753 1938 4790
rect 2006 4787 2106 4790
rect 2006 4783 2073 4787
rect 2006 4757 2018 4783
rect 2044 4761 2073 4783
rect 2099 4761 2106 4787
rect 2044 4757 2106 4761
rect 2006 4753 2106 4757
rect 126 4693 163 4699
rect 206 4693 232 4752
rect 739 4733 760 4752
rect 126 4690 232 4693
rect 126 4672 135 4690
rect 153 4676 232 4690
rect 317 4708 567 4732
rect 153 4674 229 4676
rect 153 4672 163 4674
rect 126 4662 163 4672
rect 131 4597 162 4662
rect 317 4637 354 4708
rect 469 4647 500 4648
rect 317 4617 326 4637
rect 346 4617 354 4637
rect 317 4607 354 4617
rect 413 4637 500 4647
rect 413 4617 422 4637
rect 442 4617 500 4637
rect 413 4608 500 4617
rect 413 4607 450 4608
rect 130 4588 167 4597
rect 130 4570 140 4588
rect 158 4570 167 4588
rect 130 4560 167 4570
rect 469 4555 500 4608
rect 530 4637 567 4708
rect 738 4713 1131 4733
rect 1151 4713 1154 4733
rect 1482 4732 1513 4753
rect 1903 4732 1939 4753
rect 1325 4731 1362 4732
rect 738 4708 1154 4713
rect 1324 4722 1362 4731
rect 738 4707 1079 4708
rect 682 4647 713 4648
rect 530 4617 539 4637
rect 559 4617 567 4637
rect 530 4607 567 4617
rect 626 4640 713 4647
rect 626 4637 687 4640
rect 626 4617 635 4637
rect 655 4620 687 4637
rect 708 4620 713 4640
rect 655 4617 713 4620
rect 626 4610 713 4617
rect 738 4637 775 4707
rect 1041 4706 1078 4707
rect 1324 4702 1333 4722
rect 1353 4702 1362 4722
rect 1324 4694 1362 4702
rect 1428 4726 1513 4732
rect 1538 4731 1575 4732
rect 1428 4706 1436 4726
rect 1456 4706 1513 4726
rect 1428 4698 1513 4706
rect 1537 4722 1575 4731
rect 1537 4702 1546 4722
rect 1566 4702 1575 4722
rect 1428 4697 1464 4698
rect 1537 4694 1575 4702
rect 1641 4726 1726 4732
rect 1746 4731 1783 4732
rect 1641 4706 1649 4726
rect 1669 4725 1726 4726
rect 1669 4706 1698 4725
rect 1641 4705 1698 4706
rect 1719 4705 1726 4725
rect 1641 4698 1726 4705
rect 1745 4722 1783 4731
rect 1745 4702 1754 4722
rect 1774 4702 1783 4722
rect 1641 4697 1677 4698
rect 1745 4694 1783 4702
rect 1849 4727 1993 4732
rect 1849 4726 1908 4727
rect 1849 4706 1857 4726
rect 1877 4707 1908 4726
rect 1932 4726 1993 4727
rect 1932 4707 1965 4726
rect 1877 4706 1965 4707
rect 1985 4706 1993 4726
rect 1849 4698 1993 4706
rect 1849 4697 1885 4698
rect 1957 4697 1993 4698
rect 2059 4731 2096 4732
rect 2059 4730 2097 4731
rect 2059 4722 2123 4730
rect 2059 4702 2068 4722
rect 2088 4708 2123 4722
rect 2143 4708 2146 4728
rect 2088 4703 2146 4708
rect 2088 4702 2123 4703
rect 1325 4665 1362 4694
rect 1326 4663 1362 4665
rect 1538 4663 1575 4694
rect 890 4647 926 4648
rect 738 4617 747 4637
rect 767 4617 775 4637
rect 626 4608 682 4610
rect 626 4607 663 4608
rect 738 4607 775 4617
rect 834 4637 982 4647
rect 1082 4644 1178 4646
rect 834 4617 843 4637
rect 863 4617 953 4637
rect 973 4617 982 4637
rect 834 4608 982 4617
rect 1040 4637 1178 4644
rect 1326 4641 1575 4663
rect 1746 4662 1783 4694
rect 2059 4690 2123 4702
rect 2163 4664 2190 4842
rect 2022 4662 2190 4664
rect 1746 4658 2190 4662
rect 1040 4617 1049 4637
rect 1069 4617 1178 4637
rect 1746 4639 1795 4658
rect 1815 4639 2190 4658
rect 1746 4636 2190 4639
rect 2022 4635 2190 4636
rect 2211 4661 2242 5055
rect 2303 5059 2308 5077
rect 2328 5059 2335 5077
rect 2303 5054 2335 5059
rect 2306 5052 2335 5054
rect 2211 4635 2216 4661
rect 2235 4635 2242 4661
rect 2749 4636 2787 6467
rect 2815 6354 2842 6532
rect 2882 6494 2946 6506
rect 3222 6502 3259 6534
rect 3430 6533 3679 6555
rect 4134 6541 4171 6542
rect 4437 6541 4474 6611
rect 4499 6631 4586 6638
rect 4499 6628 4557 6631
rect 4499 6608 4504 6628
rect 4525 6611 4557 6628
rect 4577 6611 4586 6631
rect 4525 6608 4586 6611
rect 4499 6601 4586 6608
rect 4645 6631 4682 6641
rect 4645 6611 4653 6631
rect 4673 6611 4682 6631
rect 4499 6600 4530 6601
rect 4133 6540 4474 6541
rect 3430 6502 3467 6533
rect 3643 6531 3679 6533
rect 4058 6535 4474 6540
rect 3643 6502 3680 6531
rect 4058 6515 4061 6535
rect 4081 6515 4474 6535
rect 4645 6540 4682 6611
rect 4712 6640 4743 6693
rect 5050 6691 5060 6709
rect 5078 6691 5089 6709
rect 5392 6728 6025 6737
rect 6751 6728 6782 6781
rect 6812 6810 6849 6881
rect 7020 6886 7413 6906
rect 7433 6886 7436 6906
rect 7020 6881 7436 6886
rect 7020 6880 7361 6881
rect 6964 6820 6995 6821
rect 6812 6790 6821 6810
rect 6841 6790 6849 6810
rect 6812 6780 6849 6790
rect 6908 6813 6995 6820
rect 6908 6810 6969 6813
rect 6908 6790 6917 6810
rect 6937 6793 6969 6810
rect 6990 6793 6995 6813
rect 6937 6790 6995 6793
rect 6908 6783 6995 6790
rect 7020 6810 7057 6880
rect 7323 6879 7360 6880
rect 7172 6820 7208 6821
rect 7020 6790 7029 6810
rect 7049 6790 7057 6810
rect 6908 6781 6964 6783
rect 6908 6780 6945 6781
rect 7020 6780 7057 6790
rect 7116 6810 7264 6820
rect 7364 6817 7460 6819
rect 7116 6790 7125 6810
rect 7145 6790 7235 6810
rect 7255 6790 7264 6810
rect 7116 6781 7264 6790
rect 7322 6810 7460 6817
rect 7322 6790 7331 6810
rect 7351 6790 7460 6810
rect 7322 6781 7460 6790
rect 7116 6780 7153 6781
rect 7172 6729 7208 6781
rect 7227 6780 7264 6781
rect 7323 6780 7360 6781
rect 5392 6710 5402 6728
rect 5420 6727 6025 6728
rect 6643 6727 6684 6728
rect 5420 6722 5441 6727
rect 5420 6710 5432 6722
rect 6535 6720 6684 6727
rect 5392 6702 5432 6710
rect 5475 6709 5501 6710
rect 5392 6700 5429 6702
rect 5475 6691 6029 6709
rect 6535 6700 6653 6720
rect 6673 6700 6684 6720
rect 6535 6692 6684 6700
rect 6751 6724 7110 6728
rect 6751 6719 7073 6724
rect 6751 6695 6864 6719
rect 6888 6700 7073 6719
rect 7097 6700 7110 6724
rect 6888 6695 7110 6700
rect 6751 6692 7110 6695
rect 7172 6692 7207 6729
rect 7275 6726 7375 6729
rect 7275 6722 7342 6726
rect 7275 6696 7287 6722
rect 7313 6700 7342 6722
rect 7368 6700 7375 6726
rect 7313 6696 7375 6700
rect 7275 6692 7375 6696
rect 5050 6682 5087 6691
rect 4762 6640 4799 6641
rect 4712 6631 4799 6640
rect 4712 6611 4770 6631
rect 4790 6611 4799 6631
rect 4712 6601 4799 6611
rect 4858 6631 4895 6641
rect 4858 6611 4866 6631
rect 4886 6611 4895 6631
rect 5395 6632 5432 6638
rect 5475 6632 5501 6691
rect 6008 6672 6029 6691
rect 5395 6629 5501 6632
rect 5053 6616 5090 6620
rect 4712 6600 4743 6601
rect 4858 6540 4895 6611
rect 4645 6516 4895 6540
rect 5051 6610 5090 6616
rect 5051 6592 5062 6610
rect 5080 6592 5090 6610
rect 5395 6611 5404 6629
rect 5422 6615 5501 6629
rect 5586 6647 5836 6671
rect 5422 6613 5498 6615
rect 5422 6611 5432 6613
rect 5395 6601 5432 6611
rect 5051 6583 5090 6592
rect 2882 6493 2917 6494
rect 2859 6488 2917 6493
rect 2859 6468 2862 6488
rect 2882 6474 2917 6488
rect 2937 6474 2946 6494
rect 2882 6466 2946 6474
rect 2908 6465 2946 6466
rect 2909 6464 2946 6465
rect 3012 6498 3048 6499
rect 3120 6498 3156 6499
rect 3012 6490 3156 6498
rect 3012 6470 3020 6490
rect 3040 6489 3128 6490
rect 3040 6470 3069 6489
rect 3092 6470 3128 6489
rect 3148 6470 3156 6490
rect 3012 6464 3156 6470
rect 3222 6494 3260 6502
rect 3328 6498 3364 6499
rect 3222 6474 3231 6494
rect 3251 6474 3260 6494
rect 3222 6465 3260 6474
rect 3279 6491 3364 6498
rect 3279 6471 3286 6491
rect 3307 6490 3364 6491
rect 3307 6471 3336 6490
rect 3279 6470 3336 6471
rect 3356 6470 3364 6490
rect 3222 6464 3259 6465
rect 3279 6464 3364 6470
rect 3430 6494 3468 6502
rect 3541 6498 3577 6499
rect 3430 6474 3439 6494
rect 3459 6474 3468 6494
rect 3430 6465 3468 6474
rect 3492 6490 3577 6498
rect 3492 6470 3549 6490
rect 3569 6470 3577 6490
rect 3430 6464 3467 6465
rect 3492 6464 3577 6470
rect 3643 6494 3681 6502
rect 3643 6474 3652 6494
rect 3672 6474 3681 6494
rect 3643 6465 3681 6474
rect 4437 6492 4474 6515
rect 5051 6505 5086 6583
rect 5400 6536 5431 6601
rect 5586 6576 5623 6647
rect 5738 6586 5769 6587
rect 5586 6556 5595 6576
rect 5615 6556 5623 6576
rect 5586 6546 5623 6556
rect 5682 6576 5769 6586
rect 5682 6556 5691 6576
rect 5711 6556 5769 6576
rect 5682 6547 5769 6556
rect 5682 6546 5719 6547
rect 5048 6495 5086 6505
rect 5399 6527 5436 6536
rect 5399 6509 5409 6527
rect 5427 6509 5436 6527
rect 5399 6499 5436 6509
rect 4437 6491 4607 6492
rect 5048 6491 5058 6495
rect 4437 6477 5058 6491
rect 5076 6477 5086 6495
rect 5738 6494 5769 6547
rect 5799 6576 5836 6647
rect 6007 6652 6400 6672
rect 6420 6652 6423 6672
rect 6751 6671 6782 6692
rect 7172 6671 7208 6692
rect 6594 6670 6631 6671
rect 6007 6647 6423 6652
rect 6593 6661 6631 6670
rect 6007 6646 6348 6647
rect 5951 6586 5982 6587
rect 5799 6556 5808 6576
rect 5828 6556 5836 6576
rect 5799 6546 5836 6556
rect 5895 6579 5982 6586
rect 5895 6576 5956 6579
rect 5895 6556 5904 6576
rect 5924 6559 5956 6576
rect 5977 6559 5982 6579
rect 5924 6556 5982 6559
rect 5895 6549 5982 6556
rect 6007 6576 6044 6646
rect 6310 6645 6347 6646
rect 6593 6641 6602 6661
rect 6622 6641 6631 6661
rect 6593 6633 6631 6641
rect 6697 6665 6782 6671
rect 6807 6670 6844 6671
rect 6697 6645 6705 6665
rect 6725 6645 6782 6665
rect 6697 6637 6782 6645
rect 6806 6661 6844 6670
rect 6806 6641 6815 6661
rect 6835 6641 6844 6661
rect 6697 6636 6733 6637
rect 6806 6633 6844 6641
rect 6910 6665 6995 6671
rect 7015 6670 7052 6671
rect 6910 6645 6918 6665
rect 6938 6664 6995 6665
rect 6938 6645 6967 6664
rect 6910 6644 6967 6645
rect 6988 6644 6995 6664
rect 6910 6637 6995 6644
rect 7014 6661 7052 6670
rect 7014 6641 7023 6661
rect 7043 6641 7052 6661
rect 6910 6636 6946 6637
rect 7014 6633 7052 6641
rect 7118 6666 7262 6671
rect 7118 6665 7177 6666
rect 7118 6645 7126 6665
rect 7146 6646 7177 6665
rect 7201 6665 7262 6666
rect 7201 6646 7234 6665
rect 7146 6645 7234 6646
rect 7254 6645 7262 6665
rect 7118 6637 7262 6645
rect 7118 6636 7154 6637
rect 7226 6636 7262 6637
rect 7328 6670 7365 6671
rect 7328 6669 7366 6670
rect 7328 6661 7392 6669
rect 7328 6641 7337 6661
rect 7357 6647 7392 6661
rect 7412 6647 7415 6667
rect 7357 6642 7415 6647
rect 7357 6641 7392 6642
rect 6594 6604 6631 6633
rect 6595 6602 6631 6604
rect 6807 6602 6844 6633
rect 6159 6586 6195 6587
rect 6007 6556 6016 6576
rect 6036 6556 6044 6576
rect 5895 6547 5951 6549
rect 5895 6546 5932 6547
rect 6007 6546 6044 6556
rect 6103 6576 6251 6586
rect 6351 6583 6447 6585
rect 6103 6556 6112 6576
rect 6132 6556 6222 6576
rect 6242 6556 6251 6576
rect 6103 6547 6251 6556
rect 6309 6576 6447 6583
rect 6595 6580 6844 6602
rect 7015 6601 7052 6633
rect 7328 6629 7392 6641
rect 7432 6603 7459 6781
rect 7291 6601 7459 6603
rect 7015 6597 7459 6601
rect 6309 6556 6318 6576
rect 6338 6556 6447 6576
rect 7015 6578 7064 6597
rect 7084 6578 7459 6597
rect 7015 6575 7459 6578
rect 7291 6574 7459 6575
rect 7480 6600 7511 6994
rect 7480 6574 7485 6600
rect 7504 6574 7511 6600
rect 7480 6571 7511 6574
rect 6309 6547 6447 6556
rect 6103 6546 6140 6547
rect 6159 6495 6195 6547
rect 6214 6546 6251 6547
rect 6310 6546 6347 6547
rect 5630 6493 5671 6494
rect 4437 6471 5086 6477
rect 5522 6486 5671 6493
rect 4437 6470 5085 6471
rect 5048 6468 5085 6470
rect 5522 6466 5640 6486
rect 5660 6466 5671 6486
rect 3643 6464 3680 6465
rect 3066 6443 3102 6464
rect 3492 6443 3523 6464
rect 5522 6458 5671 6466
rect 5738 6490 6097 6494
rect 5738 6485 6060 6490
rect 5738 6461 5851 6485
rect 5875 6466 6060 6485
rect 6084 6466 6097 6490
rect 5875 6461 6097 6466
rect 5738 6458 6097 6461
rect 6159 6458 6194 6495
rect 6262 6492 6362 6495
rect 6262 6488 6329 6492
rect 6262 6462 6274 6488
rect 6300 6466 6329 6488
rect 6355 6466 6362 6492
rect 6300 6462 6362 6466
rect 6262 6458 6362 6462
rect 2899 6439 2999 6443
rect 2899 6435 2961 6439
rect 2899 6409 2906 6435
rect 2932 6413 2961 6435
rect 2987 6413 2999 6439
rect 2932 6409 2999 6413
rect 2899 6406 2999 6409
rect 3067 6406 3102 6443
rect 3164 6440 3523 6443
rect 3164 6435 3386 6440
rect 3164 6411 3177 6435
rect 3201 6416 3386 6435
rect 3410 6416 3523 6440
rect 3201 6411 3523 6416
rect 3164 6407 3523 6411
rect 3590 6435 3739 6443
rect 5738 6437 5769 6458
rect 6159 6437 6195 6458
rect 3590 6415 3601 6435
rect 3621 6415 3739 6435
rect 3590 6408 3739 6415
rect 5402 6428 5439 6437
rect 5581 6436 5618 6437
rect 5402 6410 5411 6428
rect 5429 6410 5439 6428
rect 3590 6407 3631 6408
rect 2914 6354 2951 6355
rect 3010 6354 3047 6355
rect 3066 6354 3102 6406
rect 3121 6354 3158 6355
rect 2814 6345 2952 6354
rect 2814 6325 2923 6345
rect 2943 6325 2952 6345
rect 2814 6318 2952 6325
rect 3010 6345 3158 6354
rect 3010 6325 3019 6345
rect 3039 6325 3129 6345
rect 3149 6325 3158 6345
rect 2814 6316 2910 6318
rect 3010 6315 3158 6325
rect 3217 6345 3254 6355
rect 3329 6354 3366 6355
rect 3310 6352 3366 6354
rect 3217 6325 3225 6345
rect 3245 6325 3254 6345
rect 3066 6314 3102 6315
rect 2914 6255 2951 6256
rect 3217 6255 3254 6325
rect 3279 6345 3366 6352
rect 3279 6342 3337 6345
rect 3279 6322 3284 6342
rect 3305 6325 3337 6342
rect 3357 6325 3366 6345
rect 3305 6322 3366 6325
rect 3279 6315 3366 6322
rect 3425 6345 3462 6355
rect 3425 6325 3433 6345
rect 3453 6325 3462 6345
rect 3279 6314 3310 6315
rect 2913 6254 3254 6255
rect 2838 6249 3254 6254
rect 2838 6229 2841 6249
rect 2861 6229 3254 6249
rect 3425 6254 3462 6325
rect 3492 6354 3523 6407
rect 5051 6396 5088 6406
rect 5402 6400 5439 6410
rect 5051 6378 5060 6396
rect 5078 6378 5088 6396
rect 5051 6369 5088 6378
rect 3542 6354 3579 6355
rect 3492 6345 3579 6354
rect 3492 6325 3550 6345
rect 3570 6325 3579 6345
rect 3492 6315 3579 6325
rect 3638 6345 3675 6355
rect 3638 6325 3646 6345
rect 3666 6325 3675 6345
rect 3492 6314 3523 6315
rect 3638 6254 3675 6325
rect 5051 6323 5086 6369
rect 5403 6365 5439 6400
rect 5580 6427 5618 6436
rect 5580 6407 5589 6427
rect 5609 6407 5618 6427
rect 5580 6399 5618 6407
rect 5684 6431 5769 6437
rect 5794 6436 5831 6437
rect 5684 6411 5692 6431
rect 5712 6411 5769 6431
rect 5684 6403 5769 6411
rect 5793 6427 5831 6436
rect 5793 6407 5802 6427
rect 5822 6407 5831 6427
rect 5684 6402 5720 6403
rect 5793 6399 5831 6407
rect 5897 6431 5982 6437
rect 6002 6436 6039 6437
rect 5897 6411 5905 6431
rect 5925 6430 5982 6431
rect 5925 6411 5954 6430
rect 5897 6410 5954 6411
rect 5975 6410 5982 6430
rect 5897 6403 5982 6410
rect 6001 6427 6039 6436
rect 6001 6407 6010 6427
rect 6030 6407 6039 6427
rect 5897 6402 5933 6403
rect 6001 6399 6039 6407
rect 6105 6431 6249 6437
rect 6105 6411 6113 6431
rect 6133 6430 6221 6431
rect 6133 6411 6161 6430
rect 6105 6409 6161 6411
rect 6183 6411 6221 6430
rect 6241 6411 6249 6431
rect 6183 6409 6249 6411
rect 6105 6403 6249 6409
rect 6105 6402 6141 6403
rect 6213 6402 6249 6403
rect 6315 6436 6352 6437
rect 6315 6435 6353 6436
rect 6315 6427 6379 6435
rect 6315 6407 6324 6427
rect 6344 6413 6379 6427
rect 6399 6413 6402 6433
rect 6344 6408 6402 6413
rect 6344 6407 6379 6408
rect 5581 6370 5618 6399
rect 5401 6324 5439 6365
rect 5582 6368 5618 6370
rect 5794 6368 5831 6399
rect 5582 6346 5831 6368
rect 6002 6367 6039 6399
rect 6315 6395 6379 6407
rect 6419 6369 6446 6547
rect 8030 6536 8067 6547
rect 8156 6540 8186 7541
rect 8249 7541 8693 7552
rect 8249 7539 8417 7541
rect 8249 7361 8276 7539
rect 8316 7501 8380 7513
rect 8656 7509 8693 7541
rect 8864 7540 9113 7562
rect 9506 7561 9654 7571
rect 9713 7591 9750 7601
rect 9825 7600 9862 7601
rect 9806 7598 9862 7600
rect 9713 7571 9721 7591
rect 9741 7571 9750 7591
rect 9562 7560 9598 7561
rect 8864 7509 8901 7540
rect 9077 7538 9113 7540
rect 9077 7509 9114 7538
rect 8316 7500 8351 7501
rect 8293 7495 8351 7500
rect 8293 7475 8296 7495
rect 8316 7481 8351 7495
rect 8371 7481 8380 7501
rect 8316 7473 8380 7481
rect 8342 7472 8380 7473
rect 8343 7471 8380 7472
rect 8446 7505 8482 7506
rect 8554 7505 8590 7506
rect 8446 7497 8590 7505
rect 8446 7477 8454 7497
rect 8474 7478 8506 7497
rect 8529 7478 8562 7497
rect 8474 7477 8562 7478
rect 8582 7477 8590 7497
rect 8446 7471 8590 7477
rect 8656 7501 8694 7509
rect 8762 7505 8798 7506
rect 8656 7481 8665 7501
rect 8685 7481 8694 7501
rect 8656 7472 8694 7481
rect 8713 7498 8798 7505
rect 8713 7478 8720 7498
rect 8741 7497 8798 7498
rect 8741 7478 8770 7497
rect 8713 7477 8770 7478
rect 8790 7477 8798 7497
rect 8656 7471 8693 7472
rect 8713 7471 8798 7477
rect 8864 7501 8902 7509
rect 8975 7505 9011 7506
rect 8864 7481 8873 7501
rect 8893 7481 8902 7501
rect 8864 7472 8902 7481
rect 8926 7497 9011 7505
rect 8926 7477 8983 7497
rect 9003 7477 9011 7497
rect 8864 7471 8901 7472
rect 8926 7471 9011 7477
rect 9077 7501 9115 7509
rect 9410 7501 9447 7502
rect 9713 7501 9750 7571
rect 9775 7591 9862 7598
rect 9775 7588 9833 7591
rect 9775 7568 9780 7588
rect 9801 7571 9833 7588
rect 9853 7571 9862 7591
rect 9801 7568 9862 7571
rect 9775 7561 9862 7568
rect 9921 7591 9958 7601
rect 9921 7571 9929 7591
rect 9949 7571 9958 7591
rect 9775 7560 9806 7561
rect 9077 7481 9086 7501
rect 9106 7481 9115 7501
rect 9409 7500 9750 7501
rect 9077 7472 9115 7481
rect 9334 7495 9750 7500
rect 9334 7475 9337 7495
rect 9357 7475 9750 7495
rect 9921 7500 9958 7571
rect 9988 7600 10019 7653
rect 10326 7651 10336 7669
rect 10354 7651 10365 7669
rect 10326 7642 10363 7651
rect 10038 7600 10075 7601
rect 9988 7591 10075 7600
rect 9988 7571 10046 7591
rect 10066 7571 10075 7591
rect 9988 7561 10075 7571
rect 10134 7591 10171 7601
rect 10134 7571 10142 7591
rect 10162 7571 10171 7591
rect 10329 7576 10366 7580
rect 9988 7560 10019 7561
rect 10134 7500 10171 7571
rect 9921 7476 10171 7500
rect 10327 7570 10366 7576
rect 10327 7552 10338 7570
rect 10356 7552 10366 7570
rect 10327 7543 10366 7552
rect 9077 7471 9114 7472
rect 8500 7450 8536 7471
rect 8926 7450 8957 7471
rect 9713 7452 9750 7475
rect 10327 7465 10362 7543
rect 10324 7455 10362 7465
rect 9713 7451 9883 7452
rect 10324 7451 10334 7455
rect 8333 7446 8433 7450
rect 8333 7442 8395 7446
rect 8333 7416 8340 7442
rect 8366 7420 8395 7442
rect 8421 7420 8433 7446
rect 8366 7416 8433 7420
rect 8333 7413 8433 7416
rect 8501 7413 8536 7450
rect 8598 7447 8957 7450
rect 8598 7442 8820 7447
rect 8598 7418 8611 7442
rect 8635 7423 8820 7442
rect 8844 7423 8957 7447
rect 8635 7418 8957 7423
rect 8598 7414 8957 7418
rect 9024 7442 9173 7450
rect 9024 7422 9035 7442
rect 9055 7422 9173 7442
rect 9713 7437 10334 7451
rect 10352 7437 10362 7455
rect 9713 7431 10362 7437
rect 9713 7430 10361 7431
rect 10324 7428 10361 7430
rect 9024 7415 9173 7422
rect 9024 7414 9065 7415
rect 8348 7361 8385 7362
rect 8444 7361 8481 7362
rect 8500 7361 8536 7413
rect 8555 7361 8592 7362
rect 8248 7352 8386 7361
rect 8248 7332 8357 7352
rect 8377 7332 8386 7352
rect 8248 7325 8386 7332
rect 8444 7352 8592 7361
rect 8444 7332 8453 7352
rect 8473 7332 8563 7352
rect 8583 7332 8592 7352
rect 8248 7323 8344 7325
rect 8444 7322 8592 7332
rect 8651 7352 8688 7362
rect 8763 7361 8800 7362
rect 8744 7359 8800 7361
rect 8651 7332 8659 7352
rect 8679 7332 8688 7352
rect 8500 7321 8536 7322
rect 8348 7262 8385 7263
rect 8651 7262 8688 7332
rect 8713 7352 8800 7359
rect 8713 7349 8771 7352
rect 8713 7329 8718 7349
rect 8739 7332 8771 7349
rect 8791 7332 8800 7352
rect 8739 7329 8800 7332
rect 8713 7322 8800 7329
rect 8859 7352 8896 7362
rect 8859 7332 8867 7352
rect 8887 7332 8896 7352
rect 8713 7321 8744 7322
rect 8347 7261 8688 7262
rect 8272 7256 8688 7261
rect 8272 7236 8275 7256
rect 8295 7236 8688 7256
rect 8859 7261 8896 7332
rect 8926 7361 8957 7414
rect 8976 7361 9013 7362
rect 8926 7352 9013 7361
rect 8926 7332 8984 7352
rect 9004 7332 9013 7352
rect 8926 7322 9013 7332
rect 9072 7352 9109 7362
rect 9072 7332 9080 7352
rect 9100 7332 9109 7352
rect 8926 7321 8957 7322
rect 9072 7261 9109 7332
rect 10327 7356 10364 7366
rect 10327 7338 10336 7356
rect 10354 7338 10364 7356
rect 10327 7329 10364 7338
rect 10327 7305 10362 7329
rect 10325 7281 10362 7305
rect 10324 7275 10362 7281
rect 8859 7237 9109 7261
rect 9735 7257 10362 7275
rect 9317 7240 9485 7241
rect 9736 7240 9760 7257
rect 9317 7214 9761 7240
rect 9317 7212 9485 7214
rect 9317 7034 9344 7212
rect 9384 7174 9448 7186
rect 9724 7182 9761 7214
rect 9932 7213 10181 7235
rect 9932 7182 9969 7213
rect 10145 7211 10181 7213
rect 10324 7216 10362 7257
rect 10145 7182 10182 7211
rect 9384 7173 9419 7174
rect 9361 7168 9419 7173
rect 9361 7148 9364 7168
rect 9384 7154 9419 7168
rect 9439 7154 9448 7174
rect 9384 7146 9448 7154
rect 9410 7145 9448 7146
rect 9411 7144 9448 7145
rect 9514 7178 9550 7179
rect 9622 7178 9658 7179
rect 9514 7172 9658 7178
rect 9514 7170 9580 7172
rect 9514 7150 9522 7170
rect 9542 7151 9580 7170
rect 9602 7170 9658 7172
rect 9602 7151 9630 7170
rect 9542 7150 9630 7151
rect 9650 7150 9658 7170
rect 9514 7144 9658 7150
rect 9724 7174 9762 7182
rect 9830 7178 9866 7179
rect 9724 7154 9733 7174
rect 9753 7154 9762 7174
rect 9724 7145 9762 7154
rect 9781 7171 9866 7178
rect 9781 7151 9788 7171
rect 9809 7170 9866 7171
rect 9809 7151 9838 7170
rect 9781 7150 9838 7151
rect 9858 7150 9866 7170
rect 9724 7144 9761 7145
rect 9781 7144 9866 7150
rect 9932 7174 9970 7182
rect 10043 7178 10079 7179
rect 9932 7154 9941 7174
rect 9961 7154 9970 7174
rect 9932 7145 9970 7154
rect 9994 7170 10079 7178
rect 9994 7150 10051 7170
rect 10071 7150 10079 7170
rect 9932 7144 9969 7145
rect 9994 7144 10079 7150
rect 10145 7174 10183 7182
rect 10145 7154 10154 7174
rect 10174 7154 10183 7174
rect 10145 7145 10183 7154
rect 10324 7181 10360 7216
rect 10324 7171 10361 7181
rect 10324 7153 10334 7171
rect 10352 7153 10361 7171
rect 10145 7144 10182 7145
rect 10324 7144 10361 7153
rect 9568 7123 9604 7144
rect 9994 7123 10025 7144
rect 9401 7119 9501 7123
rect 9401 7115 9463 7119
rect 9401 7089 9408 7115
rect 9434 7093 9463 7115
rect 9489 7093 9501 7119
rect 9434 7089 9501 7093
rect 9401 7086 9501 7089
rect 9569 7086 9604 7123
rect 9666 7120 10025 7123
rect 9666 7115 9888 7120
rect 9666 7091 9679 7115
rect 9703 7096 9888 7115
rect 9912 7096 10025 7120
rect 9703 7091 10025 7096
rect 9666 7087 10025 7091
rect 10092 7115 10241 7123
rect 10092 7095 10103 7115
rect 10123 7095 10241 7115
rect 10092 7088 10241 7095
rect 10092 7087 10133 7088
rect 9416 7034 9453 7035
rect 9512 7034 9549 7035
rect 9568 7034 9604 7086
rect 9623 7034 9660 7035
rect 9316 7025 9454 7034
rect 8304 7006 8472 7007
rect 8304 7003 8748 7006
rect 8304 6984 8679 7003
rect 8699 6984 8748 7003
rect 9316 7005 9425 7025
rect 9445 7005 9454 7025
rect 8304 6980 8748 6984
rect 8304 6978 8472 6980
rect 8304 6800 8331 6978
rect 8371 6940 8435 6952
rect 8711 6948 8748 6980
rect 8919 6979 9168 7001
rect 9316 6998 9454 7005
rect 9512 7025 9660 7034
rect 9512 7005 9521 7025
rect 9541 7005 9631 7025
rect 9651 7005 9660 7025
rect 9316 6996 9412 6998
rect 9512 6995 9660 7005
rect 9719 7025 9756 7035
rect 9831 7034 9868 7035
rect 9812 7032 9868 7034
rect 9719 7005 9727 7025
rect 9747 7005 9756 7025
rect 9568 6994 9604 6995
rect 8919 6948 8956 6979
rect 9132 6977 9168 6979
rect 9132 6948 9169 6977
rect 8371 6939 8406 6940
rect 8348 6934 8406 6939
rect 8348 6914 8351 6934
rect 8371 6920 8406 6934
rect 8426 6920 8435 6940
rect 8371 6912 8435 6920
rect 8397 6911 8435 6912
rect 8398 6910 8435 6911
rect 8501 6944 8537 6945
rect 8609 6944 8645 6945
rect 8501 6936 8645 6944
rect 8501 6916 8509 6936
rect 8529 6916 8561 6936
rect 8585 6916 8617 6936
rect 8637 6916 8645 6936
rect 8501 6910 8645 6916
rect 8711 6940 8749 6948
rect 8817 6944 8853 6945
rect 8711 6920 8720 6940
rect 8740 6920 8749 6940
rect 8711 6911 8749 6920
rect 8768 6937 8853 6944
rect 8768 6917 8775 6937
rect 8796 6936 8853 6937
rect 8796 6917 8825 6936
rect 8768 6916 8825 6917
rect 8845 6916 8853 6936
rect 8711 6910 8748 6911
rect 8768 6910 8853 6916
rect 8919 6940 8957 6948
rect 9030 6944 9066 6945
rect 8919 6920 8928 6940
rect 8948 6920 8957 6940
rect 8919 6911 8957 6920
rect 8981 6936 9066 6944
rect 8981 6916 9038 6936
rect 9058 6916 9066 6936
rect 8919 6910 8956 6911
rect 8981 6910 9066 6916
rect 9132 6940 9170 6948
rect 9132 6920 9141 6940
rect 9161 6920 9170 6940
rect 9416 6935 9453 6936
rect 9719 6935 9756 7005
rect 9781 7025 9868 7032
rect 9781 7022 9839 7025
rect 9781 7002 9786 7022
rect 9807 7005 9839 7022
rect 9859 7005 9868 7025
rect 9807 7002 9868 7005
rect 9781 6995 9868 7002
rect 9927 7025 9964 7035
rect 9927 7005 9935 7025
rect 9955 7005 9964 7025
rect 9781 6994 9812 6995
rect 9415 6934 9756 6935
rect 9132 6911 9170 6920
rect 9340 6929 9756 6934
rect 9132 6910 9169 6911
rect 8555 6889 8591 6910
rect 8981 6889 9012 6910
rect 9340 6909 9343 6929
rect 9363 6909 9756 6929
rect 9927 6934 9964 7005
rect 9994 7034 10025 7087
rect 10327 7072 10364 7082
rect 10327 7054 10336 7072
rect 10354 7054 10364 7072
rect 10327 7045 10364 7054
rect 10044 7034 10081 7035
rect 9994 7025 10081 7034
rect 9994 7005 10052 7025
rect 10072 7005 10081 7025
rect 9994 6995 10081 7005
rect 10140 7025 10177 7035
rect 10140 7005 10148 7025
rect 10168 7005 10177 7025
rect 9994 6994 10025 6995
rect 10140 6934 10177 7005
rect 10332 6980 10363 7045
rect 10331 6970 10368 6980
rect 10331 6968 10341 6970
rect 10265 6966 10341 6968
rect 9927 6910 10177 6934
rect 10262 6952 10341 6966
rect 10359 6952 10368 6970
rect 10262 6949 10368 6952
rect 9734 6890 9755 6909
rect 10262 6890 10288 6949
rect 10331 6943 10368 6949
rect 8388 6885 8488 6889
rect 8388 6881 8450 6885
rect 8388 6855 8395 6881
rect 8421 6859 8450 6881
rect 8476 6859 8488 6885
rect 8421 6855 8488 6859
rect 8388 6852 8488 6855
rect 8556 6852 8591 6889
rect 8653 6886 9012 6889
rect 8653 6881 8875 6886
rect 8653 6857 8666 6881
rect 8690 6862 8875 6881
rect 8899 6862 9012 6886
rect 8690 6857 9012 6862
rect 8653 6853 9012 6857
rect 9079 6881 9228 6889
rect 9079 6861 9090 6881
rect 9110 6861 9228 6881
rect 9734 6872 10288 6890
rect 10334 6879 10371 6881
rect 10262 6871 10288 6872
rect 10331 6871 10371 6879
rect 9079 6854 9228 6861
rect 10331 6859 10343 6871
rect 10322 6854 10343 6859
rect 9079 6853 9120 6854
rect 9738 6853 10343 6854
rect 10361 6853 10371 6871
rect 8403 6800 8440 6801
rect 8499 6800 8536 6801
rect 8555 6800 8591 6852
rect 8610 6800 8647 6801
rect 8303 6791 8441 6800
rect 8303 6771 8412 6791
rect 8432 6771 8441 6791
rect 8303 6764 8441 6771
rect 8499 6791 8647 6800
rect 8499 6771 8508 6791
rect 8528 6771 8618 6791
rect 8638 6771 8647 6791
rect 8303 6762 8399 6764
rect 8499 6761 8647 6771
rect 8706 6791 8743 6801
rect 8818 6800 8855 6801
rect 8799 6798 8855 6800
rect 8706 6771 8714 6791
rect 8734 6771 8743 6791
rect 8555 6760 8591 6761
rect 8403 6701 8440 6702
rect 8706 6701 8743 6771
rect 8768 6791 8855 6798
rect 8768 6788 8826 6791
rect 8768 6768 8773 6788
rect 8794 6771 8826 6788
rect 8846 6771 8855 6791
rect 8794 6768 8855 6771
rect 8768 6761 8855 6768
rect 8914 6791 8951 6801
rect 8914 6771 8922 6791
rect 8942 6771 8951 6791
rect 8768 6760 8799 6761
rect 8402 6700 8743 6701
rect 8327 6695 8743 6700
rect 8327 6675 8330 6695
rect 8350 6675 8743 6695
rect 8914 6700 8951 6771
rect 8981 6800 9012 6853
rect 9738 6844 10371 6853
rect 9738 6837 10370 6844
rect 9738 6835 9800 6837
rect 9316 6825 9484 6826
rect 9738 6825 9760 6835
rect 9031 6800 9068 6801
rect 8981 6791 9068 6800
rect 8981 6771 9039 6791
rect 9059 6771 9068 6791
rect 8981 6761 9068 6771
rect 9127 6791 9164 6801
rect 9127 6771 9135 6791
rect 9155 6771 9164 6791
rect 8981 6760 9012 6761
rect 9127 6700 9164 6771
rect 8914 6676 9164 6700
rect 9316 6799 9760 6825
rect 9316 6797 9484 6799
rect 9316 6619 9343 6797
rect 9383 6759 9447 6771
rect 9723 6767 9760 6799
rect 9931 6798 10180 6820
rect 9931 6767 9968 6798
rect 10144 6796 10180 6798
rect 10144 6767 10181 6796
rect 9383 6758 9418 6759
rect 9360 6753 9418 6758
rect 9360 6733 9363 6753
rect 9383 6739 9418 6753
rect 9438 6739 9447 6759
rect 9383 6731 9447 6739
rect 9409 6730 9447 6731
rect 9410 6729 9447 6730
rect 9513 6763 9549 6764
rect 9621 6763 9657 6764
rect 9513 6755 9657 6763
rect 9513 6735 9521 6755
rect 9541 6735 9570 6755
rect 9513 6734 9570 6735
rect 9592 6735 9629 6755
rect 9649 6735 9657 6755
rect 9592 6734 9657 6735
rect 9513 6729 9657 6734
rect 9723 6759 9761 6767
rect 9829 6763 9865 6764
rect 9723 6739 9732 6759
rect 9752 6739 9761 6759
rect 9723 6730 9761 6739
rect 9780 6756 9865 6763
rect 9780 6736 9787 6756
rect 9808 6755 9865 6756
rect 9808 6736 9837 6755
rect 9780 6735 9837 6736
rect 9857 6735 9865 6755
rect 9723 6729 9760 6730
rect 9780 6729 9865 6735
rect 9931 6759 9969 6767
rect 10042 6763 10078 6764
rect 9931 6739 9940 6759
rect 9960 6739 9969 6759
rect 9931 6730 9969 6739
rect 9993 6755 10078 6763
rect 9993 6735 10050 6755
rect 10070 6735 10078 6755
rect 9931 6729 9968 6730
rect 9993 6729 10078 6735
rect 10144 6759 10182 6767
rect 10144 6739 10153 6759
rect 10173 6739 10182 6759
rect 10144 6730 10182 6739
rect 10144 6729 10181 6730
rect 9567 6708 9603 6729
rect 9993 6708 10024 6729
rect 9400 6704 9500 6708
rect 9400 6700 9462 6704
rect 9400 6674 9407 6700
rect 9433 6678 9462 6700
rect 9488 6678 9500 6704
rect 9433 6674 9500 6678
rect 9400 6671 9500 6674
rect 9568 6671 9603 6708
rect 9665 6705 10024 6708
rect 9665 6700 9887 6705
rect 9665 6676 9678 6700
rect 9702 6681 9887 6700
rect 9911 6681 10024 6705
rect 9702 6676 10024 6681
rect 9665 6672 10024 6676
rect 10091 6700 10240 6708
rect 10091 6680 10102 6700
rect 10122 6680 10240 6700
rect 10091 6673 10240 6680
rect 10331 6688 10370 6837
rect 10091 6672 10132 6673
rect 9415 6619 9452 6620
rect 9511 6619 9548 6620
rect 9567 6619 9603 6671
rect 9622 6619 9659 6620
rect 9315 6610 9453 6619
rect 9315 6590 9424 6610
rect 9444 6590 9453 6610
rect 9315 6583 9453 6590
rect 9511 6610 9659 6619
rect 9511 6590 9520 6610
rect 9540 6590 9630 6610
rect 9650 6590 9659 6610
rect 9315 6581 9411 6583
rect 9511 6580 9659 6590
rect 9718 6610 9755 6620
rect 9830 6619 9867 6620
rect 9811 6617 9867 6619
rect 9718 6590 9726 6610
rect 9746 6590 9755 6610
rect 9567 6579 9603 6580
rect 8030 6517 8038 6536
rect 8061 6517 8067 6536
rect 8030 6506 8067 6517
rect 8096 6539 8264 6540
rect 8096 6513 8540 6539
rect 8096 6511 8264 6513
rect 8033 6446 8066 6506
rect 6278 6367 6446 6369
rect 6002 6341 6446 6367
rect 6003 6324 6027 6341
rect 6278 6340 6446 6341
rect 6814 6369 7064 6393
rect 5050 6317 5088 6323
rect 4461 6299 5088 6317
rect 5401 6306 6028 6324
rect 5401 6300 5439 6306
rect 3425 6230 3675 6254
rect 4043 6282 4211 6283
rect 4462 6282 4486 6299
rect 4043 6256 4487 6282
rect 4043 6254 4211 6256
rect 4043 6076 4070 6254
rect 4110 6216 4174 6228
rect 4450 6224 4487 6256
rect 4658 6255 4907 6277
rect 4658 6224 4695 6255
rect 4871 6253 4907 6255
rect 5050 6258 5088 6299
rect 4871 6224 4908 6253
rect 4110 6215 4145 6216
rect 4087 6210 4145 6215
rect 4087 6190 4090 6210
rect 4110 6196 4145 6210
rect 4165 6196 4174 6216
rect 4110 6188 4174 6196
rect 4136 6187 4174 6188
rect 4137 6186 4174 6187
rect 4240 6220 4276 6221
rect 4348 6220 4384 6221
rect 4240 6214 4384 6220
rect 4240 6212 4306 6214
rect 4240 6192 4248 6212
rect 4268 6193 4306 6212
rect 4328 6212 4384 6214
rect 4328 6193 4356 6212
rect 4268 6192 4356 6193
rect 4376 6192 4384 6212
rect 4240 6186 4384 6192
rect 4450 6216 4488 6224
rect 4556 6220 4592 6221
rect 4450 6196 4459 6216
rect 4479 6196 4488 6216
rect 4450 6187 4488 6196
rect 4507 6213 4592 6220
rect 4507 6193 4514 6213
rect 4535 6212 4592 6213
rect 4535 6193 4564 6212
rect 4507 6192 4564 6193
rect 4584 6192 4592 6212
rect 4450 6186 4487 6187
rect 4507 6186 4592 6192
rect 4658 6216 4696 6224
rect 4769 6220 4805 6221
rect 4658 6196 4667 6216
rect 4687 6196 4696 6216
rect 4658 6187 4696 6196
rect 4720 6212 4805 6220
rect 4720 6192 4777 6212
rect 4797 6192 4805 6212
rect 4658 6186 4695 6187
rect 4720 6186 4805 6192
rect 4871 6216 4909 6224
rect 4871 6196 4880 6216
rect 4900 6196 4909 6216
rect 4871 6187 4909 6196
rect 5050 6223 5086 6258
rect 5403 6254 5438 6300
rect 6814 6298 6851 6369
rect 6966 6308 6997 6309
rect 6814 6278 6823 6298
rect 6843 6278 6851 6298
rect 6814 6268 6851 6278
rect 6910 6298 6997 6308
rect 6910 6278 6919 6298
rect 6939 6278 6997 6298
rect 6910 6269 6997 6278
rect 6910 6268 6947 6269
rect 5401 6245 5438 6254
rect 5401 6227 5411 6245
rect 5429 6227 5438 6245
rect 5050 6213 5087 6223
rect 5401 6217 5438 6227
rect 6966 6216 6997 6269
rect 7027 6298 7064 6369
rect 7235 6374 7628 6394
rect 7648 6374 7651 6394
rect 7235 6369 7651 6374
rect 7235 6368 7576 6369
rect 7179 6308 7210 6309
rect 7027 6278 7036 6298
rect 7056 6278 7064 6298
rect 7027 6268 7064 6278
rect 7123 6301 7210 6308
rect 7123 6298 7184 6301
rect 7123 6278 7132 6298
rect 7152 6281 7184 6298
rect 7205 6281 7210 6301
rect 7152 6278 7210 6281
rect 7123 6271 7210 6278
rect 7235 6298 7272 6368
rect 7538 6367 7575 6368
rect 7387 6308 7423 6309
rect 7235 6278 7244 6298
rect 7264 6278 7272 6298
rect 7123 6269 7179 6271
rect 7123 6268 7160 6269
rect 7235 6268 7272 6278
rect 7331 6298 7479 6308
rect 7579 6305 7675 6307
rect 7331 6278 7340 6298
rect 7360 6278 7450 6298
rect 7470 6278 7479 6298
rect 7331 6269 7479 6278
rect 7537 6298 7675 6305
rect 7537 6278 7546 6298
rect 7566 6278 7675 6298
rect 7537 6269 7675 6278
rect 7331 6268 7368 6269
rect 7387 6217 7423 6269
rect 7442 6268 7479 6269
rect 7538 6268 7575 6269
rect 6858 6215 6899 6216
rect 5050 6195 5060 6213
rect 5078 6195 5087 6213
rect 4871 6186 4908 6187
rect 5050 6186 5087 6195
rect 6750 6208 6899 6215
rect 6750 6188 6868 6208
rect 6888 6188 6899 6208
rect 4294 6165 4330 6186
rect 4720 6165 4751 6186
rect 6750 6180 6899 6188
rect 6966 6212 7325 6216
rect 6966 6207 7288 6212
rect 6966 6183 7079 6207
rect 7103 6188 7288 6207
rect 7312 6188 7325 6212
rect 7103 6183 7325 6188
rect 6966 6180 7325 6183
rect 7387 6180 7422 6217
rect 7490 6214 7590 6217
rect 7490 6210 7557 6214
rect 7490 6184 7502 6210
rect 7528 6188 7557 6210
rect 7583 6188 7590 6214
rect 7528 6184 7590 6188
rect 7490 6180 7590 6184
rect 4127 6161 4227 6165
rect 4127 6157 4189 6161
rect 4127 6131 4134 6157
rect 4160 6135 4189 6157
rect 4215 6135 4227 6161
rect 4160 6131 4227 6135
rect 4127 6128 4227 6131
rect 4295 6128 4330 6165
rect 4392 6162 4751 6165
rect 4392 6157 4614 6162
rect 4392 6133 4405 6157
rect 4429 6138 4614 6157
rect 4638 6138 4751 6162
rect 4429 6133 4751 6138
rect 4392 6129 4751 6133
rect 4818 6157 4967 6165
rect 6966 6159 6997 6180
rect 7387 6159 7423 6180
rect 6809 6158 6846 6159
rect 4818 6137 4829 6157
rect 4849 6137 4967 6157
rect 5404 6153 5441 6155
rect 5404 6152 6052 6153
rect 4818 6130 4967 6137
rect 5403 6146 6052 6152
rect 4818 6129 4859 6130
rect 4142 6076 4179 6077
rect 4238 6076 4275 6077
rect 4294 6076 4330 6128
rect 4349 6076 4386 6077
rect 4042 6067 4180 6076
rect 2978 6049 3009 6052
rect 2978 6023 2985 6049
rect 3004 6023 3009 6049
rect 2978 5629 3009 6023
rect 3030 6048 3198 6049
rect 3030 6045 3474 6048
rect 3030 6026 3405 6045
rect 3425 6026 3474 6045
rect 4042 6047 4151 6067
rect 4171 6047 4180 6067
rect 3030 6022 3474 6026
rect 3030 6020 3198 6022
rect 3030 5842 3057 6020
rect 3097 5982 3161 5994
rect 3437 5990 3474 6022
rect 3645 6021 3894 6043
rect 4042 6040 4180 6047
rect 4238 6067 4386 6076
rect 4238 6047 4247 6067
rect 4267 6047 4357 6067
rect 4377 6047 4386 6067
rect 4042 6038 4138 6040
rect 4238 6037 4386 6047
rect 4445 6067 4482 6077
rect 4557 6076 4594 6077
rect 4538 6074 4594 6076
rect 4445 6047 4453 6067
rect 4473 6047 4482 6067
rect 4294 6036 4330 6037
rect 3645 5990 3682 6021
rect 3858 6019 3894 6021
rect 3858 5990 3895 6019
rect 3097 5981 3132 5982
rect 3074 5976 3132 5981
rect 3074 5956 3077 5976
rect 3097 5962 3132 5976
rect 3152 5962 3161 5982
rect 3097 5954 3161 5962
rect 3123 5953 3161 5954
rect 3124 5952 3161 5953
rect 3227 5986 3263 5987
rect 3335 5986 3371 5987
rect 3227 5978 3371 5986
rect 3227 5958 3235 5978
rect 3255 5977 3343 5978
rect 3255 5958 3288 5977
rect 3227 5957 3288 5958
rect 3312 5958 3343 5977
rect 3363 5958 3371 5978
rect 3312 5957 3371 5958
rect 3227 5952 3371 5957
rect 3437 5982 3475 5990
rect 3543 5986 3579 5987
rect 3437 5962 3446 5982
rect 3466 5962 3475 5982
rect 3437 5953 3475 5962
rect 3494 5979 3579 5986
rect 3494 5959 3501 5979
rect 3522 5978 3579 5979
rect 3522 5959 3551 5978
rect 3494 5958 3551 5959
rect 3571 5958 3579 5978
rect 3437 5952 3474 5953
rect 3494 5952 3579 5958
rect 3645 5982 3683 5990
rect 3756 5986 3792 5987
rect 3645 5962 3654 5982
rect 3674 5962 3683 5982
rect 3645 5953 3683 5962
rect 3707 5978 3792 5986
rect 3707 5958 3764 5978
rect 3784 5958 3792 5978
rect 3645 5952 3682 5953
rect 3707 5952 3792 5958
rect 3858 5982 3896 5990
rect 3858 5962 3867 5982
rect 3887 5962 3896 5982
rect 4142 5977 4179 5978
rect 4445 5977 4482 6047
rect 4507 6067 4594 6074
rect 4507 6064 4565 6067
rect 4507 6044 4512 6064
rect 4533 6047 4565 6064
rect 4585 6047 4594 6067
rect 4533 6044 4594 6047
rect 4507 6037 4594 6044
rect 4653 6067 4690 6077
rect 4653 6047 4661 6067
rect 4681 6047 4690 6067
rect 4507 6036 4538 6037
rect 4141 5976 4482 5977
rect 3858 5953 3896 5962
rect 4066 5971 4482 5976
rect 3858 5952 3895 5953
rect 3281 5931 3317 5952
rect 3707 5931 3738 5952
rect 4066 5951 4069 5971
rect 4089 5951 4482 5971
rect 4653 5976 4690 6047
rect 4720 6076 4751 6129
rect 5403 6128 5413 6146
rect 5431 6132 6052 6146
rect 5431 6128 5441 6132
rect 5882 6131 6052 6132
rect 5053 6114 5090 6124
rect 5053 6096 5062 6114
rect 5080 6096 5090 6114
rect 5053 6087 5090 6096
rect 5403 6118 5441 6128
rect 4770 6076 4807 6077
rect 4720 6067 4807 6076
rect 4720 6047 4778 6067
rect 4798 6047 4807 6067
rect 4720 6037 4807 6047
rect 4866 6067 4903 6077
rect 4866 6047 4874 6067
rect 4894 6047 4903 6067
rect 4720 6036 4751 6037
rect 4866 5976 4903 6047
rect 5058 6022 5089 6087
rect 5403 6040 5438 6118
rect 6015 6108 6052 6131
rect 6808 6149 6846 6158
rect 6808 6129 6817 6149
rect 6837 6129 6846 6149
rect 6808 6121 6846 6129
rect 6912 6153 6997 6159
rect 7022 6158 7059 6159
rect 6912 6133 6920 6153
rect 6940 6133 6997 6153
rect 6912 6125 6997 6133
rect 7021 6149 7059 6158
rect 7021 6129 7030 6149
rect 7050 6129 7059 6149
rect 6912 6124 6948 6125
rect 7021 6121 7059 6129
rect 7125 6153 7210 6159
rect 7230 6158 7267 6159
rect 7125 6133 7133 6153
rect 7153 6152 7210 6153
rect 7153 6133 7182 6152
rect 7125 6132 7182 6133
rect 7203 6132 7210 6152
rect 7125 6125 7210 6132
rect 7229 6149 7267 6158
rect 7229 6129 7238 6149
rect 7258 6129 7267 6149
rect 7125 6124 7161 6125
rect 7229 6121 7267 6129
rect 7333 6157 7477 6159
rect 7333 6153 7391 6157
rect 7333 6133 7341 6153
rect 7361 6133 7391 6153
rect 7333 6131 7391 6133
rect 7416 6153 7477 6157
rect 7416 6133 7449 6153
rect 7469 6133 7477 6153
rect 7416 6131 7477 6133
rect 7333 6125 7477 6131
rect 7333 6124 7369 6125
rect 7441 6124 7477 6125
rect 7543 6158 7580 6159
rect 7543 6157 7581 6158
rect 7543 6149 7607 6157
rect 7543 6129 7552 6149
rect 7572 6135 7607 6149
rect 7627 6135 7630 6155
rect 7572 6130 7630 6135
rect 7572 6129 7607 6130
rect 5399 6031 5438 6040
rect 5057 6012 5094 6022
rect 5057 6010 5067 6012
rect 4991 6008 5067 6010
rect 4653 5952 4903 5976
rect 4988 5994 5067 6008
rect 5085 5994 5094 6012
rect 5399 6013 5409 6031
rect 5427 6013 5438 6031
rect 5399 6007 5438 6013
rect 5594 6083 5844 6107
rect 5594 6012 5631 6083
rect 5746 6022 5777 6023
rect 5399 6003 5436 6007
rect 4988 5991 5094 5994
rect 4460 5932 4481 5951
rect 4988 5932 5014 5991
rect 5057 5985 5094 5991
rect 5594 5992 5603 6012
rect 5623 5992 5631 6012
rect 5594 5982 5631 5992
rect 5690 6012 5777 6022
rect 5690 5992 5699 6012
rect 5719 5992 5777 6012
rect 5690 5983 5777 5992
rect 5690 5982 5727 5983
rect 5402 5932 5439 5941
rect 3114 5927 3214 5931
rect 3114 5923 3176 5927
rect 3114 5897 3121 5923
rect 3147 5901 3176 5923
rect 3202 5901 3214 5927
rect 3147 5897 3214 5901
rect 3114 5894 3214 5897
rect 3282 5894 3317 5931
rect 3379 5928 3738 5931
rect 3379 5923 3601 5928
rect 3379 5899 3392 5923
rect 3416 5904 3601 5923
rect 3625 5904 3738 5928
rect 3416 5899 3738 5904
rect 3379 5895 3738 5899
rect 3805 5923 3954 5931
rect 3805 5903 3816 5923
rect 3836 5903 3954 5923
rect 4460 5914 5014 5932
rect 5060 5921 5097 5923
rect 4988 5913 5014 5914
rect 5057 5913 5097 5921
rect 3805 5896 3954 5903
rect 5057 5901 5069 5913
rect 5048 5896 5069 5901
rect 3805 5895 3846 5896
rect 4464 5895 5069 5896
rect 5087 5895 5097 5913
rect 3129 5842 3166 5843
rect 3225 5842 3262 5843
rect 3281 5842 3317 5894
rect 3336 5842 3373 5843
rect 3029 5833 3167 5842
rect 3029 5813 3138 5833
rect 3158 5813 3167 5833
rect 3029 5806 3167 5813
rect 3225 5833 3373 5842
rect 3225 5813 3234 5833
rect 3254 5813 3344 5833
rect 3364 5813 3373 5833
rect 3029 5804 3125 5806
rect 3225 5803 3373 5813
rect 3432 5833 3469 5843
rect 3544 5842 3581 5843
rect 3525 5840 3581 5842
rect 3432 5813 3440 5833
rect 3460 5813 3469 5833
rect 3281 5802 3317 5803
rect 3129 5743 3166 5744
rect 3432 5743 3469 5813
rect 3494 5833 3581 5840
rect 3494 5830 3552 5833
rect 3494 5810 3499 5830
rect 3520 5813 3552 5830
rect 3572 5813 3581 5833
rect 3520 5810 3581 5813
rect 3494 5803 3581 5810
rect 3640 5833 3677 5843
rect 3640 5813 3648 5833
rect 3668 5813 3677 5833
rect 3494 5802 3525 5803
rect 3128 5742 3469 5743
rect 3053 5737 3469 5742
rect 3053 5717 3056 5737
rect 3076 5717 3469 5737
rect 3640 5742 3677 5813
rect 3707 5842 3738 5895
rect 4464 5886 5097 5895
rect 5400 5914 5411 5932
rect 5429 5914 5439 5932
rect 5746 5930 5777 5983
rect 5807 6012 5844 6083
rect 6015 6088 6408 6108
rect 6428 6088 6431 6108
rect 6809 6092 6846 6121
rect 6015 6083 6431 6088
rect 6810 6090 6846 6092
rect 7022 6090 7059 6121
rect 6015 6082 6356 6083
rect 5959 6022 5990 6023
rect 5807 5992 5816 6012
rect 5836 5992 5844 6012
rect 5807 5982 5844 5992
rect 5903 6015 5990 6022
rect 5903 6012 5964 6015
rect 5903 5992 5912 6012
rect 5932 5995 5964 6012
rect 5985 5995 5990 6015
rect 5932 5992 5990 5995
rect 5903 5985 5990 5992
rect 6015 6012 6052 6082
rect 6318 6081 6355 6082
rect 6810 6068 7059 6090
rect 7230 6089 7267 6121
rect 7543 6117 7607 6129
rect 7647 6091 7674 6269
rect 7506 6089 7674 6091
rect 7230 6063 7674 6089
rect 7506 6062 7674 6063
rect 6167 6022 6203 6023
rect 6015 5992 6024 6012
rect 6044 5992 6052 6012
rect 5903 5983 5959 5985
rect 5903 5982 5940 5983
rect 6015 5982 6052 5992
rect 6111 6012 6259 6022
rect 6359 6019 6455 6021
rect 6111 5992 6120 6012
rect 6140 5992 6230 6012
rect 6250 5992 6259 6012
rect 6111 5983 6259 5992
rect 6317 6012 6455 6019
rect 6317 5992 6326 6012
rect 6346 5992 6455 6012
rect 6317 5983 6455 5992
rect 6111 5982 6148 5983
rect 6167 5931 6203 5983
rect 6222 5982 6259 5983
rect 6318 5982 6355 5983
rect 5638 5929 5679 5930
rect 4464 5879 5096 5886
rect 4464 5877 4526 5879
rect 4042 5867 4210 5868
rect 4464 5867 4486 5877
rect 3757 5842 3794 5843
rect 3707 5833 3794 5842
rect 3707 5813 3765 5833
rect 3785 5813 3794 5833
rect 3707 5803 3794 5813
rect 3853 5833 3890 5843
rect 3853 5813 3861 5833
rect 3881 5813 3890 5833
rect 3707 5802 3738 5803
rect 3853 5742 3890 5813
rect 3640 5718 3890 5742
rect 4042 5841 4486 5867
rect 4042 5839 4210 5841
rect 4042 5661 4069 5839
rect 4109 5801 4173 5813
rect 4449 5809 4486 5841
rect 4657 5840 4906 5862
rect 4657 5809 4694 5840
rect 4870 5838 4906 5840
rect 4870 5809 4907 5838
rect 4109 5800 4144 5801
rect 4086 5795 4144 5800
rect 4086 5775 4089 5795
rect 4109 5781 4144 5795
rect 4164 5781 4173 5801
rect 4109 5773 4173 5781
rect 4135 5772 4173 5773
rect 4136 5771 4173 5772
rect 4239 5805 4275 5806
rect 4347 5805 4383 5806
rect 4239 5797 4383 5805
rect 4239 5777 4247 5797
rect 4267 5777 4296 5797
rect 4239 5776 4296 5777
rect 4318 5777 4355 5797
rect 4375 5777 4383 5797
rect 4318 5776 4383 5777
rect 4239 5771 4383 5776
rect 4449 5801 4487 5809
rect 4555 5805 4591 5806
rect 4449 5781 4458 5801
rect 4478 5781 4487 5801
rect 4449 5772 4487 5781
rect 4506 5798 4591 5805
rect 4506 5778 4513 5798
rect 4534 5797 4591 5798
rect 4534 5778 4563 5797
rect 4506 5777 4563 5778
rect 4583 5777 4591 5797
rect 4449 5771 4486 5772
rect 4506 5771 4591 5777
rect 4657 5801 4695 5809
rect 4768 5805 4804 5806
rect 4657 5781 4666 5801
rect 4686 5781 4695 5801
rect 4657 5772 4695 5781
rect 4719 5797 4804 5805
rect 4719 5777 4776 5797
rect 4796 5777 4804 5797
rect 4657 5771 4694 5772
rect 4719 5771 4804 5777
rect 4870 5801 4908 5809
rect 4870 5781 4879 5801
rect 4899 5781 4908 5801
rect 4870 5772 4908 5781
rect 4870 5771 4907 5772
rect 4293 5750 4329 5771
rect 4719 5750 4750 5771
rect 4126 5746 4226 5750
rect 4126 5742 4188 5746
rect 4126 5716 4133 5742
rect 4159 5720 4188 5742
rect 4214 5720 4226 5746
rect 4159 5716 4226 5720
rect 4126 5713 4226 5716
rect 4294 5713 4329 5750
rect 4391 5747 4750 5750
rect 4391 5742 4613 5747
rect 4391 5718 4404 5742
rect 4428 5723 4613 5742
rect 4637 5723 4750 5747
rect 4428 5718 4750 5723
rect 4391 5714 4750 5718
rect 4817 5742 4966 5750
rect 4817 5722 4828 5742
rect 4848 5722 4966 5742
rect 4817 5715 4966 5722
rect 5057 5730 5096 5879
rect 5400 5765 5439 5914
rect 5530 5922 5679 5929
rect 5530 5902 5648 5922
rect 5668 5902 5679 5922
rect 5530 5894 5679 5902
rect 5746 5926 6105 5930
rect 5746 5921 6068 5926
rect 5746 5897 5859 5921
rect 5883 5902 6068 5921
rect 6092 5902 6105 5926
rect 5883 5897 6105 5902
rect 5746 5894 6105 5897
rect 6167 5894 6202 5931
rect 6270 5928 6370 5931
rect 6270 5924 6337 5928
rect 6270 5898 6282 5924
rect 6308 5902 6337 5924
rect 6363 5902 6370 5928
rect 6308 5898 6370 5902
rect 6270 5894 6370 5898
rect 5746 5873 5777 5894
rect 6167 5873 6203 5894
rect 5589 5872 5626 5873
rect 5588 5863 5626 5872
rect 5588 5843 5597 5863
rect 5617 5843 5626 5863
rect 5588 5835 5626 5843
rect 5692 5867 5777 5873
rect 5802 5872 5839 5873
rect 5692 5847 5700 5867
rect 5720 5847 5777 5867
rect 5692 5839 5777 5847
rect 5801 5863 5839 5872
rect 5801 5843 5810 5863
rect 5830 5843 5839 5863
rect 5692 5838 5728 5839
rect 5801 5835 5839 5843
rect 5905 5867 5990 5873
rect 6010 5872 6047 5873
rect 5905 5847 5913 5867
rect 5933 5866 5990 5867
rect 5933 5847 5962 5866
rect 5905 5846 5962 5847
rect 5983 5846 5990 5866
rect 5905 5839 5990 5846
rect 6009 5863 6047 5872
rect 6009 5843 6018 5863
rect 6038 5843 6047 5863
rect 5905 5838 5941 5839
rect 6009 5835 6047 5843
rect 6113 5868 6257 5873
rect 6113 5867 6178 5868
rect 6113 5847 6121 5867
rect 6141 5847 6178 5867
rect 6200 5867 6257 5868
rect 6200 5847 6229 5867
rect 6249 5847 6257 5867
rect 6113 5839 6257 5847
rect 6113 5838 6149 5839
rect 6221 5838 6257 5839
rect 6323 5872 6360 5873
rect 6323 5871 6361 5872
rect 6323 5863 6387 5871
rect 6323 5843 6332 5863
rect 6352 5849 6387 5863
rect 6407 5849 6410 5869
rect 6352 5844 6410 5849
rect 6352 5843 6387 5844
rect 5589 5806 5626 5835
rect 5590 5804 5626 5806
rect 5802 5804 5839 5835
rect 5590 5782 5839 5804
rect 6010 5803 6047 5835
rect 6323 5831 6387 5843
rect 6427 5805 6454 5983
rect 6286 5803 6454 5805
rect 6010 5777 6454 5803
rect 6606 5902 6856 5926
rect 6606 5831 6643 5902
rect 6758 5841 6789 5842
rect 6606 5811 6615 5831
rect 6635 5811 6643 5831
rect 6606 5801 6643 5811
rect 6702 5831 6789 5841
rect 6702 5811 6711 5831
rect 6731 5811 6789 5831
rect 6702 5802 6789 5811
rect 6702 5801 6739 5802
rect 6010 5767 6032 5777
rect 6286 5776 6454 5777
rect 5970 5765 6032 5767
rect 5400 5758 6032 5765
rect 4817 5714 4858 5715
rect 4141 5661 4178 5662
rect 4237 5661 4274 5662
rect 4293 5661 4329 5713
rect 4348 5661 4385 5662
rect 4041 5652 4179 5661
rect 4041 5632 4150 5652
rect 4170 5632 4179 5652
rect 2978 5628 3148 5629
rect 2978 5613 3424 5628
rect 4041 5625 4179 5632
rect 4237 5652 4385 5661
rect 4237 5632 4246 5652
rect 4266 5632 4356 5652
rect 4376 5632 4385 5652
rect 4041 5623 4137 5625
rect 2980 5602 3424 5613
rect 2980 5600 3148 5602
rect 2980 5422 3007 5600
rect 3047 5562 3111 5574
rect 3387 5570 3424 5602
rect 3595 5601 3844 5623
rect 4237 5622 4385 5632
rect 4444 5652 4481 5662
rect 4556 5661 4593 5662
rect 4537 5659 4593 5661
rect 4444 5632 4452 5652
rect 4472 5632 4481 5652
rect 4293 5621 4329 5622
rect 3595 5570 3632 5601
rect 3808 5599 3844 5601
rect 3808 5570 3845 5599
rect 3047 5561 3082 5562
rect 3024 5556 3082 5561
rect 3024 5536 3027 5556
rect 3047 5542 3082 5556
rect 3102 5542 3111 5562
rect 3047 5534 3111 5542
rect 3073 5533 3111 5534
rect 3074 5532 3111 5533
rect 3177 5566 3213 5567
rect 3285 5566 3321 5567
rect 3177 5558 3321 5566
rect 3177 5538 3185 5558
rect 3205 5557 3293 5558
rect 3205 5540 3233 5557
rect 3257 5540 3293 5557
rect 3205 5538 3293 5540
rect 3313 5538 3321 5558
rect 3177 5532 3321 5538
rect 3387 5562 3425 5570
rect 3493 5566 3529 5567
rect 3387 5542 3396 5562
rect 3416 5542 3425 5562
rect 3387 5533 3425 5542
rect 3444 5559 3529 5566
rect 3444 5539 3451 5559
rect 3472 5558 3529 5559
rect 3472 5539 3501 5558
rect 3444 5538 3501 5539
rect 3521 5538 3529 5558
rect 3387 5532 3424 5533
rect 3444 5532 3529 5538
rect 3595 5562 3633 5570
rect 3706 5566 3742 5567
rect 3595 5542 3604 5562
rect 3624 5542 3633 5562
rect 3595 5533 3633 5542
rect 3657 5558 3742 5566
rect 3657 5538 3714 5558
rect 3734 5538 3742 5558
rect 3595 5532 3632 5533
rect 3657 5532 3742 5538
rect 3808 5562 3846 5570
rect 4141 5562 4178 5563
rect 4444 5562 4481 5632
rect 4506 5652 4593 5659
rect 4506 5649 4564 5652
rect 4506 5629 4511 5649
rect 4532 5632 4564 5649
rect 4584 5632 4593 5652
rect 4532 5629 4593 5632
rect 4506 5622 4593 5629
rect 4652 5652 4689 5662
rect 4652 5632 4660 5652
rect 4680 5632 4689 5652
rect 4506 5621 4537 5622
rect 3808 5542 3817 5562
rect 3837 5542 3846 5562
rect 4140 5561 4481 5562
rect 3808 5533 3846 5542
rect 4065 5556 4481 5561
rect 4065 5536 4068 5556
rect 4088 5536 4481 5556
rect 4652 5561 4689 5632
rect 4719 5661 4750 5714
rect 5057 5712 5067 5730
rect 5085 5712 5096 5730
rect 5399 5749 6032 5758
rect 6758 5749 6789 5802
rect 6819 5831 6856 5902
rect 7027 5907 7420 5927
rect 7440 5907 7443 5927
rect 7027 5902 7443 5907
rect 7027 5901 7368 5902
rect 6971 5841 7002 5842
rect 6819 5811 6828 5831
rect 6848 5811 6856 5831
rect 6819 5801 6856 5811
rect 6915 5834 7002 5841
rect 6915 5831 6976 5834
rect 6915 5811 6924 5831
rect 6944 5814 6976 5831
rect 6997 5814 7002 5834
rect 6944 5811 7002 5814
rect 6915 5804 7002 5811
rect 7027 5831 7064 5901
rect 7330 5900 7367 5901
rect 7179 5841 7215 5842
rect 7027 5811 7036 5831
rect 7056 5811 7064 5831
rect 6915 5802 6971 5804
rect 6915 5801 6952 5802
rect 7027 5801 7064 5811
rect 7123 5831 7271 5841
rect 7371 5838 7467 5840
rect 7123 5811 7132 5831
rect 7152 5811 7242 5831
rect 7262 5811 7271 5831
rect 7123 5802 7271 5811
rect 7329 5831 7467 5838
rect 7329 5811 7338 5831
rect 7358 5811 7467 5831
rect 7329 5802 7467 5811
rect 7123 5801 7160 5802
rect 7179 5750 7215 5802
rect 7234 5801 7271 5802
rect 7330 5801 7367 5802
rect 5399 5731 5409 5749
rect 5427 5748 6032 5749
rect 6650 5748 6691 5749
rect 5427 5743 5448 5748
rect 5427 5731 5439 5743
rect 6542 5741 6691 5748
rect 5399 5723 5439 5731
rect 5482 5730 5508 5731
rect 5399 5721 5436 5723
rect 5482 5712 6036 5730
rect 6542 5721 6660 5741
rect 6680 5721 6691 5741
rect 6542 5713 6691 5721
rect 6758 5745 7117 5749
rect 6758 5740 7080 5745
rect 6758 5716 6871 5740
rect 6895 5721 7080 5740
rect 7104 5721 7117 5745
rect 6895 5716 7117 5721
rect 6758 5713 7117 5716
rect 7179 5713 7214 5750
rect 7282 5747 7382 5750
rect 7282 5743 7349 5747
rect 7282 5717 7294 5743
rect 7320 5721 7349 5743
rect 7375 5721 7382 5747
rect 7320 5717 7382 5721
rect 7282 5713 7382 5717
rect 5057 5703 5094 5712
rect 4769 5661 4806 5662
rect 4719 5652 4806 5661
rect 4719 5632 4777 5652
rect 4797 5632 4806 5652
rect 4719 5622 4806 5632
rect 4865 5652 4902 5662
rect 4865 5632 4873 5652
rect 4893 5632 4902 5652
rect 5402 5653 5439 5659
rect 5482 5653 5508 5712
rect 6015 5693 6036 5712
rect 5402 5650 5508 5653
rect 5060 5637 5097 5641
rect 4719 5621 4750 5622
rect 4865 5561 4902 5632
rect 4652 5537 4902 5561
rect 5058 5631 5097 5637
rect 5058 5613 5069 5631
rect 5087 5613 5097 5631
rect 5402 5632 5411 5650
rect 5429 5636 5508 5650
rect 5593 5668 5843 5692
rect 5429 5634 5505 5636
rect 5429 5632 5439 5634
rect 5402 5622 5439 5632
rect 5058 5604 5097 5613
rect 3808 5532 3845 5533
rect 3231 5511 3267 5532
rect 3657 5511 3688 5532
rect 4444 5513 4481 5536
rect 5058 5526 5093 5604
rect 5407 5557 5438 5622
rect 5593 5597 5630 5668
rect 5745 5607 5776 5608
rect 5593 5577 5602 5597
rect 5622 5577 5630 5597
rect 5593 5567 5630 5577
rect 5689 5597 5776 5607
rect 5689 5577 5698 5597
rect 5718 5577 5776 5597
rect 5689 5568 5776 5577
rect 5689 5567 5726 5568
rect 5055 5516 5093 5526
rect 5406 5548 5443 5557
rect 5406 5530 5416 5548
rect 5434 5530 5443 5548
rect 5406 5520 5443 5530
rect 4444 5512 4614 5513
rect 5055 5512 5065 5516
rect 3064 5507 3164 5511
rect 3064 5503 3126 5507
rect 3064 5477 3071 5503
rect 3097 5481 3126 5503
rect 3152 5481 3164 5507
rect 3097 5477 3164 5481
rect 3064 5474 3164 5477
rect 3232 5474 3267 5511
rect 3329 5508 3688 5511
rect 3329 5503 3551 5508
rect 3329 5479 3342 5503
rect 3366 5484 3551 5503
rect 3575 5484 3688 5508
rect 3366 5479 3688 5484
rect 3329 5475 3688 5479
rect 3755 5503 3904 5511
rect 3755 5483 3766 5503
rect 3786 5483 3904 5503
rect 4444 5498 5065 5512
rect 5083 5498 5093 5516
rect 5745 5515 5776 5568
rect 5806 5597 5843 5668
rect 6014 5673 6407 5693
rect 6427 5673 6430 5693
rect 6758 5692 6789 5713
rect 7179 5692 7215 5713
rect 6601 5691 6638 5692
rect 6014 5668 6430 5673
rect 6600 5682 6638 5691
rect 6014 5667 6355 5668
rect 5958 5607 5989 5608
rect 5806 5577 5815 5597
rect 5835 5577 5843 5597
rect 5806 5567 5843 5577
rect 5902 5600 5989 5607
rect 5902 5597 5963 5600
rect 5902 5577 5911 5597
rect 5931 5580 5963 5597
rect 5984 5580 5989 5600
rect 5931 5577 5989 5580
rect 5902 5570 5989 5577
rect 6014 5597 6051 5667
rect 6317 5666 6354 5667
rect 6600 5662 6609 5682
rect 6629 5662 6638 5682
rect 6600 5654 6638 5662
rect 6704 5686 6789 5692
rect 6814 5691 6851 5692
rect 6704 5666 6712 5686
rect 6732 5666 6789 5686
rect 6704 5658 6789 5666
rect 6813 5682 6851 5691
rect 6813 5662 6822 5682
rect 6842 5662 6851 5682
rect 6704 5657 6740 5658
rect 6813 5654 6851 5662
rect 6917 5686 7002 5692
rect 7022 5691 7059 5692
rect 6917 5666 6925 5686
rect 6945 5685 7002 5686
rect 6945 5666 6974 5685
rect 6917 5665 6974 5666
rect 6995 5665 7002 5685
rect 6917 5658 7002 5665
rect 7021 5682 7059 5691
rect 7021 5662 7030 5682
rect 7050 5662 7059 5682
rect 6917 5657 6953 5658
rect 7021 5654 7059 5662
rect 7125 5686 7269 5692
rect 7125 5666 7133 5686
rect 7153 5666 7185 5686
rect 7209 5666 7241 5686
rect 7261 5666 7269 5686
rect 7125 5658 7269 5666
rect 7125 5657 7161 5658
rect 7233 5657 7269 5658
rect 7335 5691 7372 5692
rect 7335 5690 7373 5691
rect 7335 5682 7399 5690
rect 7335 5662 7344 5682
rect 7364 5668 7399 5682
rect 7419 5668 7422 5688
rect 7364 5663 7422 5668
rect 7364 5662 7399 5663
rect 6601 5625 6638 5654
rect 6602 5623 6638 5625
rect 6814 5623 6851 5654
rect 6166 5607 6202 5608
rect 6014 5577 6023 5597
rect 6043 5577 6051 5597
rect 5902 5568 5958 5570
rect 5902 5567 5939 5568
rect 6014 5567 6051 5577
rect 6110 5597 6258 5607
rect 6358 5604 6454 5606
rect 6110 5577 6119 5597
rect 6139 5577 6229 5597
rect 6249 5577 6258 5597
rect 6110 5568 6258 5577
rect 6316 5597 6454 5604
rect 6602 5601 6851 5623
rect 7022 5622 7059 5654
rect 7335 5650 7399 5662
rect 7439 5624 7466 5802
rect 7298 5622 7466 5624
rect 7022 5618 7466 5622
rect 6316 5577 6325 5597
rect 6345 5577 6454 5597
rect 7022 5599 7071 5618
rect 7091 5599 7466 5618
rect 7022 5596 7466 5599
rect 7298 5595 7466 5596
rect 6316 5568 6454 5577
rect 6110 5567 6147 5568
rect 6166 5516 6202 5568
rect 6221 5567 6258 5568
rect 6317 5567 6354 5568
rect 5637 5514 5678 5515
rect 4444 5492 5093 5498
rect 5529 5507 5678 5514
rect 4444 5491 5092 5492
rect 5055 5489 5092 5491
rect 3755 5476 3904 5483
rect 5529 5487 5647 5507
rect 5667 5487 5678 5507
rect 5529 5479 5678 5487
rect 5745 5511 6104 5515
rect 5745 5506 6067 5511
rect 5745 5482 5858 5506
rect 5882 5487 6067 5506
rect 6091 5487 6104 5511
rect 5882 5482 6104 5487
rect 5745 5479 6104 5482
rect 6166 5479 6201 5516
rect 6269 5513 6369 5516
rect 6269 5509 6336 5513
rect 6269 5483 6281 5509
rect 6307 5487 6336 5509
rect 6362 5487 6369 5513
rect 6307 5483 6369 5487
rect 6269 5479 6369 5483
rect 3755 5475 3796 5476
rect 3079 5422 3116 5423
rect 3175 5422 3212 5423
rect 3231 5422 3267 5474
rect 3286 5422 3323 5423
rect 2979 5413 3117 5422
rect 2979 5393 3088 5413
rect 3108 5393 3117 5413
rect 2979 5386 3117 5393
rect 3175 5413 3323 5422
rect 3175 5393 3184 5413
rect 3204 5393 3294 5413
rect 3314 5393 3323 5413
rect 2979 5384 3075 5386
rect 3175 5383 3323 5393
rect 3382 5413 3419 5423
rect 3494 5422 3531 5423
rect 3475 5420 3531 5422
rect 3382 5393 3390 5413
rect 3410 5393 3419 5413
rect 3231 5382 3267 5383
rect 3079 5323 3116 5324
rect 3382 5323 3419 5393
rect 3444 5413 3531 5420
rect 3444 5410 3502 5413
rect 3444 5390 3449 5410
rect 3470 5393 3502 5410
rect 3522 5393 3531 5413
rect 3470 5390 3531 5393
rect 3444 5383 3531 5390
rect 3590 5413 3627 5423
rect 3590 5393 3598 5413
rect 3618 5393 3627 5413
rect 3444 5382 3475 5383
rect 3078 5322 3419 5323
rect 3003 5317 3419 5322
rect 3003 5297 3006 5317
rect 3026 5297 3419 5317
rect 3590 5322 3627 5393
rect 3657 5422 3688 5475
rect 5745 5458 5776 5479
rect 6166 5458 6202 5479
rect 5409 5449 5446 5458
rect 5588 5457 5625 5458
rect 5409 5431 5418 5449
rect 5436 5431 5446 5449
rect 3707 5422 3744 5423
rect 3657 5413 3744 5422
rect 3657 5393 3715 5413
rect 3735 5393 3744 5413
rect 3657 5383 3744 5393
rect 3803 5413 3840 5423
rect 3803 5393 3811 5413
rect 3831 5393 3840 5413
rect 3657 5382 3688 5383
rect 3803 5322 3840 5393
rect 5058 5417 5095 5427
rect 5409 5421 5446 5431
rect 5058 5399 5067 5417
rect 5085 5399 5095 5417
rect 5058 5390 5095 5399
rect 5058 5366 5093 5390
rect 5410 5386 5446 5421
rect 5587 5448 5625 5457
rect 5587 5428 5596 5448
rect 5616 5428 5625 5448
rect 5587 5420 5625 5428
rect 5691 5452 5776 5458
rect 5801 5457 5838 5458
rect 5691 5432 5699 5452
rect 5719 5432 5776 5452
rect 5691 5424 5776 5432
rect 5800 5448 5838 5457
rect 5800 5428 5809 5448
rect 5829 5428 5838 5448
rect 5691 5423 5727 5424
rect 5800 5420 5838 5428
rect 5904 5452 5989 5458
rect 6009 5457 6046 5458
rect 5904 5432 5912 5452
rect 5932 5451 5989 5452
rect 5932 5432 5961 5451
rect 5904 5431 5961 5432
rect 5982 5431 5989 5451
rect 5904 5424 5989 5431
rect 6008 5448 6046 5457
rect 6008 5428 6017 5448
rect 6037 5428 6046 5448
rect 5904 5423 5940 5424
rect 6008 5420 6046 5428
rect 6112 5452 6256 5458
rect 6112 5432 6120 5452
rect 6140 5451 6228 5452
rect 6140 5432 6168 5451
rect 6112 5430 6168 5432
rect 6190 5432 6228 5451
rect 6248 5432 6256 5452
rect 6190 5430 6256 5432
rect 6112 5424 6256 5430
rect 6112 5423 6148 5424
rect 6220 5423 6256 5424
rect 6322 5457 6359 5458
rect 6322 5456 6360 5457
rect 6322 5448 6386 5456
rect 6322 5428 6331 5448
rect 6351 5434 6386 5448
rect 6406 5434 6409 5454
rect 6351 5429 6409 5434
rect 6351 5428 6386 5429
rect 5588 5391 5625 5420
rect 5056 5342 5093 5366
rect 5055 5336 5093 5342
rect 3590 5298 3840 5322
rect 4466 5318 5093 5336
rect 4048 5301 4216 5302
rect 4467 5301 4491 5318
rect 4048 5275 4492 5301
rect 4048 5273 4216 5275
rect 4048 5095 4075 5273
rect 4115 5235 4179 5247
rect 4455 5243 4492 5275
rect 4663 5274 4912 5296
rect 4663 5243 4700 5274
rect 4876 5272 4912 5274
rect 5055 5277 5093 5318
rect 5408 5345 5446 5386
rect 5589 5389 5625 5391
rect 5801 5389 5838 5420
rect 5589 5367 5838 5389
rect 6009 5388 6046 5420
rect 6322 5416 6386 5428
rect 6426 5390 6453 5568
rect 6285 5388 6453 5390
rect 6009 5362 6453 5388
rect 6010 5345 6034 5362
rect 6285 5361 6453 5362
rect 5408 5327 6035 5345
rect 6661 5341 6911 5365
rect 5408 5321 5446 5327
rect 5408 5297 5445 5321
rect 4876 5243 4913 5272
rect 4115 5234 4150 5235
rect 4092 5229 4150 5234
rect 4092 5209 4095 5229
rect 4115 5215 4150 5229
rect 4170 5215 4179 5235
rect 4115 5207 4179 5215
rect 4141 5206 4179 5207
rect 4142 5205 4179 5206
rect 4245 5239 4281 5240
rect 4353 5239 4389 5240
rect 4245 5233 4389 5239
rect 4245 5231 4311 5233
rect 4245 5211 4253 5231
rect 4273 5212 4311 5231
rect 4333 5231 4389 5233
rect 4333 5212 4361 5231
rect 4273 5211 4361 5212
rect 4381 5211 4389 5231
rect 4245 5205 4389 5211
rect 4455 5235 4493 5243
rect 4561 5239 4597 5240
rect 4455 5215 4464 5235
rect 4484 5215 4493 5235
rect 4455 5206 4493 5215
rect 4512 5232 4597 5239
rect 4512 5212 4519 5232
rect 4540 5231 4597 5232
rect 4540 5212 4569 5231
rect 4512 5211 4569 5212
rect 4589 5211 4597 5231
rect 4455 5205 4492 5206
rect 4512 5205 4597 5211
rect 4663 5235 4701 5243
rect 4774 5239 4810 5240
rect 4663 5215 4672 5235
rect 4692 5215 4701 5235
rect 4663 5206 4701 5215
rect 4725 5231 4810 5239
rect 4725 5211 4782 5231
rect 4802 5211 4810 5231
rect 4663 5205 4700 5206
rect 4725 5205 4810 5211
rect 4876 5235 4914 5243
rect 4876 5215 4885 5235
rect 4905 5215 4914 5235
rect 4876 5206 4914 5215
rect 5055 5242 5091 5277
rect 5408 5273 5443 5297
rect 5406 5264 5443 5273
rect 5406 5246 5416 5264
rect 5434 5246 5443 5264
rect 5055 5232 5092 5242
rect 5406 5236 5443 5246
rect 6661 5270 6698 5341
rect 6813 5280 6844 5281
rect 6661 5250 6670 5270
rect 6690 5250 6698 5270
rect 6661 5240 6698 5250
rect 6757 5270 6844 5280
rect 6757 5250 6766 5270
rect 6786 5250 6844 5270
rect 6757 5241 6844 5250
rect 6757 5240 6794 5241
rect 5055 5214 5065 5232
rect 5083 5214 5092 5232
rect 4876 5205 4913 5206
rect 5055 5205 5092 5214
rect 4299 5184 4335 5205
rect 4725 5184 4756 5205
rect 6813 5188 6844 5241
rect 6874 5270 6911 5341
rect 7082 5346 7475 5366
rect 7495 5346 7498 5366
rect 7082 5341 7498 5346
rect 7082 5340 7423 5341
rect 7026 5280 7057 5281
rect 6874 5250 6883 5270
rect 6903 5250 6911 5270
rect 6874 5240 6911 5250
rect 6970 5273 7057 5280
rect 6970 5270 7031 5273
rect 6970 5250 6979 5270
rect 6999 5253 7031 5270
rect 7052 5253 7057 5273
rect 6999 5250 7057 5253
rect 6970 5243 7057 5250
rect 7082 5270 7119 5340
rect 7385 5339 7422 5340
rect 7234 5280 7270 5281
rect 7082 5250 7091 5270
rect 7111 5250 7119 5270
rect 6970 5241 7026 5243
rect 6970 5240 7007 5241
rect 7082 5240 7119 5250
rect 7178 5270 7326 5280
rect 7426 5277 7522 5279
rect 7178 5250 7187 5270
rect 7207 5250 7297 5270
rect 7317 5250 7326 5270
rect 7178 5241 7326 5250
rect 7384 5270 7522 5277
rect 7384 5250 7393 5270
rect 7413 5250 7522 5270
rect 7384 5241 7522 5250
rect 7178 5240 7215 5241
rect 7234 5189 7270 5241
rect 7289 5240 7326 5241
rect 7385 5240 7422 5241
rect 6705 5187 6746 5188
rect 4132 5180 4232 5184
rect 4132 5176 4194 5180
rect 4132 5150 4139 5176
rect 4165 5154 4194 5176
rect 4220 5154 4232 5180
rect 4165 5150 4232 5154
rect 4132 5147 4232 5150
rect 4300 5147 4335 5184
rect 4397 5181 4756 5184
rect 4397 5176 4619 5181
rect 4397 5152 4410 5176
rect 4434 5157 4619 5176
rect 4643 5157 4756 5181
rect 4434 5152 4756 5157
rect 4397 5148 4756 5152
rect 4823 5176 4972 5184
rect 4823 5156 4834 5176
rect 4854 5156 4972 5176
rect 6597 5180 6746 5187
rect 5409 5172 5446 5174
rect 5409 5171 6057 5172
rect 4823 5149 4972 5156
rect 5408 5165 6057 5171
rect 4823 5148 4864 5149
rect 4147 5095 4184 5096
rect 4243 5095 4280 5096
rect 4299 5095 4335 5147
rect 4354 5095 4391 5096
rect 4047 5086 4185 5095
rect 3035 5067 3203 5068
rect 3035 5064 3479 5067
rect 3035 5045 3410 5064
rect 3430 5045 3479 5064
rect 4047 5066 4156 5086
rect 4176 5066 4185 5086
rect 3035 5041 3479 5045
rect 3035 5039 3203 5041
rect 3035 4861 3062 5039
rect 3102 5001 3166 5013
rect 3442 5009 3479 5041
rect 3650 5040 3899 5062
rect 4047 5059 4185 5066
rect 4243 5086 4391 5095
rect 4243 5066 4252 5086
rect 4272 5066 4362 5086
rect 4382 5066 4391 5086
rect 4047 5057 4143 5059
rect 4243 5056 4391 5066
rect 4450 5086 4487 5096
rect 4562 5095 4599 5096
rect 4543 5093 4599 5095
rect 4450 5066 4458 5086
rect 4478 5066 4487 5086
rect 4299 5055 4335 5056
rect 3650 5009 3687 5040
rect 3863 5038 3899 5040
rect 3863 5009 3900 5038
rect 3102 5000 3137 5001
rect 3079 4995 3137 5000
rect 3079 4975 3082 4995
rect 3102 4981 3137 4995
rect 3157 4981 3166 5001
rect 3102 4973 3166 4981
rect 3128 4972 3166 4973
rect 3129 4971 3166 4972
rect 3232 5005 3268 5006
rect 3340 5005 3376 5006
rect 3232 4997 3376 5005
rect 3232 4977 3240 4997
rect 3260 4977 3292 4997
rect 3316 4977 3348 4997
rect 3368 4977 3376 4997
rect 3232 4971 3376 4977
rect 3442 5001 3480 5009
rect 3548 5005 3584 5006
rect 3442 4981 3451 5001
rect 3471 4981 3480 5001
rect 3442 4972 3480 4981
rect 3499 4998 3584 5005
rect 3499 4978 3506 4998
rect 3527 4997 3584 4998
rect 3527 4978 3556 4997
rect 3499 4977 3556 4978
rect 3576 4977 3584 4997
rect 3442 4971 3479 4972
rect 3499 4971 3584 4977
rect 3650 5001 3688 5009
rect 3761 5005 3797 5006
rect 3650 4981 3659 5001
rect 3679 4981 3688 5001
rect 3650 4972 3688 4981
rect 3712 4997 3797 5005
rect 3712 4977 3769 4997
rect 3789 4977 3797 4997
rect 3650 4971 3687 4972
rect 3712 4971 3797 4977
rect 3863 5001 3901 5009
rect 3863 4981 3872 5001
rect 3892 4981 3901 5001
rect 4147 4996 4184 4997
rect 4450 4996 4487 5066
rect 4512 5086 4599 5093
rect 4512 5083 4570 5086
rect 4512 5063 4517 5083
rect 4538 5066 4570 5083
rect 4590 5066 4599 5086
rect 4538 5063 4599 5066
rect 4512 5056 4599 5063
rect 4658 5086 4695 5096
rect 4658 5066 4666 5086
rect 4686 5066 4695 5086
rect 4512 5055 4543 5056
rect 4146 4995 4487 4996
rect 3863 4972 3901 4981
rect 4071 4990 4487 4995
rect 3863 4971 3900 4972
rect 3286 4950 3322 4971
rect 3712 4950 3743 4971
rect 4071 4970 4074 4990
rect 4094 4970 4487 4990
rect 4658 4995 4695 5066
rect 4725 5095 4756 5148
rect 5408 5147 5418 5165
rect 5436 5151 6057 5165
rect 6597 5160 6715 5180
rect 6735 5160 6746 5180
rect 6597 5152 6746 5160
rect 6813 5184 7172 5188
rect 6813 5179 7135 5184
rect 6813 5155 6926 5179
rect 6950 5160 7135 5179
rect 7159 5160 7172 5184
rect 6950 5155 7172 5160
rect 6813 5152 7172 5155
rect 7234 5152 7269 5189
rect 7337 5186 7437 5189
rect 7337 5182 7404 5186
rect 7337 5156 7349 5182
rect 7375 5160 7404 5182
rect 7430 5160 7437 5186
rect 7375 5156 7437 5160
rect 7337 5152 7437 5156
rect 5436 5147 5446 5151
rect 5887 5150 6057 5151
rect 5058 5133 5095 5143
rect 5058 5115 5067 5133
rect 5085 5115 5095 5133
rect 5058 5106 5095 5115
rect 5408 5137 5446 5147
rect 4775 5095 4812 5096
rect 4725 5086 4812 5095
rect 4725 5066 4783 5086
rect 4803 5066 4812 5086
rect 4725 5056 4812 5066
rect 4871 5086 4908 5096
rect 4871 5066 4879 5086
rect 4899 5066 4908 5086
rect 4725 5055 4756 5056
rect 4871 4995 4908 5066
rect 5063 5041 5094 5106
rect 5408 5059 5443 5137
rect 6020 5127 6057 5150
rect 6813 5131 6844 5152
rect 7234 5131 7270 5152
rect 6656 5130 6693 5131
rect 5404 5050 5443 5059
rect 5062 5031 5099 5041
rect 5062 5029 5072 5031
rect 4996 5027 5072 5029
rect 4658 4971 4908 4995
rect 4993 5013 5072 5027
rect 5090 5013 5099 5031
rect 5404 5032 5414 5050
rect 5432 5032 5443 5050
rect 5404 5026 5443 5032
rect 5599 5102 5849 5126
rect 5599 5031 5636 5102
rect 5751 5041 5782 5042
rect 5404 5022 5441 5026
rect 4993 5010 5099 5013
rect 4465 4951 4486 4970
rect 4993 4951 5019 5010
rect 5062 5004 5099 5010
rect 5599 5011 5608 5031
rect 5628 5011 5636 5031
rect 5599 5001 5636 5011
rect 5695 5031 5782 5041
rect 5695 5011 5704 5031
rect 5724 5011 5782 5031
rect 5695 5002 5782 5011
rect 5695 5001 5732 5002
rect 5407 4951 5444 4960
rect 3119 4946 3219 4950
rect 3119 4942 3181 4946
rect 3119 4916 3126 4942
rect 3152 4920 3181 4942
rect 3207 4920 3219 4946
rect 3152 4916 3219 4920
rect 3119 4913 3219 4916
rect 3287 4913 3322 4950
rect 3384 4947 3743 4950
rect 3384 4942 3606 4947
rect 3384 4918 3397 4942
rect 3421 4923 3606 4942
rect 3630 4923 3743 4947
rect 3421 4918 3743 4923
rect 3384 4914 3743 4918
rect 3810 4942 3959 4950
rect 3810 4922 3821 4942
rect 3841 4922 3959 4942
rect 4465 4933 5019 4951
rect 5065 4940 5102 4942
rect 4993 4932 5019 4933
rect 5062 4932 5102 4940
rect 3810 4915 3959 4922
rect 5062 4920 5074 4932
rect 5053 4915 5074 4920
rect 3810 4914 3851 4915
rect 4469 4914 5074 4915
rect 5092 4914 5102 4932
rect 3134 4861 3171 4862
rect 3230 4861 3267 4862
rect 3286 4861 3322 4913
rect 3341 4861 3378 4862
rect 3034 4852 3172 4861
rect 3034 4832 3143 4852
rect 3163 4832 3172 4852
rect 3034 4825 3172 4832
rect 3230 4852 3378 4861
rect 3230 4832 3239 4852
rect 3259 4832 3349 4852
rect 3369 4832 3378 4852
rect 3034 4823 3130 4825
rect 3230 4822 3378 4832
rect 3437 4852 3474 4862
rect 3549 4861 3586 4862
rect 3530 4859 3586 4861
rect 3437 4832 3445 4852
rect 3465 4832 3474 4852
rect 3286 4821 3322 4822
rect 3134 4762 3171 4763
rect 3437 4762 3474 4832
rect 3499 4852 3586 4859
rect 3499 4849 3557 4852
rect 3499 4829 3504 4849
rect 3525 4832 3557 4849
rect 3577 4832 3586 4852
rect 3525 4829 3586 4832
rect 3499 4822 3586 4829
rect 3645 4852 3682 4862
rect 3645 4832 3653 4852
rect 3673 4832 3682 4852
rect 3499 4821 3530 4822
rect 3133 4761 3474 4762
rect 3058 4756 3474 4761
rect 3058 4736 3061 4756
rect 3081 4736 3474 4756
rect 3645 4761 3682 4832
rect 3712 4861 3743 4914
rect 4469 4905 5102 4914
rect 5405 4933 5416 4951
rect 5434 4933 5444 4951
rect 5751 4949 5782 5002
rect 5812 5031 5849 5102
rect 6020 5107 6413 5127
rect 6433 5107 6436 5127
rect 6020 5102 6436 5107
rect 6655 5121 6693 5130
rect 6020 5101 6361 5102
rect 6655 5101 6664 5121
rect 6684 5101 6693 5121
rect 5964 5041 5995 5042
rect 5812 5011 5821 5031
rect 5841 5011 5849 5031
rect 5812 5001 5849 5011
rect 5908 5034 5995 5041
rect 5908 5031 5969 5034
rect 5908 5011 5917 5031
rect 5937 5014 5969 5031
rect 5990 5014 5995 5034
rect 5937 5011 5995 5014
rect 5908 5004 5995 5011
rect 6020 5031 6057 5101
rect 6323 5100 6360 5101
rect 6655 5093 6693 5101
rect 6759 5125 6844 5131
rect 6869 5130 6906 5131
rect 6759 5105 6767 5125
rect 6787 5105 6844 5125
rect 6759 5097 6844 5105
rect 6868 5121 6906 5130
rect 6868 5101 6877 5121
rect 6897 5101 6906 5121
rect 6759 5096 6795 5097
rect 6868 5093 6906 5101
rect 6972 5125 7057 5131
rect 7077 5130 7114 5131
rect 6972 5105 6980 5125
rect 7000 5124 7057 5125
rect 7000 5105 7029 5124
rect 6972 5104 7029 5105
rect 7050 5104 7057 5124
rect 6972 5097 7057 5104
rect 7076 5121 7114 5130
rect 7076 5101 7085 5121
rect 7105 5101 7114 5121
rect 6972 5096 7008 5097
rect 7076 5093 7114 5101
rect 7180 5125 7324 5131
rect 7180 5105 7188 5125
rect 7208 5124 7296 5125
rect 7208 5105 7241 5124
rect 7264 5105 7296 5124
rect 7316 5105 7324 5125
rect 7180 5097 7324 5105
rect 7180 5096 7216 5097
rect 7288 5096 7324 5097
rect 7390 5130 7427 5131
rect 7390 5129 7428 5130
rect 7390 5121 7454 5129
rect 7390 5101 7399 5121
rect 7419 5107 7454 5121
rect 7474 5107 7477 5127
rect 7419 5102 7477 5107
rect 7419 5101 7454 5102
rect 6656 5064 6693 5093
rect 6657 5062 6693 5064
rect 6869 5062 6906 5093
rect 6172 5041 6208 5042
rect 6020 5011 6029 5031
rect 6049 5011 6057 5031
rect 5908 5002 5964 5004
rect 5908 5001 5945 5002
rect 6020 5001 6057 5011
rect 6116 5031 6264 5041
rect 6657 5040 6906 5062
rect 7077 5061 7114 5093
rect 7390 5089 7454 5101
rect 7494 5063 7521 5241
rect 7353 5061 7521 5063
rect 7077 5050 7521 5061
rect 7584 5061 7614 6062
rect 7584 5056 7616 5061
rect 6364 5038 6460 5040
rect 6116 5011 6125 5031
rect 6145 5011 6235 5031
rect 6255 5011 6264 5031
rect 6116 5002 6264 5011
rect 6322 5031 6460 5038
rect 7077 5035 7523 5050
rect 7353 5034 7523 5035
rect 6322 5011 6331 5031
rect 6351 5011 6460 5031
rect 6322 5002 6460 5011
rect 6116 5001 6153 5002
rect 6172 4950 6208 5002
rect 6227 5001 6264 5002
rect 6323 5001 6360 5002
rect 5643 4948 5684 4949
rect 4469 4898 5101 4905
rect 4469 4896 4531 4898
rect 4047 4886 4215 4887
rect 4469 4886 4491 4896
rect 3762 4861 3799 4862
rect 3712 4852 3799 4861
rect 3712 4832 3770 4852
rect 3790 4832 3799 4852
rect 3712 4822 3799 4832
rect 3858 4852 3895 4862
rect 3858 4832 3866 4852
rect 3886 4832 3895 4852
rect 3712 4821 3743 4822
rect 3858 4761 3895 4832
rect 3645 4737 3895 4761
rect 4047 4860 4491 4886
rect 4047 4858 4215 4860
rect 4047 4680 4074 4858
rect 4114 4820 4178 4832
rect 4454 4828 4491 4860
rect 4662 4859 4911 4881
rect 4662 4828 4699 4859
rect 4875 4857 4911 4859
rect 4875 4828 4912 4857
rect 4114 4819 4149 4820
rect 4091 4814 4149 4819
rect 4091 4794 4094 4814
rect 4114 4800 4149 4814
rect 4169 4800 4178 4820
rect 4114 4792 4178 4800
rect 4140 4791 4178 4792
rect 4141 4790 4178 4791
rect 4244 4824 4280 4825
rect 4352 4824 4388 4825
rect 4244 4816 4388 4824
rect 4244 4796 4252 4816
rect 4272 4796 4301 4816
rect 4244 4795 4301 4796
rect 4323 4796 4360 4816
rect 4380 4796 4388 4816
rect 4323 4795 4388 4796
rect 4244 4790 4388 4795
rect 4454 4820 4492 4828
rect 4560 4824 4596 4825
rect 4454 4800 4463 4820
rect 4483 4800 4492 4820
rect 4454 4791 4492 4800
rect 4511 4817 4596 4824
rect 4511 4797 4518 4817
rect 4539 4816 4596 4817
rect 4539 4797 4568 4816
rect 4511 4796 4568 4797
rect 4588 4796 4596 4816
rect 4454 4790 4491 4791
rect 4511 4790 4596 4796
rect 4662 4820 4700 4828
rect 4773 4824 4809 4825
rect 4662 4800 4671 4820
rect 4691 4800 4700 4820
rect 4662 4791 4700 4800
rect 4724 4816 4809 4824
rect 4724 4796 4781 4816
rect 4801 4796 4809 4816
rect 4662 4790 4699 4791
rect 4724 4790 4809 4796
rect 4875 4820 4913 4828
rect 4875 4800 4884 4820
rect 4904 4800 4913 4820
rect 4875 4791 4913 4800
rect 4875 4790 4912 4791
rect 4298 4769 4334 4790
rect 4724 4769 4755 4790
rect 4131 4765 4231 4769
rect 4131 4761 4193 4765
rect 4131 4735 4138 4761
rect 4164 4739 4193 4761
rect 4219 4739 4231 4765
rect 4164 4735 4231 4739
rect 4131 4732 4231 4735
rect 4299 4732 4334 4769
rect 4396 4766 4755 4769
rect 4396 4761 4618 4766
rect 4396 4737 4409 4761
rect 4433 4742 4618 4761
rect 4642 4742 4755 4766
rect 4433 4737 4755 4742
rect 4396 4733 4755 4737
rect 4822 4761 4971 4769
rect 4822 4741 4833 4761
rect 4853 4741 4971 4761
rect 4822 4734 4971 4741
rect 5062 4749 5101 4898
rect 5405 4784 5444 4933
rect 5535 4941 5684 4948
rect 5535 4921 5653 4941
rect 5673 4921 5684 4941
rect 5535 4913 5684 4921
rect 5751 4945 6110 4949
rect 5751 4940 6073 4945
rect 5751 4916 5864 4940
rect 5888 4921 6073 4940
rect 6097 4921 6110 4945
rect 5888 4916 6110 4921
rect 5751 4913 6110 4916
rect 6172 4913 6207 4950
rect 6275 4947 6375 4950
rect 6275 4943 6342 4947
rect 6275 4917 6287 4943
rect 6313 4921 6342 4943
rect 6368 4921 6375 4947
rect 6313 4917 6375 4921
rect 6275 4913 6375 4917
rect 5751 4892 5782 4913
rect 6172 4892 6208 4913
rect 5594 4891 5631 4892
rect 5593 4882 5631 4891
rect 5593 4862 5602 4882
rect 5622 4862 5631 4882
rect 5593 4854 5631 4862
rect 5697 4886 5782 4892
rect 5807 4891 5844 4892
rect 5697 4866 5705 4886
rect 5725 4866 5782 4886
rect 5697 4858 5782 4866
rect 5806 4882 5844 4891
rect 5806 4862 5815 4882
rect 5835 4862 5844 4882
rect 5697 4857 5733 4858
rect 5806 4854 5844 4862
rect 5910 4886 5995 4892
rect 6015 4891 6052 4892
rect 5910 4866 5918 4886
rect 5938 4885 5995 4886
rect 5938 4866 5967 4885
rect 5910 4865 5967 4866
rect 5988 4865 5995 4885
rect 5910 4858 5995 4865
rect 6014 4882 6052 4891
rect 6014 4862 6023 4882
rect 6043 4862 6052 4882
rect 5910 4857 5946 4858
rect 6014 4854 6052 4862
rect 6118 4887 6262 4892
rect 6118 4886 6183 4887
rect 6118 4866 6126 4886
rect 6146 4866 6183 4886
rect 6205 4886 6262 4887
rect 6205 4866 6234 4886
rect 6254 4866 6262 4886
rect 6118 4858 6262 4866
rect 6118 4857 6154 4858
rect 6226 4857 6262 4858
rect 6328 4891 6365 4892
rect 6328 4890 6366 4891
rect 6328 4882 6392 4890
rect 6328 4862 6337 4882
rect 6357 4868 6392 4882
rect 6412 4868 6415 4888
rect 6357 4863 6415 4868
rect 6357 4862 6392 4863
rect 5594 4825 5631 4854
rect 5595 4823 5631 4825
rect 5807 4823 5844 4854
rect 5595 4801 5844 4823
rect 6015 4822 6052 4854
rect 6328 4850 6392 4862
rect 6432 4824 6459 5002
rect 6291 4822 6459 4824
rect 6015 4796 6459 4822
rect 6611 4921 6861 4945
rect 6611 4850 6648 4921
rect 6763 4860 6794 4861
rect 6611 4830 6620 4850
rect 6640 4830 6648 4850
rect 6611 4820 6648 4830
rect 6707 4850 6794 4860
rect 6707 4830 6716 4850
rect 6736 4830 6794 4850
rect 6707 4821 6794 4830
rect 6707 4820 6744 4821
rect 6015 4786 6037 4796
rect 6291 4795 6459 4796
rect 5975 4784 6037 4786
rect 5405 4777 6037 4784
rect 4822 4733 4863 4734
rect 4146 4680 4183 4681
rect 4242 4680 4279 4681
rect 4298 4680 4334 4732
rect 4353 4680 4390 4681
rect 4046 4671 4184 4680
rect 4046 4651 4155 4671
rect 4175 4651 4184 4671
rect 4046 4644 4184 4651
rect 4242 4671 4390 4680
rect 4242 4651 4251 4671
rect 4271 4651 4361 4671
rect 4381 4651 4390 4671
rect 4046 4642 4142 4644
rect 4242 4641 4390 4651
rect 4449 4671 4486 4681
rect 4561 4680 4598 4681
rect 4542 4678 4598 4680
rect 4449 4651 4457 4671
rect 4477 4651 4486 4671
rect 4298 4640 4334 4641
rect 2211 4632 2242 4635
rect 2740 4635 2908 4636
rect 1040 4608 1178 4617
rect 2740 4609 3184 4635
rect 834 4607 871 4608
rect 890 4556 926 4608
rect 945 4607 982 4608
rect 1041 4607 1078 4608
rect 361 4554 402 4555
rect 253 4547 402 4554
rect 253 4527 371 4547
rect 391 4527 402 4547
rect 253 4519 402 4527
rect 469 4551 828 4555
rect 469 4546 791 4551
rect 469 4522 582 4546
rect 606 4527 791 4546
rect 815 4527 828 4551
rect 606 4522 828 4527
rect 469 4519 828 4522
rect 890 4519 925 4556
rect 993 4553 1093 4556
rect 993 4549 1060 4553
rect 993 4523 1005 4549
rect 1031 4527 1060 4549
rect 1086 4527 1093 4553
rect 1031 4523 1093 4527
rect 993 4519 1093 4523
rect 469 4498 500 4519
rect 890 4498 926 4519
rect 133 4489 170 4498
rect 312 4497 349 4498
rect 133 4471 142 4489
rect 160 4471 170 4489
rect 133 4461 170 4471
rect 134 4426 170 4461
rect 311 4488 349 4497
rect 311 4468 320 4488
rect 340 4468 349 4488
rect 311 4460 349 4468
rect 415 4492 500 4498
rect 525 4497 562 4498
rect 415 4472 423 4492
rect 443 4472 500 4492
rect 415 4464 500 4472
rect 524 4488 562 4497
rect 524 4468 533 4488
rect 553 4468 562 4488
rect 415 4463 451 4464
rect 524 4460 562 4468
rect 628 4492 713 4498
rect 733 4497 770 4498
rect 628 4472 636 4492
rect 656 4491 713 4492
rect 656 4472 685 4491
rect 628 4471 685 4472
rect 706 4471 713 4491
rect 628 4464 713 4471
rect 732 4488 770 4497
rect 732 4468 741 4488
rect 761 4468 770 4488
rect 628 4463 664 4464
rect 732 4460 770 4468
rect 836 4492 980 4498
rect 836 4472 844 4492
rect 864 4491 952 4492
rect 864 4472 892 4491
rect 836 4470 892 4472
rect 914 4472 952 4491
rect 972 4472 980 4492
rect 914 4470 980 4472
rect 836 4464 980 4470
rect 836 4463 872 4464
rect 944 4463 980 4464
rect 1046 4497 1083 4498
rect 1046 4496 1084 4497
rect 1046 4488 1110 4496
rect 1046 4468 1055 4488
rect 1075 4474 1110 4488
rect 1130 4474 1133 4494
rect 1075 4469 1133 4474
rect 1075 4468 1110 4469
rect 312 4431 349 4460
rect 132 4385 170 4426
rect 313 4429 349 4431
rect 525 4429 562 4460
rect 313 4407 562 4429
rect 733 4428 770 4460
rect 1046 4456 1110 4468
rect 1150 4430 1177 4608
rect 1009 4428 1177 4430
rect 2740 4607 2908 4609
rect 2740 4604 2787 4607
rect 2740 4429 2767 4604
rect 2807 4569 2871 4581
rect 3147 4577 3184 4609
rect 3355 4608 3604 4630
rect 3355 4577 3392 4608
rect 3568 4606 3604 4608
rect 3568 4577 3605 4606
rect 4146 4581 4183 4582
rect 4449 4581 4486 4651
rect 4511 4671 4598 4678
rect 4511 4668 4569 4671
rect 4511 4648 4516 4668
rect 4537 4651 4569 4668
rect 4589 4651 4598 4671
rect 4537 4648 4598 4651
rect 4511 4641 4598 4648
rect 4657 4671 4694 4681
rect 4657 4651 4665 4671
rect 4685 4651 4694 4671
rect 4511 4640 4542 4641
rect 4145 4580 4486 4581
rect 2807 4568 2842 4569
rect 2784 4563 2842 4568
rect 2784 4543 2787 4563
rect 2807 4549 2842 4563
rect 2862 4549 2871 4569
rect 2807 4541 2871 4549
rect 2833 4540 2871 4541
rect 2834 4539 2871 4540
rect 2937 4573 2973 4574
rect 3045 4573 3081 4574
rect 2937 4565 3081 4573
rect 2937 4545 2945 4565
rect 2965 4563 3053 4565
rect 2965 4545 2991 4563
rect 2937 4544 2991 4545
rect 3017 4545 3053 4563
rect 3073 4545 3081 4565
rect 3017 4544 3081 4545
rect 2937 4539 3081 4544
rect 3147 4569 3185 4577
rect 3253 4573 3289 4574
rect 3147 4549 3156 4569
rect 3176 4549 3185 4569
rect 3147 4540 3185 4549
rect 3204 4566 3289 4573
rect 3204 4546 3211 4566
rect 3232 4565 3289 4566
rect 3232 4546 3261 4565
rect 3204 4545 3261 4546
rect 3281 4545 3289 4565
rect 3147 4539 3184 4540
rect 3204 4539 3289 4545
rect 3355 4569 3393 4577
rect 3466 4573 3502 4574
rect 3355 4549 3364 4569
rect 3384 4549 3393 4569
rect 3355 4540 3393 4549
rect 3417 4565 3502 4573
rect 3417 4545 3474 4565
rect 3494 4545 3502 4565
rect 3355 4539 3392 4540
rect 3417 4539 3502 4545
rect 3568 4569 3606 4577
rect 3568 4549 3577 4569
rect 3597 4549 3606 4569
rect 4070 4575 4486 4580
rect 4070 4555 4073 4575
rect 4093 4555 4486 4575
rect 4657 4580 4694 4651
rect 4724 4680 4755 4733
rect 5062 4731 5072 4749
rect 5090 4731 5101 4749
rect 5404 4768 6037 4777
rect 6763 4768 6794 4821
rect 6824 4850 6861 4921
rect 7032 4926 7425 4946
rect 7445 4926 7448 4946
rect 7032 4921 7448 4926
rect 7032 4920 7373 4921
rect 6976 4860 7007 4861
rect 6824 4830 6833 4850
rect 6853 4830 6861 4850
rect 6824 4820 6861 4830
rect 6920 4853 7007 4860
rect 6920 4850 6981 4853
rect 6920 4830 6929 4850
rect 6949 4833 6981 4850
rect 7002 4833 7007 4853
rect 6949 4830 7007 4833
rect 6920 4823 7007 4830
rect 7032 4850 7069 4920
rect 7335 4919 7372 4920
rect 7184 4860 7220 4861
rect 7032 4830 7041 4850
rect 7061 4830 7069 4850
rect 6920 4821 6976 4823
rect 6920 4820 6957 4821
rect 7032 4820 7069 4830
rect 7128 4850 7276 4860
rect 7376 4857 7472 4859
rect 7128 4830 7137 4850
rect 7157 4830 7247 4850
rect 7267 4830 7276 4850
rect 7128 4821 7276 4830
rect 7334 4850 7472 4857
rect 7334 4830 7343 4850
rect 7363 4830 7472 4850
rect 7334 4821 7472 4830
rect 7128 4820 7165 4821
rect 7184 4769 7220 4821
rect 7239 4820 7276 4821
rect 7335 4820 7372 4821
rect 5404 4750 5414 4768
rect 5432 4767 6037 4768
rect 6655 4767 6696 4768
rect 5432 4762 5453 4767
rect 5432 4750 5444 4762
rect 6547 4760 6696 4767
rect 5404 4742 5444 4750
rect 5487 4749 5513 4750
rect 5404 4740 5441 4742
rect 5487 4731 6041 4749
rect 6547 4740 6665 4760
rect 6685 4740 6696 4760
rect 6547 4732 6696 4740
rect 6763 4764 7122 4768
rect 6763 4759 7085 4764
rect 6763 4735 6876 4759
rect 6900 4740 7085 4759
rect 7109 4740 7122 4764
rect 6900 4735 7122 4740
rect 6763 4732 7122 4735
rect 7184 4732 7219 4769
rect 7287 4766 7387 4769
rect 7287 4762 7354 4766
rect 7287 4736 7299 4762
rect 7325 4740 7354 4762
rect 7380 4740 7387 4766
rect 7325 4736 7387 4740
rect 7287 4732 7387 4736
rect 5062 4722 5099 4731
rect 4774 4680 4811 4681
rect 4724 4671 4811 4680
rect 4724 4651 4782 4671
rect 4802 4651 4811 4671
rect 4724 4641 4811 4651
rect 4870 4671 4907 4681
rect 4870 4651 4878 4671
rect 4898 4651 4907 4671
rect 5407 4672 5444 4678
rect 5487 4672 5513 4731
rect 6020 4712 6041 4731
rect 5407 4669 5513 4672
rect 5065 4656 5102 4660
rect 4724 4640 4755 4641
rect 4870 4580 4907 4651
rect 4657 4556 4907 4580
rect 5063 4650 5102 4656
rect 5063 4632 5074 4650
rect 5092 4632 5102 4650
rect 5407 4651 5416 4669
rect 5434 4655 5513 4669
rect 5598 4687 5848 4711
rect 5434 4653 5510 4655
rect 5434 4651 5444 4653
rect 5407 4641 5444 4651
rect 5063 4623 5102 4632
rect 3568 4540 3606 4549
rect 3568 4539 3605 4540
rect 2991 4518 3027 4539
rect 3417 4518 3448 4539
rect 4449 4532 4486 4555
rect 5063 4545 5098 4623
rect 5412 4576 5443 4641
rect 5598 4616 5635 4687
rect 5750 4626 5781 4627
rect 5598 4596 5607 4616
rect 5627 4596 5635 4616
rect 5598 4586 5635 4596
rect 5694 4616 5781 4626
rect 5694 4596 5703 4616
rect 5723 4596 5781 4616
rect 5694 4587 5781 4596
rect 5694 4586 5731 4587
rect 5060 4535 5098 4545
rect 5411 4567 5448 4576
rect 5411 4549 5421 4567
rect 5439 4549 5448 4567
rect 5411 4539 5448 4549
rect 4449 4531 4619 4532
rect 5060 4531 5070 4535
rect 2824 4514 2924 4518
rect 2824 4510 2886 4514
rect 2824 4484 2831 4510
rect 2857 4488 2886 4510
rect 2912 4488 2924 4514
rect 2857 4484 2924 4488
rect 2824 4481 2924 4484
rect 2992 4481 3027 4518
rect 3089 4515 3448 4518
rect 3089 4510 3311 4515
rect 3089 4486 3102 4510
rect 3126 4491 3311 4510
rect 3335 4491 3448 4515
rect 3126 4486 3448 4491
rect 3089 4482 3448 4486
rect 3515 4510 3664 4518
rect 4449 4517 5070 4531
rect 5088 4517 5098 4535
rect 5750 4534 5781 4587
rect 5811 4616 5848 4687
rect 6019 4692 6412 4712
rect 6432 4692 6435 4712
rect 6763 4711 6794 4732
rect 7184 4711 7220 4732
rect 6606 4710 6643 4711
rect 6019 4687 6435 4692
rect 6605 4701 6643 4710
rect 6019 4686 6360 4687
rect 5963 4626 5994 4627
rect 5811 4596 5820 4616
rect 5840 4596 5848 4616
rect 5811 4586 5848 4596
rect 5907 4619 5994 4626
rect 5907 4616 5968 4619
rect 5907 4596 5916 4616
rect 5936 4599 5968 4616
rect 5989 4599 5994 4619
rect 5936 4596 5994 4599
rect 5907 4589 5994 4596
rect 6019 4616 6056 4686
rect 6322 4685 6359 4686
rect 6605 4681 6614 4701
rect 6634 4681 6643 4701
rect 6605 4673 6643 4681
rect 6709 4705 6794 4711
rect 6819 4710 6856 4711
rect 6709 4685 6717 4705
rect 6737 4685 6794 4705
rect 6709 4677 6794 4685
rect 6818 4701 6856 4710
rect 6818 4681 6827 4701
rect 6847 4681 6856 4701
rect 6709 4676 6745 4677
rect 6818 4673 6856 4681
rect 6922 4705 7007 4711
rect 7027 4710 7064 4711
rect 6922 4685 6930 4705
rect 6950 4704 7007 4705
rect 6950 4685 6979 4704
rect 6922 4684 6979 4685
rect 7000 4684 7007 4704
rect 6922 4677 7007 4684
rect 7026 4701 7064 4710
rect 7026 4681 7035 4701
rect 7055 4681 7064 4701
rect 6922 4676 6958 4677
rect 7026 4673 7064 4681
rect 7130 4706 7274 4711
rect 7130 4705 7189 4706
rect 7130 4685 7138 4705
rect 7158 4686 7189 4705
rect 7213 4705 7274 4706
rect 7213 4686 7246 4705
rect 7158 4685 7246 4686
rect 7266 4685 7274 4705
rect 7130 4677 7274 4685
rect 7130 4676 7166 4677
rect 7238 4676 7274 4677
rect 7340 4710 7377 4711
rect 7340 4709 7378 4710
rect 7340 4701 7404 4709
rect 7340 4681 7349 4701
rect 7369 4687 7404 4701
rect 7424 4687 7427 4707
rect 7369 4682 7427 4687
rect 7369 4681 7404 4682
rect 6606 4644 6643 4673
rect 6607 4642 6643 4644
rect 6819 4642 6856 4673
rect 6171 4626 6207 4627
rect 6019 4596 6028 4616
rect 6048 4596 6056 4616
rect 5907 4587 5963 4589
rect 5907 4586 5944 4587
rect 6019 4586 6056 4596
rect 6115 4616 6263 4626
rect 6363 4623 6459 4625
rect 6115 4596 6124 4616
rect 6144 4596 6234 4616
rect 6254 4596 6263 4616
rect 6115 4587 6263 4596
rect 6321 4616 6459 4623
rect 6607 4620 6856 4642
rect 7027 4641 7064 4673
rect 7340 4669 7404 4681
rect 7444 4643 7471 4821
rect 7303 4641 7471 4643
rect 7027 4637 7471 4641
rect 6321 4596 6330 4616
rect 6350 4596 6459 4616
rect 7027 4618 7076 4637
rect 7096 4618 7471 4637
rect 7027 4615 7471 4618
rect 7303 4614 7471 4615
rect 7492 4640 7523 5034
rect 7584 5038 7589 5056
rect 7609 5038 7616 5056
rect 7584 5033 7616 5038
rect 7587 5031 7616 5033
rect 7492 4614 7497 4640
rect 7516 4614 7523 4640
rect 8030 4615 8068 6446
rect 8096 6333 8123 6511
rect 8163 6473 8227 6485
rect 8503 6481 8540 6513
rect 8711 6512 8960 6534
rect 9415 6520 9452 6521
rect 9718 6520 9755 6590
rect 9780 6610 9867 6617
rect 9780 6607 9838 6610
rect 9780 6587 9785 6607
rect 9806 6590 9838 6607
rect 9858 6590 9867 6610
rect 9806 6587 9867 6590
rect 9780 6580 9867 6587
rect 9926 6610 9963 6620
rect 9926 6590 9934 6610
rect 9954 6590 9963 6610
rect 9780 6579 9811 6580
rect 9414 6519 9755 6520
rect 8711 6481 8748 6512
rect 8924 6510 8960 6512
rect 9339 6514 9755 6519
rect 8924 6481 8961 6510
rect 9339 6494 9342 6514
rect 9362 6494 9755 6514
rect 9926 6519 9963 6590
rect 9993 6619 10024 6672
rect 10331 6670 10341 6688
rect 10359 6670 10370 6688
rect 10331 6661 10368 6670
rect 10043 6619 10080 6620
rect 9993 6610 10080 6619
rect 9993 6590 10051 6610
rect 10071 6590 10080 6610
rect 9993 6580 10080 6590
rect 10139 6610 10176 6620
rect 10139 6590 10147 6610
rect 10167 6590 10176 6610
rect 10334 6595 10371 6599
rect 9993 6579 10024 6580
rect 10139 6519 10176 6590
rect 9926 6495 10176 6519
rect 10332 6589 10371 6595
rect 10332 6571 10343 6589
rect 10361 6571 10371 6589
rect 10332 6562 10371 6571
rect 8163 6472 8198 6473
rect 8140 6467 8198 6472
rect 8140 6447 8143 6467
rect 8163 6453 8198 6467
rect 8218 6453 8227 6473
rect 8163 6445 8227 6453
rect 8189 6444 8227 6445
rect 8190 6443 8227 6444
rect 8293 6477 8329 6478
rect 8401 6477 8437 6478
rect 8293 6469 8437 6477
rect 8293 6449 8301 6469
rect 8321 6468 8409 6469
rect 8321 6449 8350 6468
rect 8373 6449 8409 6468
rect 8429 6449 8437 6469
rect 8293 6443 8437 6449
rect 8503 6473 8541 6481
rect 8609 6477 8645 6478
rect 8503 6453 8512 6473
rect 8532 6453 8541 6473
rect 8503 6444 8541 6453
rect 8560 6470 8645 6477
rect 8560 6450 8567 6470
rect 8588 6469 8645 6470
rect 8588 6450 8617 6469
rect 8560 6449 8617 6450
rect 8637 6449 8645 6469
rect 8503 6443 8540 6444
rect 8560 6443 8645 6449
rect 8711 6473 8749 6481
rect 8822 6477 8858 6478
rect 8711 6453 8720 6473
rect 8740 6453 8749 6473
rect 8711 6444 8749 6453
rect 8773 6469 8858 6477
rect 8773 6449 8830 6469
rect 8850 6449 8858 6469
rect 8711 6443 8748 6444
rect 8773 6443 8858 6449
rect 8924 6473 8962 6481
rect 8924 6453 8933 6473
rect 8953 6453 8962 6473
rect 8924 6444 8962 6453
rect 9718 6471 9755 6494
rect 10332 6484 10367 6562
rect 10329 6474 10367 6484
rect 9718 6470 9888 6471
rect 10329 6470 10339 6474
rect 9718 6456 10339 6470
rect 10357 6456 10367 6474
rect 9718 6450 10367 6456
rect 9718 6449 10366 6450
rect 10329 6447 10366 6449
rect 8924 6443 8961 6444
rect 8347 6422 8383 6443
rect 8773 6422 8804 6443
rect 8180 6418 8280 6422
rect 8180 6414 8242 6418
rect 8180 6388 8187 6414
rect 8213 6392 8242 6414
rect 8268 6392 8280 6418
rect 8213 6388 8280 6392
rect 8180 6385 8280 6388
rect 8348 6385 8383 6422
rect 8445 6419 8804 6422
rect 8445 6414 8667 6419
rect 8445 6390 8458 6414
rect 8482 6395 8667 6414
rect 8691 6395 8804 6419
rect 8482 6390 8804 6395
rect 8445 6386 8804 6390
rect 8871 6414 9020 6422
rect 8871 6394 8882 6414
rect 8902 6394 9020 6414
rect 8871 6387 9020 6394
rect 8871 6386 8912 6387
rect 8195 6333 8232 6334
rect 8291 6333 8328 6334
rect 8347 6333 8383 6385
rect 8402 6333 8439 6334
rect 8095 6324 8233 6333
rect 8095 6304 8204 6324
rect 8224 6304 8233 6324
rect 8095 6297 8233 6304
rect 8291 6324 8439 6333
rect 8291 6304 8300 6324
rect 8320 6304 8410 6324
rect 8430 6304 8439 6324
rect 8095 6295 8191 6297
rect 8291 6294 8439 6304
rect 8498 6324 8535 6334
rect 8610 6333 8647 6334
rect 8591 6331 8647 6333
rect 8498 6304 8506 6324
rect 8526 6304 8535 6324
rect 8347 6293 8383 6294
rect 8195 6234 8232 6235
rect 8498 6234 8535 6304
rect 8560 6324 8647 6331
rect 8560 6321 8618 6324
rect 8560 6301 8565 6321
rect 8586 6304 8618 6321
rect 8638 6304 8647 6324
rect 8586 6301 8647 6304
rect 8560 6294 8647 6301
rect 8706 6324 8743 6334
rect 8706 6304 8714 6324
rect 8734 6304 8743 6324
rect 8560 6293 8591 6294
rect 8194 6233 8535 6234
rect 8119 6228 8535 6233
rect 8119 6208 8122 6228
rect 8142 6208 8535 6228
rect 8706 6233 8743 6304
rect 8773 6333 8804 6386
rect 10332 6375 10369 6385
rect 10332 6357 10341 6375
rect 10359 6357 10369 6375
rect 10332 6348 10369 6357
rect 8823 6333 8860 6334
rect 8773 6324 8860 6333
rect 8773 6304 8831 6324
rect 8851 6304 8860 6324
rect 8773 6294 8860 6304
rect 8919 6324 8956 6334
rect 8919 6304 8927 6324
rect 8947 6304 8956 6324
rect 8773 6293 8804 6294
rect 8919 6233 8956 6304
rect 10332 6302 10367 6348
rect 10331 6296 10369 6302
rect 9742 6278 10369 6296
rect 8706 6209 8956 6233
rect 9324 6261 9492 6262
rect 9743 6261 9767 6278
rect 9324 6235 9768 6261
rect 9324 6233 9492 6235
rect 9324 6055 9351 6233
rect 9391 6195 9455 6207
rect 9731 6203 9768 6235
rect 9939 6234 10188 6256
rect 9939 6203 9976 6234
rect 10152 6232 10188 6234
rect 10331 6237 10369 6278
rect 10152 6203 10189 6232
rect 9391 6194 9426 6195
rect 9368 6189 9426 6194
rect 9368 6169 9371 6189
rect 9391 6175 9426 6189
rect 9446 6175 9455 6195
rect 9391 6167 9455 6175
rect 9417 6166 9455 6167
rect 9418 6165 9455 6166
rect 9521 6199 9557 6200
rect 9629 6199 9665 6200
rect 9521 6193 9665 6199
rect 9521 6191 9587 6193
rect 9521 6171 9529 6191
rect 9549 6172 9587 6191
rect 9609 6191 9665 6193
rect 9609 6172 9637 6191
rect 9549 6171 9637 6172
rect 9657 6171 9665 6191
rect 9521 6165 9665 6171
rect 9731 6195 9769 6203
rect 9837 6199 9873 6200
rect 9731 6175 9740 6195
rect 9760 6175 9769 6195
rect 9731 6166 9769 6175
rect 9788 6192 9873 6199
rect 9788 6172 9795 6192
rect 9816 6191 9873 6192
rect 9816 6172 9845 6191
rect 9788 6171 9845 6172
rect 9865 6171 9873 6191
rect 9731 6165 9768 6166
rect 9788 6165 9873 6171
rect 9939 6195 9977 6203
rect 10050 6199 10086 6200
rect 9939 6175 9948 6195
rect 9968 6175 9977 6195
rect 9939 6166 9977 6175
rect 10001 6191 10086 6199
rect 10001 6171 10058 6191
rect 10078 6171 10086 6191
rect 9939 6165 9976 6166
rect 10001 6165 10086 6171
rect 10152 6195 10190 6203
rect 10152 6175 10161 6195
rect 10181 6175 10190 6195
rect 10152 6166 10190 6175
rect 10331 6202 10367 6237
rect 10331 6192 10368 6202
rect 10331 6174 10341 6192
rect 10359 6174 10368 6192
rect 10152 6165 10189 6166
rect 10331 6165 10368 6174
rect 9575 6144 9611 6165
rect 10001 6144 10032 6165
rect 9408 6140 9508 6144
rect 9408 6136 9470 6140
rect 9408 6110 9415 6136
rect 9441 6114 9470 6136
rect 9496 6114 9508 6140
rect 9441 6110 9508 6114
rect 9408 6107 9508 6110
rect 9576 6107 9611 6144
rect 9673 6141 10032 6144
rect 9673 6136 9895 6141
rect 9673 6112 9686 6136
rect 9710 6117 9895 6136
rect 9919 6117 10032 6141
rect 9710 6112 10032 6117
rect 9673 6108 10032 6112
rect 10099 6136 10248 6144
rect 10099 6116 10110 6136
rect 10130 6116 10248 6136
rect 10099 6109 10248 6116
rect 10099 6108 10140 6109
rect 9423 6055 9460 6056
rect 9519 6055 9556 6056
rect 9575 6055 9611 6107
rect 9630 6055 9667 6056
rect 9323 6046 9461 6055
rect 8259 6028 8290 6031
rect 8259 6002 8266 6028
rect 8285 6002 8290 6028
rect 8259 5608 8290 6002
rect 8311 6027 8479 6028
rect 8311 6024 8755 6027
rect 8311 6005 8686 6024
rect 8706 6005 8755 6024
rect 9323 6026 9432 6046
rect 9452 6026 9461 6046
rect 8311 6001 8755 6005
rect 8311 5999 8479 6001
rect 8311 5821 8338 5999
rect 8378 5961 8442 5973
rect 8718 5969 8755 6001
rect 8926 6000 9175 6022
rect 9323 6019 9461 6026
rect 9519 6046 9667 6055
rect 9519 6026 9528 6046
rect 9548 6026 9638 6046
rect 9658 6026 9667 6046
rect 9323 6017 9419 6019
rect 9519 6016 9667 6026
rect 9726 6046 9763 6056
rect 9838 6055 9875 6056
rect 9819 6053 9875 6055
rect 9726 6026 9734 6046
rect 9754 6026 9763 6046
rect 9575 6015 9611 6016
rect 8926 5969 8963 6000
rect 9139 5998 9175 6000
rect 9139 5969 9176 5998
rect 8378 5960 8413 5961
rect 8355 5955 8413 5960
rect 8355 5935 8358 5955
rect 8378 5941 8413 5955
rect 8433 5941 8442 5961
rect 8378 5933 8442 5941
rect 8404 5932 8442 5933
rect 8405 5931 8442 5932
rect 8508 5965 8544 5966
rect 8616 5965 8652 5966
rect 8508 5957 8652 5965
rect 8508 5937 8516 5957
rect 8536 5956 8624 5957
rect 8536 5937 8569 5956
rect 8508 5936 8569 5937
rect 8593 5937 8624 5956
rect 8644 5937 8652 5957
rect 8593 5936 8652 5937
rect 8508 5931 8652 5936
rect 8718 5961 8756 5969
rect 8824 5965 8860 5966
rect 8718 5941 8727 5961
rect 8747 5941 8756 5961
rect 8718 5932 8756 5941
rect 8775 5958 8860 5965
rect 8775 5938 8782 5958
rect 8803 5957 8860 5958
rect 8803 5938 8832 5957
rect 8775 5937 8832 5938
rect 8852 5937 8860 5957
rect 8718 5931 8755 5932
rect 8775 5931 8860 5937
rect 8926 5961 8964 5969
rect 9037 5965 9073 5966
rect 8926 5941 8935 5961
rect 8955 5941 8964 5961
rect 8926 5932 8964 5941
rect 8988 5957 9073 5965
rect 8988 5937 9045 5957
rect 9065 5937 9073 5957
rect 8926 5931 8963 5932
rect 8988 5931 9073 5937
rect 9139 5961 9177 5969
rect 9139 5941 9148 5961
rect 9168 5941 9177 5961
rect 9423 5956 9460 5957
rect 9726 5956 9763 6026
rect 9788 6046 9875 6053
rect 9788 6043 9846 6046
rect 9788 6023 9793 6043
rect 9814 6026 9846 6043
rect 9866 6026 9875 6046
rect 9814 6023 9875 6026
rect 9788 6016 9875 6023
rect 9934 6046 9971 6056
rect 9934 6026 9942 6046
rect 9962 6026 9971 6046
rect 9788 6015 9819 6016
rect 9422 5955 9763 5956
rect 9139 5932 9177 5941
rect 9347 5950 9763 5955
rect 9139 5931 9176 5932
rect 8562 5910 8598 5931
rect 8988 5910 9019 5931
rect 9347 5930 9350 5950
rect 9370 5930 9763 5950
rect 9934 5955 9971 6026
rect 10001 6055 10032 6108
rect 10334 6093 10371 6103
rect 10334 6075 10343 6093
rect 10361 6075 10371 6093
rect 10334 6066 10371 6075
rect 10051 6055 10088 6056
rect 10001 6046 10088 6055
rect 10001 6026 10059 6046
rect 10079 6026 10088 6046
rect 10001 6016 10088 6026
rect 10147 6046 10184 6056
rect 10147 6026 10155 6046
rect 10175 6026 10184 6046
rect 10001 6015 10032 6016
rect 10147 5955 10184 6026
rect 10339 6001 10370 6066
rect 10338 5991 10375 6001
rect 10338 5989 10348 5991
rect 10272 5987 10348 5989
rect 9934 5931 10184 5955
rect 10269 5973 10348 5987
rect 10366 5973 10375 5991
rect 10269 5970 10375 5973
rect 9741 5911 9762 5930
rect 10269 5911 10295 5970
rect 10338 5964 10375 5970
rect 8395 5906 8495 5910
rect 8395 5902 8457 5906
rect 8395 5876 8402 5902
rect 8428 5880 8457 5902
rect 8483 5880 8495 5906
rect 8428 5876 8495 5880
rect 8395 5873 8495 5876
rect 8563 5873 8598 5910
rect 8660 5907 9019 5910
rect 8660 5902 8882 5907
rect 8660 5878 8673 5902
rect 8697 5883 8882 5902
rect 8906 5883 9019 5907
rect 8697 5878 9019 5883
rect 8660 5874 9019 5878
rect 9086 5902 9235 5910
rect 9086 5882 9097 5902
rect 9117 5882 9235 5902
rect 9741 5893 10295 5911
rect 10341 5900 10378 5902
rect 10269 5892 10295 5893
rect 10338 5892 10378 5900
rect 9086 5875 9235 5882
rect 10338 5880 10350 5892
rect 10329 5875 10350 5880
rect 9086 5874 9127 5875
rect 9745 5874 10350 5875
rect 10368 5874 10378 5892
rect 8410 5821 8447 5822
rect 8506 5821 8543 5822
rect 8562 5821 8598 5873
rect 8617 5821 8654 5822
rect 8310 5812 8448 5821
rect 8310 5792 8419 5812
rect 8439 5792 8448 5812
rect 8310 5785 8448 5792
rect 8506 5812 8654 5821
rect 8506 5792 8515 5812
rect 8535 5792 8625 5812
rect 8645 5792 8654 5812
rect 8310 5783 8406 5785
rect 8506 5782 8654 5792
rect 8713 5812 8750 5822
rect 8825 5821 8862 5822
rect 8806 5819 8862 5821
rect 8713 5792 8721 5812
rect 8741 5792 8750 5812
rect 8562 5781 8598 5782
rect 8410 5722 8447 5723
rect 8713 5722 8750 5792
rect 8775 5812 8862 5819
rect 8775 5809 8833 5812
rect 8775 5789 8780 5809
rect 8801 5792 8833 5809
rect 8853 5792 8862 5812
rect 8801 5789 8862 5792
rect 8775 5782 8862 5789
rect 8921 5812 8958 5822
rect 8921 5792 8929 5812
rect 8949 5792 8958 5812
rect 8775 5781 8806 5782
rect 8409 5721 8750 5722
rect 8334 5716 8750 5721
rect 8334 5696 8337 5716
rect 8357 5696 8750 5716
rect 8921 5721 8958 5792
rect 8988 5821 9019 5874
rect 9745 5865 10378 5874
rect 9745 5858 10377 5865
rect 9745 5856 9807 5858
rect 9323 5846 9491 5847
rect 9745 5846 9767 5856
rect 9038 5821 9075 5822
rect 8988 5812 9075 5821
rect 8988 5792 9046 5812
rect 9066 5792 9075 5812
rect 8988 5782 9075 5792
rect 9134 5812 9171 5822
rect 9134 5792 9142 5812
rect 9162 5792 9171 5812
rect 8988 5781 9019 5782
rect 9134 5721 9171 5792
rect 8921 5697 9171 5721
rect 9323 5820 9767 5846
rect 9323 5818 9491 5820
rect 9323 5640 9350 5818
rect 9390 5780 9454 5792
rect 9730 5788 9767 5820
rect 9938 5819 10187 5841
rect 9938 5788 9975 5819
rect 10151 5817 10187 5819
rect 10151 5788 10188 5817
rect 9390 5779 9425 5780
rect 9367 5774 9425 5779
rect 9367 5754 9370 5774
rect 9390 5760 9425 5774
rect 9445 5760 9454 5780
rect 9390 5752 9454 5760
rect 9416 5751 9454 5752
rect 9417 5750 9454 5751
rect 9520 5784 9556 5785
rect 9628 5784 9664 5785
rect 9520 5776 9664 5784
rect 9520 5756 9528 5776
rect 9548 5756 9577 5776
rect 9520 5755 9577 5756
rect 9599 5756 9636 5776
rect 9656 5756 9664 5776
rect 9599 5755 9664 5756
rect 9520 5750 9664 5755
rect 9730 5780 9768 5788
rect 9836 5784 9872 5785
rect 9730 5760 9739 5780
rect 9759 5760 9768 5780
rect 9730 5751 9768 5760
rect 9787 5777 9872 5784
rect 9787 5757 9794 5777
rect 9815 5776 9872 5777
rect 9815 5757 9844 5776
rect 9787 5756 9844 5757
rect 9864 5756 9872 5776
rect 9730 5750 9767 5751
rect 9787 5750 9872 5756
rect 9938 5780 9976 5788
rect 10049 5784 10085 5785
rect 9938 5760 9947 5780
rect 9967 5760 9976 5780
rect 9938 5751 9976 5760
rect 10000 5776 10085 5784
rect 10000 5756 10057 5776
rect 10077 5756 10085 5776
rect 9938 5750 9975 5751
rect 10000 5750 10085 5756
rect 10151 5780 10189 5788
rect 10151 5760 10160 5780
rect 10180 5760 10189 5780
rect 10151 5751 10189 5760
rect 10151 5750 10188 5751
rect 9574 5729 9610 5750
rect 10000 5729 10031 5750
rect 9407 5725 9507 5729
rect 9407 5721 9469 5725
rect 9407 5695 9414 5721
rect 9440 5699 9469 5721
rect 9495 5699 9507 5725
rect 9440 5695 9507 5699
rect 9407 5692 9507 5695
rect 9575 5692 9610 5729
rect 9672 5726 10031 5729
rect 9672 5721 9894 5726
rect 9672 5697 9685 5721
rect 9709 5702 9894 5721
rect 9918 5702 10031 5726
rect 9709 5697 10031 5702
rect 9672 5693 10031 5697
rect 10098 5721 10247 5729
rect 10098 5701 10109 5721
rect 10129 5701 10247 5721
rect 10098 5694 10247 5701
rect 10338 5709 10377 5858
rect 10098 5693 10139 5694
rect 9422 5640 9459 5641
rect 9518 5640 9555 5641
rect 9574 5640 9610 5692
rect 9629 5640 9666 5641
rect 9322 5631 9460 5640
rect 9322 5611 9431 5631
rect 9451 5611 9460 5631
rect 8259 5607 8429 5608
rect 8259 5592 8705 5607
rect 9322 5604 9460 5611
rect 9518 5631 9666 5640
rect 9518 5611 9527 5631
rect 9547 5611 9637 5631
rect 9657 5611 9666 5631
rect 9322 5602 9418 5604
rect 8261 5581 8705 5592
rect 8261 5579 8429 5581
rect 8261 5401 8288 5579
rect 8328 5541 8392 5553
rect 8668 5549 8705 5581
rect 8876 5580 9125 5602
rect 9518 5601 9666 5611
rect 9725 5631 9762 5641
rect 9837 5640 9874 5641
rect 9818 5638 9874 5640
rect 9725 5611 9733 5631
rect 9753 5611 9762 5631
rect 9574 5600 9610 5601
rect 8876 5549 8913 5580
rect 9089 5578 9125 5580
rect 9089 5549 9126 5578
rect 8328 5540 8363 5541
rect 8305 5535 8363 5540
rect 8305 5515 8308 5535
rect 8328 5521 8363 5535
rect 8383 5521 8392 5541
rect 8328 5513 8392 5521
rect 8354 5512 8392 5513
rect 8355 5511 8392 5512
rect 8458 5545 8494 5546
rect 8566 5545 8602 5546
rect 8458 5537 8602 5545
rect 8458 5517 8466 5537
rect 8486 5536 8574 5537
rect 8486 5519 8514 5536
rect 8538 5519 8574 5536
rect 8486 5517 8574 5519
rect 8594 5517 8602 5537
rect 8458 5511 8602 5517
rect 8668 5541 8706 5549
rect 8774 5545 8810 5546
rect 8668 5521 8677 5541
rect 8697 5521 8706 5541
rect 8668 5512 8706 5521
rect 8725 5538 8810 5545
rect 8725 5518 8732 5538
rect 8753 5537 8810 5538
rect 8753 5518 8782 5537
rect 8725 5517 8782 5518
rect 8802 5517 8810 5537
rect 8668 5511 8705 5512
rect 8725 5511 8810 5517
rect 8876 5541 8914 5549
rect 8987 5545 9023 5546
rect 8876 5521 8885 5541
rect 8905 5521 8914 5541
rect 8876 5512 8914 5521
rect 8938 5537 9023 5545
rect 8938 5517 8995 5537
rect 9015 5517 9023 5537
rect 8876 5511 8913 5512
rect 8938 5511 9023 5517
rect 9089 5541 9127 5549
rect 9422 5541 9459 5542
rect 9725 5541 9762 5611
rect 9787 5631 9874 5638
rect 9787 5628 9845 5631
rect 9787 5608 9792 5628
rect 9813 5611 9845 5628
rect 9865 5611 9874 5631
rect 9813 5608 9874 5611
rect 9787 5601 9874 5608
rect 9933 5631 9970 5641
rect 9933 5611 9941 5631
rect 9961 5611 9970 5631
rect 9787 5600 9818 5601
rect 9089 5521 9098 5541
rect 9118 5521 9127 5541
rect 9421 5540 9762 5541
rect 9089 5512 9127 5521
rect 9346 5535 9762 5540
rect 9346 5515 9349 5535
rect 9369 5515 9762 5535
rect 9933 5540 9970 5611
rect 10000 5640 10031 5693
rect 10338 5691 10348 5709
rect 10366 5691 10377 5709
rect 10338 5682 10375 5691
rect 10050 5640 10087 5641
rect 10000 5631 10087 5640
rect 10000 5611 10058 5631
rect 10078 5611 10087 5631
rect 10000 5601 10087 5611
rect 10146 5631 10183 5641
rect 10146 5611 10154 5631
rect 10174 5611 10183 5631
rect 10341 5616 10378 5620
rect 10000 5600 10031 5601
rect 10146 5540 10183 5611
rect 9933 5516 10183 5540
rect 10339 5610 10378 5616
rect 10339 5592 10350 5610
rect 10368 5592 10378 5610
rect 10339 5583 10378 5592
rect 9089 5511 9126 5512
rect 8512 5490 8548 5511
rect 8938 5490 8969 5511
rect 9725 5492 9762 5515
rect 10339 5505 10374 5583
rect 10336 5495 10374 5505
rect 9725 5491 9895 5492
rect 10336 5491 10346 5495
rect 8345 5486 8445 5490
rect 8345 5482 8407 5486
rect 8345 5456 8352 5482
rect 8378 5460 8407 5482
rect 8433 5460 8445 5486
rect 8378 5456 8445 5460
rect 8345 5453 8445 5456
rect 8513 5453 8548 5490
rect 8610 5487 8969 5490
rect 8610 5482 8832 5487
rect 8610 5458 8623 5482
rect 8647 5463 8832 5482
rect 8856 5463 8969 5487
rect 8647 5458 8969 5463
rect 8610 5454 8969 5458
rect 9036 5482 9185 5490
rect 9036 5462 9047 5482
rect 9067 5462 9185 5482
rect 9725 5477 10346 5491
rect 10364 5477 10374 5495
rect 9725 5471 10374 5477
rect 9725 5470 10373 5471
rect 10336 5468 10373 5470
rect 9036 5455 9185 5462
rect 9036 5454 9077 5455
rect 8360 5401 8397 5402
rect 8456 5401 8493 5402
rect 8512 5401 8548 5453
rect 8567 5401 8604 5402
rect 8260 5392 8398 5401
rect 8260 5372 8369 5392
rect 8389 5372 8398 5392
rect 8260 5365 8398 5372
rect 8456 5392 8604 5401
rect 8456 5372 8465 5392
rect 8485 5372 8575 5392
rect 8595 5372 8604 5392
rect 8260 5363 8356 5365
rect 8456 5362 8604 5372
rect 8663 5392 8700 5402
rect 8775 5401 8812 5402
rect 8756 5399 8812 5401
rect 8663 5372 8671 5392
rect 8691 5372 8700 5392
rect 8512 5361 8548 5362
rect 8360 5302 8397 5303
rect 8663 5302 8700 5372
rect 8725 5392 8812 5399
rect 8725 5389 8783 5392
rect 8725 5369 8730 5389
rect 8751 5372 8783 5389
rect 8803 5372 8812 5392
rect 8751 5369 8812 5372
rect 8725 5362 8812 5369
rect 8871 5392 8908 5402
rect 8871 5372 8879 5392
rect 8899 5372 8908 5392
rect 8725 5361 8756 5362
rect 8359 5301 8700 5302
rect 8284 5296 8700 5301
rect 8284 5276 8287 5296
rect 8307 5276 8700 5296
rect 8871 5301 8908 5372
rect 8938 5401 8969 5454
rect 8988 5401 9025 5402
rect 8938 5392 9025 5401
rect 8938 5372 8996 5392
rect 9016 5372 9025 5392
rect 8938 5362 9025 5372
rect 9084 5392 9121 5402
rect 9084 5372 9092 5392
rect 9112 5372 9121 5392
rect 8938 5361 8969 5362
rect 9084 5301 9121 5372
rect 10339 5396 10376 5406
rect 10339 5378 10348 5396
rect 10366 5378 10376 5396
rect 10339 5369 10376 5378
rect 10339 5345 10374 5369
rect 10337 5321 10374 5345
rect 10336 5315 10374 5321
rect 8871 5277 9121 5301
rect 9747 5297 10374 5315
rect 9329 5280 9497 5281
rect 9748 5280 9772 5297
rect 9329 5254 9773 5280
rect 9329 5252 9497 5254
rect 9329 5074 9356 5252
rect 9396 5214 9460 5226
rect 9736 5222 9773 5254
rect 9944 5253 10193 5275
rect 9944 5222 9981 5253
rect 10157 5251 10193 5253
rect 10336 5256 10374 5297
rect 10157 5222 10194 5251
rect 9396 5213 9431 5214
rect 9373 5208 9431 5213
rect 9373 5188 9376 5208
rect 9396 5194 9431 5208
rect 9451 5194 9460 5214
rect 9396 5186 9460 5194
rect 9422 5185 9460 5186
rect 9423 5184 9460 5185
rect 9526 5218 9562 5219
rect 9634 5218 9670 5219
rect 9526 5212 9670 5218
rect 9526 5210 9592 5212
rect 9526 5190 9534 5210
rect 9554 5191 9592 5210
rect 9614 5210 9670 5212
rect 9614 5191 9642 5210
rect 9554 5190 9642 5191
rect 9662 5190 9670 5210
rect 9526 5184 9670 5190
rect 9736 5214 9774 5222
rect 9842 5218 9878 5219
rect 9736 5194 9745 5214
rect 9765 5194 9774 5214
rect 9736 5185 9774 5194
rect 9793 5211 9878 5218
rect 9793 5191 9800 5211
rect 9821 5210 9878 5211
rect 9821 5191 9850 5210
rect 9793 5190 9850 5191
rect 9870 5190 9878 5210
rect 9736 5184 9773 5185
rect 9793 5184 9878 5190
rect 9944 5214 9982 5222
rect 10055 5218 10091 5219
rect 9944 5194 9953 5214
rect 9973 5194 9982 5214
rect 9944 5185 9982 5194
rect 10006 5210 10091 5218
rect 10006 5190 10063 5210
rect 10083 5190 10091 5210
rect 9944 5184 9981 5185
rect 10006 5184 10091 5190
rect 10157 5214 10195 5222
rect 10157 5194 10166 5214
rect 10186 5194 10195 5214
rect 10157 5185 10195 5194
rect 10336 5221 10372 5256
rect 10336 5211 10373 5221
rect 10336 5193 10346 5211
rect 10364 5193 10373 5211
rect 10157 5184 10194 5185
rect 10336 5184 10373 5193
rect 9580 5163 9616 5184
rect 10006 5163 10037 5184
rect 9413 5159 9513 5163
rect 9413 5155 9475 5159
rect 9413 5129 9420 5155
rect 9446 5133 9475 5155
rect 9501 5133 9513 5159
rect 9446 5129 9513 5133
rect 9413 5126 9513 5129
rect 9581 5126 9616 5163
rect 9678 5160 10037 5163
rect 9678 5155 9900 5160
rect 9678 5131 9691 5155
rect 9715 5136 9900 5155
rect 9924 5136 10037 5160
rect 9715 5131 10037 5136
rect 9678 5127 10037 5131
rect 10104 5155 10253 5163
rect 10104 5135 10115 5155
rect 10135 5135 10253 5155
rect 10104 5128 10253 5135
rect 10104 5127 10145 5128
rect 9428 5074 9465 5075
rect 9524 5074 9561 5075
rect 9580 5074 9616 5126
rect 9635 5074 9672 5075
rect 9328 5065 9466 5074
rect 8316 5046 8484 5047
rect 8316 5043 8760 5046
rect 8316 5024 8691 5043
rect 8711 5024 8760 5043
rect 9328 5045 9437 5065
rect 9457 5045 9466 5065
rect 8316 5020 8760 5024
rect 8316 5018 8484 5020
rect 8316 4840 8343 5018
rect 8383 4980 8447 4992
rect 8723 4988 8760 5020
rect 8931 5019 9180 5041
rect 9328 5038 9466 5045
rect 9524 5065 9672 5074
rect 9524 5045 9533 5065
rect 9553 5045 9643 5065
rect 9663 5045 9672 5065
rect 9328 5036 9424 5038
rect 9524 5035 9672 5045
rect 9731 5065 9768 5075
rect 9843 5074 9880 5075
rect 9824 5072 9880 5074
rect 9731 5045 9739 5065
rect 9759 5045 9768 5065
rect 9580 5034 9616 5035
rect 8931 4988 8968 5019
rect 9144 5017 9180 5019
rect 9144 4988 9181 5017
rect 8383 4979 8418 4980
rect 8360 4974 8418 4979
rect 8360 4954 8363 4974
rect 8383 4960 8418 4974
rect 8438 4960 8447 4980
rect 8383 4952 8447 4960
rect 8409 4951 8447 4952
rect 8410 4950 8447 4951
rect 8513 4984 8549 4985
rect 8621 4984 8657 4985
rect 8513 4976 8657 4984
rect 8513 4956 8521 4976
rect 8541 4956 8573 4976
rect 8597 4956 8629 4976
rect 8649 4956 8657 4976
rect 8513 4950 8657 4956
rect 8723 4980 8761 4988
rect 8829 4984 8865 4985
rect 8723 4960 8732 4980
rect 8752 4960 8761 4980
rect 8723 4951 8761 4960
rect 8780 4977 8865 4984
rect 8780 4957 8787 4977
rect 8808 4976 8865 4977
rect 8808 4957 8837 4976
rect 8780 4956 8837 4957
rect 8857 4956 8865 4976
rect 8723 4950 8760 4951
rect 8780 4950 8865 4956
rect 8931 4980 8969 4988
rect 9042 4984 9078 4985
rect 8931 4960 8940 4980
rect 8960 4960 8969 4980
rect 8931 4951 8969 4960
rect 8993 4976 9078 4984
rect 8993 4956 9050 4976
rect 9070 4956 9078 4976
rect 8931 4950 8968 4951
rect 8993 4950 9078 4956
rect 9144 4980 9182 4988
rect 9144 4960 9153 4980
rect 9173 4960 9182 4980
rect 9428 4975 9465 4976
rect 9731 4975 9768 5045
rect 9793 5065 9880 5072
rect 9793 5062 9851 5065
rect 9793 5042 9798 5062
rect 9819 5045 9851 5062
rect 9871 5045 9880 5065
rect 9819 5042 9880 5045
rect 9793 5035 9880 5042
rect 9939 5065 9976 5075
rect 9939 5045 9947 5065
rect 9967 5045 9976 5065
rect 9793 5034 9824 5035
rect 9427 4974 9768 4975
rect 9144 4951 9182 4960
rect 9352 4969 9768 4974
rect 9144 4950 9181 4951
rect 8567 4929 8603 4950
rect 8993 4929 9024 4950
rect 9352 4949 9355 4969
rect 9375 4949 9768 4969
rect 9939 4974 9976 5045
rect 10006 5074 10037 5127
rect 10339 5112 10376 5122
rect 10339 5094 10348 5112
rect 10366 5094 10376 5112
rect 10339 5085 10376 5094
rect 10056 5074 10093 5075
rect 10006 5065 10093 5074
rect 10006 5045 10064 5065
rect 10084 5045 10093 5065
rect 10006 5035 10093 5045
rect 10152 5065 10189 5075
rect 10152 5045 10160 5065
rect 10180 5045 10189 5065
rect 10006 5034 10037 5035
rect 10152 4974 10189 5045
rect 10344 5020 10375 5085
rect 10343 5010 10380 5020
rect 10343 5008 10353 5010
rect 10277 5006 10353 5008
rect 9939 4950 10189 4974
rect 10274 4992 10353 5006
rect 10371 4992 10380 5010
rect 10274 4989 10380 4992
rect 9746 4930 9767 4949
rect 10274 4930 10300 4989
rect 10343 4983 10380 4989
rect 8400 4925 8500 4929
rect 8400 4921 8462 4925
rect 8400 4895 8407 4921
rect 8433 4899 8462 4921
rect 8488 4899 8500 4925
rect 8433 4895 8500 4899
rect 8400 4892 8500 4895
rect 8568 4892 8603 4929
rect 8665 4926 9024 4929
rect 8665 4921 8887 4926
rect 8665 4897 8678 4921
rect 8702 4902 8887 4921
rect 8911 4902 9024 4926
rect 8702 4897 9024 4902
rect 8665 4893 9024 4897
rect 9091 4921 9240 4929
rect 9091 4901 9102 4921
rect 9122 4901 9240 4921
rect 9746 4912 10300 4930
rect 10346 4919 10383 4921
rect 10274 4911 10300 4912
rect 10343 4911 10383 4919
rect 9091 4894 9240 4901
rect 10343 4899 10355 4911
rect 10334 4894 10355 4899
rect 9091 4893 9132 4894
rect 9750 4893 10355 4894
rect 10373 4893 10383 4911
rect 8415 4840 8452 4841
rect 8511 4840 8548 4841
rect 8567 4840 8603 4892
rect 8622 4840 8659 4841
rect 8315 4831 8453 4840
rect 8315 4811 8424 4831
rect 8444 4811 8453 4831
rect 8315 4804 8453 4811
rect 8511 4831 8659 4840
rect 8511 4811 8520 4831
rect 8540 4811 8630 4831
rect 8650 4811 8659 4831
rect 8315 4802 8411 4804
rect 8511 4801 8659 4811
rect 8718 4831 8755 4841
rect 8830 4840 8867 4841
rect 8811 4838 8867 4840
rect 8718 4811 8726 4831
rect 8746 4811 8755 4831
rect 8567 4800 8603 4801
rect 8415 4741 8452 4742
rect 8718 4741 8755 4811
rect 8780 4831 8867 4838
rect 8780 4828 8838 4831
rect 8780 4808 8785 4828
rect 8806 4811 8838 4828
rect 8858 4811 8867 4831
rect 8806 4808 8867 4811
rect 8780 4801 8867 4808
rect 8926 4831 8963 4841
rect 8926 4811 8934 4831
rect 8954 4811 8963 4831
rect 8780 4800 8811 4801
rect 8414 4740 8755 4741
rect 8339 4735 8755 4740
rect 8339 4715 8342 4735
rect 8362 4715 8755 4735
rect 8926 4740 8963 4811
rect 8993 4840 9024 4893
rect 9750 4884 10383 4893
rect 9750 4877 10382 4884
rect 9750 4875 9812 4877
rect 9328 4865 9496 4866
rect 9750 4865 9772 4875
rect 9043 4840 9080 4841
rect 8993 4831 9080 4840
rect 8993 4811 9051 4831
rect 9071 4811 9080 4831
rect 8993 4801 9080 4811
rect 9139 4831 9176 4841
rect 9139 4811 9147 4831
rect 9167 4811 9176 4831
rect 8993 4800 9024 4801
rect 9139 4740 9176 4811
rect 8926 4716 9176 4740
rect 9328 4839 9772 4865
rect 9328 4837 9496 4839
rect 9328 4659 9355 4837
rect 9395 4799 9459 4811
rect 9735 4807 9772 4839
rect 9943 4838 10192 4860
rect 9943 4807 9980 4838
rect 10156 4836 10192 4838
rect 10156 4807 10193 4836
rect 9395 4798 9430 4799
rect 9372 4793 9430 4798
rect 9372 4773 9375 4793
rect 9395 4779 9430 4793
rect 9450 4779 9459 4799
rect 9395 4771 9459 4779
rect 9421 4770 9459 4771
rect 9422 4769 9459 4770
rect 9525 4803 9561 4804
rect 9633 4803 9669 4804
rect 9525 4795 9669 4803
rect 9525 4775 9533 4795
rect 9553 4775 9582 4795
rect 9525 4774 9582 4775
rect 9604 4775 9641 4795
rect 9661 4775 9669 4795
rect 9604 4774 9669 4775
rect 9525 4769 9669 4774
rect 9735 4799 9773 4807
rect 9841 4803 9877 4804
rect 9735 4779 9744 4799
rect 9764 4779 9773 4799
rect 9735 4770 9773 4779
rect 9792 4796 9877 4803
rect 9792 4776 9799 4796
rect 9820 4795 9877 4796
rect 9820 4776 9849 4795
rect 9792 4775 9849 4776
rect 9869 4775 9877 4795
rect 9735 4769 9772 4770
rect 9792 4769 9877 4775
rect 9943 4799 9981 4807
rect 10054 4803 10090 4804
rect 9943 4779 9952 4799
rect 9972 4779 9981 4799
rect 9943 4770 9981 4779
rect 10005 4795 10090 4803
rect 10005 4775 10062 4795
rect 10082 4775 10090 4795
rect 9943 4769 9980 4770
rect 10005 4769 10090 4775
rect 10156 4799 10194 4807
rect 10156 4779 10165 4799
rect 10185 4779 10194 4799
rect 10156 4770 10194 4779
rect 10156 4769 10193 4770
rect 9579 4748 9615 4769
rect 10005 4748 10036 4769
rect 9412 4744 9512 4748
rect 9412 4740 9474 4744
rect 9412 4714 9419 4740
rect 9445 4718 9474 4740
rect 9500 4718 9512 4744
rect 9445 4714 9512 4718
rect 9412 4711 9512 4714
rect 9580 4711 9615 4748
rect 9677 4745 10036 4748
rect 9677 4740 9899 4745
rect 9677 4716 9690 4740
rect 9714 4721 9899 4740
rect 9923 4721 10036 4745
rect 9714 4716 10036 4721
rect 9677 4712 10036 4716
rect 10103 4740 10252 4748
rect 10103 4720 10114 4740
rect 10134 4720 10252 4740
rect 10103 4713 10252 4720
rect 10343 4728 10382 4877
rect 10103 4712 10144 4713
rect 9427 4659 9464 4660
rect 9523 4659 9560 4660
rect 9579 4659 9615 4711
rect 9634 4659 9671 4660
rect 9327 4650 9465 4659
rect 9327 4630 9436 4650
rect 9456 4630 9465 4650
rect 9327 4623 9465 4630
rect 9523 4650 9671 4659
rect 9523 4630 9532 4650
rect 9552 4630 9642 4650
rect 9662 4630 9671 4650
rect 9327 4621 9423 4623
rect 9523 4620 9671 4630
rect 9730 4650 9767 4660
rect 9842 4659 9879 4660
rect 9823 4657 9879 4659
rect 9730 4630 9738 4650
rect 9758 4630 9767 4650
rect 9579 4619 9615 4620
rect 7492 4611 7523 4614
rect 8021 4614 8189 4615
rect 6321 4587 6459 4596
rect 8021 4588 8465 4614
rect 6115 4586 6152 4587
rect 6171 4535 6207 4587
rect 6226 4586 6263 4587
rect 6322 4586 6359 4587
rect 5642 4533 5683 4534
rect 4449 4511 5098 4517
rect 5534 4526 5683 4533
rect 4449 4510 5097 4511
rect 3515 4490 3526 4510
rect 3546 4490 3664 4510
rect 5060 4508 5097 4510
rect 5534 4506 5652 4526
rect 5672 4506 5683 4526
rect 5534 4498 5683 4506
rect 5750 4530 6109 4534
rect 5750 4525 6072 4530
rect 5750 4501 5863 4525
rect 5887 4506 6072 4525
rect 6096 4506 6109 4530
rect 5887 4501 6109 4506
rect 5750 4498 6109 4501
rect 6171 4498 6206 4535
rect 6274 4532 6374 4535
rect 6274 4528 6341 4532
rect 6274 4502 6286 4528
rect 6312 4506 6341 4528
rect 6367 4506 6374 4532
rect 6312 4502 6374 4506
rect 6274 4498 6374 4502
rect 3515 4483 3664 4490
rect 3515 4482 3556 4483
rect 2839 4429 2876 4430
rect 2935 4429 2972 4430
rect 2991 4429 3027 4481
rect 3046 4429 3083 4430
rect 733 4402 1177 4428
rect 734 4385 758 4402
rect 1009 4401 1177 4402
rect 1628 4398 1878 4422
rect 132 4367 759 4385
rect 132 4366 170 4367
rect 130 4361 170 4366
rect 130 4318 165 4361
rect 128 4309 165 4318
rect 128 4291 138 4309
rect 156 4291 165 4309
rect 1628 4327 1665 4398
rect 1780 4337 1811 4338
rect 1628 4307 1637 4327
rect 1657 4307 1665 4327
rect 1628 4297 1665 4307
rect 1724 4327 1811 4337
rect 1724 4307 1733 4327
rect 1753 4307 1811 4327
rect 1724 4298 1811 4307
rect 1724 4297 1761 4298
rect 128 4281 165 4291
rect 1780 4245 1811 4298
rect 1841 4327 1878 4398
rect 2049 4403 2442 4423
rect 2462 4403 2465 4423
rect 2049 4398 2465 4403
rect 2739 4420 2877 4429
rect 2739 4400 2848 4420
rect 2868 4400 2877 4420
rect 2049 4397 2390 4398
rect 1993 4337 2024 4338
rect 1841 4307 1850 4327
rect 1870 4307 1878 4327
rect 1841 4297 1878 4307
rect 1937 4330 2024 4337
rect 1937 4327 1998 4330
rect 1937 4307 1946 4327
rect 1966 4310 1998 4327
rect 2019 4310 2024 4330
rect 1966 4307 2024 4310
rect 1937 4300 2024 4307
rect 2049 4327 2086 4397
rect 2352 4396 2389 4397
rect 2739 4393 2877 4400
rect 2935 4420 3083 4429
rect 2935 4400 2944 4420
rect 2964 4400 3054 4420
rect 3074 4400 3083 4420
rect 2739 4391 2835 4393
rect 2935 4390 3083 4400
rect 3142 4420 3179 4430
rect 3254 4429 3291 4430
rect 3235 4427 3291 4429
rect 3142 4400 3150 4420
rect 3170 4400 3179 4420
rect 2991 4389 3027 4390
rect 2201 4337 2237 4338
rect 2049 4307 2058 4327
rect 2078 4307 2086 4327
rect 1937 4298 1993 4300
rect 1937 4297 1974 4298
rect 2049 4297 2086 4307
rect 2145 4327 2293 4337
rect 2393 4334 2489 4336
rect 2145 4307 2154 4327
rect 2174 4307 2264 4327
rect 2284 4307 2293 4327
rect 2145 4298 2293 4307
rect 2351 4327 2489 4334
rect 2839 4330 2876 4331
rect 3142 4330 3179 4400
rect 3204 4420 3291 4427
rect 3204 4417 3262 4420
rect 3204 4397 3209 4417
rect 3230 4400 3262 4417
rect 3282 4400 3291 4420
rect 3230 4397 3291 4400
rect 3204 4390 3291 4397
rect 3350 4420 3387 4430
rect 3350 4400 3358 4420
rect 3378 4400 3387 4420
rect 3204 4389 3235 4390
rect 2838 4329 3179 4330
rect 2351 4307 2360 4327
rect 2380 4307 2489 4327
rect 2351 4298 2489 4307
rect 2763 4324 3179 4329
rect 2763 4304 2766 4324
rect 2786 4304 3179 4324
rect 3350 4329 3387 4400
rect 3417 4429 3448 4482
rect 5750 4477 5781 4498
rect 6171 4477 6207 4498
rect 5414 4468 5451 4477
rect 5593 4476 5630 4477
rect 5414 4450 5423 4468
rect 5441 4450 5451 4468
rect 5063 4436 5100 4446
rect 5414 4440 5451 4450
rect 3467 4429 3504 4430
rect 3417 4420 3504 4429
rect 3417 4400 3475 4420
rect 3495 4400 3504 4420
rect 3417 4390 3504 4400
rect 3563 4420 3600 4430
rect 3563 4400 3571 4420
rect 3591 4400 3600 4420
rect 3417 4389 3448 4390
rect 3563 4329 3600 4400
rect 5063 4418 5072 4436
rect 5090 4418 5100 4436
rect 5063 4409 5100 4418
rect 5063 4366 5098 4409
rect 5415 4405 5451 4440
rect 5592 4467 5630 4476
rect 5592 4447 5601 4467
rect 5621 4447 5630 4467
rect 5592 4439 5630 4447
rect 5696 4471 5781 4477
rect 5806 4476 5843 4477
rect 5696 4451 5704 4471
rect 5724 4451 5781 4471
rect 5696 4443 5781 4451
rect 5805 4467 5843 4476
rect 5805 4447 5814 4467
rect 5834 4447 5843 4467
rect 5696 4442 5732 4443
rect 5805 4439 5843 4447
rect 5909 4471 5994 4477
rect 6014 4476 6051 4477
rect 5909 4451 5917 4471
rect 5937 4470 5994 4471
rect 5937 4451 5966 4470
rect 5909 4450 5966 4451
rect 5987 4450 5994 4470
rect 5909 4443 5994 4450
rect 6013 4467 6051 4476
rect 6013 4447 6022 4467
rect 6042 4447 6051 4467
rect 5909 4442 5945 4443
rect 6013 4439 6051 4447
rect 6117 4471 6261 4477
rect 6117 4451 6125 4471
rect 6145 4470 6233 4471
rect 6145 4451 6173 4470
rect 6117 4449 6173 4451
rect 6195 4451 6233 4470
rect 6253 4451 6261 4471
rect 6195 4449 6261 4451
rect 6117 4443 6261 4449
rect 6117 4442 6153 4443
rect 6225 4442 6261 4443
rect 6327 4476 6364 4477
rect 6327 4475 6365 4476
rect 6327 4467 6391 4475
rect 6327 4447 6336 4467
rect 6356 4453 6391 4467
rect 6411 4453 6414 4473
rect 6356 4448 6414 4453
rect 6356 4447 6391 4448
rect 5593 4410 5630 4439
rect 5058 4361 5098 4366
rect 5413 4364 5451 4405
rect 5594 4408 5630 4410
rect 5806 4408 5843 4439
rect 5594 4386 5843 4408
rect 6014 4407 6051 4439
rect 6327 4435 6391 4447
rect 6431 4409 6458 4587
rect 6290 4407 6458 4409
rect 8021 4586 8189 4588
rect 8021 4583 8068 4586
rect 8021 4408 8048 4583
rect 8088 4548 8152 4560
rect 8428 4556 8465 4588
rect 8636 4587 8885 4609
rect 8636 4556 8673 4587
rect 8849 4585 8885 4587
rect 8849 4556 8886 4585
rect 9427 4560 9464 4561
rect 9730 4560 9767 4630
rect 9792 4650 9879 4657
rect 9792 4647 9850 4650
rect 9792 4627 9797 4647
rect 9818 4630 9850 4647
rect 9870 4630 9879 4650
rect 9818 4627 9879 4630
rect 9792 4620 9879 4627
rect 9938 4650 9975 4660
rect 9938 4630 9946 4650
rect 9966 4630 9975 4650
rect 9792 4619 9823 4620
rect 9426 4559 9767 4560
rect 8088 4547 8123 4548
rect 8065 4542 8123 4547
rect 8065 4522 8068 4542
rect 8088 4528 8123 4542
rect 8143 4528 8152 4548
rect 8088 4520 8152 4528
rect 8114 4519 8152 4520
rect 8115 4518 8152 4519
rect 8218 4552 8254 4553
rect 8326 4552 8362 4553
rect 8218 4544 8362 4552
rect 8218 4524 8226 4544
rect 8246 4542 8334 4544
rect 8246 4524 8272 4542
rect 8218 4523 8272 4524
rect 8298 4524 8334 4542
rect 8354 4524 8362 4544
rect 8298 4523 8362 4524
rect 8218 4518 8362 4523
rect 8428 4548 8466 4556
rect 8534 4552 8570 4553
rect 8428 4528 8437 4548
rect 8457 4528 8466 4548
rect 8428 4519 8466 4528
rect 8485 4545 8570 4552
rect 8485 4525 8492 4545
rect 8513 4544 8570 4545
rect 8513 4525 8542 4544
rect 8485 4524 8542 4525
rect 8562 4524 8570 4544
rect 8428 4518 8465 4519
rect 8485 4518 8570 4524
rect 8636 4548 8674 4556
rect 8747 4552 8783 4553
rect 8636 4528 8645 4548
rect 8665 4528 8674 4548
rect 8636 4519 8674 4528
rect 8698 4544 8783 4552
rect 8698 4524 8755 4544
rect 8775 4524 8783 4544
rect 8636 4518 8673 4519
rect 8698 4518 8783 4524
rect 8849 4548 8887 4556
rect 8849 4528 8858 4548
rect 8878 4528 8887 4548
rect 9351 4554 9767 4559
rect 9351 4534 9354 4554
rect 9374 4534 9767 4554
rect 9938 4559 9975 4630
rect 10005 4659 10036 4712
rect 10343 4710 10353 4728
rect 10371 4710 10382 4728
rect 10343 4701 10380 4710
rect 10055 4659 10092 4660
rect 10005 4650 10092 4659
rect 10005 4630 10063 4650
rect 10083 4630 10092 4650
rect 10005 4620 10092 4630
rect 10151 4650 10188 4660
rect 10151 4630 10159 4650
rect 10179 4630 10188 4650
rect 10346 4635 10383 4639
rect 10005 4619 10036 4620
rect 10151 4559 10188 4630
rect 9938 4535 10188 4559
rect 10344 4629 10383 4635
rect 10344 4611 10355 4629
rect 10373 4611 10383 4629
rect 10344 4602 10383 4611
rect 8849 4519 8887 4528
rect 8849 4518 8886 4519
rect 8272 4497 8308 4518
rect 8698 4497 8729 4518
rect 9730 4511 9767 4534
rect 10344 4524 10379 4602
rect 10341 4514 10379 4524
rect 9730 4510 9900 4511
rect 10341 4510 10351 4514
rect 8105 4493 8205 4497
rect 8105 4489 8167 4493
rect 8105 4463 8112 4489
rect 8138 4467 8167 4489
rect 8193 4467 8205 4493
rect 8138 4463 8205 4467
rect 8105 4460 8205 4463
rect 8273 4460 8308 4497
rect 8370 4494 8729 4497
rect 8370 4489 8592 4494
rect 8370 4465 8383 4489
rect 8407 4470 8592 4489
rect 8616 4470 8729 4494
rect 8407 4465 8729 4470
rect 8370 4461 8729 4465
rect 8796 4489 8945 4497
rect 9730 4496 10351 4510
rect 10369 4496 10379 4514
rect 9730 4490 10379 4496
rect 9730 4489 10378 4490
rect 8796 4469 8807 4489
rect 8827 4469 8945 4489
rect 10341 4487 10378 4489
rect 8796 4462 8945 4469
rect 8796 4461 8837 4462
rect 8120 4408 8157 4409
rect 8216 4408 8253 4409
rect 8272 4408 8308 4460
rect 8327 4408 8364 4409
rect 6014 4381 6458 4407
rect 6015 4364 6039 4381
rect 6290 4380 6458 4381
rect 6909 4377 7159 4401
rect 5058 4360 5096 4361
rect 4469 4342 5096 4360
rect 5413 4346 6040 4364
rect 5413 4345 5451 4346
rect 3350 4305 3600 4329
rect 4051 4325 4219 4326
rect 4470 4325 4494 4342
rect 4051 4299 4495 4325
rect 2145 4297 2182 4298
rect 2201 4246 2237 4298
rect 2256 4297 2293 4298
rect 2352 4297 2389 4298
rect 1672 4244 1713 4245
rect 1564 4237 1713 4244
rect 131 4217 168 4219
rect 1564 4217 1682 4237
rect 1702 4217 1713 4237
rect 131 4216 779 4217
rect 130 4210 779 4216
rect 130 4192 140 4210
rect 158 4196 779 4210
rect 1564 4209 1713 4217
rect 1780 4241 2139 4245
rect 1780 4236 2102 4241
rect 1780 4212 1893 4236
rect 1917 4217 2102 4236
rect 2126 4217 2139 4241
rect 1917 4212 2139 4217
rect 1780 4209 2139 4212
rect 2201 4209 2236 4246
rect 2304 4243 2404 4246
rect 2304 4239 2371 4243
rect 2304 4213 2316 4239
rect 2342 4217 2371 4239
rect 2397 4217 2404 4243
rect 2342 4213 2404 4217
rect 2304 4209 2404 4213
rect 158 4192 168 4196
rect 609 4195 779 4196
rect 130 4182 168 4192
rect 130 4104 165 4182
rect 742 4172 779 4195
rect 1780 4188 1811 4209
rect 2201 4188 2237 4209
rect 1623 4187 1660 4188
rect 1622 4178 1660 4187
rect 126 4095 165 4104
rect 126 4077 136 4095
rect 154 4077 165 4095
rect 126 4071 165 4077
rect 321 4147 571 4171
rect 321 4076 358 4147
rect 473 4086 504 4087
rect 126 4067 163 4071
rect 321 4056 330 4076
rect 350 4056 358 4076
rect 321 4046 358 4056
rect 417 4076 504 4086
rect 417 4056 426 4076
rect 446 4056 504 4076
rect 417 4047 504 4056
rect 417 4046 454 4047
rect 129 3996 166 4005
rect 127 3978 138 3996
rect 156 3978 166 3996
rect 473 3994 504 4047
rect 534 4076 571 4147
rect 742 4152 1135 4172
rect 1155 4152 1158 4172
rect 742 4147 1158 4152
rect 1622 4158 1631 4178
rect 1651 4158 1660 4178
rect 1622 4150 1660 4158
rect 1726 4182 1811 4188
rect 1836 4187 1873 4188
rect 1726 4162 1734 4182
rect 1754 4162 1811 4182
rect 1726 4154 1811 4162
rect 1835 4178 1873 4187
rect 1835 4158 1844 4178
rect 1864 4158 1873 4178
rect 1726 4153 1762 4154
rect 1835 4150 1873 4158
rect 1939 4182 2024 4188
rect 2044 4187 2081 4188
rect 1939 4162 1947 4182
rect 1967 4181 2024 4182
rect 1967 4162 1996 4181
rect 1939 4161 1996 4162
rect 2017 4161 2024 4181
rect 1939 4154 2024 4161
rect 2043 4178 2081 4187
rect 2043 4158 2052 4178
rect 2072 4158 2081 4178
rect 1939 4153 1975 4154
rect 2043 4150 2081 4158
rect 2147 4183 2291 4188
rect 2147 4182 2211 4183
rect 2147 4162 2155 4182
rect 2175 4164 2211 4182
rect 2237 4182 2291 4183
rect 2237 4164 2263 4182
rect 2175 4162 2263 4164
rect 2283 4162 2291 4182
rect 2147 4154 2291 4162
rect 2147 4153 2183 4154
rect 2255 4153 2291 4154
rect 2357 4187 2394 4188
rect 2357 4186 2395 4187
rect 2357 4178 2421 4186
rect 2357 4158 2366 4178
rect 2386 4164 2421 4178
rect 2441 4164 2444 4184
rect 2386 4159 2444 4164
rect 2386 4158 2421 4159
rect 742 4146 1083 4147
rect 686 4086 717 4087
rect 534 4056 543 4076
rect 563 4056 571 4076
rect 534 4046 571 4056
rect 630 4079 717 4086
rect 630 4076 691 4079
rect 630 4056 639 4076
rect 659 4059 691 4076
rect 712 4059 717 4079
rect 659 4056 717 4059
rect 630 4049 717 4056
rect 742 4076 779 4146
rect 1045 4145 1082 4146
rect 1623 4121 1660 4150
rect 1624 4119 1660 4121
rect 1836 4119 1873 4150
rect 1624 4097 1873 4119
rect 2044 4118 2081 4150
rect 2357 4146 2421 4158
rect 2461 4123 2488 4298
rect 2441 4120 2488 4123
rect 2320 4118 2488 4120
rect 4051 4297 4219 4299
rect 4051 4119 4078 4297
rect 4118 4259 4182 4271
rect 4458 4267 4495 4299
rect 4666 4298 4915 4320
rect 4666 4267 4703 4298
rect 4879 4296 4915 4298
rect 5058 4301 5096 4342
rect 5411 4340 5451 4345
rect 4879 4267 4916 4296
rect 4118 4258 4153 4259
rect 4095 4253 4153 4258
rect 4095 4233 4098 4253
rect 4118 4239 4153 4253
rect 4173 4239 4182 4259
rect 4118 4231 4182 4239
rect 4144 4230 4182 4231
rect 4145 4229 4182 4230
rect 4248 4263 4284 4264
rect 4356 4263 4392 4264
rect 4248 4257 4392 4263
rect 4248 4255 4314 4257
rect 4248 4235 4256 4255
rect 4276 4236 4314 4255
rect 4336 4255 4392 4257
rect 4336 4236 4364 4255
rect 4276 4235 4364 4236
rect 4384 4235 4392 4255
rect 4248 4229 4392 4235
rect 4458 4259 4496 4267
rect 4564 4263 4600 4264
rect 4458 4239 4467 4259
rect 4487 4239 4496 4259
rect 4458 4230 4496 4239
rect 4515 4256 4600 4263
rect 4515 4236 4522 4256
rect 4543 4255 4600 4256
rect 4543 4236 4572 4255
rect 4515 4235 4572 4236
rect 4592 4235 4600 4255
rect 4458 4229 4495 4230
rect 4515 4229 4600 4235
rect 4666 4259 4704 4267
rect 4777 4263 4813 4264
rect 4666 4239 4675 4259
rect 4695 4239 4704 4259
rect 4666 4230 4704 4239
rect 4728 4255 4813 4263
rect 4728 4235 4785 4255
rect 4805 4235 4813 4255
rect 4666 4229 4703 4230
rect 4728 4229 4813 4235
rect 4879 4259 4917 4267
rect 4879 4239 4888 4259
rect 4908 4239 4917 4259
rect 4879 4230 4917 4239
rect 5058 4266 5094 4301
rect 5411 4297 5446 4340
rect 5409 4288 5446 4297
rect 5409 4270 5419 4288
rect 5437 4270 5446 4288
rect 6909 4306 6946 4377
rect 7061 4316 7092 4317
rect 6909 4286 6918 4306
rect 6938 4286 6946 4306
rect 6909 4276 6946 4286
rect 7005 4306 7092 4316
rect 7005 4286 7014 4306
rect 7034 4286 7092 4306
rect 7005 4277 7092 4286
rect 7005 4276 7042 4277
rect 5058 4256 5095 4266
rect 5409 4260 5446 4270
rect 5058 4238 5068 4256
rect 5086 4238 5095 4256
rect 4879 4229 4916 4230
rect 5058 4229 5095 4238
rect 4302 4208 4338 4229
rect 4728 4208 4759 4229
rect 7061 4224 7092 4277
rect 7122 4306 7159 4377
rect 7330 4382 7723 4402
rect 7743 4382 7746 4402
rect 7330 4377 7746 4382
rect 8020 4399 8158 4408
rect 8020 4379 8129 4399
rect 8149 4379 8158 4399
rect 7330 4376 7671 4377
rect 7274 4316 7305 4317
rect 7122 4286 7131 4306
rect 7151 4286 7159 4306
rect 7122 4276 7159 4286
rect 7218 4309 7305 4316
rect 7218 4306 7279 4309
rect 7218 4286 7227 4306
rect 7247 4289 7279 4306
rect 7300 4289 7305 4309
rect 7247 4286 7305 4289
rect 7218 4279 7305 4286
rect 7330 4306 7367 4376
rect 7633 4375 7670 4376
rect 8020 4372 8158 4379
rect 8216 4399 8364 4408
rect 8216 4379 8225 4399
rect 8245 4379 8335 4399
rect 8355 4379 8364 4399
rect 8020 4370 8116 4372
rect 8216 4369 8364 4379
rect 8423 4399 8460 4409
rect 8535 4408 8572 4409
rect 8516 4406 8572 4408
rect 8423 4379 8431 4399
rect 8451 4379 8460 4399
rect 8272 4368 8308 4369
rect 7482 4316 7518 4317
rect 7330 4286 7339 4306
rect 7359 4286 7367 4306
rect 7218 4277 7274 4279
rect 7218 4276 7255 4277
rect 7330 4276 7367 4286
rect 7426 4306 7574 4316
rect 7674 4313 7770 4315
rect 7426 4286 7435 4306
rect 7455 4286 7545 4306
rect 7565 4286 7574 4306
rect 7426 4277 7574 4286
rect 7632 4306 7770 4313
rect 8120 4309 8157 4310
rect 8423 4309 8460 4379
rect 8485 4399 8572 4406
rect 8485 4396 8543 4399
rect 8485 4376 8490 4396
rect 8511 4379 8543 4396
rect 8563 4379 8572 4399
rect 8511 4376 8572 4379
rect 8485 4369 8572 4376
rect 8631 4399 8668 4409
rect 8631 4379 8639 4399
rect 8659 4379 8668 4399
rect 8485 4368 8516 4369
rect 8119 4308 8460 4309
rect 7632 4286 7641 4306
rect 7661 4286 7770 4306
rect 7632 4277 7770 4286
rect 8044 4303 8460 4308
rect 8044 4283 8047 4303
rect 8067 4283 8460 4303
rect 8631 4308 8668 4379
rect 8698 4408 8729 4461
rect 10344 4415 10381 4425
rect 8748 4408 8785 4409
rect 8698 4399 8785 4408
rect 8698 4379 8756 4399
rect 8776 4379 8785 4399
rect 8698 4369 8785 4379
rect 8844 4399 8881 4409
rect 8844 4379 8852 4399
rect 8872 4379 8881 4399
rect 8698 4368 8729 4369
rect 8844 4308 8881 4379
rect 10344 4397 10353 4415
rect 10371 4397 10381 4415
rect 10344 4388 10381 4397
rect 10344 4345 10379 4388
rect 10339 4340 10379 4345
rect 10339 4339 10377 4340
rect 9750 4321 10377 4339
rect 8631 4284 8881 4308
rect 9332 4304 9500 4305
rect 9751 4304 9775 4321
rect 9332 4278 9776 4304
rect 7426 4276 7463 4277
rect 7482 4225 7518 4277
rect 7537 4276 7574 4277
rect 7633 4276 7670 4277
rect 6953 4223 6994 4224
rect 6845 4216 6994 4223
rect 4135 4204 4235 4208
rect 4135 4200 4197 4204
rect 4135 4174 4142 4200
rect 4168 4178 4197 4200
rect 4223 4178 4235 4204
rect 4168 4174 4235 4178
rect 4135 4171 4235 4174
rect 4303 4171 4338 4208
rect 4400 4205 4759 4208
rect 4400 4200 4622 4205
rect 4400 4176 4413 4200
rect 4437 4181 4622 4200
rect 4646 4181 4759 4205
rect 4437 4176 4759 4181
rect 4400 4172 4759 4176
rect 4826 4200 4975 4208
rect 4826 4180 4837 4200
rect 4857 4180 4975 4200
rect 5412 4196 5449 4198
rect 6845 4196 6963 4216
rect 6983 4196 6994 4216
rect 5412 4195 6060 4196
rect 4826 4173 4975 4180
rect 5411 4189 6060 4195
rect 4826 4172 4867 4173
rect 4150 4119 4187 4120
rect 4246 4119 4283 4120
rect 4302 4119 4338 4171
rect 4357 4119 4394 4120
rect 2044 4092 2488 4118
rect 4050 4110 4188 4119
rect 2320 4091 2488 4092
rect 2986 4092 3017 4095
rect 894 4086 930 4087
rect 742 4056 751 4076
rect 771 4056 779 4076
rect 630 4047 686 4049
rect 630 4046 667 4047
rect 742 4046 779 4056
rect 838 4076 986 4086
rect 1086 4083 1182 4085
rect 838 4056 847 4076
rect 867 4056 957 4076
rect 977 4056 986 4076
rect 838 4047 986 4056
rect 1044 4076 1182 4083
rect 1044 4056 1053 4076
rect 1073 4056 1182 4076
rect 1044 4047 1182 4056
rect 838 4046 875 4047
rect 894 3995 930 4047
rect 949 4046 986 4047
rect 1045 4046 1082 4047
rect 365 3993 406 3994
rect 127 3829 166 3978
rect 257 3986 406 3993
rect 257 3966 375 3986
rect 395 3966 406 3986
rect 257 3958 406 3966
rect 473 3990 832 3994
rect 473 3985 795 3990
rect 473 3961 586 3985
rect 610 3966 795 3985
rect 819 3966 832 3990
rect 610 3961 832 3966
rect 473 3958 832 3961
rect 894 3958 929 3995
rect 997 3992 1097 3995
rect 997 3988 1064 3992
rect 997 3962 1009 3988
rect 1035 3966 1064 3988
rect 1090 3966 1097 3992
rect 1035 3962 1097 3966
rect 997 3958 1097 3962
rect 473 3937 504 3958
rect 894 3937 930 3958
rect 316 3936 353 3937
rect 315 3927 353 3936
rect 315 3907 324 3927
rect 344 3907 353 3927
rect 315 3899 353 3907
rect 419 3931 504 3937
rect 529 3936 566 3937
rect 419 3911 427 3931
rect 447 3911 504 3931
rect 419 3903 504 3911
rect 528 3927 566 3936
rect 528 3907 537 3927
rect 557 3907 566 3927
rect 419 3902 455 3903
rect 528 3899 566 3907
rect 632 3931 717 3937
rect 737 3936 774 3937
rect 632 3911 640 3931
rect 660 3930 717 3931
rect 660 3911 689 3930
rect 632 3910 689 3911
rect 710 3910 717 3930
rect 632 3903 717 3910
rect 736 3927 774 3936
rect 736 3907 745 3927
rect 765 3907 774 3927
rect 632 3902 668 3903
rect 736 3899 774 3907
rect 840 3932 984 3937
rect 840 3931 905 3932
rect 840 3911 848 3931
rect 868 3911 905 3931
rect 927 3931 984 3932
rect 927 3911 956 3931
rect 976 3911 984 3931
rect 840 3903 984 3911
rect 840 3902 876 3903
rect 948 3902 984 3903
rect 1050 3936 1087 3937
rect 1050 3935 1088 3936
rect 1050 3927 1114 3935
rect 1050 3907 1059 3927
rect 1079 3913 1114 3927
rect 1134 3913 1137 3933
rect 1079 3908 1137 3913
rect 1079 3907 1114 3908
rect 316 3870 353 3899
rect 317 3868 353 3870
rect 529 3868 566 3899
rect 317 3846 566 3868
rect 737 3867 774 3899
rect 1050 3895 1114 3907
rect 1154 3869 1181 4047
rect 1013 3867 1181 3869
rect 737 3841 1181 3867
rect 1333 3966 1583 3990
rect 1333 3895 1370 3966
rect 1485 3905 1516 3906
rect 1333 3875 1342 3895
rect 1362 3875 1370 3895
rect 1333 3865 1370 3875
rect 1429 3895 1516 3905
rect 1429 3875 1438 3895
rect 1458 3875 1516 3895
rect 1429 3866 1516 3875
rect 1429 3865 1466 3866
rect 737 3831 759 3841
rect 1013 3840 1181 3841
rect 697 3829 759 3831
rect 127 3822 759 3829
rect 126 3813 759 3822
rect 1485 3813 1516 3866
rect 1546 3895 1583 3966
rect 1754 3971 2147 3991
rect 2167 3971 2170 3991
rect 1754 3966 2170 3971
rect 1754 3965 2095 3966
rect 1698 3905 1729 3906
rect 1546 3875 1555 3895
rect 1575 3875 1583 3895
rect 1546 3865 1583 3875
rect 1642 3898 1729 3905
rect 1642 3895 1703 3898
rect 1642 3875 1651 3895
rect 1671 3878 1703 3895
rect 1724 3878 1729 3898
rect 1671 3875 1729 3878
rect 1642 3868 1729 3875
rect 1754 3895 1791 3965
rect 2057 3964 2094 3965
rect 1906 3905 1942 3906
rect 1754 3875 1763 3895
rect 1783 3875 1791 3895
rect 1642 3866 1698 3868
rect 1642 3865 1679 3866
rect 1754 3865 1791 3875
rect 1850 3895 1998 3905
rect 2098 3902 2194 3904
rect 1850 3875 1859 3895
rect 1879 3875 1969 3895
rect 1989 3875 1998 3895
rect 1850 3866 1998 3875
rect 2056 3895 2194 3902
rect 2056 3875 2065 3895
rect 2085 3875 2194 3895
rect 2056 3866 2194 3875
rect 1850 3865 1887 3866
rect 1906 3814 1942 3866
rect 1961 3865 1998 3866
rect 2057 3865 2094 3866
rect 126 3795 136 3813
rect 154 3812 759 3813
rect 1377 3812 1418 3813
rect 154 3807 175 3812
rect 154 3795 166 3807
rect 1269 3805 1418 3812
rect 126 3787 166 3795
rect 209 3794 235 3795
rect 126 3785 163 3787
rect 209 3776 763 3794
rect 1269 3785 1387 3805
rect 1407 3785 1418 3805
rect 1269 3777 1418 3785
rect 1485 3809 1844 3813
rect 1485 3804 1807 3809
rect 1485 3780 1598 3804
rect 1622 3785 1807 3804
rect 1831 3785 1844 3809
rect 1622 3780 1844 3785
rect 1485 3777 1844 3780
rect 1906 3777 1941 3814
rect 2009 3811 2109 3814
rect 2009 3807 2076 3811
rect 2009 3781 2021 3807
rect 2047 3785 2076 3807
rect 2102 3785 2109 3811
rect 2047 3781 2109 3785
rect 2009 3777 2109 3781
rect 129 3717 166 3723
rect 209 3717 235 3776
rect 742 3757 763 3776
rect 129 3714 235 3717
rect 129 3696 138 3714
rect 156 3700 235 3714
rect 320 3732 570 3756
rect 156 3698 232 3700
rect 156 3696 166 3698
rect 129 3686 166 3696
rect 134 3621 165 3686
rect 320 3661 357 3732
rect 472 3671 503 3672
rect 320 3641 329 3661
rect 349 3641 357 3661
rect 320 3631 357 3641
rect 416 3661 503 3671
rect 416 3641 425 3661
rect 445 3641 503 3661
rect 416 3632 503 3641
rect 416 3631 453 3632
rect 133 3612 170 3621
rect 133 3594 143 3612
rect 161 3594 170 3612
rect 133 3584 170 3594
rect 472 3579 503 3632
rect 533 3661 570 3732
rect 741 3737 1134 3757
rect 1154 3737 1157 3757
rect 1485 3756 1516 3777
rect 1906 3756 1942 3777
rect 1328 3755 1365 3756
rect 741 3732 1157 3737
rect 1327 3746 1365 3755
rect 741 3731 1082 3732
rect 685 3671 716 3672
rect 533 3641 542 3661
rect 562 3641 570 3661
rect 533 3631 570 3641
rect 629 3664 716 3671
rect 629 3661 690 3664
rect 629 3641 638 3661
rect 658 3644 690 3661
rect 711 3644 716 3664
rect 658 3641 716 3644
rect 629 3634 716 3641
rect 741 3661 778 3731
rect 1044 3730 1081 3731
rect 1327 3726 1336 3746
rect 1356 3726 1365 3746
rect 1327 3718 1365 3726
rect 1431 3750 1516 3756
rect 1541 3755 1578 3756
rect 1431 3730 1439 3750
rect 1459 3730 1516 3750
rect 1431 3722 1516 3730
rect 1540 3746 1578 3755
rect 1540 3726 1549 3746
rect 1569 3726 1578 3746
rect 1431 3721 1467 3722
rect 1540 3718 1578 3726
rect 1644 3750 1729 3756
rect 1749 3755 1786 3756
rect 1644 3730 1652 3750
rect 1672 3749 1729 3750
rect 1672 3730 1701 3749
rect 1644 3729 1701 3730
rect 1722 3729 1729 3749
rect 1644 3722 1729 3729
rect 1748 3746 1786 3755
rect 1748 3726 1757 3746
rect 1777 3726 1786 3746
rect 1644 3721 1680 3722
rect 1748 3718 1786 3726
rect 1852 3750 1996 3756
rect 1852 3730 1860 3750
rect 1880 3730 1912 3750
rect 1936 3730 1968 3750
rect 1988 3730 1996 3750
rect 1852 3722 1996 3730
rect 1852 3721 1888 3722
rect 1960 3721 1996 3722
rect 2062 3755 2099 3756
rect 2062 3754 2100 3755
rect 2062 3746 2126 3754
rect 2062 3726 2071 3746
rect 2091 3732 2126 3746
rect 2146 3732 2149 3752
rect 2091 3727 2149 3732
rect 2091 3726 2126 3727
rect 1328 3689 1365 3718
rect 1329 3687 1365 3689
rect 1541 3687 1578 3718
rect 893 3671 929 3672
rect 741 3641 750 3661
rect 770 3641 778 3661
rect 629 3632 685 3634
rect 629 3631 666 3632
rect 741 3631 778 3641
rect 837 3661 985 3671
rect 1085 3668 1181 3670
rect 837 3641 846 3661
rect 866 3641 956 3661
rect 976 3641 985 3661
rect 837 3632 985 3641
rect 1043 3661 1181 3668
rect 1329 3665 1578 3687
rect 1749 3686 1786 3718
rect 2062 3714 2126 3726
rect 2166 3688 2193 3866
rect 2025 3686 2193 3688
rect 1749 3682 2193 3686
rect 1043 3641 1052 3661
rect 1072 3641 1181 3661
rect 1749 3663 1798 3682
rect 1818 3663 2193 3682
rect 1749 3660 2193 3663
rect 2025 3659 2193 3660
rect 1043 3632 1181 3641
rect 837 3631 874 3632
rect 893 3580 929 3632
rect 948 3631 985 3632
rect 1044 3631 1081 3632
rect 364 3578 405 3579
rect 256 3571 405 3578
rect 256 3551 374 3571
rect 394 3551 405 3571
rect 256 3543 405 3551
rect 472 3575 831 3579
rect 472 3570 794 3575
rect 472 3546 585 3570
rect 609 3551 794 3570
rect 818 3551 831 3575
rect 609 3546 831 3551
rect 472 3543 831 3546
rect 893 3543 928 3580
rect 996 3577 1096 3580
rect 996 3573 1063 3577
rect 996 3547 1008 3573
rect 1034 3551 1063 3573
rect 1089 3551 1096 3577
rect 1034 3547 1096 3551
rect 996 3543 1096 3547
rect 472 3522 503 3543
rect 893 3522 929 3543
rect 136 3513 173 3522
rect 315 3521 352 3522
rect 136 3495 145 3513
rect 163 3495 173 3513
rect 136 3485 173 3495
rect 137 3450 173 3485
rect 314 3512 352 3521
rect 314 3492 323 3512
rect 343 3492 352 3512
rect 314 3484 352 3492
rect 418 3516 503 3522
rect 528 3521 565 3522
rect 418 3496 426 3516
rect 446 3496 503 3516
rect 418 3488 503 3496
rect 527 3512 565 3521
rect 527 3492 536 3512
rect 556 3492 565 3512
rect 418 3487 454 3488
rect 527 3484 565 3492
rect 631 3516 716 3522
rect 736 3521 773 3522
rect 631 3496 639 3516
rect 659 3515 716 3516
rect 659 3496 688 3515
rect 631 3495 688 3496
rect 709 3495 716 3515
rect 631 3488 716 3495
rect 735 3512 773 3521
rect 735 3492 744 3512
rect 764 3492 773 3512
rect 631 3487 667 3488
rect 735 3484 773 3492
rect 839 3516 983 3522
rect 839 3496 847 3516
rect 867 3515 955 3516
rect 867 3496 895 3515
rect 839 3494 895 3496
rect 917 3496 955 3515
rect 975 3496 983 3516
rect 917 3494 983 3496
rect 839 3488 983 3494
rect 839 3487 875 3488
rect 947 3487 983 3488
rect 1049 3521 1086 3522
rect 1049 3520 1087 3521
rect 1049 3512 1113 3520
rect 1049 3492 1058 3512
rect 1078 3498 1113 3512
rect 1133 3498 1136 3518
rect 1078 3493 1136 3498
rect 1078 3492 1113 3493
rect 315 3455 352 3484
rect 135 3409 173 3450
rect 316 3453 352 3455
rect 528 3453 565 3484
rect 316 3431 565 3453
rect 736 3452 773 3484
rect 1049 3480 1113 3492
rect 1153 3454 1180 3632
rect 1012 3452 1180 3454
rect 736 3426 1180 3452
rect 737 3409 761 3426
rect 1012 3425 1180 3426
rect 135 3391 762 3409
rect 1388 3405 1638 3429
rect 135 3385 173 3391
rect 135 3361 172 3385
rect 135 3337 170 3361
rect 133 3328 170 3337
rect 133 3310 143 3328
rect 161 3310 170 3328
rect 133 3300 170 3310
rect 1388 3334 1425 3405
rect 1540 3344 1571 3345
rect 1388 3314 1397 3334
rect 1417 3314 1425 3334
rect 1388 3304 1425 3314
rect 1484 3334 1571 3344
rect 1484 3314 1493 3334
rect 1513 3314 1571 3334
rect 1484 3305 1571 3314
rect 1484 3304 1521 3305
rect 1540 3252 1571 3305
rect 1601 3334 1638 3405
rect 1809 3410 2202 3430
rect 2222 3410 2225 3430
rect 1809 3405 2225 3410
rect 1809 3404 2150 3405
rect 1753 3344 1784 3345
rect 1601 3314 1610 3334
rect 1630 3314 1638 3334
rect 1601 3304 1638 3314
rect 1697 3337 1784 3344
rect 1697 3334 1758 3337
rect 1697 3314 1706 3334
rect 1726 3317 1758 3334
rect 1779 3317 1784 3337
rect 1726 3314 1784 3317
rect 1697 3307 1784 3314
rect 1809 3334 1846 3404
rect 2112 3403 2149 3404
rect 1961 3344 1997 3345
rect 1809 3314 1818 3334
rect 1838 3314 1846 3334
rect 1697 3305 1753 3307
rect 1697 3304 1734 3305
rect 1809 3304 1846 3314
rect 1905 3334 2053 3344
rect 2153 3341 2249 3343
rect 1905 3314 1914 3334
rect 1934 3314 2024 3334
rect 2044 3314 2053 3334
rect 1905 3305 2053 3314
rect 2111 3334 2249 3341
rect 2111 3314 2120 3334
rect 2140 3314 2249 3334
rect 2111 3305 2249 3314
rect 1905 3304 1942 3305
rect 1961 3253 1997 3305
rect 2016 3304 2053 3305
rect 2112 3304 2149 3305
rect 1432 3251 1473 3252
rect 1324 3244 1473 3251
rect 136 3236 173 3238
rect 136 3235 784 3236
rect 135 3229 784 3235
rect 135 3211 145 3229
rect 163 3215 784 3229
rect 1324 3224 1442 3244
rect 1462 3224 1473 3244
rect 1324 3216 1473 3224
rect 1540 3248 1899 3252
rect 1540 3243 1862 3248
rect 1540 3219 1653 3243
rect 1677 3224 1862 3243
rect 1886 3224 1899 3248
rect 1677 3219 1899 3224
rect 1540 3216 1899 3219
rect 1961 3216 1996 3253
rect 2064 3250 2164 3253
rect 2064 3246 2131 3250
rect 2064 3220 2076 3246
rect 2102 3224 2131 3246
rect 2157 3224 2164 3250
rect 2102 3220 2164 3224
rect 2064 3216 2164 3220
rect 163 3211 173 3215
rect 614 3214 784 3215
rect 135 3201 173 3211
rect 135 3123 170 3201
rect 747 3191 784 3214
rect 1540 3195 1571 3216
rect 1961 3195 1997 3216
rect 1383 3194 1420 3195
rect 131 3114 170 3123
rect 131 3096 141 3114
rect 159 3096 170 3114
rect 131 3090 170 3096
rect 326 3166 576 3190
rect 326 3095 363 3166
rect 478 3105 509 3106
rect 131 3086 168 3090
rect 326 3075 335 3095
rect 355 3075 363 3095
rect 326 3065 363 3075
rect 422 3095 509 3105
rect 422 3075 431 3095
rect 451 3075 509 3095
rect 422 3066 509 3075
rect 422 3065 459 3066
rect 134 3015 171 3024
rect 132 2997 143 3015
rect 161 2997 171 3015
rect 478 3013 509 3066
rect 539 3095 576 3166
rect 747 3171 1140 3191
rect 1160 3171 1163 3191
rect 747 3166 1163 3171
rect 1382 3185 1420 3194
rect 747 3165 1088 3166
rect 1382 3165 1391 3185
rect 1411 3165 1420 3185
rect 691 3105 722 3106
rect 539 3075 548 3095
rect 568 3075 576 3095
rect 539 3065 576 3075
rect 635 3098 722 3105
rect 635 3095 696 3098
rect 635 3075 644 3095
rect 664 3078 696 3095
rect 717 3078 722 3098
rect 664 3075 722 3078
rect 635 3068 722 3075
rect 747 3095 784 3165
rect 1050 3164 1087 3165
rect 1382 3157 1420 3165
rect 1486 3189 1571 3195
rect 1596 3194 1633 3195
rect 1486 3169 1494 3189
rect 1514 3169 1571 3189
rect 1486 3161 1571 3169
rect 1595 3185 1633 3194
rect 1595 3165 1604 3185
rect 1624 3165 1633 3185
rect 1486 3160 1522 3161
rect 1595 3157 1633 3165
rect 1699 3189 1784 3195
rect 1804 3194 1841 3195
rect 1699 3169 1707 3189
rect 1727 3188 1784 3189
rect 1727 3169 1756 3188
rect 1699 3168 1756 3169
rect 1777 3168 1784 3188
rect 1699 3161 1784 3168
rect 1803 3185 1841 3194
rect 1803 3165 1812 3185
rect 1832 3165 1841 3185
rect 1699 3160 1735 3161
rect 1803 3157 1841 3165
rect 1907 3189 2051 3195
rect 1907 3169 1915 3189
rect 1935 3187 2023 3189
rect 1935 3170 1971 3187
rect 1995 3170 2023 3187
rect 1935 3169 2023 3170
rect 2043 3169 2051 3189
rect 1907 3161 2051 3169
rect 1907 3160 1943 3161
rect 2015 3160 2051 3161
rect 2117 3194 2154 3195
rect 2117 3193 2155 3194
rect 2117 3185 2181 3193
rect 2117 3165 2126 3185
rect 2146 3171 2181 3185
rect 2201 3171 2204 3191
rect 2146 3166 2204 3171
rect 2146 3165 2181 3166
rect 1383 3128 1420 3157
rect 1384 3126 1420 3128
rect 1596 3126 1633 3157
rect 899 3105 935 3106
rect 747 3075 756 3095
rect 776 3075 784 3095
rect 635 3066 691 3068
rect 635 3065 672 3066
rect 747 3065 784 3075
rect 843 3095 991 3105
rect 1384 3104 1633 3126
rect 1804 3125 1841 3157
rect 2117 3153 2181 3165
rect 2221 3127 2248 3305
rect 2080 3125 2248 3127
rect 1804 3114 2248 3125
rect 1091 3102 1187 3104
rect 843 3075 852 3095
rect 872 3075 962 3095
rect 982 3075 991 3095
rect 843 3066 991 3075
rect 1049 3095 1187 3102
rect 1804 3099 2250 3114
rect 2080 3098 2250 3099
rect 1049 3075 1058 3095
rect 1078 3075 1187 3095
rect 1049 3066 1187 3075
rect 843 3065 880 3066
rect 899 3014 935 3066
rect 954 3065 991 3066
rect 1050 3065 1087 3066
rect 370 3012 411 3013
rect 132 2848 171 2997
rect 262 3005 411 3012
rect 262 2985 380 3005
rect 400 2985 411 3005
rect 262 2977 411 2985
rect 478 3009 837 3013
rect 478 3004 800 3009
rect 478 2980 591 3004
rect 615 2985 800 3004
rect 824 2985 837 3009
rect 615 2980 837 2985
rect 478 2977 837 2980
rect 899 2977 934 3014
rect 1002 3011 1102 3014
rect 1002 3007 1069 3011
rect 1002 2981 1014 3007
rect 1040 2985 1069 3007
rect 1095 2985 1102 3011
rect 1040 2981 1102 2985
rect 1002 2977 1102 2981
rect 478 2956 509 2977
rect 899 2956 935 2977
rect 321 2955 358 2956
rect 320 2946 358 2955
rect 320 2926 329 2946
rect 349 2926 358 2946
rect 320 2918 358 2926
rect 424 2950 509 2956
rect 534 2955 571 2956
rect 424 2930 432 2950
rect 452 2930 509 2950
rect 424 2922 509 2930
rect 533 2946 571 2955
rect 533 2926 542 2946
rect 562 2926 571 2946
rect 424 2921 460 2922
rect 533 2918 571 2926
rect 637 2950 722 2956
rect 742 2955 779 2956
rect 637 2930 645 2950
rect 665 2949 722 2950
rect 665 2930 694 2949
rect 637 2929 694 2930
rect 715 2929 722 2949
rect 637 2922 722 2929
rect 741 2946 779 2955
rect 741 2926 750 2946
rect 770 2926 779 2946
rect 637 2921 673 2922
rect 741 2918 779 2926
rect 845 2951 989 2956
rect 845 2950 910 2951
rect 845 2930 853 2950
rect 873 2930 910 2950
rect 932 2950 989 2951
rect 932 2930 961 2950
rect 981 2930 989 2950
rect 845 2922 989 2930
rect 845 2921 881 2922
rect 953 2921 989 2922
rect 1055 2955 1092 2956
rect 1055 2954 1093 2955
rect 1055 2946 1119 2954
rect 1055 2926 1064 2946
rect 1084 2932 1119 2946
rect 1139 2932 1142 2952
rect 1084 2927 1142 2932
rect 1084 2926 1119 2927
rect 321 2889 358 2918
rect 322 2887 358 2889
rect 534 2887 571 2918
rect 322 2865 571 2887
rect 742 2886 779 2918
rect 1055 2914 1119 2926
rect 1159 2888 1186 3066
rect 1018 2886 1186 2888
rect 742 2860 1186 2886
rect 1338 2985 1588 3009
rect 1338 2914 1375 2985
rect 1490 2924 1521 2925
rect 1338 2894 1347 2914
rect 1367 2894 1375 2914
rect 1338 2884 1375 2894
rect 1434 2914 1521 2924
rect 1434 2894 1443 2914
rect 1463 2894 1521 2914
rect 1434 2885 1521 2894
rect 1434 2884 1471 2885
rect 742 2850 764 2860
rect 1018 2859 1186 2860
rect 702 2848 764 2850
rect 132 2841 764 2848
rect 131 2832 764 2841
rect 1490 2832 1521 2885
rect 1551 2914 1588 2985
rect 1759 2990 2152 3010
rect 2172 2990 2175 3010
rect 1759 2985 2175 2990
rect 1759 2984 2100 2985
rect 1703 2924 1734 2925
rect 1551 2894 1560 2914
rect 1580 2894 1588 2914
rect 1551 2884 1588 2894
rect 1647 2917 1734 2924
rect 1647 2914 1708 2917
rect 1647 2894 1656 2914
rect 1676 2897 1708 2914
rect 1729 2897 1734 2917
rect 1676 2894 1734 2897
rect 1647 2887 1734 2894
rect 1759 2914 1796 2984
rect 2062 2983 2099 2984
rect 1911 2924 1947 2925
rect 1759 2894 1768 2914
rect 1788 2894 1796 2914
rect 1647 2885 1703 2887
rect 1647 2884 1684 2885
rect 1759 2884 1796 2894
rect 1855 2914 2003 2924
rect 2103 2921 2199 2923
rect 1855 2894 1864 2914
rect 1884 2894 1974 2914
rect 1994 2894 2003 2914
rect 1855 2885 2003 2894
rect 2061 2914 2199 2921
rect 2061 2894 2070 2914
rect 2090 2894 2199 2914
rect 2061 2885 2199 2894
rect 1855 2884 1892 2885
rect 1911 2833 1947 2885
rect 1966 2884 2003 2885
rect 2062 2884 2099 2885
rect 131 2814 141 2832
rect 159 2831 764 2832
rect 1382 2831 1423 2832
rect 159 2826 180 2831
rect 159 2814 171 2826
rect 1274 2824 1423 2831
rect 131 2806 171 2814
rect 214 2813 240 2814
rect 131 2804 168 2806
rect 214 2795 768 2813
rect 1274 2804 1392 2824
rect 1412 2804 1423 2824
rect 1274 2796 1423 2804
rect 1490 2828 1849 2832
rect 1490 2823 1812 2828
rect 1490 2799 1603 2823
rect 1627 2804 1812 2823
rect 1836 2804 1849 2828
rect 1627 2799 1849 2804
rect 1490 2796 1849 2799
rect 1911 2796 1946 2833
rect 2014 2830 2114 2833
rect 2014 2826 2081 2830
rect 2014 2800 2026 2826
rect 2052 2804 2081 2826
rect 2107 2804 2114 2830
rect 2052 2800 2114 2804
rect 2014 2796 2114 2800
rect 134 2736 171 2742
rect 214 2736 240 2795
rect 747 2776 768 2795
rect 134 2733 240 2736
rect 134 2715 143 2733
rect 161 2719 240 2733
rect 325 2751 575 2775
rect 161 2717 237 2719
rect 161 2715 171 2717
rect 134 2705 171 2715
rect 139 2640 170 2705
rect 325 2680 362 2751
rect 477 2690 508 2691
rect 325 2660 334 2680
rect 354 2660 362 2680
rect 325 2650 362 2660
rect 421 2680 508 2690
rect 421 2660 430 2680
rect 450 2660 508 2680
rect 421 2651 508 2660
rect 421 2650 458 2651
rect 138 2631 175 2640
rect 138 2613 148 2631
rect 166 2613 175 2631
rect 138 2603 175 2613
rect 477 2598 508 2651
rect 538 2680 575 2751
rect 746 2756 1139 2776
rect 1159 2756 1162 2776
rect 1490 2775 1521 2796
rect 1911 2775 1947 2796
rect 1333 2774 1370 2775
rect 746 2751 1162 2756
rect 1332 2765 1370 2774
rect 746 2750 1087 2751
rect 690 2690 721 2691
rect 538 2660 547 2680
rect 567 2660 575 2680
rect 538 2650 575 2660
rect 634 2683 721 2690
rect 634 2680 695 2683
rect 634 2660 643 2680
rect 663 2663 695 2680
rect 716 2663 721 2683
rect 663 2660 721 2663
rect 634 2653 721 2660
rect 746 2680 783 2750
rect 1049 2749 1086 2750
rect 1332 2745 1341 2765
rect 1361 2745 1370 2765
rect 1332 2737 1370 2745
rect 1436 2769 1521 2775
rect 1546 2774 1583 2775
rect 1436 2749 1444 2769
rect 1464 2749 1521 2769
rect 1436 2741 1521 2749
rect 1545 2765 1583 2774
rect 1545 2745 1554 2765
rect 1574 2745 1583 2765
rect 1436 2740 1472 2741
rect 1545 2737 1583 2745
rect 1649 2769 1734 2775
rect 1754 2774 1791 2775
rect 1649 2749 1657 2769
rect 1677 2768 1734 2769
rect 1677 2749 1706 2768
rect 1649 2748 1706 2749
rect 1727 2748 1734 2768
rect 1649 2741 1734 2748
rect 1753 2765 1791 2774
rect 1753 2745 1762 2765
rect 1782 2745 1791 2765
rect 1649 2740 1685 2741
rect 1753 2737 1791 2745
rect 1857 2770 2001 2775
rect 1857 2769 1916 2770
rect 1857 2749 1865 2769
rect 1885 2750 1916 2769
rect 1940 2769 2001 2770
rect 1940 2750 1973 2769
rect 1885 2749 1973 2750
rect 1993 2749 2001 2769
rect 1857 2741 2001 2749
rect 1857 2740 1893 2741
rect 1965 2740 2001 2741
rect 2067 2774 2104 2775
rect 2067 2773 2105 2774
rect 2067 2765 2131 2773
rect 2067 2745 2076 2765
rect 2096 2751 2131 2765
rect 2151 2751 2154 2771
rect 2096 2746 2154 2751
rect 2096 2745 2131 2746
rect 1333 2708 1370 2737
rect 1334 2706 1370 2708
rect 1546 2706 1583 2737
rect 898 2690 934 2691
rect 746 2660 755 2680
rect 775 2660 783 2680
rect 634 2651 690 2653
rect 634 2650 671 2651
rect 746 2650 783 2660
rect 842 2680 990 2690
rect 1090 2687 1186 2689
rect 842 2660 851 2680
rect 871 2660 961 2680
rect 981 2660 990 2680
rect 842 2651 990 2660
rect 1048 2680 1186 2687
rect 1334 2684 1583 2706
rect 1754 2705 1791 2737
rect 2067 2733 2131 2745
rect 2171 2707 2198 2885
rect 2030 2705 2198 2707
rect 1754 2701 2198 2705
rect 1048 2660 1057 2680
rect 1077 2660 1186 2680
rect 1754 2682 1803 2701
rect 1823 2682 2198 2701
rect 1754 2679 2198 2682
rect 2030 2678 2198 2679
rect 2219 2704 2250 3098
rect 2219 2678 2224 2704
rect 2243 2678 2250 2704
rect 2219 2675 2250 2678
rect 1048 2651 1186 2660
rect 842 2650 879 2651
rect 898 2599 934 2651
rect 953 2650 990 2651
rect 1049 2650 1086 2651
rect 369 2597 410 2598
rect 261 2590 410 2597
rect 261 2570 379 2590
rect 399 2570 410 2590
rect 261 2562 410 2570
rect 477 2594 836 2598
rect 477 2589 799 2594
rect 477 2565 590 2589
rect 614 2570 799 2589
rect 823 2570 836 2594
rect 614 2565 836 2570
rect 477 2562 836 2565
rect 898 2562 933 2599
rect 1001 2596 1101 2599
rect 1001 2592 1068 2596
rect 1001 2566 1013 2592
rect 1039 2570 1068 2592
rect 1094 2570 1101 2596
rect 1039 2566 1101 2570
rect 1001 2562 1101 2566
rect 477 2541 508 2562
rect 898 2541 934 2562
rect 141 2532 178 2541
rect 320 2540 357 2541
rect 141 2514 150 2532
rect 168 2514 178 2532
rect 141 2504 178 2514
rect 142 2469 178 2504
rect 319 2531 357 2540
rect 319 2511 328 2531
rect 348 2511 357 2531
rect 319 2503 357 2511
rect 423 2535 508 2541
rect 533 2540 570 2541
rect 423 2515 431 2535
rect 451 2515 508 2535
rect 423 2507 508 2515
rect 532 2531 570 2540
rect 532 2511 541 2531
rect 561 2511 570 2531
rect 423 2506 459 2507
rect 532 2503 570 2511
rect 636 2535 721 2541
rect 741 2540 778 2541
rect 636 2515 644 2535
rect 664 2534 721 2535
rect 664 2515 693 2534
rect 636 2514 693 2515
rect 714 2514 721 2534
rect 636 2507 721 2514
rect 740 2531 778 2540
rect 740 2511 749 2531
rect 769 2511 778 2531
rect 636 2506 672 2507
rect 740 2503 778 2511
rect 844 2535 988 2541
rect 844 2515 852 2535
rect 872 2534 960 2535
rect 872 2515 900 2534
rect 844 2513 900 2515
rect 922 2515 960 2534
rect 980 2515 988 2535
rect 922 2513 988 2515
rect 844 2507 988 2513
rect 844 2506 880 2507
rect 952 2506 988 2507
rect 1054 2540 1091 2541
rect 1054 2539 1092 2540
rect 1054 2531 1118 2539
rect 1054 2511 1063 2531
rect 1083 2517 1118 2531
rect 1138 2517 1141 2537
rect 1083 2512 1141 2517
rect 1083 2511 1118 2512
rect 320 2474 357 2503
rect 140 2428 178 2469
rect 321 2472 357 2474
rect 533 2472 570 2503
rect 321 2450 570 2472
rect 741 2471 778 2503
rect 1054 2499 1118 2511
rect 1158 2473 1185 2651
rect 1017 2471 1185 2473
rect 741 2445 1185 2471
rect 742 2428 766 2445
rect 1017 2444 1185 2445
rect 1553 2473 1803 2497
rect 140 2410 767 2428
rect 140 2404 178 2410
rect 142 2358 177 2404
rect 1553 2402 1590 2473
rect 1705 2412 1736 2413
rect 1553 2382 1562 2402
rect 1582 2382 1590 2402
rect 1553 2372 1590 2382
rect 1649 2402 1736 2412
rect 1649 2382 1658 2402
rect 1678 2382 1736 2402
rect 1649 2373 1736 2382
rect 1649 2372 1686 2373
rect 140 2349 177 2358
rect 140 2331 150 2349
rect 168 2331 177 2349
rect 140 2321 177 2331
rect 1705 2320 1736 2373
rect 1766 2402 1803 2473
rect 1974 2478 2367 2498
rect 2387 2478 2390 2498
rect 1974 2473 2390 2478
rect 1974 2472 2315 2473
rect 1918 2412 1949 2413
rect 1766 2382 1775 2402
rect 1795 2382 1803 2402
rect 1766 2372 1803 2382
rect 1862 2405 1949 2412
rect 1862 2402 1923 2405
rect 1862 2382 1871 2402
rect 1891 2385 1923 2402
rect 1944 2385 1949 2405
rect 1891 2382 1949 2385
rect 1862 2375 1949 2382
rect 1974 2402 2011 2472
rect 2277 2471 2314 2472
rect 2126 2412 2162 2413
rect 1974 2382 1983 2402
rect 2003 2382 2011 2402
rect 1862 2373 1918 2375
rect 1862 2372 1899 2373
rect 1974 2372 2011 2382
rect 2070 2402 2218 2412
rect 2318 2409 2414 2411
rect 2070 2382 2079 2402
rect 2099 2382 2189 2402
rect 2209 2382 2218 2402
rect 2070 2373 2218 2382
rect 2276 2402 2414 2409
rect 2276 2382 2285 2402
rect 2305 2382 2414 2402
rect 2276 2373 2414 2382
rect 2070 2372 2107 2373
rect 2126 2321 2162 2373
rect 2181 2372 2218 2373
rect 2277 2372 2314 2373
rect 1597 2319 1638 2320
rect 1489 2312 1638 2319
rect 1489 2292 1607 2312
rect 1627 2292 1638 2312
rect 1489 2284 1638 2292
rect 1705 2316 2064 2320
rect 1705 2311 2027 2316
rect 1705 2287 1818 2311
rect 1842 2292 2027 2311
rect 2051 2292 2064 2316
rect 1842 2287 2064 2292
rect 1705 2284 2064 2287
rect 2126 2284 2161 2321
rect 2229 2318 2329 2321
rect 2229 2314 2296 2318
rect 2229 2288 2241 2314
rect 2267 2292 2296 2314
rect 2322 2292 2329 2318
rect 2267 2288 2329 2292
rect 2229 2284 2329 2288
rect 1705 2263 1736 2284
rect 2126 2263 2162 2284
rect 1548 2262 1585 2263
rect 143 2257 180 2259
rect 143 2256 791 2257
rect 142 2250 791 2256
rect 142 2232 152 2250
rect 170 2236 791 2250
rect 170 2232 180 2236
rect 621 2235 791 2236
rect 142 2222 180 2232
rect 142 2144 177 2222
rect 754 2212 791 2235
rect 1547 2253 1585 2262
rect 1547 2233 1556 2253
rect 1576 2233 1585 2253
rect 1547 2225 1585 2233
rect 1651 2257 1736 2263
rect 1761 2262 1798 2263
rect 1651 2237 1659 2257
rect 1679 2237 1736 2257
rect 1651 2229 1736 2237
rect 1760 2253 1798 2262
rect 1760 2233 1769 2253
rect 1789 2233 1798 2253
rect 1651 2228 1687 2229
rect 1760 2225 1798 2233
rect 1864 2257 1949 2263
rect 1969 2262 2006 2263
rect 1864 2237 1872 2257
rect 1892 2256 1949 2257
rect 1892 2237 1921 2256
rect 1864 2236 1921 2237
rect 1942 2236 1949 2256
rect 1864 2229 1949 2236
rect 1968 2253 2006 2262
rect 1968 2233 1977 2253
rect 1997 2233 2006 2253
rect 1864 2228 1900 2229
rect 1968 2225 2006 2233
rect 2072 2257 2216 2263
rect 2072 2237 2080 2257
rect 2100 2238 2136 2257
rect 2159 2238 2188 2257
rect 2100 2237 2188 2238
rect 2208 2237 2216 2257
rect 2072 2229 2216 2237
rect 2072 2228 2108 2229
rect 2180 2228 2216 2229
rect 2282 2262 2319 2263
rect 2282 2261 2320 2262
rect 2282 2253 2346 2261
rect 2282 2233 2291 2253
rect 2311 2239 2346 2253
rect 2366 2239 2369 2259
rect 2311 2234 2369 2239
rect 2311 2233 2346 2234
rect 138 2135 177 2144
rect 138 2117 148 2135
rect 166 2117 177 2135
rect 138 2111 177 2117
rect 333 2187 583 2211
rect 333 2116 370 2187
rect 485 2126 516 2127
rect 138 2107 175 2111
rect 333 2096 342 2116
rect 362 2096 370 2116
rect 333 2086 370 2096
rect 429 2116 516 2126
rect 429 2096 438 2116
rect 458 2096 516 2116
rect 429 2087 516 2096
rect 429 2086 466 2087
rect 141 2036 178 2045
rect 139 2018 150 2036
rect 168 2018 178 2036
rect 485 2034 516 2087
rect 546 2116 583 2187
rect 754 2192 1147 2212
rect 1167 2192 1170 2212
rect 1548 2196 1585 2225
rect 754 2187 1170 2192
rect 1549 2194 1585 2196
rect 1761 2194 1798 2225
rect 754 2186 1095 2187
rect 698 2126 729 2127
rect 546 2096 555 2116
rect 575 2096 583 2116
rect 546 2086 583 2096
rect 642 2119 729 2126
rect 642 2116 703 2119
rect 642 2096 651 2116
rect 671 2099 703 2116
rect 724 2099 729 2119
rect 671 2096 729 2099
rect 642 2089 729 2096
rect 754 2116 791 2186
rect 1057 2185 1094 2186
rect 1549 2172 1798 2194
rect 1969 2193 2006 2225
rect 2282 2221 2346 2233
rect 2386 2195 2413 2373
rect 2441 2260 2479 4091
rect 2986 4066 2993 4092
rect 3012 4066 3017 4092
rect 2893 3673 2922 3675
rect 2893 3668 2925 3673
rect 2893 3650 2900 3668
rect 2920 3650 2925 3668
rect 2986 3672 3017 4066
rect 3038 4091 3206 4092
rect 3038 4088 3482 4091
rect 3038 4069 3413 4088
rect 3433 4069 3482 4088
rect 4050 4090 4159 4110
rect 4179 4090 4188 4110
rect 3038 4065 3482 4069
rect 3038 4063 3206 4065
rect 3038 3885 3065 4063
rect 3105 4025 3169 4037
rect 3445 4033 3482 4065
rect 3653 4064 3902 4086
rect 4050 4083 4188 4090
rect 4246 4110 4394 4119
rect 4246 4090 4255 4110
rect 4275 4090 4365 4110
rect 4385 4090 4394 4110
rect 4050 4081 4146 4083
rect 4246 4080 4394 4090
rect 4453 4110 4490 4120
rect 4565 4119 4602 4120
rect 4546 4117 4602 4119
rect 4453 4090 4461 4110
rect 4481 4090 4490 4110
rect 4302 4079 4338 4080
rect 3653 4033 3690 4064
rect 3866 4062 3902 4064
rect 3866 4033 3903 4062
rect 3105 4024 3140 4025
rect 3082 4019 3140 4024
rect 3082 3999 3085 4019
rect 3105 4005 3140 4019
rect 3160 4005 3169 4025
rect 3105 3997 3169 4005
rect 3131 3996 3169 3997
rect 3132 3995 3169 3996
rect 3235 4029 3271 4030
rect 3343 4029 3379 4030
rect 3235 4021 3379 4029
rect 3235 4001 3243 4021
rect 3263 4020 3351 4021
rect 3263 4001 3296 4020
rect 3235 4000 3296 4001
rect 3320 4001 3351 4020
rect 3371 4001 3379 4021
rect 3320 4000 3379 4001
rect 3235 3995 3379 4000
rect 3445 4025 3483 4033
rect 3551 4029 3587 4030
rect 3445 4005 3454 4025
rect 3474 4005 3483 4025
rect 3445 3996 3483 4005
rect 3502 4022 3587 4029
rect 3502 4002 3509 4022
rect 3530 4021 3587 4022
rect 3530 4002 3559 4021
rect 3502 4001 3559 4002
rect 3579 4001 3587 4021
rect 3445 3995 3482 3996
rect 3502 3995 3587 4001
rect 3653 4025 3691 4033
rect 3764 4029 3800 4030
rect 3653 4005 3662 4025
rect 3682 4005 3691 4025
rect 3653 3996 3691 4005
rect 3715 4021 3800 4029
rect 3715 4001 3772 4021
rect 3792 4001 3800 4021
rect 3653 3995 3690 3996
rect 3715 3995 3800 4001
rect 3866 4025 3904 4033
rect 3866 4005 3875 4025
rect 3895 4005 3904 4025
rect 4150 4020 4187 4021
rect 4453 4020 4490 4090
rect 4515 4110 4602 4117
rect 4515 4107 4573 4110
rect 4515 4087 4520 4107
rect 4541 4090 4573 4107
rect 4593 4090 4602 4110
rect 4541 4087 4602 4090
rect 4515 4080 4602 4087
rect 4661 4110 4698 4120
rect 4661 4090 4669 4110
rect 4689 4090 4698 4110
rect 4515 4079 4546 4080
rect 4149 4019 4490 4020
rect 3866 3996 3904 4005
rect 4074 4014 4490 4019
rect 3866 3995 3903 3996
rect 3289 3974 3325 3995
rect 3715 3974 3746 3995
rect 4074 3994 4077 4014
rect 4097 3994 4490 4014
rect 4661 4019 4698 4090
rect 4728 4119 4759 4172
rect 5411 4171 5421 4189
rect 5439 4175 6060 4189
rect 6845 4188 6994 4196
rect 7061 4220 7420 4224
rect 7061 4215 7383 4220
rect 7061 4191 7174 4215
rect 7198 4196 7383 4215
rect 7407 4196 7420 4220
rect 7198 4191 7420 4196
rect 7061 4188 7420 4191
rect 7482 4188 7517 4225
rect 7585 4222 7685 4225
rect 7585 4218 7652 4222
rect 7585 4192 7597 4218
rect 7623 4196 7652 4218
rect 7678 4196 7685 4222
rect 7623 4192 7685 4196
rect 7585 4188 7685 4192
rect 5439 4171 5449 4175
rect 5890 4174 6060 4175
rect 5061 4157 5098 4167
rect 5061 4139 5070 4157
rect 5088 4139 5098 4157
rect 5061 4130 5098 4139
rect 5411 4161 5449 4171
rect 4778 4119 4815 4120
rect 4728 4110 4815 4119
rect 4728 4090 4786 4110
rect 4806 4090 4815 4110
rect 4728 4080 4815 4090
rect 4874 4110 4911 4120
rect 4874 4090 4882 4110
rect 4902 4090 4911 4110
rect 4728 4079 4759 4080
rect 4874 4019 4911 4090
rect 5066 4065 5097 4130
rect 5411 4083 5446 4161
rect 6023 4151 6060 4174
rect 7061 4167 7092 4188
rect 7482 4167 7518 4188
rect 6904 4166 6941 4167
rect 6903 4157 6941 4166
rect 5407 4074 5446 4083
rect 5065 4055 5102 4065
rect 5065 4053 5075 4055
rect 4999 4051 5075 4053
rect 4661 3995 4911 4019
rect 4996 4037 5075 4051
rect 5093 4037 5102 4055
rect 5407 4056 5417 4074
rect 5435 4056 5446 4074
rect 5407 4050 5446 4056
rect 5602 4126 5852 4150
rect 5602 4055 5639 4126
rect 5754 4065 5785 4066
rect 5407 4046 5444 4050
rect 4996 4034 5102 4037
rect 4468 3975 4489 3994
rect 4996 3975 5022 4034
rect 5065 4028 5102 4034
rect 5602 4035 5611 4055
rect 5631 4035 5639 4055
rect 5602 4025 5639 4035
rect 5698 4055 5785 4065
rect 5698 4035 5707 4055
rect 5727 4035 5785 4055
rect 5698 4026 5785 4035
rect 5698 4025 5735 4026
rect 5410 3975 5447 3984
rect 3122 3970 3222 3974
rect 3122 3966 3184 3970
rect 3122 3940 3129 3966
rect 3155 3944 3184 3966
rect 3210 3944 3222 3970
rect 3155 3940 3222 3944
rect 3122 3937 3222 3940
rect 3290 3937 3325 3974
rect 3387 3971 3746 3974
rect 3387 3966 3609 3971
rect 3387 3942 3400 3966
rect 3424 3947 3609 3966
rect 3633 3947 3746 3971
rect 3424 3942 3746 3947
rect 3387 3938 3746 3942
rect 3813 3966 3962 3974
rect 3813 3946 3824 3966
rect 3844 3946 3962 3966
rect 4468 3957 5022 3975
rect 5068 3964 5105 3966
rect 4996 3956 5022 3957
rect 5065 3956 5105 3964
rect 3813 3939 3962 3946
rect 5065 3944 5077 3956
rect 5056 3939 5077 3944
rect 3813 3938 3854 3939
rect 4472 3938 5077 3939
rect 5095 3938 5105 3956
rect 3137 3885 3174 3886
rect 3233 3885 3270 3886
rect 3289 3885 3325 3937
rect 3344 3885 3381 3886
rect 3037 3876 3175 3885
rect 3037 3856 3146 3876
rect 3166 3856 3175 3876
rect 3037 3849 3175 3856
rect 3233 3876 3381 3885
rect 3233 3856 3242 3876
rect 3262 3856 3352 3876
rect 3372 3856 3381 3876
rect 3037 3847 3133 3849
rect 3233 3846 3381 3856
rect 3440 3876 3477 3886
rect 3552 3885 3589 3886
rect 3533 3883 3589 3885
rect 3440 3856 3448 3876
rect 3468 3856 3477 3876
rect 3289 3845 3325 3846
rect 3137 3786 3174 3787
rect 3440 3786 3477 3856
rect 3502 3876 3589 3883
rect 3502 3873 3560 3876
rect 3502 3853 3507 3873
rect 3528 3856 3560 3873
rect 3580 3856 3589 3876
rect 3528 3853 3589 3856
rect 3502 3846 3589 3853
rect 3648 3876 3685 3886
rect 3648 3856 3656 3876
rect 3676 3856 3685 3876
rect 3502 3845 3533 3846
rect 3136 3785 3477 3786
rect 3061 3780 3477 3785
rect 3061 3760 3064 3780
rect 3084 3760 3477 3780
rect 3648 3785 3685 3856
rect 3715 3885 3746 3938
rect 4472 3929 5105 3938
rect 5408 3957 5419 3975
rect 5437 3957 5447 3975
rect 5754 3973 5785 4026
rect 5815 4055 5852 4126
rect 6023 4131 6416 4151
rect 6436 4131 6439 4151
rect 6023 4126 6439 4131
rect 6903 4137 6912 4157
rect 6932 4137 6941 4157
rect 6903 4129 6941 4137
rect 7007 4161 7092 4167
rect 7117 4166 7154 4167
rect 7007 4141 7015 4161
rect 7035 4141 7092 4161
rect 7007 4133 7092 4141
rect 7116 4157 7154 4166
rect 7116 4137 7125 4157
rect 7145 4137 7154 4157
rect 7007 4132 7043 4133
rect 7116 4129 7154 4137
rect 7220 4161 7305 4167
rect 7325 4166 7362 4167
rect 7220 4141 7228 4161
rect 7248 4160 7305 4161
rect 7248 4141 7277 4160
rect 7220 4140 7277 4141
rect 7298 4140 7305 4160
rect 7220 4133 7305 4140
rect 7324 4157 7362 4166
rect 7324 4137 7333 4157
rect 7353 4137 7362 4157
rect 7220 4132 7256 4133
rect 7324 4129 7362 4137
rect 7428 4162 7572 4167
rect 7428 4161 7492 4162
rect 7428 4141 7436 4161
rect 7456 4143 7492 4161
rect 7518 4161 7572 4162
rect 7518 4143 7544 4161
rect 7456 4141 7544 4143
rect 7564 4141 7572 4161
rect 7428 4133 7572 4141
rect 7428 4132 7464 4133
rect 7536 4132 7572 4133
rect 7638 4166 7675 4167
rect 7638 4165 7676 4166
rect 7638 4157 7702 4165
rect 7638 4137 7647 4157
rect 7667 4143 7702 4157
rect 7722 4143 7725 4163
rect 7667 4138 7725 4143
rect 7667 4137 7702 4138
rect 6023 4125 6364 4126
rect 5967 4065 5998 4066
rect 5815 4035 5824 4055
rect 5844 4035 5852 4055
rect 5815 4025 5852 4035
rect 5911 4058 5998 4065
rect 5911 4055 5972 4058
rect 5911 4035 5920 4055
rect 5940 4038 5972 4055
rect 5993 4038 5998 4058
rect 5940 4035 5998 4038
rect 5911 4028 5998 4035
rect 6023 4055 6060 4125
rect 6326 4124 6363 4125
rect 6904 4100 6941 4129
rect 6905 4098 6941 4100
rect 7117 4098 7154 4129
rect 6905 4076 7154 4098
rect 7325 4097 7362 4129
rect 7638 4125 7702 4137
rect 7742 4102 7769 4277
rect 7722 4099 7769 4102
rect 7601 4097 7769 4099
rect 9332 4276 9500 4278
rect 9332 4098 9359 4276
rect 9399 4238 9463 4250
rect 9739 4246 9776 4278
rect 9947 4277 10196 4299
rect 9947 4246 9984 4277
rect 10160 4275 10196 4277
rect 10339 4280 10377 4321
rect 10160 4246 10197 4275
rect 9399 4237 9434 4238
rect 9376 4232 9434 4237
rect 9376 4212 9379 4232
rect 9399 4218 9434 4232
rect 9454 4218 9463 4238
rect 9399 4210 9463 4218
rect 9425 4209 9463 4210
rect 9426 4208 9463 4209
rect 9529 4242 9565 4243
rect 9637 4242 9673 4243
rect 9529 4236 9673 4242
rect 9529 4234 9595 4236
rect 9529 4214 9537 4234
rect 9557 4215 9595 4234
rect 9617 4234 9673 4236
rect 9617 4215 9645 4234
rect 9557 4214 9645 4215
rect 9665 4214 9673 4234
rect 9529 4208 9673 4214
rect 9739 4238 9777 4246
rect 9845 4242 9881 4243
rect 9739 4218 9748 4238
rect 9768 4218 9777 4238
rect 9739 4209 9777 4218
rect 9796 4235 9881 4242
rect 9796 4215 9803 4235
rect 9824 4234 9881 4235
rect 9824 4215 9853 4234
rect 9796 4214 9853 4215
rect 9873 4214 9881 4234
rect 9739 4208 9776 4209
rect 9796 4208 9881 4214
rect 9947 4238 9985 4246
rect 10058 4242 10094 4243
rect 9947 4218 9956 4238
rect 9976 4218 9985 4238
rect 9947 4209 9985 4218
rect 10009 4234 10094 4242
rect 10009 4214 10066 4234
rect 10086 4214 10094 4234
rect 9947 4208 9984 4209
rect 10009 4208 10094 4214
rect 10160 4238 10198 4246
rect 10160 4218 10169 4238
rect 10189 4218 10198 4238
rect 10160 4209 10198 4218
rect 10339 4245 10375 4280
rect 10339 4235 10376 4245
rect 10339 4217 10349 4235
rect 10367 4217 10376 4235
rect 10160 4208 10197 4209
rect 10339 4208 10376 4217
rect 9583 4187 9619 4208
rect 10009 4187 10040 4208
rect 9416 4183 9516 4187
rect 9416 4179 9478 4183
rect 9416 4153 9423 4179
rect 9449 4157 9478 4179
rect 9504 4157 9516 4183
rect 9449 4153 9516 4157
rect 9416 4150 9516 4153
rect 9584 4150 9619 4187
rect 9681 4184 10040 4187
rect 9681 4179 9903 4184
rect 9681 4155 9694 4179
rect 9718 4160 9903 4179
rect 9927 4160 10040 4184
rect 9718 4155 10040 4160
rect 9681 4151 10040 4155
rect 10107 4179 10256 4187
rect 10107 4159 10118 4179
rect 10138 4159 10256 4179
rect 10107 4152 10256 4159
rect 10107 4151 10148 4152
rect 9431 4098 9468 4099
rect 9527 4098 9564 4099
rect 9583 4098 9619 4150
rect 9638 4098 9675 4099
rect 7325 4071 7769 4097
rect 9331 4089 9469 4098
rect 7601 4070 7769 4071
rect 8267 4071 8298 4074
rect 6175 4065 6211 4066
rect 6023 4035 6032 4055
rect 6052 4035 6060 4055
rect 5911 4026 5967 4028
rect 5911 4025 5948 4026
rect 6023 4025 6060 4035
rect 6119 4055 6267 4065
rect 6367 4062 6463 4064
rect 6119 4035 6128 4055
rect 6148 4035 6238 4055
rect 6258 4035 6267 4055
rect 6119 4026 6267 4035
rect 6325 4055 6463 4062
rect 6325 4035 6334 4055
rect 6354 4035 6463 4055
rect 6325 4026 6463 4035
rect 6119 4025 6156 4026
rect 6175 3974 6211 4026
rect 6230 4025 6267 4026
rect 6326 4025 6363 4026
rect 5646 3972 5687 3973
rect 4472 3922 5104 3929
rect 4472 3920 4534 3922
rect 4050 3910 4218 3911
rect 4472 3910 4494 3920
rect 3765 3885 3802 3886
rect 3715 3876 3802 3885
rect 3715 3856 3773 3876
rect 3793 3856 3802 3876
rect 3715 3846 3802 3856
rect 3861 3876 3898 3886
rect 3861 3856 3869 3876
rect 3889 3856 3898 3876
rect 3715 3845 3746 3846
rect 3861 3785 3898 3856
rect 3648 3761 3898 3785
rect 4050 3884 4494 3910
rect 4050 3882 4218 3884
rect 4050 3704 4077 3882
rect 4117 3844 4181 3856
rect 4457 3852 4494 3884
rect 4665 3883 4914 3905
rect 4665 3852 4702 3883
rect 4878 3881 4914 3883
rect 4878 3852 4915 3881
rect 4117 3843 4152 3844
rect 4094 3838 4152 3843
rect 4094 3818 4097 3838
rect 4117 3824 4152 3838
rect 4172 3824 4181 3844
rect 4117 3816 4181 3824
rect 4143 3815 4181 3816
rect 4144 3814 4181 3815
rect 4247 3848 4283 3849
rect 4355 3848 4391 3849
rect 4247 3840 4391 3848
rect 4247 3820 4255 3840
rect 4275 3820 4304 3840
rect 4247 3819 4304 3820
rect 4326 3820 4363 3840
rect 4383 3820 4391 3840
rect 4326 3819 4391 3820
rect 4247 3814 4391 3819
rect 4457 3844 4495 3852
rect 4563 3848 4599 3849
rect 4457 3824 4466 3844
rect 4486 3824 4495 3844
rect 4457 3815 4495 3824
rect 4514 3841 4599 3848
rect 4514 3821 4521 3841
rect 4542 3840 4599 3841
rect 4542 3821 4571 3840
rect 4514 3820 4571 3821
rect 4591 3820 4599 3840
rect 4457 3814 4494 3815
rect 4514 3814 4599 3820
rect 4665 3844 4703 3852
rect 4776 3848 4812 3849
rect 4665 3824 4674 3844
rect 4694 3824 4703 3844
rect 4665 3815 4703 3824
rect 4727 3840 4812 3848
rect 4727 3820 4784 3840
rect 4804 3820 4812 3840
rect 4665 3814 4702 3815
rect 4727 3814 4812 3820
rect 4878 3844 4916 3852
rect 4878 3824 4887 3844
rect 4907 3824 4916 3844
rect 4878 3815 4916 3824
rect 4878 3814 4915 3815
rect 4301 3793 4337 3814
rect 4727 3793 4758 3814
rect 4134 3789 4234 3793
rect 4134 3785 4196 3789
rect 4134 3759 4141 3785
rect 4167 3763 4196 3785
rect 4222 3763 4234 3789
rect 4167 3759 4234 3763
rect 4134 3756 4234 3759
rect 4302 3756 4337 3793
rect 4399 3790 4758 3793
rect 4399 3785 4621 3790
rect 4399 3761 4412 3785
rect 4436 3766 4621 3785
rect 4645 3766 4758 3790
rect 4436 3761 4758 3766
rect 4399 3757 4758 3761
rect 4825 3785 4974 3793
rect 4825 3765 4836 3785
rect 4856 3765 4974 3785
rect 4825 3758 4974 3765
rect 5065 3773 5104 3922
rect 5408 3808 5447 3957
rect 5538 3965 5687 3972
rect 5538 3945 5656 3965
rect 5676 3945 5687 3965
rect 5538 3937 5687 3945
rect 5754 3969 6113 3973
rect 5754 3964 6076 3969
rect 5754 3940 5867 3964
rect 5891 3945 6076 3964
rect 6100 3945 6113 3969
rect 5891 3940 6113 3945
rect 5754 3937 6113 3940
rect 6175 3937 6210 3974
rect 6278 3971 6378 3974
rect 6278 3967 6345 3971
rect 6278 3941 6290 3967
rect 6316 3945 6345 3967
rect 6371 3945 6378 3971
rect 6316 3941 6378 3945
rect 6278 3937 6378 3941
rect 5754 3916 5785 3937
rect 6175 3916 6211 3937
rect 5597 3915 5634 3916
rect 5596 3906 5634 3915
rect 5596 3886 5605 3906
rect 5625 3886 5634 3906
rect 5596 3878 5634 3886
rect 5700 3910 5785 3916
rect 5810 3915 5847 3916
rect 5700 3890 5708 3910
rect 5728 3890 5785 3910
rect 5700 3882 5785 3890
rect 5809 3906 5847 3915
rect 5809 3886 5818 3906
rect 5838 3886 5847 3906
rect 5700 3881 5736 3882
rect 5809 3878 5847 3886
rect 5913 3910 5998 3916
rect 6018 3915 6055 3916
rect 5913 3890 5921 3910
rect 5941 3909 5998 3910
rect 5941 3890 5970 3909
rect 5913 3889 5970 3890
rect 5991 3889 5998 3909
rect 5913 3882 5998 3889
rect 6017 3906 6055 3915
rect 6017 3886 6026 3906
rect 6046 3886 6055 3906
rect 5913 3881 5949 3882
rect 6017 3878 6055 3886
rect 6121 3911 6265 3916
rect 6121 3910 6186 3911
rect 6121 3890 6129 3910
rect 6149 3890 6186 3910
rect 6208 3910 6265 3911
rect 6208 3890 6237 3910
rect 6257 3890 6265 3910
rect 6121 3882 6265 3890
rect 6121 3881 6157 3882
rect 6229 3881 6265 3882
rect 6331 3915 6368 3916
rect 6331 3914 6369 3915
rect 6331 3906 6395 3914
rect 6331 3886 6340 3906
rect 6360 3892 6395 3906
rect 6415 3892 6418 3912
rect 6360 3887 6418 3892
rect 6360 3886 6395 3887
rect 5597 3849 5634 3878
rect 5598 3847 5634 3849
rect 5810 3847 5847 3878
rect 5598 3825 5847 3847
rect 6018 3846 6055 3878
rect 6331 3874 6395 3886
rect 6435 3848 6462 4026
rect 6294 3846 6462 3848
rect 6018 3820 6462 3846
rect 6614 3945 6864 3969
rect 6614 3874 6651 3945
rect 6766 3884 6797 3885
rect 6614 3854 6623 3874
rect 6643 3854 6651 3874
rect 6614 3844 6651 3854
rect 6710 3874 6797 3884
rect 6710 3854 6719 3874
rect 6739 3854 6797 3874
rect 6710 3845 6797 3854
rect 6710 3844 6747 3845
rect 6018 3810 6040 3820
rect 6294 3819 6462 3820
rect 5978 3808 6040 3810
rect 5408 3801 6040 3808
rect 4825 3757 4866 3758
rect 4149 3704 4186 3705
rect 4245 3704 4282 3705
rect 4301 3704 4337 3756
rect 4356 3704 4393 3705
rect 4049 3695 4187 3704
rect 4049 3675 4158 3695
rect 4178 3675 4187 3695
rect 2986 3671 3156 3672
rect 2986 3656 3432 3671
rect 4049 3668 4187 3675
rect 4245 3695 4393 3704
rect 4245 3675 4254 3695
rect 4274 3675 4364 3695
rect 4384 3675 4393 3695
rect 4049 3666 4145 3668
rect 2893 3645 2925 3650
rect 2895 2644 2925 3645
rect 2988 3645 3432 3656
rect 2988 3643 3156 3645
rect 2988 3465 3015 3643
rect 3055 3605 3119 3617
rect 3395 3613 3432 3645
rect 3603 3644 3852 3666
rect 4245 3665 4393 3675
rect 4452 3695 4489 3705
rect 4564 3704 4601 3705
rect 4545 3702 4601 3704
rect 4452 3675 4460 3695
rect 4480 3675 4489 3695
rect 4301 3664 4337 3665
rect 3603 3613 3640 3644
rect 3816 3642 3852 3644
rect 3816 3613 3853 3642
rect 3055 3604 3090 3605
rect 3032 3599 3090 3604
rect 3032 3579 3035 3599
rect 3055 3585 3090 3599
rect 3110 3585 3119 3605
rect 3055 3577 3119 3585
rect 3081 3576 3119 3577
rect 3082 3575 3119 3576
rect 3185 3609 3221 3610
rect 3293 3609 3329 3610
rect 3185 3601 3329 3609
rect 3185 3581 3193 3601
rect 3213 3582 3245 3601
rect 3268 3582 3301 3601
rect 3213 3581 3301 3582
rect 3321 3581 3329 3601
rect 3185 3575 3329 3581
rect 3395 3605 3433 3613
rect 3501 3609 3537 3610
rect 3395 3585 3404 3605
rect 3424 3585 3433 3605
rect 3395 3576 3433 3585
rect 3452 3602 3537 3609
rect 3452 3582 3459 3602
rect 3480 3601 3537 3602
rect 3480 3582 3509 3601
rect 3452 3581 3509 3582
rect 3529 3581 3537 3601
rect 3395 3575 3432 3576
rect 3452 3575 3537 3581
rect 3603 3605 3641 3613
rect 3714 3609 3750 3610
rect 3603 3585 3612 3605
rect 3632 3585 3641 3605
rect 3603 3576 3641 3585
rect 3665 3601 3750 3609
rect 3665 3581 3722 3601
rect 3742 3581 3750 3601
rect 3603 3575 3640 3576
rect 3665 3575 3750 3581
rect 3816 3605 3854 3613
rect 4149 3605 4186 3606
rect 4452 3605 4489 3675
rect 4514 3695 4601 3702
rect 4514 3692 4572 3695
rect 4514 3672 4519 3692
rect 4540 3675 4572 3692
rect 4592 3675 4601 3695
rect 4540 3672 4601 3675
rect 4514 3665 4601 3672
rect 4660 3695 4697 3705
rect 4660 3675 4668 3695
rect 4688 3675 4697 3695
rect 4514 3664 4545 3665
rect 3816 3585 3825 3605
rect 3845 3585 3854 3605
rect 4148 3604 4489 3605
rect 3816 3576 3854 3585
rect 4073 3599 4489 3604
rect 4073 3579 4076 3599
rect 4096 3579 4489 3599
rect 4660 3604 4697 3675
rect 4727 3704 4758 3757
rect 5065 3755 5075 3773
rect 5093 3755 5104 3773
rect 5407 3792 6040 3801
rect 6766 3792 6797 3845
rect 6827 3874 6864 3945
rect 7035 3950 7428 3970
rect 7448 3950 7451 3970
rect 7035 3945 7451 3950
rect 7035 3944 7376 3945
rect 6979 3884 7010 3885
rect 6827 3854 6836 3874
rect 6856 3854 6864 3874
rect 6827 3844 6864 3854
rect 6923 3877 7010 3884
rect 6923 3874 6984 3877
rect 6923 3854 6932 3874
rect 6952 3857 6984 3874
rect 7005 3857 7010 3877
rect 6952 3854 7010 3857
rect 6923 3847 7010 3854
rect 7035 3874 7072 3944
rect 7338 3943 7375 3944
rect 7187 3884 7223 3885
rect 7035 3854 7044 3874
rect 7064 3854 7072 3874
rect 6923 3845 6979 3847
rect 6923 3844 6960 3845
rect 7035 3844 7072 3854
rect 7131 3874 7279 3884
rect 7379 3881 7475 3883
rect 7131 3854 7140 3874
rect 7160 3854 7250 3874
rect 7270 3854 7279 3874
rect 7131 3845 7279 3854
rect 7337 3874 7475 3881
rect 7337 3854 7346 3874
rect 7366 3854 7475 3874
rect 7337 3845 7475 3854
rect 7131 3844 7168 3845
rect 7187 3793 7223 3845
rect 7242 3844 7279 3845
rect 7338 3844 7375 3845
rect 5407 3774 5417 3792
rect 5435 3791 6040 3792
rect 6658 3791 6699 3792
rect 5435 3786 5456 3791
rect 5435 3774 5447 3786
rect 6550 3784 6699 3791
rect 5407 3766 5447 3774
rect 5490 3773 5516 3774
rect 5407 3764 5444 3766
rect 5490 3755 6044 3773
rect 6550 3764 6668 3784
rect 6688 3764 6699 3784
rect 6550 3756 6699 3764
rect 6766 3788 7125 3792
rect 6766 3783 7088 3788
rect 6766 3759 6879 3783
rect 6903 3764 7088 3783
rect 7112 3764 7125 3788
rect 6903 3759 7125 3764
rect 6766 3756 7125 3759
rect 7187 3756 7222 3793
rect 7290 3790 7390 3793
rect 7290 3786 7357 3790
rect 7290 3760 7302 3786
rect 7328 3764 7357 3786
rect 7383 3764 7390 3790
rect 7328 3760 7390 3764
rect 7290 3756 7390 3760
rect 5065 3746 5102 3755
rect 4777 3704 4814 3705
rect 4727 3695 4814 3704
rect 4727 3675 4785 3695
rect 4805 3675 4814 3695
rect 4727 3665 4814 3675
rect 4873 3695 4910 3705
rect 4873 3675 4881 3695
rect 4901 3675 4910 3695
rect 5410 3696 5447 3702
rect 5490 3696 5516 3755
rect 6023 3736 6044 3755
rect 5410 3693 5516 3696
rect 5068 3680 5105 3684
rect 4727 3664 4758 3665
rect 4873 3604 4910 3675
rect 4660 3580 4910 3604
rect 5066 3674 5105 3680
rect 5066 3656 5077 3674
rect 5095 3656 5105 3674
rect 5410 3675 5419 3693
rect 5437 3679 5516 3693
rect 5601 3711 5851 3735
rect 5437 3677 5513 3679
rect 5437 3675 5447 3677
rect 5410 3665 5447 3675
rect 5066 3647 5105 3656
rect 3816 3575 3853 3576
rect 3239 3554 3275 3575
rect 3665 3554 3696 3575
rect 4452 3556 4489 3579
rect 5066 3569 5101 3647
rect 5415 3600 5446 3665
rect 5601 3640 5638 3711
rect 5753 3650 5784 3651
rect 5601 3620 5610 3640
rect 5630 3620 5638 3640
rect 5601 3610 5638 3620
rect 5697 3640 5784 3650
rect 5697 3620 5706 3640
rect 5726 3620 5784 3640
rect 5697 3611 5784 3620
rect 5697 3610 5734 3611
rect 5063 3559 5101 3569
rect 5414 3591 5451 3600
rect 5414 3573 5424 3591
rect 5442 3573 5451 3591
rect 5414 3563 5451 3573
rect 4452 3555 4622 3556
rect 5063 3555 5073 3559
rect 3072 3550 3172 3554
rect 3072 3546 3134 3550
rect 3072 3520 3079 3546
rect 3105 3524 3134 3546
rect 3160 3524 3172 3550
rect 3105 3520 3172 3524
rect 3072 3517 3172 3520
rect 3240 3517 3275 3554
rect 3337 3551 3696 3554
rect 3337 3546 3559 3551
rect 3337 3522 3350 3546
rect 3374 3527 3559 3546
rect 3583 3527 3696 3551
rect 3374 3522 3696 3527
rect 3337 3518 3696 3522
rect 3763 3546 3912 3554
rect 3763 3526 3774 3546
rect 3794 3526 3912 3546
rect 4452 3541 5073 3555
rect 5091 3541 5101 3559
rect 5753 3558 5784 3611
rect 5814 3640 5851 3711
rect 6022 3716 6415 3736
rect 6435 3716 6438 3736
rect 6766 3735 6797 3756
rect 7187 3735 7223 3756
rect 6609 3734 6646 3735
rect 6022 3711 6438 3716
rect 6608 3725 6646 3734
rect 6022 3710 6363 3711
rect 5966 3650 5997 3651
rect 5814 3620 5823 3640
rect 5843 3620 5851 3640
rect 5814 3610 5851 3620
rect 5910 3643 5997 3650
rect 5910 3640 5971 3643
rect 5910 3620 5919 3640
rect 5939 3623 5971 3640
rect 5992 3623 5997 3643
rect 5939 3620 5997 3623
rect 5910 3613 5997 3620
rect 6022 3640 6059 3710
rect 6325 3709 6362 3710
rect 6608 3705 6617 3725
rect 6637 3705 6646 3725
rect 6608 3697 6646 3705
rect 6712 3729 6797 3735
rect 6822 3734 6859 3735
rect 6712 3709 6720 3729
rect 6740 3709 6797 3729
rect 6712 3701 6797 3709
rect 6821 3725 6859 3734
rect 6821 3705 6830 3725
rect 6850 3705 6859 3725
rect 6712 3700 6748 3701
rect 6821 3697 6859 3705
rect 6925 3729 7010 3735
rect 7030 3734 7067 3735
rect 6925 3709 6933 3729
rect 6953 3728 7010 3729
rect 6953 3709 6982 3728
rect 6925 3708 6982 3709
rect 7003 3708 7010 3728
rect 6925 3701 7010 3708
rect 7029 3725 7067 3734
rect 7029 3705 7038 3725
rect 7058 3705 7067 3725
rect 6925 3700 6961 3701
rect 7029 3697 7067 3705
rect 7133 3729 7277 3735
rect 7133 3709 7141 3729
rect 7161 3709 7193 3729
rect 7217 3709 7249 3729
rect 7269 3709 7277 3729
rect 7133 3701 7277 3709
rect 7133 3700 7169 3701
rect 7241 3700 7277 3701
rect 7343 3734 7380 3735
rect 7343 3733 7381 3734
rect 7343 3725 7407 3733
rect 7343 3705 7352 3725
rect 7372 3711 7407 3725
rect 7427 3711 7430 3731
rect 7372 3706 7430 3711
rect 7372 3705 7407 3706
rect 6609 3668 6646 3697
rect 6610 3666 6646 3668
rect 6822 3666 6859 3697
rect 6174 3650 6210 3651
rect 6022 3620 6031 3640
rect 6051 3620 6059 3640
rect 5910 3611 5966 3613
rect 5910 3610 5947 3611
rect 6022 3610 6059 3620
rect 6118 3640 6266 3650
rect 6366 3647 6462 3649
rect 6118 3620 6127 3640
rect 6147 3620 6237 3640
rect 6257 3620 6266 3640
rect 6118 3611 6266 3620
rect 6324 3640 6462 3647
rect 6610 3644 6859 3666
rect 7030 3665 7067 3697
rect 7343 3693 7407 3705
rect 7447 3667 7474 3845
rect 7306 3665 7474 3667
rect 7030 3661 7474 3665
rect 6324 3620 6333 3640
rect 6353 3620 6462 3640
rect 7030 3642 7079 3661
rect 7099 3642 7474 3661
rect 7030 3639 7474 3642
rect 7306 3638 7474 3639
rect 6324 3611 6462 3620
rect 6118 3610 6155 3611
rect 6174 3559 6210 3611
rect 6229 3610 6266 3611
rect 6325 3610 6362 3611
rect 5645 3557 5686 3558
rect 4452 3535 5101 3541
rect 5537 3550 5686 3557
rect 4452 3534 5100 3535
rect 5063 3532 5100 3534
rect 3763 3519 3912 3526
rect 5537 3530 5655 3550
rect 5675 3530 5686 3550
rect 5537 3522 5686 3530
rect 5753 3554 6112 3558
rect 5753 3549 6075 3554
rect 5753 3525 5866 3549
rect 5890 3530 6075 3549
rect 6099 3530 6112 3554
rect 5890 3525 6112 3530
rect 5753 3522 6112 3525
rect 6174 3522 6209 3559
rect 6277 3556 6377 3559
rect 6277 3552 6344 3556
rect 6277 3526 6289 3552
rect 6315 3530 6344 3552
rect 6370 3530 6377 3556
rect 6315 3526 6377 3530
rect 6277 3522 6377 3526
rect 3763 3518 3804 3519
rect 3087 3465 3124 3466
rect 3183 3465 3220 3466
rect 3239 3465 3275 3517
rect 3294 3465 3331 3466
rect 2987 3456 3125 3465
rect 2987 3436 3096 3456
rect 3116 3436 3125 3456
rect 2987 3429 3125 3436
rect 3183 3456 3331 3465
rect 3183 3436 3192 3456
rect 3212 3436 3302 3456
rect 3322 3436 3331 3456
rect 2987 3427 3083 3429
rect 3183 3426 3331 3436
rect 3390 3456 3427 3466
rect 3502 3465 3539 3466
rect 3483 3463 3539 3465
rect 3390 3436 3398 3456
rect 3418 3436 3427 3456
rect 3239 3425 3275 3426
rect 3087 3366 3124 3367
rect 3390 3366 3427 3436
rect 3452 3456 3539 3463
rect 3452 3453 3510 3456
rect 3452 3433 3457 3453
rect 3478 3436 3510 3453
rect 3530 3436 3539 3456
rect 3478 3433 3539 3436
rect 3452 3426 3539 3433
rect 3598 3456 3635 3466
rect 3598 3436 3606 3456
rect 3626 3436 3635 3456
rect 3452 3425 3483 3426
rect 3086 3365 3427 3366
rect 3011 3360 3427 3365
rect 3011 3340 3014 3360
rect 3034 3340 3427 3360
rect 3598 3365 3635 3436
rect 3665 3465 3696 3518
rect 5753 3501 5784 3522
rect 6174 3501 6210 3522
rect 5417 3492 5454 3501
rect 5596 3500 5633 3501
rect 5417 3474 5426 3492
rect 5444 3474 5454 3492
rect 3715 3465 3752 3466
rect 3665 3456 3752 3465
rect 3665 3436 3723 3456
rect 3743 3436 3752 3456
rect 3665 3426 3752 3436
rect 3811 3456 3848 3466
rect 3811 3436 3819 3456
rect 3839 3436 3848 3456
rect 3665 3425 3696 3426
rect 3811 3365 3848 3436
rect 5066 3460 5103 3470
rect 5417 3464 5454 3474
rect 5066 3442 5075 3460
rect 5093 3442 5103 3460
rect 5066 3433 5103 3442
rect 5066 3409 5101 3433
rect 5418 3429 5454 3464
rect 5595 3491 5633 3500
rect 5595 3471 5604 3491
rect 5624 3471 5633 3491
rect 5595 3463 5633 3471
rect 5699 3495 5784 3501
rect 5809 3500 5846 3501
rect 5699 3475 5707 3495
rect 5727 3475 5784 3495
rect 5699 3467 5784 3475
rect 5808 3491 5846 3500
rect 5808 3471 5817 3491
rect 5837 3471 5846 3491
rect 5699 3466 5735 3467
rect 5808 3463 5846 3471
rect 5912 3495 5997 3501
rect 6017 3500 6054 3501
rect 5912 3475 5920 3495
rect 5940 3494 5997 3495
rect 5940 3475 5969 3494
rect 5912 3474 5969 3475
rect 5990 3474 5997 3494
rect 5912 3467 5997 3474
rect 6016 3491 6054 3500
rect 6016 3471 6025 3491
rect 6045 3471 6054 3491
rect 5912 3466 5948 3467
rect 6016 3463 6054 3471
rect 6120 3495 6264 3501
rect 6120 3475 6128 3495
rect 6148 3494 6236 3495
rect 6148 3475 6176 3494
rect 6120 3473 6176 3475
rect 6198 3475 6236 3494
rect 6256 3475 6264 3495
rect 6198 3473 6264 3475
rect 6120 3467 6264 3473
rect 6120 3466 6156 3467
rect 6228 3466 6264 3467
rect 6330 3500 6367 3501
rect 6330 3499 6368 3500
rect 6330 3491 6394 3499
rect 6330 3471 6339 3491
rect 6359 3477 6394 3491
rect 6414 3477 6417 3497
rect 6359 3472 6417 3477
rect 6359 3471 6394 3472
rect 5596 3434 5633 3463
rect 5064 3385 5101 3409
rect 5063 3379 5101 3385
rect 3598 3341 3848 3365
rect 4474 3361 5101 3379
rect 4056 3344 4224 3345
rect 4475 3344 4499 3361
rect 4056 3318 4500 3344
rect 4056 3316 4224 3318
rect 4056 3138 4083 3316
rect 4123 3278 4187 3290
rect 4463 3286 4500 3318
rect 4671 3317 4920 3339
rect 4671 3286 4708 3317
rect 4884 3315 4920 3317
rect 5063 3320 5101 3361
rect 5416 3388 5454 3429
rect 5597 3432 5633 3434
rect 5809 3432 5846 3463
rect 5597 3410 5846 3432
rect 6017 3431 6054 3463
rect 6330 3459 6394 3471
rect 6434 3433 6461 3611
rect 6293 3431 6461 3433
rect 6017 3405 6461 3431
rect 6018 3388 6042 3405
rect 6293 3404 6461 3405
rect 5416 3370 6043 3388
rect 6669 3384 6919 3408
rect 5416 3364 5454 3370
rect 5416 3340 5453 3364
rect 4884 3286 4921 3315
rect 4123 3277 4158 3278
rect 4100 3272 4158 3277
rect 4100 3252 4103 3272
rect 4123 3258 4158 3272
rect 4178 3258 4187 3278
rect 4123 3250 4187 3258
rect 4149 3249 4187 3250
rect 4150 3248 4187 3249
rect 4253 3282 4289 3283
rect 4361 3282 4397 3283
rect 4253 3276 4397 3282
rect 4253 3274 4319 3276
rect 4253 3254 4261 3274
rect 4281 3255 4319 3274
rect 4341 3274 4397 3276
rect 4341 3255 4369 3274
rect 4281 3254 4369 3255
rect 4389 3254 4397 3274
rect 4253 3248 4397 3254
rect 4463 3278 4501 3286
rect 4569 3282 4605 3283
rect 4463 3258 4472 3278
rect 4492 3258 4501 3278
rect 4463 3249 4501 3258
rect 4520 3275 4605 3282
rect 4520 3255 4527 3275
rect 4548 3274 4605 3275
rect 4548 3255 4577 3274
rect 4520 3254 4577 3255
rect 4597 3254 4605 3274
rect 4463 3248 4500 3249
rect 4520 3248 4605 3254
rect 4671 3278 4709 3286
rect 4782 3282 4818 3283
rect 4671 3258 4680 3278
rect 4700 3258 4709 3278
rect 4671 3249 4709 3258
rect 4733 3274 4818 3282
rect 4733 3254 4790 3274
rect 4810 3254 4818 3274
rect 4671 3248 4708 3249
rect 4733 3248 4818 3254
rect 4884 3278 4922 3286
rect 4884 3258 4893 3278
rect 4913 3258 4922 3278
rect 4884 3249 4922 3258
rect 5063 3285 5099 3320
rect 5416 3316 5451 3340
rect 5414 3307 5451 3316
rect 5414 3289 5424 3307
rect 5442 3289 5451 3307
rect 5063 3275 5100 3285
rect 5414 3279 5451 3289
rect 6669 3313 6706 3384
rect 6821 3323 6852 3324
rect 6669 3293 6678 3313
rect 6698 3293 6706 3313
rect 6669 3283 6706 3293
rect 6765 3313 6852 3323
rect 6765 3293 6774 3313
rect 6794 3293 6852 3313
rect 6765 3284 6852 3293
rect 6765 3283 6802 3284
rect 5063 3257 5073 3275
rect 5091 3257 5100 3275
rect 4884 3248 4921 3249
rect 5063 3248 5100 3257
rect 4307 3227 4343 3248
rect 4733 3227 4764 3248
rect 6821 3231 6852 3284
rect 6882 3313 6919 3384
rect 7090 3389 7483 3409
rect 7503 3389 7506 3409
rect 7090 3384 7506 3389
rect 7090 3383 7431 3384
rect 7034 3323 7065 3324
rect 6882 3293 6891 3313
rect 6911 3293 6919 3313
rect 6882 3283 6919 3293
rect 6978 3316 7065 3323
rect 6978 3313 7039 3316
rect 6978 3293 6987 3313
rect 7007 3296 7039 3313
rect 7060 3296 7065 3316
rect 7007 3293 7065 3296
rect 6978 3286 7065 3293
rect 7090 3313 7127 3383
rect 7393 3382 7430 3383
rect 7242 3323 7278 3324
rect 7090 3293 7099 3313
rect 7119 3293 7127 3313
rect 6978 3284 7034 3286
rect 6978 3283 7015 3284
rect 7090 3283 7127 3293
rect 7186 3313 7334 3323
rect 7434 3320 7530 3322
rect 7186 3293 7195 3313
rect 7215 3293 7305 3313
rect 7325 3293 7334 3313
rect 7186 3284 7334 3293
rect 7392 3313 7530 3320
rect 7392 3293 7401 3313
rect 7421 3293 7530 3313
rect 7392 3284 7530 3293
rect 7186 3283 7223 3284
rect 7242 3232 7278 3284
rect 7297 3283 7334 3284
rect 7393 3283 7430 3284
rect 6713 3230 6754 3231
rect 4140 3223 4240 3227
rect 4140 3219 4202 3223
rect 4140 3193 4147 3219
rect 4173 3197 4202 3219
rect 4228 3197 4240 3223
rect 4173 3193 4240 3197
rect 4140 3190 4240 3193
rect 4308 3190 4343 3227
rect 4405 3224 4764 3227
rect 4405 3219 4627 3224
rect 4405 3195 4418 3219
rect 4442 3200 4627 3219
rect 4651 3200 4764 3224
rect 4442 3195 4764 3200
rect 4405 3191 4764 3195
rect 4831 3219 4980 3227
rect 4831 3199 4842 3219
rect 4862 3199 4980 3219
rect 6605 3223 6754 3230
rect 5417 3215 5454 3217
rect 5417 3214 6065 3215
rect 4831 3192 4980 3199
rect 5416 3208 6065 3214
rect 4831 3191 4872 3192
rect 4155 3138 4192 3139
rect 4251 3138 4288 3139
rect 4307 3138 4343 3190
rect 4362 3138 4399 3139
rect 4055 3129 4193 3138
rect 3043 3110 3211 3111
rect 3043 3107 3487 3110
rect 3043 3088 3418 3107
rect 3438 3088 3487 3107
rect 4055 3109 4164 3129
rect 4184 3109 4193 3129
rect 3043 3084 3487 3088
rect 3043 3082 3211 3084
rect 3043 2904 3070 3082
rect 3110 3044 3174 3056
rect 3450 3052 3487 3084
rect 3658 3083 3907 3105
rect 4055 3102 4193 3109
rect 4251 3129 4399 3138
rect 4251 3109 4260 3129
rect 4280 3109 4370 3129
rect 4390 3109 4399 3129
rect 4055 3100 4151 3102
rect 4251 3099 4399 3109
rect 4458 3129 4495 3139
rect 4570 3138 4607 3139
rect 4551 3136 4607 3138
rect 4458 3109 4466 3129
rect 4486 3109 4495 3129
rect 4307 3098 4343 3099
rect 3658 3052 3695 3083
rect 3871 3081 3907 3083
rect 3871 3052 3908 3081
rect 3110 3043 3145 3044
rect 3087 3038 3145 3043
rect 3087 3018 3090 3038
rect 3110 3024 3145 3038
rect 3165 3024 3174 3044
rect 3110 3016 3174 3024
rect 3136 3015 3174 3016
rect 3137 3014 3174 3015
rect 3240 3048 3276 3049
rect 3348 3048 3384 3049
rect 3240 3040 3384 3048
rect 3240 3020 3248 3040
rect 3268 3020 3300 3040
rect 3324 3020 3356 3040
rect 3376 3020 3384 3040
rect 3240 3014 3384 3020
rect 3450 3044 3488 3052
rect 3556 3048 3592 3049
rect 3450 3024 3459 3044
rect 3479 3024 3488 3044
rect 3450 3015 3488 3024
rect 3507 3041 3592 3048
rect 3507 3021 3514 3041
rect 3535 3040 3592 3041
rect 3535 3021 3564 3040
rect 3507 3020 3564 3021
rect 3584 3020 3592 3040
rect 3450 3014 3487 3015
rect 3507 3014 3592 3020
rect 3658 3044 3696 3052
rect 3769 3048 3805 3049
rect 3658 3024 3667 3044
rect 3687 3024 3696 3044
rect 3658 3015 3696 3024
rect 3720 3040 3805 3048
rect 3720 3020 3777 3040
rect 3797 3020 3805 3040
rect 3658 3014 3695 3015
rect 3720 3014 3805 3020
rect 3871 3044 3909 3052
rect 3871 3024 3880 3044
rect 3900 3024 3909 3044
rect 4155 3039 4192 3040
rect 4458 3039 4495 3109
rect 4520 3129 4607 3136
rect 4520 3126 4578 3129
rect 4520 3106 4525 3126
rect 4546 3109 4578 3126
rect 4598 3109 4607 3129
rect 4546 3106 4607 3109
rect 4520 3099 4607 3106
rect 4666 3129 4703 3139
rect 4666 3109 4674 3129
rect 4694 3109 4703 3129
rect 4520 3098 4551 3099
rect 4154 3038 4495 3039
rect 3871 3015 3909 3024
rect 4079 3033 4495 3038
rect 3871 3014 3908 3015
rect 3294 2993 3330 3014
rect 3720 2993 3751 3014
rect 4079 3013 4082 3033
rect 4102 3013 4495 3033
rect 4666 3038 4703 3109
rect 4733 3138 4764 3191
rect 5416 3190 5426 3208
rect 5444 3194 6065 3208
rect 6605 3203 6723 3223
rect 6743 3203 6754 3223
rect 6605 3195 6754 3203
rect 6821 3227 7180 3231
rect 6821 3222 7143 3227
rect 6821 3198 6934 3222
rect 6958 3203 7143 3222
rect 7167 3203 7180 3227
rect 6958 3198 7180 3203
rect 6821 3195 7180 3198
rect 7242 3195 7277 3232
rect 7345 3229 7445 3232
rect 7345 3225 7412 3229
rect 7345 3199 7357 3225
rect 7383 3203 7412 3225
rect 7438 3203 7445 3229
rect 7383 3199 7445 3203
rect 7345 3195 7445 3199
rect 5444 3190 5454 3194
rect 5895 3193 6065 3194
rect 5066 3176 5103 3186
rect 5066 3158 5075 3176
rect 5093 3158 5103 3176
rect 5066 3149 5103 3158
rect 5416 3180 5454 3190
rect 4783 3138 4820 3139
rect 4733 3129 4820 3138
rect 4733 3109 4791 3129
rect 4811 3109 4820 3129
rect 4733 3099 4820 3109
rect 4879 3129 4916 3139
rect 4879 3109 4887 3129
rect 4907 3109 4916 3129
rect 4733 3098 4764 3099
rect 4879 3038 4916 3109
rect 5071 3084 5102 3149
rect 5416 3102 5451 3180
rect 6028 3170 6065 3193
rect 6821 3174 6852 3195
rect 7242 3174 7278 3195
rect 6664 3173 6701 3174
rect 5412 3093 5451 3102
rect 5070 3074 5107 3084
rect 5070 3072 5080 3074
rect 5004 3070 5080 3072
rect 4666 3014 4916 3038
rect 5001 3056 5080 3070
rect 5098 3056 5107 3074
rect 5412 3075 5422 3093
rect 5440 3075 5451 3093
rect 5412 3069 5451 3075
rect 5607 3145 5857 3169
rect 5607 3074 5644 3145
rect 5759 3084 5790 3085
rect 5412 3065 5449 3069
rect 5001 3053 5107 3056
rect 4473 2994 4494 3013
rect 5001 2994 5027 3053
rect 5070 3047 5107 3053
rect 5607 3054 5616 3074
rect 5636 3054 5644 3074
rect 5607 3044 5644 3054
rect 5703 3074 5790 3084
rect 5703 3054 5712 3074
rect 5732 3054 5790 3074
rect 5703 3045 5790 3054
rect 5703 3044 5740 3045
rect 5415 2994 5452 3003
rect 3127 2989 3227 2993
rect 3127 2985 3189 2989
rect 3127 2959 3134 2985
rect 3160 2963 3189 2985
rect 3215 2963 3227 2989
rect 3160 2959 3227 2963
rect 3127 2956 3227 2959
rect 3295 2956 3330 2993
rect 3392 2990 3751 2993
rect 3392 2985 3614 2990
rect 3392 2961 3405 2985
rect 3429 2966 3614 2985
rect 3638 2966 3751 2990
rect 3429 2961 3751 2966
rect 3392 2957 3751 2961
rect 3818 2985 3967 2993
rect 3818 2965 3829 2985
rect 3849 2965 3967 2985
rect 4473 2976 5027 2994
rect 5073 2983 5110 2985
rect 5001 2975 5027 2976
rect 5070 2975 5110 2983
rect 3818 2958 3967 2965
rect 5070 2963 5082 2975
rect 5061 2958 5082 2963
rect 3818 2957 3859 2958
rect 4477 2957 5082 2958
rect 5100 2957 5110 2975
rect 3142 2904 3179 2905
rect 3238 2904 3275 2905
rect 3294 2904 3330 2956
rect 3349 2904 3386 2905
rect 3042 2895 3180 2904
rect 3042 2875 3151 2895
rect 3171 2875 3180 2895
rect 3042 2868 3180 2875
rect 3238 2895 3386 2904
rect 3238 2875 3247 2895
rect 3267 2875 3357 2895
rect 3377 2875 3386 2895
rect 3042 2866 3138 2868
rect 3238 2865 3386 2875
rect 3445 2895 3482 2905
rect 3557 2904 3594 2905
rect 3538 2902 3594 2904
rect 3445 2875 3453 2895
rect 3473 2875 3482 2895
rect 3294 2864 3330 2865
rect 3142 2805 3179 2806
rect 3445 2805 3482 2875
rect 3507 2895 3594 2902
rect 3507 2892 3565 2895
rect 3507 2872 3512 2892
rect 3533 2875 3565 2892
rect 3585 2875 3594 2895
rect 3533 2872 3594 2875
rect 3507 2865 3594 2872
rect 3653 2895 3690 2905
rect 3653 2875 3661 2895
rect 3681 2875 3690 2895
rect 3507 2864 3538 2865
rect 3141 2804 3482 2805
rect 3066 2799 3482 2804
rect 3066 2779 3069 2799
rect 3089 2779 3482 2799
rect 3653 2804 3690 2875
rect 3720 2904 3751 2957
rect 4477 2948 5110 2957
rect 5413 2976 5424 2994
rect 5442 2976 5452 2994
rect 5759 2992 5790 3045
rect 5820 3074 5857 3145
rect 6028 3150 6421 3170
rect 6441 3150 6444 3170
rect 6028 3145 6444 3150
rect 6663 3164 6701 3173
rect 6028 3144 6369 3145
rect 6663 3144 6672 3164
rect 6692 3144 6701 3164
rect 5972 3084 6003 3085
rect 5820 3054 5829 3074
rect 5849 3054 5857 3074
rect 5820 3044 5857 3054
rect 5916 3077 6003 3084
rect 5916 3074 5977 3077
rect 5916 3054 5925 3074
rect 5945 3057 5977 3074
rect 5998 3057 6003 3077
rect 5945 3054 6003 3057
rect 5916 3047 6003 3054
rect 6028 3074 6065 3144
rect 6331 3143 6368 3144
rect 6663 3136 6701 3144
rect 6767 3168 6852 3174
rect 6877 3173 6914 3174
rect 6767 3148 6775 3168
rect 6795 3148 6852 3168
rect 6767 3140 6852 3148
rect 6876 3164 6914 3173
rect 6876 3144 6885 3164
rect 6905 3144 6914 3164
rect 6767 3139 6803 3140
rect 6876 3136 6914 3144
rect 6980 3168 7065 3174
rect 7085 3173 7122 3174
rect 6980 3148 6988 3168
rect 7008 3167 7065 3168
rect 7008 3148 7037 3167
rect 6980 3147 7037 3148
rect 7058 3147 7065 3167
rect 6980 3140 7065 3147
rect 7084 3164 7122 3173
rect 7084 3144 7093 3164
rect 7113 3144 7122 3164
rect 6980 3139 7016 3140
rect 7084 3136 7122 3144
rect 7188 3168 7332 3174
rect 7188 3148 7196 3168
rect 7216 3166 7304 3168
rect 7216 3149 7252 3166
rect 7276 3149 7304 3166
rect 7216 3148 7304 3149
rect 7324 3148 7332 3168
rect 7188 3140 7332 3148
rect 7188 3139 7224 3140
rect 7296 3139 7332 3140
rect 7398 3173 7435 3174
rect 7398 3172 7436 3173
rect 7398 3164 7462 3172
rect 7398 3144 7407 3164
rect 7427 3150 7462 3164
rect 7482 3150 7485 3170
rect 7427 3145 7485 3150
rect 7427 3144 7462 3145
rect 6664 3107 6701 3136
rect 6665 3105 6701 3107
rect 6877 3105 6914 3136
rect 6180 3084 6216 3085
rect 6028 3054 6037 3074
rect 6057 3054 6065 3074
rect 5916 3045 5972 3047
rect 5916 3044 5953 3045
rect 6028 3044 6065 3054
rect 6124 3074 6272 3084
rect 6665 3083 6914 3105
rect 7085 3104 7122 3136
rect 7398 3132 7462 3144
rect 7502 3106 7529 3284
rect 7361 3104 7529 3106
rect 7085 3093 7529 3104
rect 6372 3081 6468 3083
rect 6124 3054 6133 3074
rect 6153 3054 6243 3074
rect 6263 3054 6272 3074
rect 6124 3045 6272 3054
rect 6330 3074 6468 3081
rect 7085 3078 7531 3093
rect 7361 3077 7531 3078
rect 6330 3054 6339 3074
rect 6359 3054 6468 3074
rect 6330 3045 6468 3054
rect 6124 3044 6161 3045
rect 6180 2993 6216 3045
rect 6235 3044 6272 3045
rect 6331 3044 6368 3045
rect 5651 2991 5692 2992
rect 4477 2941 5109 2948
rect 4477 2939 4539 2941
rect 4055 2929 4223 2930
rect 4477 2929 4499 2939
rect 3770 2904 3807 2905
rect 3720 2895 3807 2904
rect 3720 2875 3778 2895
rect 3798 2875 3807 2895
rect 3720 2865 3807 2875
rect 3866 2895 3903 2905
rect 3866 2875 3874 2895
rect 3894 2875 3903 2895
rect 3720 2864 3751 2865
rect 3866 2804 3903 2875
rect 3653 2780 3903 2804
rect 4055 2903 4499 2929
rect 4055 2901 4223 2903
rect 4055 2723 4082 2901
rect 4122 2863 4186 2875
rect 4462 2871 4499 2903
rect 4670 2902 4919 2924
rect 4670 2871 4707 2902
rect 4883 2900 4919 2902
rect 4883 2871 4920 2900
rect 4122 2862 4157 2863
rect 4099 2857 4157 2862
rect 4099 2837 4102 2857
rect 4122 2843 4157 2857
rect 4177 2843 4186 2863
rect 4122 2835 4186 2843
rect 4148 2834 4186 2835
rect 4149 2833 4186 2834
rect 4252 2867 4288 2868
rect 4360 2867 4396 2868
rect 4252 2859 4396 2867
rect 4252 2839 4260 2859
rect 4280 2839 4309 2859
rect 4252 2838 4309 2839
rect 4331 2839 4368 2859
rect 4388 2839 4396 2859
rect 4331 2838 4396 2839
rect 4252 2833 4396 2838
rect 4462 2863 4500 2871
rect 4568 2867 4604 2868
rect 4462 2843 4471 2863
rect 4491 2843 4500 2863
rect 4462 2834 4500 2843
rect 4519 2860 4604 2867
rect 4519 2840 4526 2860
rect 4547 2859 4604 2860
rect 4547 2840 4576 2859
rect 4519 2839 4576 2840
rect 4596 2839 4604 2859
rect 4462 2833 4499 2834
rect 4519 2833 4604 2839
rect 4670 2863 4708 2871
rect 4781 2867 4817 2868
rect 4670 2843 4679 2863
rect 4699 2843 4708 2863
rect 4670 2834 4708 2843
rect 4732 2859 4817 2867
rect 4732 2839 4789 2859
rect 4809 2839 4817 2859
rect 4670 2833 4707 2834
rect 4732 2833 4817 2839
rect 4883 2863 4921 2871
rect 4883 2843 4892 2863
rect 4912 2843 4921 2863
rect 4883 2834 4921 2843
rect 4883 2833 4920 2834
rect 4306 2812 4342 2833
rect 4732 2812 4763 2833
rect 4139 2808 4239 2812
rect 4139 2804 4201 2808
rect 4139 2778 4146 2804
rect 4172 2782 4201 2804
rect 4227 2782 4239 2808
rect 4172 2778 4239 2782
rect 4139 2775 4239 2778
rect 4307 2775 4342 2812
rect 4404 2809 4763 2812
rect 4404 2804 4626 2809
rect 4404 2780 4417 2804
rect 4441 2785 4626 2804
rect 4650 2785 4763 2809
rect 4441 2780 4763 2785
rect 4404 2776 4763 2780
rect 4830 2804 4979 2812
rect 4830 2784 4841 2804
rect 4861 2784 4979 2804
rect 4830 2777 4979 2784
rect 5070 2792 5109 2941
rect 5413 2827 5452 2976
rect 5543 2984 5692 2991
rect 5543 2964 5661 2984
rect 5681 2964 5692 2984
rect 5543 2956 5692 2964
rect 5759 2988 6118 2992
rect 5759 2983 6081 2988
rect 5759 2959 5872 2983
rect 5896 2964 6081 2983
rect 6105 2964 6118 2988
rect 5896 2959 6118 2964
rect 5759 2956 6118 2959
rect 6180 2956 6215 2993
rect 6283 2990 6383 2993
rect 6283 2986 6350 2990
rect 6283 2960 6295 2986
rect 6321 2964 6350 2986
rect 6376 2964 6383 2990
rect 6321 2960 6383 2964
rect 6283 2956 6383 2960
rect 5759 2935 5790 2956
rect 6180 2935 6216 2956
rect 5602 2934 5639 2935
rect 5601 2925 5639 2934
rect 5601 2905 5610 2925
rect 5630 2905 5639 2925
rect 5601 2897 5639 2905
rect 5705 2929 5790 2935
rect 5815 2934 5852 2935
rect 5705 2909 5713 2929
rect 5733 2909 5790 2929
rect 5705 2901 5790 2909
rect 5814 2925 5852 2934
rect 5814 2905 5823 2925
rect 5843 2905 5852 2925
rect 5705 2900 5741 2901
rect 5814 2897 5852 2905
rect 5918 2929 6003 2935
rect 6023 2934 6060 2935
rect 5918 2909 5926 2929
rect 5946 2928 6003 2929
rect 5946 2909 5975 2928
rect 5918 2908 5975 2909
rect 5996 2908 6003 2928
rect 5918 2901 6003 2908
rect 6022 2925 6060 2934
rect 6022 2905 6031 2925
rect 6051 2905 6060 2925
rect 5918 2900 5954 2901
rect 6022 2897 6060 2905
rect 6126 2930 6270 2935
rect 6126 2929 6191 2930
rect 6126 2909 6134 2929
rect 6154 2909 6191 2929
rect 6213 2929 6270 2930
rect 6213 2909 6242 2929
rect 6262 2909 6270 2929
rect 6126 2901 6270 2909
rect 6126 2900 6162 2901
rect 6234 2900 6270 2901
rect 6336 2934 6373 2935
rect 6336 2933 6374 2934
rect 6336 2925 6400 2933
rect 6336 2905 6345 2925
rect 6365 2911 6400 2925
rect 6420 2911 6423 2931
rect 6365 2906 6423 2911
rect 6365 2905 6400 2906
rect 5602 2868 5639 2897
rect 5603 2866 5639 2868
rect 5815 2866 5852 2897
rect 5603 2844 5852 2866
rect 6023 2865 6060 2897
rect 6336 2893 6400 2905
rect 6440 2867 6467 3045
rect 6299 2865 6467 2867
rect 6023 2839 6467 2865
rect 6619 2964 6869 2988
rect 6619 2893 6656 2964
rect 6771 2903 6802 2904
rect 6619 2873 6628 2893
rect 6648 2873 6656 2893
rect 6619 2863 6656 2873
rect 6715 2893 6802 2903
rect 6715 2873 6724 2893
rect 6744 2873 6802 2893
rect 6715 2864 6802 2873
rect 6715 2863 6752 2864
rect 6023 2829 6045 2839
rect 6299 2838 6467 2839
rect 5983 2827 6045 2829
rect 5413 2820 6045 2827
rect 4830 2776 4871 2777
rect 4154 2723 4191 2724
rect 4250 2723 4287 2724
rect 4306 2723 4342 2775
rect 4361 2723 4398 2724
rect 4054 2714 4192 2723
rect 4054 2694 4163 2714
rect 4183 2694 4192 2714
rect 4054 2687 4192 2694
rect 4250 2714 4398 2723
rect 4250 2694 4259 2714
rect 4279 2694 4369 2714
rect 4389 2694 4398 2714
rect 4054 2685 4150 2687
rect 4250 2684 4398 2694
rect 4457 2714 4494 2724
rect 4569 2723 4606 2724
rect 4550 2721 4606 2723
rect 4457 2694 4465 2714
rect 4485 2694 4494 2714
rect 4306 2683 4342 2684
rect 2835 2643 3003 2644
rect 2835 2617 3279 2643
rect 2835 2615 3003 2617
rect 2835 2437 2862 2615
rect 2902 2577 2966 2589
rect 3242 2585 3279 2617
rect 3450 2616 3699 2638
rect 4154 2624 4191 2625
rect 4457 2624 4494 2694
rect 4519 2714 4606 2721
rect 4519 2711 4577 2714
rect 4519 2691 4524 2711
rect 4545 2694 4577 2711
rect 4597 2694 4606 2714
rect 4545 2691 4606 2694
rect 4519 2684 4606 2691
rect 4665 2714 4702 2724
rect 4665 2694 4673 2714
rect 4693 2694 4702 2714
rect 4519 2683 4550 2684
rect 4153 2623 4494 2624
rect 3450 2585 3487 2616
rect 3663 2614 3699 2616
rect 4078 2618 4494 2623
rect 3663 2585 3700 2614
rect 4078 2598 4081 2618
rect 4101 2598 4494 2618
rect 4665 2623 4702 2694
rect 4732 2723 4763 2776
rect 5070 2774 5080 2792
rect 5098 2774 5109 2792
rect 5412 2811 6045 2820
rect 6771 2811 6802 2864
rect 6832 2893 6869 2964
rect 7040 2969 7433 2989
rect 7453 2969 7456 2989
rect 7040 2964 7456 2969
rect 7040 2963 7381 2964
rect 6984 2903 7015 2904
rect 6832 2873 6841 2893
rect 6861 2873 6869 2893
rect 6832 2863 6869 2873
rect 6928 2896 7015 2903
rect 6928 2893 6989 2896
rect 6928 2873 6937 2893
rect 6957 2876 6989 2893
rect 7010 2876 7015 2896
rect 6957 2873 7015 2876
rect 6928 2866 7015 2873
rect 7040 2893 7077 2963
rect 7343 2962 7380 2963
rect 7192 2903 7228 2904
rect 7040 2873 7049 2893
rect 7069 2873 7077 2893
rect 6928 2864 6984 2866
rect 6928 2863 6965 2864
rect 7040 2863 7077 2873
rect 7136 2893 7284 2903
rect 7384 2900 7480 2902
rect 7136 2873 7145 2893
rect 7165 2873 7255 2893
rect 7275 2873 7284 2893
rect 7136 2864 7284 2873
rect 7342 2893 7480 2900
rect 7342 2873 7351 2893
rect 7371 2873 7480 2893
rect 7342 2864 7480 2873
rect 7136 2863 7173 2864
rect 7192 2812 7228 2864
rect 7247 2863 7284 2864
rect 7343 2863 7380 2864
rect 5412 2793 5422 2811
rect 5440 2810 6045 2811
rect 6663 2810 6704 2811
rect 5440 2805 5461 2810
rect 5440 2793 5452 2805
rect 6555 2803 6704 2810
rect 5412 2785 5452 2793
rect 5495 2792 5521 2793
rect 5412 2783 5449 2785
rect 5495 2774 6049 2792
rect 6555 2783 6673 2803
rect 6693 2783 6704 2803
rect 6555 2775 6704 2783
rect 6771 2807 7130 2811
rect 6771 2802 7093 2807
rect 6771 2778 6884 2802
rect 6908 2783 7093 2802
rect 7117 2783 7130 2807
rect 6908 2778 7130 2783
rect 6771 2775 7130 2778
rect 7192 2775 7227 2812
rect 7295 2809 7395 2812
rect 7295 2805 7362 2809
rect 7295 2779 7307 2805
rect 7333 2783 7362 2805
rect 7388 2783 7395 2809
rect 7333 2779 7395 2783
rect 7295 2775 7395 2779
rect 5070 2765 5107 2774
rect 4782 2723 4819 2724
rect 4732 2714 4819 2723
rect 4732 2694 4790 2714
rect 4810 2694 4819 2714
rect 4732 2684 4819 2694
rect 4878 2714 4915 2724
rect 4878 2694 4886 2714
rect 4906 2694 4915 2714
rect 5415 2715 5452 2721
rect 5495 2715 5521 2774
rect 6028 2755 6049 2774
rect 5415 2712 5521 2715
rect 5073 2699 5110 2703
rect 4732 2683 4763 2684
rect 4878 2623 4915 2694
rect 4665 2599 4915 2623
rect 5071 2693 5110 2699
rect 5071 2675 5082 2693
rect 5100 2675 5110 2693
rect 5415 2694 5424 2712
rect 5442 2698 5521 2712
rect 5606 2730 5856 2754
rect 5442 2696 5518 2698
rect 5442 2694 5452 2696
rect 5415 2684 5452 2694
rect 5071 2666 5110 2675
rect 2902 2576 2937 2577
rect 2879 2571 2937 2576
rect 2879 2551 2882 2571
rect 2902 2557 2937 2571
rect 2957 2557 2966 2577
rect 2902 2549 2966 2557
rect 2928 2548 2966 2549
rect 2929 2547 2966 2548
rect 3032 2581 3068 2582
rect 3140 2581 3176 2582
rect 3032 2575 3176 2581
rect 3032 2573 3093 2575
rect 3032 2553 3040 2573
rect 3060 2553 3093 2573
rect 3032 2549 3093 2553
rect 3118 2573 3176 2575
rect 3118 2553 3148 2573
rect 3168 2553 3176 2573
rect 3118 2549 3176 2553
rect 3032 2547 3176 2549
rect 3242 2577 3280 2585
rect 3348 2581 3384 2582
rect 3242 2557 3251 2577
rect 3271 2557 3280 2577
rect 3242 2548 3280 2557
rect 3299 2574 3384 2581
rect 3299 2554 3306 2574
rect 3327 2573 3384 2574
rect 3327 2554 3356 2573
rect 3299 2553 3356 2554
rect 3376 2553 3384 2573
rect 3242 2547 3279 2548
rect 3299 2547 3384 2553
rect 3450 2577 3488 2585
rect 3561 2581 3597 2582
rect 3450 2557 3459 2577
rect 3479 2557 3488 2577
rect 3450 2548 3488 2557
rect 3512 2573 3597 2581
rect 3512 2553 3569 2573
rect 3589 2553 3597 2573
rect 3450 2547 3487 2548
rect 3512 2547 3597 2553
rect 3663 2577 3701 2585
rect 3663 2557 3672 2577
rect 3692 2557 3701 2577
rect 3663 2548 3701 2557
rect 4457 2575 4494 2598
rect 5071 2588 5106 2666
rect 5420 2619 5451 2684
rect 5606 2659 5643 2730
rect 5758 2669 5789 2670
rect 5606 2639 5615 2659
rect 5635 2639 5643 2659
rect 5606 2629 5643 2639
rect 5702 2659 5789 2669
rect 5702 2639 5711 2659
rect 5731 2639 5789 2659
rect 5702 2630 5789 2639
rect 5702 2629 5739 2630
rect 5068 2578 5106 2588
rect 5419 2610 5456 2619
rect 5419 2592 5429 2610
rect 5447 2592 5456 2610
rect 5419 2582 5456 2592
rect 4457 2574 4627 2575
rect 5068 2574 5078 2578
rect 4457 2560 5078 2574
rect 5096 2560 5106 2578
rect 5758 2577 5789 2630
rect 5819 2659 5856 2730
rect 6027 2735 6420 2755
rect 6440 2735 6443 2755
rect 6771 2754 6802 2775
rect 7192 2754 7228 2775
rect 6614 2753 6651 2754
rect 6027 2730 6443 2735
rect 6613 2744 6651 2753
rect 6027 2729 6368 2730
rect 5971 2669 6002 2670
rect 5819 2639 5828 2659
rect 5848 2639 5856 2659
rect 5819 2629 5856 2639
rect 5915 2662 6002 2669
rect 5915 2659 5976 2662
rect 5915 2639 5924 2659
rect 5944 2642 5976 2659
rect 5997 2642 6002 2662
rect 5944 2639 6002 2642
rect 5915 2632 6002 2639
rect 6027 2659 6064 2729
rect 6330 2728 6367 2729
rect 6613 2724 6622 2744
rect 6642 2724 6651 2744
rect 6613 2716 6651 2724
rect 6717 2748 6802 2754
rect 6827 2753 6864 2754
rect 6717 2728 6725 2748
rect 6745 2728 6802 2748
rect 6717 2720 6802 2728
rect 6826 2744 6864 2753
rect 6826 2724 6835 2744
rect 6855 2724 6864 2744
rect 6717 2719 6753 2720
rect 6826 2716 6864 2724
rect 6930 2748 7015 2754
rect 7035 2753 7072 2754
rect 6930 2728 6938 2748
rect 6958 2747 7015 2748
rect 6958 2728 6987 2747
rect 6930 2727 6987 2728
rect 7008 2727 7015 2747
rect 6930 2720 7015 2727
rect 7034 2744 7072 2753
rect 7034 2724 7043 2744
rect 7063 2724 7072 2744
rect 6930 2719 6966 2720
rect 7034 2716 7072 2724
rect 7138 2749 7282 2754
rect 7138 2748 7197 2749
rect 7138 2728 7146 2748
rect 7166 2729 7197 2748
rect 7221 2748 7282 2749
rect 7221 2729 7254 2748
rect 7166 2728 7254 2729
rect 7274 2728 7282 2748
rect 7138 2720 7282 2728
rect 7138 2719 7174 2720
rect 7246 2719 7282 2720
rect 7348 2753 7385 2754
rect 7348 2752 7386 2753
rect 7348 2744 7412 2752
rect 7348 2724 7357 2744
rect 7377 2730 7412 2744
rect 7432 2730 7435 2750
rect 7377 2725 7435 2730
rect 7377 2724 7412 2725
rect 6614 2687 6651 2716
rect 6615 2685 6651 2687
rect 6827 2685 6864 2716
rect 6179 2669 6215 2670
rect 6027 2639 6036 2659
rect 6056 2639 6064 2659
rect 5915 2630 5971 2632
rect 5915 2629 5952 2630
rect 6027 2629 6064 2639
rect 6123 2659 6271 2669
rect 6371 2666 6467 2668
rect 6123 2639 6132 2659
rect 6152 2639 6242 2659
rect 6262 2639 6271 2659
rect 6123 2630 6271 2639
rect 6329 2659 6467 2666
rect 6615 2663 6864 2685
rect 7035 2684 7072 2716
rect 7348 2712 7412 2724
rect 7452 2686 7479 2864
rect 7311 2684 7479 2686
rect 7035 2680 7479 2684
rect 6329 2639 6338 2659
rect 6358 2639 6467 2659
rect 7035 2661 7084 2680
rect 7104 2661 7479 2680
rect 7035 2658 7479 2661
rect 7311 2657 7479 2658
rect 7500 2683 7531 3077
rect 7500 2657 7505 2683
rect 7524 2657 7531 2683
rect 7500 2654 7531 2657
rect 6329 2630 6467 2639
rect 6123 2629 6160 2630
rect 6179 2578 6215 2630
rect 6234 2629 6271 2630
rect 6330 2629 6367 2630
rect 5650 2576 5691 2577
rect 4457 2554 5106 2560
rect 5542 2569 5691 2576
rect 4457 2553 5105 2554
rect 5068 2551 5105 2553
rect 5542 2549 5660 2569
rect 5680 2549 5691 2569
rect 3663 2547 3700 2548
rect 3086 2526 3122 2547
rect 3512 2526 3543 2547
rect 5542 2541 5691 2549
rect 5758 2573 6117 2577
rect 5758 2568 6080 2573
rect 5758 2544 5871 2568
rect 5895 2549 6080 2568
rect 6104 2549 6117 2573
rect 5895 2544 6117 2549
rect 5758 2541 6117 2544
rect 6179 2541 6214 2578
rect 6282 2575 6382 2578
rect 6282 2571 6349 2575
rect 6282 2545 6294 2571
rect 6320 2549 6349 2571
rect 6375 2549 6382 2575
rect 6320 2545 6382 2549
rect 6282 2541 6382 2545
rect 2919 2522 3019 2526
rect 2919 2518 2981 2522
rect 2919 2492 2926 2518
rect 2952 2496 2981 2518
rect 3007 2496 3019 2522
rect 2952 2492 3019 2496
rect 2919 2489 3019 2492
rect 3087 2489 3122 2526
rect 3184 2523 3543 2526
rect 3184 2518 3406 2523
rect 3184 2494 3197 2518
rect 3221 2499 3406 2518
rect 3430 2499 3543 2523
rect 3221 2494 3543 2499
rect 3184 2490 3543 2494
rect 3610 2518 3759 2526
rect 5758 2520 5789 2541
rect 6179 2520 6215 2541
rect 3610 2498 3621 2518
rect 3641 2498 3759 2518
rect 3610 2491 3759 2498
rect 5422 2511 5459 2520
rect 5601 2519 5638 2520
rect 5422 2493 5431 2511
rect 5449 2493 5459 2511
rect 3610 2490 3651 2491
rect 2934 2437 2971 2438
rect 3030 2437 3067 2438
rect 3086 2437 3122 2489
rect 3141 2437 3178 2438
rect 2834 2428 2972 2437
rect 2834 2408 2943 2428
rect 2963 2408 2972 2428
rect 2834 2401 2972 2408
rect 3030 2428 3178 2437
rect 3030 2408 3039 2428
rect 3059 2408 3149 2428
rect 3169 2408 3178 2428
rect 2834 2399 2930 2401
rect 3030 2398 3178 2408
rect 3237 2428 3274 2438
rect 3349 2437 3386 2438
rect 3330 2435 3386 2437
rect 3237 2408 3245 2428
rect 3265 2408 3274 2428
rect 3086 2397 3122 2398
rect 2934 2338 2971 2339
rect 3237 2338 3274 2408
rect 3299 2428 3386 2435
rect 3299 2425 3357 2428
rect 3299 2405 3304 2425
rect 3325 2408 3357 2425
rect 3377 2408 3386 2428
rect 3325 2405 3386 2408
rect 3299 2398 3386 2405
rect 3445 2428 3482 2438
rect 3445 2408 3453 2428
rect 3473 2408 3482 2428
rect 3299 2397 3330 2398
rect 2933 2337 3274 2338
rect 2858 2332 3274 2337
rect 2858 2312 2861 2332
rect 2881 2312 3274 2332
rect 3445 2337 3482 2408
rect 3512 2437 3543 2490
rect 5071 2479 5108 2489
rect 5422 2483 5459 2493
rect 5071 2461 5080 2479
rect 5098 2461 5108 2479
rect 5071 2452 5108 2461
rect 3562 2437 3599 2438
rect 3512 2428 3599 2437
rect 3512 2408 3570 2428
rect 3590 2408 3599 2428
rect 3512 2398 3599 2408
rect 3658 2428 3695 2438
rect 3658 2408 3666 2428
rect 3686 2408 3695 2428
rect 3512 2397 3543 2398
rect 3658 2337 3695 2408
rect 5071 2406 5106 2452
rect 5423 2448 5459 2483
rect 5600 2510 5638 2519
rect 5600 2490 5609 2510
rect 5629 2490 5638 2510
rect 5600 2482 5638 2490
rect 5704 2514 5789 2520
rect 5814 2519 5851 2520
rect 5704 2494 5712 2514
rect 5732 2494 5789 2514
rect 5704 2486 5789 2494
rect 5813 2510 5851 2519
rect 5813 2490 5822 2510
rect 5842 2490 5851 2510
rect 5704 2485 5740 2486
rect 5813 2482 5851 2490
rect 5917 2514 6002 2520
rect 6022 2519 6059 2520
rect 5917 2494 5925 2514
rect 5945 2513 6002 2514
rect 5945 2494 5974 2513
rect 5917 2493 5974 2494
rect 5995 2493 6002 2513
rect 5917 2486 6002 2493
rect 6021 2510 6059 2519
rect 6021 2490 6030 2510
rect 6050 2490 6059 2510
rect 5917 2485 5953 2486
rect 6021 2482 6059 2490
rect 6125 2514 6269 2520
rect 6125 2494 6133 2514
rect 6153 2513 6241 2514
rect 6153 2494 6181 2513
rect 6125 2492 6181 2494
rect 6203 2494 6241 2513
rect 6261 2494 6269 2514
rect 6203 2492 6269 2494
rect 6125 2486 6269 2492
rect 6125 2485 6161 2486
rect 6233 2485 6269 2486
rect 6335 2519 6372 2520
rect 6335 2518 6373 2519
rect 6335 2510 6399 2518
rect 6335 2490 6344 2510
rect 6364 2496 6399 2510
rect 6419 2496 6422 2516
rect 6364 2491 6422 2496
rect 6364 2490 6399 2491
rect 5601 2453 5638 2482
rect 5421 2407 5459 2448
rect 5602 2451 5638 2453
rect 5814 2451 5851 2482
rect 5602 2429 5851 2451
rect 6022 2450 6059 2482
rect 6335 2478 6399 2490
rect 6439 2452 6466 2630
rect 6298 2450 6466 2452
rect 6022 2424 6466 2450
rect 6023 2407 6047 2424
rect 6298 2423 6466 2424
rect 6834 2452 7084 2476
rect 5070 2400 5108 2406
rect 4481 2382 5108 2400
rect 5421 2389 6048 2407
rect 5421 2383 5459 2389
rect 3445 2313 3695 2337
rect 4063 2365 4231 2366
rect 4482 2365 4506 2382
rect 4063 2339 4507 2365
rect 4063 2337 4231 2339
rect 2443 2200 2476 2260
rect 2245 2193 2413 2195
rect 1969 2167 2413 2193
rect 2245 2166 2413 2167
rect 2442 2189 2479 2200
rect 2442 2170 2448 2189
rect 2471 2170 2479 2189
rect 906 2126 942 2127
rect 754 2096 763 2116
rect 783 2096 791 2116
rect 642 2087 698 2089
rect 642 2086 679 2087
rect 754 2086 791 2096
rect 850 2116 998 2126
rect 1098 2123 1194 2125
rect 850 2096 859 2116
rect 879 2096 969 2116
rect 989 2096 998 2116
rect 850 2087 998 2096
rect 1056 2116 1194 2123
rect 1056 2096 1065 2116
rect 1085 2096 1194 2116
rect 1056 2087 1194 2096
rect 850 2086 887 2087
rect 906 2035 942 2087
rect 961 2086 998 2087
rect 1057 2086 1094 2087
rect 377 2033 418 2034
rect 139 1869 178 2018
rect 269 2026 418 2033
rect 269 2006 387 2026
rect 407 2006 418 2026
rect 269 1998 418 2006
rect 485 2030 844 2034
rect 485 2025 807 2030
rect 485 2001 598 2025
rect 622 2006 807 2025
rect 831 2006 844 2030
rect 622 2001 844 2006
rect 485 1998 844 2001
rect 906 1998 941 2035
rect 1009 2032 1109 2035
rect 1009 2028 1076 2032
rect 1009 2002 1021 2028
rect 1047 2006 1076 2028
rect 1102 2006 1109 2032
rect 1047 2002 1109 2006
rect 1009 1998 1109 2002
rect 485 1977 516 1998
rect 906 1977 942 1998
rect 328 1976 365 1977
rect 327 1967 365 1976
rect 327 1947 336 1967
rect 356 1947 365 1967
rect 327 1939 365 1947
rect 431 1971 516 1977
rect 541 1976 578 1977
rect 431 1951 439 1971
rect 459 1951 516 1971
rect 431 1943 516 1951
rect 540 1967 578 1976
rect 540 1947 549 1967
rect 569 1947 578 1967
rect 431 1942 467 1943
rect 540 1939 578 1947
rect 644 1971 729 1977
rect 749 1976 786 1977
rect 644 1951 652 1971
rect 672 1970 729 1971
rect 672 1951 701 1970
rect 644 1950 701 1951
rect 722 1950 729 1970
rect 644 1943 729 1950
rect 748 1967 786 1976
rect 748 1947 757 1967
rect 777 1947 786 1967
rect 644 1942 680 1943
rect 748 1939 786 1947
rect 852 1972 996 1977
rect 852 1971 917 1972
rect 852 1951 860 1971
rect 880 1951 917 1971
rect 939 1971 996 1972
rect 939 1951 968 1971
rect 988 1951 996 1971
rect 852 1943 996 1951
rect 852 1942 888 1943
rect 960 1942 996 1943
rect 1062 1976 1099 1977
rect 1062 1975 1100 1976
rect 1062 1967 1126 1975
rect 1062 1947 1071 1967
rect 1091 1953 1126 1967
rect 1146 1953 1149 1973
rect 1091 1948 1149 1953
rect 1091 1947 1126 1948
rect 328 1910 365 1939
rect 329 1908 365 1910
rect 541 1908 578 1939
rect 329 1886 578 1908
rect 749 1907 786 1939
rect 1062 1935 1126 1947
rect 1166 1909 1193 2087
rect 1025 1907 1193 1909
rect 749 1881 1193 1907
rect 1345 2006 1595 2030
rect 1345 1935 1382 2006
rect 1497 1945 1528 1946
rect 1345 1915 1354 1935
rect 1374 1915 1382 1935
rect 1345 1905 1382 1915
rect 1441 1935 1528 1945
rect 1441 1915 1450 1935
rect 1470 1915 1528 1935
rect 1441 1906 1528 1915
rect 1441 1905 1478 1906
rect 749 1871 771 1881
rect 1025 1880 1193 1881
rect 709 1869 771 1871
rect 139 1862 771 1869
rect 138 1853 771 1862
rect 1497 1853 1528 1906
rect 1558 1935 1595 2006
rect 1766 2011 2159 2031
rect 2179 2011 2182 2031
rect 1766 2006 2182 2011
rect 1766 2005 2107 2006
rect 1710 1945 1741 1946
rect 1558 1915 1567 1935
rect 1587 1915 1595 1935
rect 1558 1905 1595 1915
rect 1654 1938 1741 1945
rect 1654 1935 1715 1938
rect 1654 1915 1663 1935
rect 1683 1918 1715 1935
rect 1736 1918 1741 1938
rect 1683 1915 1741 1918
rect 1654 1908 1741 1915
rect 1766 1935 1803 2005
rect 2069 2004 2106 2005
rect 1918 1945 1954 1946
rect 1766 1915 1775 1935
rect 1795 1915 1803 1935
rect 1654 1906 1710 1908
rect 1654 1905 1691 1906
rect 1766 1905 1803 1915
rect 1862 1935 2010 1945
rect 2110 1942 2206 1944
rect 1862 1915 1871 1935
rect 1891 1915 1981 1935
rect 2001 1915 2010 1935
rect 1862 1906 2010 1915
rect 2068 1935 2206 1942
rect 2068 1915 2077 1935
rect 2097 1915 2206 1935
rect 2068 1906 2206 1915
rect 1862 1905 1899 1906
rect 1918 1854 1954 1906
rect 1973 1905 2010 1906
rect 2069 1905 2106 1906
rect 138 1835 148 1853
rect 166 1852 771 1853
rect 1389 1852 1430 1853
rect 166 1847 187 1852
rect 166 1835 178 1847
rect 1281 1845 1430 1852
rect 138 1827 178 1835
rect 221 1834 247 1835
rect 138 1825 175 1827
rect 221 1816 775 1834
rect 1281 1825 1399 1845
rect 1419 1825 1430 1845
rect 1281 1817 1430 1825
rect 1497 1849 1856 1853
rect 1497 1844 1819 1849
rect 1497 1820 1610 1844
rect 1634 1825 1819 1844
rect 1843 1825 1856 1849
rect 1634 1820 1856 1825
rect 1497 1817 1856 1820
rect 1918 1817 1953 1854
rect 2021 1851 2121 1854
rect 2021 1847 2088 1851
rect 2021 1821 2033 1847
rect 2059 1825 2088 1847
rect 2114 1825 2121 1851
rect 2059 1821 2121 1825
rect 2021 1817 2121 1821
rect 141 1757 178 1763
rect 221 1757 247 1816
rect 754 1797 775 1816
rect 141 1754 247 1757
rect 141 1736 150 1754
rect 168 1740 247 1754
rect 332 1772 582 1796
rect 168 1738 244 1740
rect 168 1736 178 1738
rect 141 1726 178 1736
rect 146 1661 177 1726
rect 332 1701 369 1772
rect 484 1711 515 1712
rect 332 1681 341 1701
rect 361 1681 369 1701
rect 332 1671 369 1681
rect 428 1701 515 1711
rect 428 1681 437 1701
rect 457 1681 515 1701
rect 428 1672 515 1681
rect 428 1671 465 1672
rect 145 1652 182 1661
rect 145 1634 155 1652
rect 173 1634 182 1652
rect 145 1624 182 1634
rect 484 1619 515 1672
rect 545 1701 582 1772
rect 753 1777 1146 1797
rect 1166 1777 1169 1797
rect 1497 1796 1528 1817
rect 1918 1796 1954 1817
rect 1340 1795 1377 1796
rect 753 1772 1169 1777
rect 1339 1786 1377 1795
rect 753 1771 1094 1772
rect 697 1711 728 1712
rect 545 1681 554 1701
rect 574 1681 582 1701
rect 545 1671 582 1681
rect 641 1704 728 1711
rect 641 1701 702 1704
rect 641 1681 650 1701
rect 670 1684 702 1701
rect 723 1684 728 1704
rect 670 1681 728 1684
rect 641 1674 728 1681
rect 753 1701 790 1771
rect 1056 1770 1093 1771
rect 1339 1766 1348 1786
rect 1368 1766 1377 1786
rect 1339 1758 1377 1766
rect 1443 1790 1528 1796
rect 1553 1795 1590 1796
rect 1443 1770 1451 1790
rect 1471 1770 1528 1790
rect 1443 1762 1528 1770
rect 1552 1786 1590 1795
rect 1552 1766 1561 1786
rect 1581 1766 1590 1786
rect 1443 1761 1479 1762
rect 1552 1758 1590 1766
rect 1656 1790 1741 1796
rect 1761 1795 1798 1796
rect 1656 1770 1664 1790
rect 1684 1789 1741 1790
rect 1684 1770 1713 1789
rect 1656 1769 1713 1770
rect 1734 1769 1741 1789
rect 1656 1762 1741 1769
rect 1760 1786 1798 1795
rect 1760 1766 1769 1786
rect 1789 1766 1798 1786
rect 1656 1761 1692 1762
rect 1760 1758 1798 1766
rect 1864 1790 2008 1796
rect 1864 1770 1872 1790
rect 1892 1770 1924 1790
rect 1948 1770 1980 1790
rect 2000 1770 2008 1790
rect 1864 1762 2008 1770
rect 1864 1761 1900 1762
rect 1972 1761 2008 1762
rect 2074 1795 2111 1796
rect 2074 1794 2112 1795
rect 2074 1786 2138 1794
rect 2074 1766 2083 1786
rect 2103 1772 2138 1786
rect 2158 1772 2161 1792
rect 2103 1767 2161 1772
rect 2103 1766 2138 1767
rect 1340 1729 1377 1758
rect 1341 1727 1377 1729
rect 1553 1727 1590 1758
rect 905 1711 941 1712
rect 753 1681 762 1701
rect 782 1681 790 1701
rect 641 1672 697 1674
rect 641 1671 678 1672
rect 753 1671 790 1681
rect 849 1701 997 1711
rect 1097 1708 1193 1710
rect 849 1681 858 1701
rect 878 1681 968 1701
rect 988 1681 997 1701
rect 849 1672 997 1681
rect 1055 1701 1193 1708
rect 1341 1705 1590 1727
rect 1761 1726 1798 1758
rect 2074 1754 2138 1766
rect 2178 1728 2205 1906
rect 2037 1726 2205 1728
rect 1761 1722 2205 1726
rect 1055 1681 1064 1701
rect 1084 1681 1193 1701
rect 1761 1703 1810 1722
rect 1830 1703 2205 1722
rect 1761 1700 2205 1703
rect 2037 1699 2205 1700
rect 1055 1672 1193 1681
rect 849 1671 886 1672
rect 905 1620 941 1672
rect 960 1671 997 1672
rect 1056 1671 1093 1672
rect 376 1618 417 1619
rect 268 1611 417 1618
rect 268 1591 386 1611
rect 406 1591 417 1611
rect 268 1583 417 1591
rect 484 1615 843 1619
rect 484 1610 806 1615
rect 484 1586 597 1610
rect 621 1591 806 1610
rect 830 1591 843 1615
rect 621 1586 843 1591
rect 484 1583 843 1586
rect 905 1583 940 1620
rect 1008 1617 1108 1620
rect 1008 1613 1075 1617
rect 1008 1587 1020 1613
rect 1046 1591 1075 1613
rect 1101 1591 1108 1617
rect 1046 1587 1108 1591
rect 1008 1583 1108 1587
rect 484 1562 515 1583
rect 905 1562 941 1583
rect 148 1553 185 1562
rect 327 1561 364 1562
rect 148 1535 157 1553
rect 175 1535 185 1553
rect 148 1525 185 1535
rect 149 1490 185 1525
rect 326 1552 364 1561
rect 326 1532 335 1552
rect 355 1532 364 1552
rect 326 1524 364 1532
rect 430 1556 515 1562
rect 540 1561 577 1562
rect 430 1536 438 1556
rect 458 1536 515 1556
rect 430 1528 515 1536
rect 539 1552 577 1561
rect 539 1532 548 1552
rect 568 1532 577 1552
rect 430 1527 466 1528
rect 539 1524 577 1532
rect 643 1556 728 1562
rect 748 1561 785 1562
rect 643 1536 651 1556
rect 671 1555 728 1556
rect 671 1536 700 1555
rect 643 1535 700 1536
rect 721 1535 728 1555
rect 643 1528 728 1535
rect 747 1552 785 1561
rect 747 1532 756 1552
rect 776 1532 785 1552
rect 643 1527 679 1528
rect 747 1524 785 1532
rect 851 1556 995 1562
rect 851 1536 859 1556
rect 879 1555 967 1556
rect 879 1536 907 1555
rect 851 1534 907 1536
rect 929 1536 967 1555
rect 987 1536 995 1556
rect 929 1534 995 1536
rect 851 1528 995 1534
rect 851 1527 887 1528
rect 959 1527 995 1528
rect 1061 1561 1098 1562
rect 1061 1560 1099 1561
rect 1061 1552 1125 1560
rect 1061 1532 1070 1552
rect 1090 1538 1125 1552
rect 1145 1538 1148 1558
rect 1090 1533 1148 1538
rect 1090 1532 1125 1533
rect 327 1495 364 1524
rect 147 1449 185 1490
rect 328 1493 364 1495
rect 540 1493 577 1524
rect 328 1471 577 1493
rect 748 1492 785 1524
rect 1061 1520 1125 1532
rect 1165 1494 1192 1672
rect 1024 1492 1192 1494
rect 748 1466 1192 1492
rect 749 1449 773 1466
rect 1024 1465 1192 1466
rect 147 1431 774 1449
rect 1400 1445 1650 1469
rect 147 1425 185 1431
rect 147 1401 184 1425
rect 147 1377 182 1401
rect 145 1368 182 1377
rect 145 1350 155 1368
rect 173 1350 182 1368
rect 145 1340 182 1350
rect 1400 1374 1437 1445
rect 1552 1384 1583 1385
rect 1400 1354 1409 1374
rect 1429 1354 1437 1374
rect 1400 1344 1437 1354
rect 1496 1374 1583 1384
rect 1496 1354 1505 1374
rect 1525 1354 1583 1374
rect 1496 1345 1583 1354
rect 1496 1344 1533 1345
rect 1552 1292 1583 1345
rect 1613 1374 1650 1445
rect 1821 1450 2214 1470
rect 2234 1450 2237 1470
rect 1821 1445 2237 1450
rect 1821 1444 2162 1445
rect 1765 1384 1796 1385
rect 1613 1354 1622 1374
rect 1642 1354 1650 1374
rect 1613 1344 1650 1354
rect 1709 1377 1796 1384
rect 1709 1374 1770 1377
rect 1709 1354 1718 1374
rect 1738 1357 1770 1374
rect 1791 1357 1796 1377
rect 1738 1354 1796 1357
rect 1709 1347 1796 1354
rect 1821 1374 1858 1444
rect 2124 1443 2161 1444
rect 1973 1384 2009 1385
rect 1821 1354 1830 1374
rect 1850 1354 1858 1374
rect 1709 1345 1765 1347
rect 1709 1344 1746 1345
rect 1821 1344 1858 1354
rect 1917 1374 2065 1384
rect 2165 1381 2261 1383
rect 1917 1354 1926 1374
rect 1946 1354 2036 1374
rect 2056 1354 2065 1374
rect 1917 1345 2065 1354
rect 2123 1374 2261 1381
rect 2123 1354 2132 1374
rect 2152 1354 2261 1374
rect 2123 1345 2261 1354
rect 1917 1344 1954 1345
rect 1973 1293 2009 1345
rect 2028 1344 2065 1345
rect 2124 1344 2161 1345
rect 1444 1291 1485 1292
rect 1336 1284 1485 1291
rect 148 1276 185 1278
rect 148 1275 796 1276
rect 147 1269 796 1275
rect 147 1251 157 1269
rect 175 1255 796 1269
rect 1336 1264 1454 1284
rect 1474 1264 1485 1284
rect 1336 1256 1485 1264
rect 1552 1288 1911 1292
rect 1552 1283 1874 1288
rect 1552 1259 1665 1283
rect 1689 1264 1874 1283
rect 1898 1264 1911 1288
rect 1689 1259 1911 1264
rect 1552 1256 1911 1259
rect 1973 1256 2008 1293
rect 2076 1290 2176 1293
rect 2076 1286 2143 1290
rect 2076 1260 2088 1286
rect 2114 1264 2143 1286
rect 2169 1264 2176 1290
rect 2114 1260 2176 1264
rect 2076 1256 2176 1260
rect 175 1251 185 1255
rect 626 1254 796 1255
rect 147 1241 185 1251
rect 147 1163 182 1241
rect 759 1231 796 1254
rect 1552 1235 1583 1256
rect 1973 1235 2009 1256
rect 1395 1234 1432 1235
rect 143 1154 182 1163
rect 143 1136 153 1154
rect 171 1136 182 1154
rect 143 1130 182 1136
rect 338 1206 588 1230
rect 338 1135 375 1206
rect 490 1145 521 1146
rect 143 1126 180 1130
rect 338 1115 347 1135
rect 367 1115 375 1135
rect 338 1105 375 1115
rect 434 1135 521 1145
rect 434 1115 443 1135
rect 463 1115 521 1135
rect 434 1106 521 1115
rect 434 1105 471 1106
rect 146 1055 183 1064
rect 144 1037 155 1055
rect 173 1037 183 1055
rect 490 1053 521 1106
rect 551 1135 588 1206
rect 759 1211 1152 1231
rect 1172 1211 1175 1231
rect 759 1206 1175 1211
rect 1394 1225 1432 1234
rect 759 1205 1100 1206
rect 1394 1205 1403 1225
rect 1423 1205 1432 1225
rect 703 1145 734 1146
rect 551 1115 560 1135
rect 580 1115 588 1135
rect 551 1105 588 1115
rect 647 1138 734 1145
rect 647 1135 708 1138
rect 647 1115 656 1135
rect 676 1118 708 1135
rect 729 1118 734 1138
rect 676 1115 734 1118
rect 647 1108 734 1115
rect 759 1135 796 1205
rect 1062 1204 1099 1205
rect 1394 1197 1432 1205
rect 1498 1229 1583 1235
rect 1608 1234 1645 1235
rect 1498 1209 1506 1229
rect 1526 1209 1583 1229
rect 1498 1201 1583 1209
rect 1607 1225 1645 1234
rect 1607 1205 1616 1225
rect 1636 1205 1645 1225
rect 1498 1200 1534 1201
rect 1607 1197 1645 1205
rect 1711 1229 1796 1235
rect 1816 1234 1853 1235
rect 1711 1209 1719 1229
rect 1739 1228 1796 1229
rect 1739 1209 1768 1228
rect 1711 1208 1768 1209
rect 1789 1208 1796 1228
rect 1711 1201 1796 1208
rect 1815 1225 1853 1234
rect 1815 1205 1824 1225
rect 1844 1205 1853 1225
rect 1711 1200 1747 1201
rect 1815 1197 1853 1205
rect 1919 1229 2063 1235
rect 1919 1209 1927 1229
rect 1947 1228 2035 1229
rect 1947 1209 1980 1228
rect 2003 1209 2035 1228
rect 2055 1209 2063 1229
rect 1919 1201 2063 1209
rect 1919 1200 1955 1201
rect 2027 1200 2063 1201
rect 2129 1234 2166 1235
rect 2129 1233 2167 1234
rect 2129 1225 2193 1233
rect 2129 1205 2138 1225
rect 2158 1211 2193 1225
rect 2213 1211 2216 1231
rect 2158 1206 2216 1211
rect 2158 1205 2193 1206
rect 1395 1168 1432 1197
rect 1396 1166 1432 1168
rect 1608 1166 1645 1197
rect 911 1145 947 1146
rect 759 1115 768 1135
rect 788 1115 796 1135
rect 647 1106 703 1108
rect 647 1105 684 1106
rect 759 1105 796 1115
rect 855 1135 1003 1145
rect 1396 1144 1645 1166
rect 1816 1165 1853 1197
rect 2129 1193 2193 1205
rect 2233 1167 2260 1345
rect 2092 1165 2260 1167
rect 1816 1154 2260 1165
rect 2323 1165 2353 2166
rect 2442 2159 2479 2170
rect 4063 2159 4090 2337
rect 4130 2299 4194 2311
rect 4470 2307 4507 2339
rect 4678 2338 4927 2360
rect 4678 2307 4715 2338
rect 4891 2336 4927 2338
rect 5070 2341 5108 2382
rect 4891 2307 4928 2336
rect 4130 2298 4165 2299
rect 4107 2293 4165 2298
rect 4107 2273 4110 2293
rect 4130 2279 4165 2293
rect 4185 2279 4194 2299
rect 4130 2271 4194 2279
rect 4156 2270 4194 2271
rect 4157 2269 4194 2270
rect 4260 2303 4296 2304
rect 4368 2303 4404 2304
rect 4260 2297 4404 2303
rect 4260 2295 4326 2297
rect 4260 2275 4268 2295
rect 4288 2276 4326 2295
rect 4348 2295 4404 2297
rect 4348 2276 4376 2295
rect 4288 2275 4376 2276
rect 4396 2275 4404 2295
rect 4260 2269 4404 2275
rect 4470 2299 4508 2307
rect 4576 2303 4612 2304
rect 4470 2279 4479 2299
rect 4499 2279 4508 2299
rect 4470 2270 4508 2279
rect 4527 2296 4612 2303
rect 4527 2276 4534 2296
rect 4555 2295 4612 2296
rect 4555 2276 4584 2295
rect 4527 2275 4584 2276
rect 4604 2275 4612 2295
rect 4470 2269 4507 2270
rect 4527 2269 4612 2275
rect 4678 2299 4716 2307
rect 4789 2303 4825 2304
rect 4678 2279 4687 2299
rect 4707 2279 4716 2299
rect 4678 2270 4716 2279
rect 4740 2295 4825 2303
rect 4740 2275 4797 2295
rect 4817 2275 4825 2295
rect 4678 2269 4715 2270
rect 4740 2269 4825 2275
rect 4891 2299 4929 2307
rect 4891 2279 4900 2299
rect 4920 2279 4929 2299
rect 4891 2270 4929 2279
rect 5070 2306 5106 2341
rect 5423 2337 5458 2383
rect 6834 2381 6871 2452
rect 6986 2391 7017 2392
rect 6834 2361 6843 2381
rect 6863 2361 6871 2381
rect 6834 2351 6871 2361
rect 6930 2381 7017 2391
rect 6930 2361 6939 2381
rect 6959 2361 7017 2381
rect 6930 2352 7017 2361
rect 6930 2351 6967 2352
rect 5421 2328 5458 2337
rect 5421 2310 5431 2328
rect 5449 2310 5458 2328
rect 5070 2296 5107 2306
rect 5421 2300 5458 2310
rect 6986 2299 7017 2352
rect 7047 2381 7084 2452
rect 7255 2457 7648 2477
rect 7668 2457 7671 2477
rect 7255 2452 7671 2457
rect 7255 2451 7596 2452
rect 7199 2391 7230 2392
rect 7047 2361 7056 2381
rect 7076 2361 7084 2381
rect 7047 2351 7084 2361
rect 7143 2384 7230 2391
rect 7143 2381 7204 2384
rect 7143 2361 7152 2381
rect 7172 2364 7204 2381
rect 7225 2364 7230 2384
rect 7172 2361 7230 2364
rect 7143 2354 7230 2361
rect 7255 2381 7292 2451
rect 7558 2450 7595 2451
rect 7407 2391 7443 2392
rect 7255 2361 7264 2381
rect 7284 2361 7292 2381
rect 7143 2352 7199 2354
rect 7143 2351 7180 2352
rect 7255 2351 7292 2361
rect 7351 2381 7499 2391
rect 7599 2388 7695 2390
rect 7351 2361 7360 2381
rect 7380 2361 7470 2381
rect 7490 2361 7499 2381
rect 7351 2352 7499 2361
rect 7557 2381 7695 2388
rect 7557 2361 7566 2381
rect 7586 2361 7695 2381
rect 7557 2352 7695 2361
rect 7351 2351 7388 2352
rect 7407 2300 7443 2352
rect 7462 2351 7499 2352
rect 7558 2351 7595 2352
rect 6878 2298 6919 2299
rect 5070 2278 5080 2296
rect 5098 2278 5107 2296
rect 4891 2269 4928 2270
rect 5070 2269 5107 2278
rect 6770 2291 6919 2298
rect 6770 2271 6888 2291
rect 6908 2271 6919 2291
rect 4314 2248 4350 2269
rect 4740 2248 4771 2269
rect 6770 2263 6919 2271
rect 6986 2295 7345 2299
rect 6986 2290 7308 2295
rect 6986 2266 7099 2290
rect 7123 2271 7308 2290
rect 7332 2271 7345 2295
rect 7123 2266 7345 2271
rect 6986 2263 7345 2266
rect 7407 2263 7442 2300
rect 7510 2297 7610 2300
rect 7510 2293 7577 2297
rect 7510 2267 7522 2293
rect 7548 2271 7577 2293
rect 7603 2271 7610 2297
rect 7548 2267 7610 2271
rect 7510 2263 7610 2267
rect 4147 2244 4247 2248
rect 4147 2240 4209 2244
rect 4147 2214 4154 2240
rect 4180 2218 4209 2240
rect 4235 2218 4247 2244
rect 4180 2214 4247 2218
rect 4147 2211 4247 2214
rect 4315 2211 4350 2248
rect 4412 2245 4771 2248
rect 4412 2240 4634 2245
rect 4412 2216 4425 2240
rect 4449 2221 4634 2240
rect 4658 2221 4771 2245
rect 4449 2216 4771 2221
rect 4412 2212 4771 2216
rect 4838 2240 4987 2248
rect 6986 2242 7017 2263
rect 7407 2242 7443 2263
rect 6829 2241 6866 2242
rect 4838 2220 4849 2240
rect 4869 2220 4987 2240
rect 5424 2236 5461 2238
rect 5424 2235 6072 2236
rect 4838 2213 4987 2220
rect 5423 2229 6072 2235
rect 4838 2212 4879 2213
rect 4162 2159 4199 2160
rect 4258 2159 4295 2160
rect 4314 2159 4350 2211
rect 4369 2159 4406 2160
rect 4062 2150 4200 2159
rect 2998 2132 3029 2135
rect 2998 2106 3005 2132
rect 3024 2106 3029 2132
rect 2998 1712 3029 2106
rect 3050 2131 3218 2132
rect 3050 2128 3494 2131
rect 3050 2109 3425 2128
rect 3445 2109 3494 2128
rect 4062 2130 4171 2150
rect 4191 2130 4200 2150
rect 3050 2105 3494 2109
rect 3050 2103 3218 2105
rect 3050 1925 3077 2103
rect 3117 2065 3181 2077
rect 3457 2073 3494 2105
rect 3665 2104 3914 2126
rect 4062 2123 4200 2130
rect 4258 2150 4406 2159
rect 4258 2130 4267 2150
rect 4287 2130 4377 2150
rect 4397 2130 4406 2150
rect 4062 2121 4158 2123
rect 4258 2120 4406 2130
rect 4465 2150 4502 2160
rect 4577 2159 4614 2160
rect 4558 2157 4614 2159
rect 4465 2130 4473 2150
rect 4493 2130 4502 2150
rect 4314 2119 4350 2120
rect 3665 2073 3702 2104
rect 3878 2102 3914 2104
rect 3878 2073 3915 2102
rect 3117 2064 3152 2065
rect 3094 2059 3152 2064
rect 3094 2039 3097 2059
rect 3117 2045 3152 2059
rect 3172 2045 3181 2065
rect 3117 2037 3181 2045
rect 3143 2036 3181 2037
rect 3144 2035 3181 2036
rect 3247 2069 3283 2070
rect 3355 2069 3391 2070
rect 3247 2061 3391 2069
rect 3247 2041 3255 2061
rect 3275 2060 3363 2061
rect 3275 2041 3308 2060
rect 3247 2040 3308 2041
rect 3332 2041 3363 2060
rect 3383 2041 3391 2061
rect 3332 2040 3391 2041
rect 3247 2035 3391 2040
rect 3457 2065 3495 2073
rect 3563 2069 3599 2070
rect 3457 2045 3466 2065
rect 3486 2045 3495 2065
rect 3457 2036 3495 2045
rect 3514 2062 3599 2069
rect 3514 2042 3521 2062
rect 3542 2061 3599 2062
rect 3542 2042 3571 2061
rect 3514 2041 3571 2042
rect 3591 2041 3599 2061
rect 3457 2035 3494 2036
rect 3514 2035 3599 2041
rect 3665 2065 3703 2073
rect 3776 2069 3812 2070
rect 3665 2045 3674 2065
rect 3694 2045 3703 2065
rect 3665 2036 3703 2045
rect 3727 2061 3812 2069
rect 3727 2041 3784 2061
rect 3804 2041 3812 2061
rect 3665 2035 3702 2036
rect 3727 2035 3812 2041
rect 3878 2065 3916 2073
rect 3878 2045 3887 2065
rect 3907 2045 3916 2065
rect 4162 2060 4199 2061
rect 4465 2060 4502 2130
rect 4527 2150 4614 2157
rect 4527 2147 4585 2150
rect 4527 2127 4532 2147
rect 4553 2130 4585 2147
rect 4605 2130 4614 2150
rect 4553 2127 4614 2130
rect 4527 2120 4614 2127
rect 4673 2150 4710 2160
rect 4673 2130 4681 2150
rect 4701 2130 4710 2150
rect 4527 2119 4558 2120
rect 4161 2059 4502 2060
rect 3878 2036 3916 2045
rect 4086 2054 4502 2059
rect 3878 2035 3915 2036
rect 3301 2014 3337 2035
rect 3727 2014 3758 2035
rect 4086 2034 4089 2054
rect 4109 2034 4502 2054
rect 4673 2059 4710 2130
rect 4740 2159 4771 2212
rect 5423 2211 5433 2229
rect 5451 2215 6072 2229
rect 5451 2211 5461 2215
rect 5902 2214 6072 2215
rect 5073 2197 5110 2207
rect 5073 2179 5082 2197
rect 5100 2179 5110 2197
rect 5073 2170 5110 2179
rect 5423 2201 5461 2211
rect 4790 2159 4827 2160
rect 4740 2150 4827 2159
rect 4740 2130 4798 2150
rect 4818 2130 4827 2150
rect 4740 2120 4827 2130
rect 4886 2150 4923 2160
rect 4886 2130 4894 2150
rect 4914 2130 4923 2150
rect 4740 2119 4771 2120
rect 4886 2059 4923 2130
rect 5078 2105 5109 2170
rect 5423 2123 5458 2201
rect 6035 2191 6072 2214
rect 6828 2232 6866 2241
rect 6828 2212 6837 2232
rect 6857 2212 6866 2232
rect 6828 2204 6866 2212
rect 6932 2236 7017 2242
rect 7042 2241 7079 2242
rect 6932 2216 6940 2236
rect 6960 2216 7017 2236
rect 6932 2208 7017 2216
rect 7041 2232 7079 2241
rect 7041 2212 7050 2232
rect 7070 2212 7079 2232
rect 6932 2207 6968 2208
rect 7041 2204 7079 2212
rect 7145 2236 7230 2242
rect 7250 2241 7287 2242
rect 7145 2216 7153 2236
rect 7173 2235 7230 2236
rect 7173 2216 7202 2235
rect 7145 2215 7202 2216
rect 7223 2215 7230 2235
rect 7145 2208 7230 2215
rect 7249 2232 7287 2241
rect 7249 2212 7258 2232
rect 7278 2212 7287 2232
rect 7145 2207 7181 2208
rect 7249 2204 7287 2212
rect 7353 2236 7497 2242
rect 7353 2216 7361 2236
rect 7381 2217 7417 2236
rect 7440 2217 7469 2236
rect 7381 2216 7469 2217
rect 7489 2216 7497 2236
rect 7353 2208 7497 2216
rect 7353 2207 7389 2208
rect 7461 2207 7497 2208
rect 7563 2241 7600 2242
rect 7563 2240 7601 2241
rect 7563 2232 7627 2240
rect 7563 2212 7572 2232
rect 7592 2218 7627 2232
rect 7647 2218 7650 2238
rect 7592 2213 7650 2218
rect 7592 2212 7627 2213
rect 5419 2114 5458 2123
rect 5077 2095 5114 2105
rect 5077 2093 5087 2095
rect 5011 2091 5087 2093
rect 4673 2035 4923 2059
rect 5008 2077 5087 2091
rect 5105 2077 5114 2095
rect 5419 2096 5429 2114
rect 5447 2096 5458 2114
rect 5419 2090 5458 2096
rect 5614 2166 5864 2190
rect 5614 2095 5651 2166
rect 5766 2105 5797 2106
rect 5419 2086 5456 2090
rect 5008 2074 5114 2077
rect 4480 2015 4501 2034
rect 5008 2015 5034 2074
rect 5077 2068 5114 2074
rect 5614 2075 5623 2095
rect 5643 2075 5651 2095
rect 5614 2065 5651 2075
rect 5710 2095 5797 2105
rect 5710 2075 5719 2095
rect 5739 2075 5797 2095
rect 5710 2066 5797 2075
rect 5710 2065 5747 2066
rect 5422 2015 5459 2024
rect 3134 2010 3234 2014
rect 3134 2006 3196 2010
rect 3134 1980 3141 2006
rect 3167 1984 3196 2006
rect 3222 1984 3234 2010
rect 3167 1980 3234 1984
rect 3134 1977 3234 1980
rect 3302 1977 3337 2014
rect 3399 2011 3758 2014
rect 3399 2006 3621 2011
rect 3399 1982 3412 2006
rect 3436 1987 3621 2006
rect 3645 1987 3758 2011
rect 3436 1982 3758 1987
rect 3399 1978 3758 1982
rect 3825 2006 3974 2014
rect 3825 1986 3836 2006
rect 3856 1986 3974 2006
rect 4480 1997 5034 2015
rect 5080 2004 5117 2006
rect 5008 1996 5034 1997
rect 5077 1996 5117 2004
rect 3825 1979 3974 1986
rect 5077 1984 5089 1996
rect 5068 1979 5089 1984
rect 3825 1978 3866 1979
rect 4484 1978 5089 1979
rect 5107 1978 5117 1996
rect 3149 1925 3186 1926
rect 3245 1925 3282 1926
rect 3301 1925 3337 1977
rect 3356 1925 3393 1926
rect 3049 1916 3187 1925
rect 3049 1896 3158 1916
rect 3178 1896 3187 1916
rect 3049 1889 3187 1896
rect 3245 1916 3393 1925
rect 3245 1896 3254 1916
rect 3274 1896 3364 1916
rect 3384 1896 3393 1916
rect 3049 1887 3145 1889
rect 3245 1886 3393 1896
rect 3452 1916 3489 1926
rect 3564 1925 3601 1926
rect 3545 1923 3601 1925
rect 3452 1896 3460 1916
rect 3480 1896 3489 1916
rect 3301 1885 3337 1886
rect 3149 1826 3186 1827
rect 3452 1826 3489 1896
rect 3514 1916 3601 1923
rect 3514 1913 3572 1916
rect 3514 1893 3519 1913
rect 3540 1896 3572 1913
rect 3592 1896 3601 1916
rect 3540 1893 3601 1896
rect 3514 1886 3601 1893
rect 3660 1916 3697 1926
rect 3660 1896 3668 1916
rect 3688 1896 3697 1916
rect 3514 1885 3545 1886
rect 3148 1825 3489 1826
rect 3073 1820 3489 1825
rect 3073 1800 3076 1820
rect 3096 1800 3489 1820
rect 3660 1825 3697 1896
rect 3727 1925 3758 1978
rect 4484 1969 5117 1978
rect 5420 1997 5431 2015
rect 5449 1997 5459 2015
rect 5766 2013 5797 2066
rect 5827 2095 5864 2166
rect 6035 2171 6428 2191
rect 6448 2171 6451 2191
rect 6829 2175 6866 2204
rect 6035 2166 6451 2171
rect 6830 2173 6866 2175
rect 7042 2173 7079 2204
rect 6035 2165 6376 2166
rect 5979 2105 6010 2106
rect 5827 2075 5836 2095
rect 5856 2075 5864 2095
rect 5827 2065 5864 2075
rect 5923 2098 6010 2105
rect 5923 2095 5984 2098
rect 5923 2075 5932 2095
rect 5952 2078 5984 2095
rect 6005 2078 6010 2098
rect 5952 2075 6010 2078
rect 5923 2068 6010 2075
rect 6035 2095 6072 2165
rect 6338 2164 6375 2165
rect 6830 2151 7079 2173
rect 7250 2172 7287 2204
rect 7563 2200 7627 2212
rect 7667 2174 7694 2352
rect 7722 2239 7760 4070
rect 8267 4045 8274 4071
rect 8293 4045 8298 4071
rect 8174 3652 8203 3654
rect 8174 3647 8206 3652
rect 8174 3629 8181 3647
rect 8201 3629 8206 3647
rect 8267 3651 8298 4045
rect 8319 4070 8487 4071
rect 8319 4067 8763 4070
rect 8319 4048 8694 4067
rect 8714 4048 8763 4067
rect 9331 4069 9440 4089
rect 9460 4069 9469 4089
rect 8319 4044 8763 4048
rect 8319 4042 8487 4044
rect 8319 3864 8346 4042
rect 8386 4004 8450 4016
rect 8726 4012 8763 4044
rect 8934 4043 9183 4065
rect 9331 4062 9469 4069
rect 9527 4089 9675 4098
rect 9527 4069 9536 4089
rect 9556 4069 9646 4089
rect 9666 4069 9675 4089
rect 9331 4060 9427 4062
rect 9527 4059 9675 4069
rect 9734 4089 9771 4099
rect 9846 4098 9883 4099
rect 9827 4096 9883 4098
rect 9734 4069 9742 4089
rect 9762 4069 9771 4089
rect 9583 4058 9619 4059
rect 8934 4012 8971 4043
rect 9147 4041 9183 4043
rect 9147 4012 9184 4041
rect 8386 4003 8421 4004
rect 8363 3998 8421 4003
rect 8363 3978 8366 3998
rect 8386 3984 8421 3998
rect 8441 3984 8450 4004
rect 8386 3976 8450 3984
rect 8412 3975 8450 3976
rect 8413 3974 8450 3975
rect 8516 4008 8552 4009
rect 8624 4008 8660 4009
rect 8516 4000 8660 4008
rect 8516 3980 8524 4000
rect 8544 3999 8632 4000
rect 8544 3980 8577 3999
rect 8516 3979 8577 3980
rect 8601 3980 8632 3999
rect 8652 3980 8660 4000
rect 8601 3979 8660 3980
rect 8516 3974 8660 3979
rect 8726 4004 8764 4012
rect 8832 4008 8868 4009
rect 8726 3984 8735 4004
rect 8755 3984 8764 4004
rect 8726 3975 8764 3984
rect 8783 4001 8868 4008
rect 8783 3981 8790 4001
rect 8811 4000 8868 4001
rect 8811 3981 8840 4000
rect 8783 3980 8840 3981
rect 8860 3980 8868 4000
rect 8726 3974 8763 3975
rect 8783 3974 8868 3980
rect 8934 4004 8972 4012
rect 9045 4008 9081 4009
rect 8934 3984 8943 4004
rect 8963 3984 8972 4004
rect 8934 3975 8972 3984
rect 8996 4000 9081 4008
rect 8996 3980 9053 4000
rect 9073 3980 9081 4000
rect 8934 3974 8971 3975
rect 8996 3974 9081 3980
rect 9147 4004 9185 4012
rect 9147 3984 9156 4004
rect 9176 3984 9185 4004
rect 9431 3999 9468 4000
rect 9734 3999 9771 4069
rect 9796 4089 9883 4096
rect 9796 4086 9854 4089
rect 9796 4066 9801 4086
rect 9822 4069 9854 4086
rect 9874 4069 9883 4089
rect 9822 4066 9883 4069
rect 9796 4059 9883 4066
rect 9942 4089 9979 4099
rect 9942 4069 9950 4089
rect 9970 4069 9979 4089
rect 9796 4058 9827 4059
rect 9430 3998 9771 3999
rect 9147 3975 9185 3984
rect 9355 3993 9771 3998
rect 9147 3974 9184 3975
rect 8570 3953 8606 3974
rect 8996 3953 9027 3974
rect 9355 3973 9358 3993
rect 9378 3973 9771 3993
rect 9942 3998 9979 4069
rect 10009 4098 10040 4151
rect 10342 4136 10379 4146
rect 10342 4118 10351 4136
rect 10369 4118 10379 4136
rect 10342 4109 10379 4118
rect 10059 4098 10096 4099
rect 10009 4089 10096 4098
rect 10009 4069 10067 4089
rect 10087 4069 10096 4089
rect 10009 4059 10096 4069
rect 10155 4089 10192 4099
rect 10155 4069 10163 4089
rect 10183 4069 10192 4089
rect 10009 4058 10040 4059
rect 10155 3998 10192 4069
rect 10347 4044 10378 4109
rect 10346 4034 10383 4044
rect 10346 4032 10356 4034
rect 10280 4030 10356 4032
rect 9942 3974 10192 3998
rect 10277 4016 10356 4030
rect 10374 4016 10383 4034
rect 10277 4013 10383 4016
rect 9749 3954 9770 3973
rect 10277 3954 10303 4013
rect 10346 4007 10383 4013
rect 8403 3949 8503 3953
rect 8403 3945 8465 3949
rect 8403 3919 8410 3945
rect 8436 3923 8465 3945
rect 8491 3923 8503 3949
rect 8436 3919 8503 3923
rect 8403 3916 8503 3919
rect 8571 3916 8606 3953
rect 8668 3950 9027 3953
rect 8668 3945 8890 3950
rect 8668 3921 8681 3945
rect 8705 3926 8890 3945
rect 8914 3926 9027 3950
rect 8705 3921 9027 3926
rect 8668 3917 9027 3921
rect 9094 3945 9243 3953
rect 9094 3925 9105 3945
rect 9125 3925 9243 3945
rect 9749 3936 10303 3954
rect 10349 3943 10386 3945
rect 10277 3935 10303 3936
rect 10346 3935 10386 3943
rect 9094 3918 9243 3925
rect 10346 3923 10358 3935
rect 10337 3918 10358 3923
rect 9094 3917 9135 3918
rect 9753 3917 10358 3918
rect 10376 3917 10386 3935
rect 8418 3864 8455 3865
rect 8514 3864 8551 3865
rect 8570 3864 8606 3916
rect 8625 3864 8662 3865
rect 8318 3855 8456 3864
rect 8318 3835 8427 3855
rect 8447 3835 8456 3855
rect 8318 3828 8456 3835
rect 8514 3855 8662 3864
rect 8514 3835 8523 3855
rect 8543 3835 8633 3855
rect 8653 3835 8662 3855
rect 8318 3826 8414 3828
rect 8514 3825 8662 3835
rect 8721 3855 8758 3865
rect 8833 3864 8870 3865
rect 8814 3862 8870 3864
rect 8721 3835 8729 3855
rect 8749 3835 8758 3855
rect 8570 3824 8606 3825
rect 8418 3765 8455 3766
rect 8721 3765 8758 3835
rect 8783 3855 8870 3862
rect 8783 3852 8841 3855
rect 8783 3832 8788 3852
rect 8809 3835 8841 3852
rect 8861 3835 8870 3855
rect 8809 3832 8870 3835
rect 8783 3825 8870 3832
rect 8929 3855 8966 3865
rect 8929 3835 8937 3855
rect 8957 3835 8966 3855
rect 8783 3824 8814 3825
rect 8417 3764 8758 3765
rect 8342 3759 8758 3764
rect 8342 3739 8345 3759
rect 8365 3739 8758 3759
rect 8929 3764 8966 3835
rect 8996 3864 9027 3917
rect 9753 3908 10386 3917
rect 9753 3901 10385 3908
rect 9753 3899 9815 3901
rect 9331 3889 9499 3890
rect 9753 3889 9775 3899
rect 9046 3864 9083 3865
rect 8996 3855 9083 3864
rect 8996 3835 9054 3855
rect 9074 3835 9083 3855
rect 8996 3825 9083 3835
rect 9142 3855 9179 3865
rect 9142 3835 9150 3855
rect 9170 3835 9179 3855
rect 8996 3824 9027 3825
rect 9142 3764 9179 3835
rect 8929 3740 9179 3764
rect 9331 3863 9775 3889
rect 9331 3861 9499 3863
rect 9331 3683 9358 3861
rect 9398 3823 9462 3835
rect 9738 3831 9775 3863
rect 9946 3862 10195 3884
rect 9946 3831 9983 3862
rect 10159 3860 10195 3862
rect 10159 3831 10196 3860
rect 9398 3822 9433 3823
rect 9375 3817 9433 3822
rect 9375 3797 9378 3817
rect 9398 3803 9433 3817
rect 9453 3803 9462 3823
rect 9398 3795 9462 3803
rect 9424 3794 9462 3795
rect 9425 3793 9462 3794
rect 9528 3827 9564 3828
rect 9636 3827 9672 3828
rect 9528 3819 9672 3827
rect 9528 3799 9536 3819
rect 9556 3799 9585 3819
rect 9528 3798 9585 3799
rect 9607 3799 9644 3819
rect 9664 3799 9672 3819
rect 9607 3798 9672 3799
rect 9528 3793 9672 3798
rect 9738 3823 9776 3831
rect 9844 3827 9880 3828
rect 9738 3803 9747 3823
rect 9767 3803 9776 3823
rect 9738 3794 9776 3803
rect 9795 3820 9880 3827
rect 9795 3800 9802 3820
rect 9823 3819 9880 3820
rect 9823 3800 9852 3819
rect 9795 3799 9852 3800
rect 9872 3799 9880 3819
rect 9738 3793 9775 3794
rect 9795 3793 9880 3799
rect 9946 3823 9984 3831
rect 10057 3827 10093 3828
rect 9946 3803 9955 3823
rect 9975 3803 9984 3823
rect 9946 3794 9984 3803
rect 10008 3819 10093 3827
rect 10008 3799 10065 3819
rect 10085 3799 10093 3819
rect 9946 3793 9983 3794
rect 10008 3793 10093 3799
rect 10159 3823 10197 3831
rect 10159 3803 10168 3823
rect 10188 3803 10197 3823
rect 10159 3794 10197 3803
rect 10159 3793 10196 3794
rect 9582 3772 9618 3793
rect 10008 3772 10039 3793
rect 9415 3768 9515 3772
rect 9415 3764 9477 3768
rect 9415 3738 9422 3764
rect 9448 3742 9477 3764
rect 9503 3742 9515 3768
rect 9448 3738 9515 3742
rect 9415 3735 9515 3738
rect 9583 3735 9618 3772
rect 9680 3769 10039 3772
rect 9680 3764 9902 3769
rect 9680 3740 9693 3764
rect 9717 3745 9902 3764
rect 9926 3745 10039 3769
rect 9717 3740 10039 3745
rect 9680 3736 10039 3740
rect 10106 3764 10255 3772
rect 10106 3744 10117 3764
rect 10137 3744 10255 3764
rect 10106 3737 10255 3744
rect 10346 3752 10385 3901
rect 10106 3736 10147 3737
rect 9430 3683 9467 3684
rect 9526 3683 9563 3684
rect 9582 3683 9618 3735
rect 9637 3683 9674 3684
rect 9330 3674 9468 3683
rect 9330 3654 9439 3674
rect 9459 3654 9468 3674
rect 8267 3650 8437 3651
rect 8267 3635 8713 3650
rect 9330 3647 9468 3654
rect 9526 3674 9674 3683
rect 9526 3654 9535 3674
rect 9555 3654 9645 3674
rect 9665 3654 9674 3674
rect 9330 3645 9426 3647
rect 8174 3624 8206 3629
rect 8176 2623 8206 3624
rect 8269 3624 8713 3635
rect 8269 3622 8437 3624
rect 8269 3444 8296 3622
rect 8336 3584 8400 3596
rect 8676 3592 8713 3624
rect 8884 3623 9133 3645
rect 9526 3644 9674 3654
rect 9733 3674 9770 3684
rect 9845 3683 9882 3684
rect 9826 3681 9882 3683
rect 9733 3654 9741 3674
rect 9761 3654 9770 3674
rect 9582 3643 9618 3644
rect 8884 3592 8921 3623
rect 9097 3621 9133 3623
rect 9097 3592 9134 3621
rect 8336 3583 8371 3584
rect 8313 3578 8371 3583
rect 8313 3558 8316 3578
rect 8336 3564 8371 3578
rect 8391 3564 8400 3584
rect 8336 3556 8400 3564
rect 8362 3555 8400 3556
rect 8363 3554 8400 3555
rect 8466 3588 8502 3589
rect 8574 3588 8610 3589
rect 8466 3580 8610 3588
rect 8466 3560 8474 3580
rect 8494 3561 8526 3580
rect 8549 3561 8582 3580
rect 8494 3560 8582 3561
rect 8602 3560 8610 3580
rect 8466 3554 8610 3560
rect 8676 3584 8714 3592
rect 8782 3588 8818 3589
rect 8676 3564 8685 3584
rect 8705 3564 8714 3584
rect 8676 3555 8714 3564
rect 8733 3581 8818 3588
rect 8733 3561 8740 3581
rect 8761 3580 8818 3581
rect 8761 3561 8790 3580
rect 8733 3560 8790 3561
rect 8810 3560 8818 3580
rect 8676 3554 8713 3555
rect 8733 3554 8818 3560
rect 8884 3584 8922 3592
rect 8995 3588 9031 3589
rect 8884 3564 8893 3584
rect 8913 3564 8922 3584
rect 8884 3555 8922 3564
rect 8946 3580 9031 3588
rect 8946 3560 9003 3580
rect 9023 3560 9031 3580
rect 8884 3554 8921 3555
rect 8946 3554 9031 3560
rect 9097 3584 9135 3592
rect 9430 3584 9467 3585
rect 9733 3584 9770 3654
rect 9795 3674 9882 3681
rect 9795 3671 9853 3674
rect 9795 3651 9800 3671
rect 9821 3654 9853 3671
rect 9873 3654 9882 3674
rect 9821 3651 9882 3654
rect 9795 3644 9882 3651
rect 9941 3674 9978 3684
rect 9941 3654 9949 3674
rect 9969 3654 9978 3674
rect 9795 3643 9826 3644
rect 9097 3564 9106 3584
rect 9126 3564 9135 3584
rect 9429 3583 9770 3584
rect 9097 3555 9135 3564
rect 9354 3578 9770 3583
rect 9354 3558 9357 3578
rect 9377 3558 9770 3578
rect 9941 3583 9978 3654
rect 10008 3683 10039 3736
rect 10346 3734 10356 3752
rect 10374 3734 10385 3752
rect 10346 3725 10383 3734
rect 10058 3683 10095 3684
rect 10008 3674 10095 3683
rect 10008 3654 10066 3674
rect 10086 3654 10095 3674
rect 10008 3644 10095 3654
rect 10154 3674 10191 3684
rect 10154 3654 10162 3674
rect 10182 3654 10191 3674
rect 10349 3659 10386 3663
rect 10008 3643 10039 3644
rect 10154 3583 10191 3654
rect 9941 3559 10191 3583
rect 10347 3653 10386 3659
rect 10347 3635 10358 3653
rect 10376 3635 10386 3653
rect 10347 3626 10386 3635
rect 9097 3554 9134 3555
rect 8520 3533 8556 3554
rect 8946 3533 8977 3554
rect 9733 3535 9770 3558
rect 10347 3548 10382 3626
rect 10344 3538 10382 3548
rect 9733 3534 9903 3535
rect 10344 3534 10354 3538
rect 8353 3529 8453 3533
rect 8353 3525 8415 3529
rect 8353 3499 8360 3525
rect 8386 3503 8415 3525
rect 8441 3503 8453 3529
rect 8386 3499 8453 3503
rect 8353 3496 8453 3499
rect 8521 3496 8556 3533
rect 8618 3530 8977 3533
rect 8618 3525 8840 3530
rect 8618 3501 8631 3525
rect 8655 3506 8840 3525
rect 8864 3506 8977 3530
rect 8655 3501 8977 3506
rect 8618 3497 8977 3501
rect 9044 3525 9193 3533
rect 9044 3505 9055 3525
rect 9075 3505 9193 3525
rect 9733 3520 10354 3534
rect 10372 3520 10382 3538
rect 9733 3514 10382 3520
rect 9733 3513 10381 3514
rect 10344 3511 10381 3513
rect 9044 3498 9193 3505
rect 9044 3497 9085 3498
rect 8368 3444 8405 3445
rect 8464 3444 8501 3445
rect 8520 3444 8556 3496
rect 8575 3444 8612 3445
rect 8268 3435 8406 3444
rect 8268 3415 8377 3435
rect 8397 3415 8406 3435
rect 8268 3408 8406 3415
rect 8464 3435 8612 3444
rect 8464 3415 8473 3435
rect 8493 3415 8583 3435
rect 8603 3415 8612 3435
rect 8268 3406 8364 3408
rect 8464 3405 8612 3415
rect 8671 3435 8708 3445
rect 8783 3444 8820 3445
rect 8764 3442 8820 3444
rect 8671 3415 8679 3435
rect 8699 3415 8708 3435
rect 8520 3404 8556 3405
rect 8368 3345 8405 3346
rect 8671 3345 8708 3415
rect 8733 3435 8820 3442
rect 8733 3432 8791 3435
rect 8733 3412 8738 3432
rect 8759 3415 8791 3432
rect 8811 3415 8820 3435
rect 8759 3412 8820 3415
rect 8733 3405 8820 3412
rect 8879 3435 8916 3445
rect 8879 3415 8887 3435
rect 8907 3415 8916 3435
rect 8733 3404 8764 3405
rect 8367 3344 8708 3345
rect 8292 3339 8708 3344
rect 8292 3319 8295 3339
rect 8315 3319 8708 3339
rect 8879 3344 8916 3415
rect 8946 3444 8977 3497
rect 8996 3444 9033 3445
rect 8946 3435 9033 3444
rect 8946 3415 9004 3435
rect 9024 3415 9033 3435
rect 8946 3405 9033 3415
rect 9092 3435 9129 3445
rect 9092 3415 9100 3435
rect 9120 3415 9129 3435
rect 8946 3404 8977 3405
rect 9092 3344 9129 3415
rect 10347 3439 10384 3449
rect 10347 3421 10356 3439
rect 10374 3421 10384 3439
rect 10347 3412 10384 3421
rect 10347 3388 10382 3412
rect 10345 3364 10382 3388
rect 10344 3358 10382 3364
rect 8879 3320 9129 3344
rect 9755 3340 10382 3358
rect 9337 3323 9505 3324
rect 9756 3323 9780 3340
rect 9337 3297 9781 3323
rect 9337 3295 9505 3297
rect 9337 3117 9364 3295
rect 9404 3257 9468 3269
rect 9744 3265 9781 3297
rect 9952 3296 10201 3318
rect 9952 3265 9989 3296
rect 10165 3294 10201 3296
rect 10344 3299 10382 3340
rect 10165 3265 10202 3294
rect 9404 3256 9439 3257
rect 9381 3251 9439 3256
rect 9381 3231 9384 3251
rect 9404 3237 9439 3251
rect 9459 3237 9468 3257
rect 9404 3229 9468 3237
rect 9430 3228 9468 3229
rect 9431 3227 9468 3228
rect 9534 3261 9570 3262
rect 9642 3261 9678 3262
rect 9534 3255 9678 3261
rect 9534 3253 9600 3255
rect 9534 3233 9542 3253
rect 9562 3234 9600 3253
rect 9622 3253 9678 3255
rect 9622 3234 9650 3253
rect 9562 3233 9650 3234
rect 9670 3233 9678 3253
rect 9534 3227 9678 3233
rect 9744 3257 9782 3265
rect 9850 3261 9886 3262
rect 9744 3237 9753 3257
rect 9773 3237 9782 3257
rect 9744 3228 9782 3237
rect 9801 3254 9886 3261
rect 9801 3234 9808 3254
rect 9829 3253 9886 3254
rect 9829 3234 9858 3253
rect 9801 3233 9858 3234
rect 9878 3233 9886 3253
rect 9744 3227 9781 3228
rect 9801 3227 9886 3233
rect 9952 3257 9990 3265
rect 10063 3261 10099 3262
rect 9952 3237 9961 3257
rect 9981 3237 9990 3257
rect 9952 3228 9990 3237
rect 10014 3253 10099 3261
rect 10014 3233 10071 3253
rect 10091 3233 10099 3253
rect 9952 3227 9989 3228
rect 10014 3227 10099 3233
rect 10165 3257 10203 3265
rect 10165 3237 10174 3257
rect 10194 3237 10203 3257
rect 10165 3228 10203 3237
rect 10344 3264 10380 3299
rect 10344 3254 10381 3264
rect 10344 3236 10354 3254
rect 10372 3236 10381 3254
rect 10165 3227 10202 3228
rect 10344 3227 10381 3236
rect 9588 3206 9624 3227
rect 10014 3206 10045 3227
rect 9421 3202 9521 3206
rect 9421 3198 9483 3202
rect 9421 3172 9428 3198
rect 9454 3176 9483 3198
rect 9509 3176 9521 3202
rect 9454 3172 9521 3176
rect 9421 3169 9521 3172
rect 9589 3169 9624 3206
rect 9686 3203 10045 3206
rect 9686 3198 9908 3203
rect 9686 3174 9699 3198
rect 9723 3179 9908 3198
rect 9932 3179 10045 3203
rect 9723 3174 10045 3179
rect 9686 3170 10045 3174
rect 10112 3198 10261 3206
rect 10112 3178 10123 3198
rect 10143 3178 10261 3198
rect 10112 3171 10261 3178
rect 10112 3170 10153 3171
rect 9436 3117 9473 3118
rect 9532 3117 9569 3118
rect 9588 3117 9624 3169
rect 9643 3117 9680 3118
rect 9336 3108 9474 3117
rect 8324 3089 8492 3090
rect 8324 3086 8768 3089
rect 8324 3067 8699 3086
rect 8719 3067 8768 3086
rect 9336 3088 9445 3108
rect 9465 3088 9474 3108
rect 8324 3063 8768 3067
rect 8324 3061 8492 3063
rect 8324 2883 8351 3061
rect 8391 3023 8455 3035
rect 8731 3031 8768 3063
rect 8939 3062 9188 3084
rect 9336 3081 9474 3088
rect 9532 3108 9680 3117
rect 9532 3088 9541 3108
rect 9561 3088 9651 3108
rect 9671 3088 9680 3108
rect 9336 3079 9432 3081
rect 9532 3078 9680 3088
rect 9739 3108 9776 3118
rect 9851 3117 9888 3118
rect 9832 3115 9888 3117
rect 9739 3088 9747 3108
rect 9767 3088 9776 3108
rect 9588 3077 9624 3078
rect 8939 3031 8976 3062
rect 9152 3060 9188 3062
rect 9152 3031 9189 3060
rect 8391 3022 8426 3023
rect 8368 3017 8426 3022
rect 8368 2997 8371 3017
rect 8391 3003 8426 3017
rect 8446 3003 8455 3023
rect 8391 2995 8455 3003
rect 8417 2994 8455 2995
rect 8418 2993 8455 2994
rect 8521 3027 8557 3028
rect 8629 3027 8665 3028
rect 8521 3019 8665 3027
rect 8521 2999 8529 3019
rect 8549 2999 8581 3019
rect 8605 2999 8637 3019
rect 8657 2999 8665 3019
rect 8521 2993 8665 2999
rect 8731 3023 8769 3031
rect 8837 3027 8873 3028
rect 8731 3003 8740 3023
rect 8760 3003 8769 3023
rect 8731 2994 8769 3003
rect 8788 3020 8873 3027
rect 8788 3000 8795 3020
rect 8816 3019 8873 3020
rect 8816 3000 8845 3019
rect 8788 2999 8845 3000
rect 8865 2999 8873 3019
rect 8731 2993 8768 2994
rect 8788 2993 8873 2999
rect 8939 3023 8977 3031
rect 9050 3027 9086 3028
rect 8939 3003 8948 3023
rect 8968 3003 8977 3023
rect 8939 2994 8977 3003
rect 9001 3019 9086 3027
rect 9001 2999 9058 3019
rect 9078 2999 9086 3019
rect 8939 2993 8976 2994
rect 9001 2993 9086 2999
rect 9152 3023 9190 3031
rect 9152 3003 9161 3023
rect 9181 3003 9190 3023
rect 9436 3018 9473 3019
rect 9739 3018 9776 3088
rect 9801 3108 9888 3115
rect 9801 3105 9859 3108
rect 9801 3085 9806 3105
rect 9827 3088 9859 3105
rect 9879 3088 9888 3108
rect 9827 3085 9888 3088
rect 9801 3078 9888 3085
rect 9947 3108 9984 3118
rect 9947 3088 9955 3108
rect 9975 3088 9984 3108
rect 9801 3077 9832 3078
rect 9435 3017 9776 3018
rect 9152 2994 9190 3003
rect 9360 3012 9776 3017
rect 9152 2993 9189 2994
rect 8575 2972 8611 2993
rect 9001 2972 9032 2993
rect 9360 2992 9363 3012
rect 9383 2992 9776 3012
rect 9947 3017 9984 3088
rect 10014 3117 10045 3170
rect 10347 3155 10384 3165
rect 10347 3137 10356 3155
rect 10374 3137 10384 3155
rect 10347 3128 10384 3137
rect 10064 3117 10101 3118
rect 10014 3108 10101 3117
rect 10014 3088 10072 3108
rect 10092 3088 10101 3108
rect 10014 3078 10101 3088
rect 10160 3108 10197 3118
rect 10160 3088 10168 3108
rect 10188 3088 10197 3108
rect 10014 3077 10045 3078
rect 10160 3017 10197 3088
rect 10352 3063 10383 3128
rect 10351 3053 10388 3063
rect 10351 3051 10361 3053
rect 10285 3049 10361 3051
rect 9947 2993 10197 3017
rect 10282 3035 10361 3049
rect 10379 3035 10388 3053
rect 10282 3032 10388 3035
rect 9754 2973 9775 2992
rect 10282 2973 10308 3032
rect 10351 3026 10388 3032
rect 8408 2968 8508 2972
rect 8408 2964 8470 2968
rect 8408 2938 8415 2964
rect 8441 2942 8470 2964
rect 8496 2942 8508 2968
rect 8441 2938 8508 2942
rect 8408 2935 8508 2938
rect 8576 2935 8611 2972
rect 8673 2969 9032 2972
rect 8673 2964 8895 2969
rect 8673 2940 8686 2964
rect 8710 2945 8895 2964
rect 8919 2945 9032 2969
rect 8710 2940 9032 2945
rect 8673 2936 9032 2940
rect 9099 2964 9248 2972
rect 9099 2944 9110 2964
rect 9130 2944 9248 2964
rect 9754 2955 10308 2973
rect 10354 2962 10391 2964
rect 10282 2954 10308 2955
rect 10351 2954 10391 2962
rect 9099 2937 9248 2944
rect 10351 2942 10363 2954
rect 10342 2937 10363 2942
rect 9099 2936 9140 2937
rect 9758 2936 10363 2937
rect 10381 2936 10391 2954
rect 8423 2883 8460 2884
rect 8519 2883 8556 2884
rect 8575 2883 8611 2935
rect 8630 2883 8667 2884
rect 8323 2874 8461 2883
rect 8323 2854 8432 2874
rect 8452 2854 8461 2874
rect 8323 2847 8461 2854
rect 8519 2874 8667 2883
rect 8519 2854 8528 2874
rect 8548 2854 8638 2874
rect 8658 2854 8667 2874
rect 8323 2845 8419 2847
rect 8519 2844 8667 2854
rect 8726 2874 8763 2884
rect 8838 2883 8875 2884
rect 8819 2881 8875 2883
rect 8726 2854 8734 2874
rect 8754 2854 8763 2874
rect 8575 2843 8611 2844
rect 8423 2784 8460 2785
rect 8726 2784 8763 2854
rect 8788 2874 8875 2881
rect 8788 2871 8846 2874
rect 8788 2851 8793 2871
rect 8814 2854 8846 2871
rect 8866 2854 8875 2874
rect 8814 2851 8875 2854
rect 8788 2844 8875 2851
rect 8934 2874 8971 2884
rect 8934 2854 8942 2874
rect 8962 2854 8971 2874
rect 8788 2843 8819 2844
rect 8422 2783 8763 2784
rect 8347 2778 8763 2783
rect 8347 2758 8350 2778
rect 8370 2758 8763 2778
rect 8934 2783 8971 2854
rect 9001 2883 9032 2936
rect 9758 2927 10391 2936
rect 9758 2920 10390 2927
rect 9758 2918 9820 2920
rect 9336 2908 9504 2909
rect 9758 2908 9780 2918
rect 9051 2883 9088 2884
rect 9001 2874 9088 2883
rect 9001 2854 9059 2874
rect 9079 2854 9088 2874
rect 9001 2844 9088 2854
rect 9147 2874 9184 2884
rect 9147 2854 9155 2874
rect 9175 2854 9184 2874
rect 9001 2843 9032 2844
rect 9147 2783 9184 2854
rect 8934 2759 9184 2783
rect 9336 2882 9780 2908
rect 9336 2880 9504 2882
rect 9336 2702 9363 2880
rect 9403 2842 9467 2854
rect 9743 2850 9780 2882
rect 9951 2881 10200 2903
rect 9951 2850 9988 2881
rect 10164 2879 10200 2881
rect 10164 2850 10201 2879
rect 9403 2841 9438 2842
rect 9380 2836 9438 2841
rect 9380 2816 9383 2836
rect 9403 2822 9438 2836
rect 9458 2822 9467 2842
rect 9403 2814 9467 2822
rect 9429 2813 9467 2814
rect 9430 2812 9467 2813
rect 9533 2846 9569 2847
rect 9641 2846 9677 2847
rect 9533 2838 9677 2846
rect 9533 2818 9541 2838
rect 9561 2818 9590 2838
rect 9533 2817 9590 2818
rect 9612 2818 9649 2838
rect 9669 2818 9677 2838
rect 9612 2817 9677 2818
rect 9533 2812 9677 2817
rect 9743 2842 9781 2850
rect 9849 2846 9885 2847
rect 9743 2822 9752 2842
rect 9772 2822 9781 2842
rect 9743 2813 9781 2822
rect 9800 2839 9885 2846
rect 9800 2819 9807 2839
rect 9828 2838 9885 2839
rect 9828 2819 9857 2838
rect 9800 2818 9857 2819
rect 9877 2818 9885 2838
rect 9743 2812 9780 2813
rect 9800 2812 9885 2818
rect 9951 2842 9989 2850
rect 10062 2846 10098 2847
rect 9951 2822 9960 2842
rect 9980 2822 9989 2842
rect 9951 2813 9989 2822
rect 10013 2838 10098 2846
rect 10013 2818 10070 2838
rect 10090 2818 10098 2838
rect 9951 2812 9988 2813
rect 10013 2812 10098 2818
rect 10164 2842 10202 2850
rect 10164 2822 10173 2842
rect 10193 2822 10202 2842
rect 10164 2813 10202 2822
rect 10164 2812 10201 2813
rect 9587 2791 9623 2812
rect 10013 2791 10044 2812
rect 9420 2787 9520 2791
rect 9420 2783 9482 2787
rect 9420 2757 9427 2783
rect 9453 2761 9482 2783
rect 9508 2761 9520 2787
rect 9453 2757 9520 2761
rect 9420 2754 9520 2757
rect 9588 2754 9623 2791
rect 9685 2788 10044 2791
rect 9685 2783 9907 2788
rect 9685 2759 9698 2783
rect 9722 2764 9907 2783
rect 9931 2764 10044 2788
rect 9722 2759 10044 2764
rect 9685 2755 10044 2759
rect 10111 2783 10260 2791
rect 10111 2763 10122 2783
rect 10142 2763 10260 2783
rect 10111 2756 10260 2763
rect 10351 2771 10390 2920
rect 10111 2755 10152 2756
rect 9435 2702 9472 2703
rect 9531 2702 9568 2703
rect 9587 2702 9623 2754
rect 9642 2702 9679 2703
rect 9335 2693 9473 2702
rect 9335 2673 9444 2693
rect 9464 2673 9473 2693
rect 9335 2666 9473 2673
rect 9531 2693 9679 2702
rect 9531 2673 9540 2693
rect 9560 2673 9650 2693
rect 9670 2673 9679 2693
rect 9335 2664 9431 2666
rect 9531 2663 9679 2673
rect 9738 2693 9775 2703
rect 9850 2702 9887 2703
rect 9831 2700 9887 2702
rect 9738 2673 9746 2693
rect 9766 2673 9775 2693
rect 9587 2662 9623 2663
rect 8116 2622 8284 2623
rect 8116 2596 8560 2622
rect 8116 2594 8284 2596
rect 8116 2416 8143 2594
rect 8183 2556 8247 2568
rect 8523 2564 8560 2596
rect 8731 2595 8980 2617
rect 9435 2603 9472 2604
rect 9738 2603 9775 2673
rect 9800 2693 9887 2700
rect 9800 2690 9858 2693
rect 9800 2670 9805 2690
rect 9826 2673 9858 2690
rect 9878 2673 9887 2693
rect 9826 2670 9887 2673
rect 9800 2663 9887 2670
rect 9946 2693 9983 2703
rect 9946 2673 9954 2693
rect 9974 2673 9983 2693
rect 9800 2662 9831 2663
rect 9434 2602 9775 2603
rect 8731 2564 8768 2595
rect 8944 2593 8980 2595
rect 9359 2597 9775 2602
rect 8944 2564 8981 2593
rect 9359 2577 9362 2597
rect 9382 2577 9775 2597
rect 9946 2602 9983 2673
rect 10013 2702 10044 2755
rect 10351 2753 10361 2771
rect 10379 2753 10390 2771
rect 10351 2744 10388 2753
rect 10063 2702 10100 2703
rect 10013 2693 10100 2702
rect 10013 2673 10071 2693
rect 10091 2673 10100 2693
rect 10013 2663 10100 2673
rect 10159 2693 10196 2703
rect 10159 2673 10167 2693
rect 10187 2673 10196 2693
rect 10354 2678 10391 2682
rect 10013 2662 10044 2663
rect 10159 2602 10196 2673
rect 9946 2578 10196 2602
rect 10352 2672 10391 2678
rect 10352 2654 10363 2672
rect 10381 2654 10391 2672
rect 10352 2645 10391 2654
rect 8183 2555 8218 2556
rect 8160 2550 8218 2555
rect 8160 2530 8163 2550
rect 8183 2536 8218 2550
rect 8238 2536 8247 2556
rect 8183 2528 8247 2536
rect 8209 2527 8247 2528
rect 8210 2526 8247 2527
rect 8313 2560 8349 2561
rect 8421 2560 8457 2561
rect 8313 2554 8457 2560
rect 8313 2552 8374 2554
rect 8313 2532 8321 2552
rect 8341 2532 8374 2552
rect 8313 2528 8374 2532
rect 8399 2552 8457 2554
rect 8399 2532 8429 2552
rect 8449 2532 8457 2552
rect 8399 2528 8457 2532
rect 8313 2526 8457 2528
rect 8523 2556 8561 2564
rect 8629 2560 8665 2561
rect 8523 2536 8532 2556
rect 8552 2536 8561 2556
rect 8523 2527 8561 2536
rect 8580 2553 8665 2560
rect 8580 2533 8587 2553
rect 8608 2552 8665 2553
rect 8608 2533 8637 2552
rect 8580 2532 8637 2533
rect 8657 2532 8665 2552
rect 8523 2526 8560 2527
rect 8580 2526 8665 2532
rect 8731 2556 8769 2564
rect 8842 2560 8878 2561
rect 8731 2536 8740 2556
rect 8760 2536 8769 2556
rect 8731 2527 8769 2536
rect 8793 2552 8878 2560
rect 8793 2532 8850 2552
rect 8870 2532 8878 2552
rect 8731 2526 8768 2527
rect 8793 2526 8878 2532
rect 8944 2556 8982 2564
rect 8944 2536 8953 2556
rect 8973 2536 8982 2556
rect 8944 2527 8982 2536
rect 9738 2554 9775 2577
rect 10352 2567 10387 2645
rect 10349 2557 10387 2567
rect 9738 2553 9908 2554
rect 10349 2553 10359 2557
rect 9738 2539 10359 2553
rect 10377 2539 10387 2557
rect 9738 2533 10387 2539
rect 9738 2532 10386 2533
rect 10349 2530 10386 2532
rect 8944 2526 8981 2527
rect 8367 2505 8403 2526
rect 8793 2505 8824 2526
rect 8200 2501 8300 2505
rect 8200 2497 8262 2501
rect 8200 2471 8207 2497
rect 8233 2475 8262 2497
rect 8288 2475 8300 2501
rect 8233 2471 8300 2475
rect 8200 2468 8300 2471
rect 8368 2468 8403 2505
rect 8465 2502 8824 2505
rect 8465 2497 8687 2502
rect 8465 2473 8478 2497
rect 8502 2478 8687 2497
rect 8711 2478 8824 2502
rect 8502 2473 8824 2478
rect 8465 2469 8824 2473
rect 8891 2497 9040 2505
rect 8891 2477 8902 2497
rect 8922 2477 9040 2497
rect 8891 2470 9040 2477
rect 8891 2469 8932 2470
rect 8215 2416 8252 2417
rect 8311 2416 8348 2417
rect 8367 2416 8403 2468
rect 8422 2416 8459 2417
rect 8115 2407 8253 2416
rect 8115 2387 8224 2407
rect 8244 2387 8253 2407
rect 8115 2380 8253 2387
rect 8311 2407 8459 2416
rect 8311 2387 8320 2407
rect 8340 2387 8430 2407
rect 8450 2387 8459 2407
rect 8115 2378 8211 2380
rect 8311 2377 8459 2387
rect 8518 2407 8555 2417
rect 8630 2416 8667 2417
rect 8611 2414 8667 2416
rect 8518 2387 8526 2407
rect 8546 2387 8555 2407
rect 8367 2376 8403 2377
rect 8215 2317 8252 2318
rect 8518 2317 8555 2387
rect 8580 2407 8667 2414
rect 8580 2404 8638 2407
rect 8580 2384 8585 2404
rect 8606 2387 8638 2404
rect 8658 2387 8667 2407
rect 8606 2384 8667 2387
rect 8580 2377 8667 2384
rect 8726 2407 8763 2417
rect 8726 2387 8734 2407
rect 8754 2387 8763 2407
rect 8580 2376 8611 2377
rect 8214 2316 8555 2317
rect 8139 2311 8555 2316
rect 8139 2291 8142 2311
rect 8162 2291 8555 2311
rect 8726 2316 8763 2387
rect 8793 2416 8824 2469
rect 10352 2458 10389 2468
rect 10352 2440 10361 2458
rect 10379 2440 10389 2458
rect 10352 2431 10389 2440
rect 8843 2416 8880 2417
rect 8793 2407 8880 2416
rect 8793 2387 8851 2407
rect 8871 2387 8880 2407
rect 8793 2377 8880 2387
rect 8939 2407 8976 2417
rect 8939 2387 8947 2407
rect 8967 2387 8976 2407
rect 8793 2376 8824 2377
rect 8939 2316 8976 2387
rect 10352 2385 10387 2431
rect 10351 2379 10389 2385
rect 9762 2361 10389 2379
rect 8726 2292 8976 2316
rect 9344 2344 9512 2345
rect 9763 2344 9787 2361
rect 9344 2318 9788 2344
rect 9344 2316 9512 2318
rect 7724 2179 7757 2239
rect 7526 2172 7694 2174
rect 7250 2146 7694 2172
rect 7526 2145 7694 2146
rect 7723 2168 7760 2179
rect 7723 2149 7729 2168
rect 7752 2149 7760 2168
rect 6187 2105 6223 2106
rect 6035 2075 6044 2095
rect 6064 2075 6072 2095
rect 5923 2066 5979 2068
rect 5923 2065 5960 2066
rect 6035 2065 6072 2075
rect 6131 2095 6279 2105
rect 6379 2102 6475 2104
rect 6131 2075 6140 2095
rect 6160 2075 6250 2095
rect 6270 2075 6279 2095
rect 6131 2066 6279 2075
rect 6337 2095 6475 2102
rect 6337 2075 6346 2095
rect 6366 2075 6475 2095
rect 6337 2066 6475 2075
rect 6131 2065 6168 2066
rect 6187 2014 6223 2066
rect 6242 2065 6279 2066
rect 6338 2065 6375 2066
rect 5658 2012 5699 2013
rect 4484 1962 5116 1969
rect 4484 1960 4546 1962
rect 4062 1950 4230 1951
rect 4484 1950 4506 1960
rect 3777 1925 3814 1926
rect 3727 1916 3814 1925
rect 3727 1896 3785 1916
rect 3805 1896 3814 1916
rect 3727 1886 3814 1896
rect 3873 1916 3910 1926
rect 3873 1896 3881 1916
rect 3901 1896 3910 1916
rect 3727 1885 3758 1886
rect 3873 1825 3910 1896
rect 3660 1801 3910 1825
rect 4062 1924 4506 1950
rect 4062 1922 4230 1924
rect 4062 1744 4089 1922
rect 4129 1884 4193 1896
rect 4469 1892 4506 1924
rect 4677 1923 4926 1945
rect 4677 1892 4714 1923
rect 4890 1921 4926 1923
rect 4890 1892 4927 1921
rect 4129 1883 4164 1884
rect 4106 1878 4164 1883
rect 4106 1858 4109 1878
rect 4129 1864 4164 1878
rect 4184 1864 4193 1884
rect 4129 1856 4193 1864
rect 4155 1855 4193 1856
rect 4156 1854 4193 1855
rect 4259 1888 4295 1889
rect 4367 1888 4403 1889
rect 4259 1880 4403 1888
rect 4259 1860 4267 1880
rect 4287 1860 4316 1880
rect 4259 1859 4316 1860
rect 4338 1860 4375 1880
rect 4395 1860 4403 1880
rect 4338 1859 4403 1860
rect 4259 1854 4403 1859
rect 4469 1884 4507 1892
rect 4575 1888 4611 1889
rect 4469 1864 4478 1884
rect 4498 1864 4507 1884
rect 4469 1855 4507 1864
rect 4526 1881 4611 1888
rect 4526 1861 4533 1881
rect 4554 1880 4611 1881
rect 4554 1861 4583 1880
rect 4526 1860 4583 1861
rect 4603 1860 4611 1880
rect 4469 1854 4506 1855
rect 4526 1854 4611 1860
rect 4677 1884 4715 1892
rect 4788 1888 4824 1889
rect 4677 1864 4686 1884
rect 4706 1864 4715 1884
rect 4677 1855 4715 1864
rect 4739 1880 4824 1888
rect 4739 1860 4796 1880
rect 4816 1860 4824 1880
rect 4677 1854 4714 1855
rect 4739 1854 4824 1860
rect 4890 1884 4928 1892
rect 4890 1864 4899 1884
rect 4919 1864 4928 1884
rect 4890 1855 4928 1864
rect 4890 1854 4927 1855
rect 4313 1833 4349 1854
rect 4739 1833 4770 1854
rect 4146 1829 4246 1833
rect 4146 1825 4208 1829
rect 4146 1799 4153 1825
rect 4179 1803 4208 1825
rect 4234 1803 4246 1829
rect 4179 1799 4246 1803
rect 4146 1796 4246 1799
rect 4314 1796 4349 1833
rect 4411 1830 4770 1833
rect 4411 1825 4633 1830
rect 4411 1801 4424 1825
rect 4448 1806 4633 1825
rect 4657 1806 4770 1830
rect 4448 1801 4770 1806
rect 4411 1797 4770 1801
rect 4837 1825 4986 1833
rect 4837 1805 4848 1825
rect 4868 1805 4986 1825
rect 4837 1798 4986 1805
rect 5077 1813 5116 1962
rect 5420 1848 5459 1997
rect 5550 2005 5699 2012
rect 5550 1985 5668 2005
rect 5688 1985 5699 2005
rect 5550 1977 5699 1985
rect 5766 2009 6125 2013
rect 5766 2004 6088 2009
rect 5766 1980 5879 2004
rect 5903 1985 6088 2004
rect 6112 1985 6125 2009
rect 5903 1980 6125 1985
rect 5766 1977 6125 1980
rect 6187 1977 6222 2014
rect 6290 2011 6390 2014
rect 6290 2007 6357 2011
rect 6290 1981 6302 2007
rect 6328 1985 6357 2007
rect 6383 1985 6390 2011
rect 6328 1981 6390 1985
rect 6290 1977 6390 1981
rect 5766 1956 5797 1977
rect 6187 1956 6223 1977
rect 5609 1955 5646 1956
rect 5608 1946 5646 1955
rect 5608 1926 5617 1946
rect 5637 1926 5646 1946
rect 5608 1918 5646 1926
rect 5712 1950 5797 1956
rect 5822 1955 5859 1956
rect 5712 1930 5720 1950
rect 5740 1930 5797 1950
rect 5712 1922 5797 1930
rect 5821 1946 5859 1955
rect 5821 1926 5830 1946
rect 5850 1926 5859 1946
rect 5712 1921 5748 1922
rect 5821 1918 5859 1926
rect 5925 1950 6010 1956
rect 6030 1955 6067 1956
rect 5925 1930 5933 1950
rect 5953 1949 6010 1950
rect 5953 1930 5982 1949
rect 5925 1929 5982 1930
rect 6003 1929 6010 1949
rect 5925 1922 6010 1929
rect 6029 1946 6067 1955
rect 6029 1926 6038 1946
rect 6058 1926 6067 1946
rect 5925 1921 5961 1922
rect 6029 1918 6067 1926
rect 6133 1951 6277 1956
rect 6133 1950 6198 1951
rect 6133 1930 6141 1950
rect 6161 1930 6198 1950
rect 6220 1950 6277 1951
rect 6220 1930 6249 1950
rect 6269 1930 6277 1950
rect 6133 1922 6277 1930
rect 6133 1921 6169 1922
rect 6241 1921 6277 1922
rect 6343 1955 6380 1956
rect 6343 1954 6381 1955
rect 6343 1946 6407 1954
rect 6343 1926 6352 1946
rect 6372 1932 6407 1946
rect 6427 1932 6430 1952
rect 6372 1927 6430 1932
rect 6372 1926 6407 1927
rect 5609 1889 5646 1918
rect 5610 1887 5646 1889
rect 5822 1887 5859 1918
rect 5610 1865 5859 1887
rect 6030 1886 6067 1918
rect 6343 1914 6407 1926
rect 6447 1888 6474 2066
rect 6306 1886 6474 1888
rect 6030 1860 6474 1886
rect 6626 1985 6876 2009
rect 6626 1914 6663 1985
rect 6778 1924 6809 1925
rect 6626 1894 6635 1914
rect 6655 1894 6663 1914
rect 6626 1884 6663 1894
rect 6722 1914 6809 1924
rect 6722 1894 6731 1914
rect 6751 1894 6809 1914
rect 6722 1885 6809 1894
rect 6722 1884 6759 1885
rect 6030 1850 6052 1860
rect 6306 1859 6474 1860
rect 5990 1848 6052 1850
rect 5420 1841 6052 1848
rect 4837 1797 4878 1798
rect 4161 1744 4198 1745
rect 4257 1744 4294 1745
rect 4313 1744 4349 1796
rect 4368 1744 4405 1745
rect 4061 1735 4199 1744
rect 4061 1715 4170 1735
rect 4190 1715 4199 1735
rect 2998 1711 3168 1712
rect 2998 1696 3444 1711
rect 4061 1708 4199 1715
rect 4257 1735 4405 1744
rect 4257 1715 4266 1735
rect 4286 1715 4376 1735
rect 4396 1715 4405 1735
rect 4061 1706 4157 1708
rect 3000 1685 3444 1696
rect 3000 1683 3168 1685
rect 3000 1505 3027 1683
rect 3067 1645 3131 1657
rect 3407 1653 3444 1685
rect 3615 1684 3864 1706
rect 4257 1705 4405 1715
rect 4464 1735 4501 1745
rect 4576 1744 4613 1745
rect 4557 1742 4613 1744
rect 4464 1715 4472 1735
rect 4492 1715 4501 1735
rect 4313 1704 4349 1705
rect 3615 1653 3652 1684
rect 3828 1682 3864 1684
rect 3828 1653 3865 1682
rect 3067 1644 3102 1645
rect 3044 1639 3102 1644
rect 3044 1619 3047 1639
rect 3067 1625 3102 1639
rect 3122 1625 3131 1645
rect 3067 1617 3131 1625
rect 3093 1616 3131 1617
rect 3094 1615 3131 1616
rect 3197 1649 3233 1650
rect 3305 1649 3341 1650
rect 3197 1641 3341 1649
rect 3197 1621 3205 1641
rect 3225 1640 3313 1641
rect 3225 1623 3253 1640
rect 3277 1623 3313 1640
rect 3225 1621 3313 1623
rect 3333 1621 3341 1641
rect 3197 1615 3341 1621
rect 3407 1645 3445 1653
rect 3513 1649 3549 1650
rect 3407 1625 3416 1645
rect 3436 1625 3445 1645
rect 3407 1616 3445 1625
rect 3464 1642 3549 1649
rect 3464 1622 3471 1642
rect 3492 1641 3549 1642
rect 3492 1622 3521 1641
rect 3464 1621 3521 1622
rect 3541 1621 3549 1641
rect 3407 1615 3444 1616
rect 3464 1615 3549 1621
rect 3615 1645 3653 1653
rect 3726 1649 3762 1650
rect 3615 1625 3624 1645
rect 3644 1625 3653 1645
rect 3615 1616 3653 1625
rect 3677 1641 3762 1649
rect 3677 1621 3734 1641
rect 3754 1621 3762 1641
rect 3615 1615 3652 1616
rect 3677 1615 3762 1621
rect 3828 1645 3866 1653
rect 4161 1645 4198 1646
rect 4464 1645 4501 1715
rect 4526 1735 4613 1742
rect 4526 1732 4584 1735
rect 4526 1712 4531 1732
rect 4552 1715 4584 1732
rect 4604 1715 4613 1735
rect 4552 1712 4613 1715
rect 4526 1705 4613 1712
rect 4672 1735 4709 1745
rect 4672 1715 4680 1735
rect 4700 1715 4709 1735
rect 4526 1704 4557 1705
rect 3828 1625 3837 1645
rect 3857 1625 3866 1645
rect 4160 1644 4501 1645
rect 3828 1616 3866 1625
rect 4085 1639 4501 1644
rect 4085 1619 4088 1639
rect 4108 1619 4501 1639
rect 4672 1644 4709 1715
rect 4739 1744 4770 1797
rect 5077 1795 5087 1813
rect 5105 1795 5116 1813
rect 5419 1832 6052 1841
rect 6778 1832 6809 1885
rect 6839 1914 6876 1985
rect 7047 1990 7440 2010
rect 7460 1990 7463 2010
rect 7047 1985 7463 1990
rect 7047 1984 7388 1985
rect 6991 1924 7022 1925
rect 6839 1894 6848 1914
rect 6868 1894 6876 1914
rect 6839 1884 6876 1894
rect 6935 1917 7022 1924
rect 6935 1914 6996 1917
rect 6935 1894 6944 1914
rect 6964 1897 6996 1914
rect 7017 1897 7022 1917
rect 6964 1894 7022 1897
rect 6935 1887 7022 1894
rect 7047 1914 7084 1984
rect 7350 1983 7387 1984
rect 7199 1924 7235 1925
rect 7047 1894 7056 1914
rect 7076 1894 7084 1914
rect 6935 1885 6991 1887
rect 6935 1884 6972 1885
rect 7047 1884 7084 1894
rect 7143 1914 7291 1924
rect 7391 1921 7487 1923
rect 7143 1894 7152 1914
rect 7172 1894 7262 1914
rect 7282 1894 7291 1914
rect 7143 1885 7291 1894
rect 7349 1914 7487 1921
rect 7349 1894 7358 1914
rect 7378 1894 7487 1914
rect 7349 1885 7487 1894
rect 7143 1884 7180 1885
rect 7199 1833 7235 1885
rect 7254 1884 7291 1885
rect 7350 1884 7387 1885
rect 5419 1814 5429 1832
rect 5447 1831 6052 1832
rect 6670 1831 6711 1832
rect 5447 1826 5468 1831
rect 5447 1814 5459 1826
rect 6562 1824 6711 1831
rect 5419 1806 5459 1814
rect 5502 1813 5528 1814
rect 5419 1804 5456 1806
rect 5502 1795 6056 1813
rect 6562 1804 6680 1824
rect 6700 1804 6711 1824
rect 6562 1796 6711 1804
rect 6778 1828 7137 1832
rect 6778 1823 7100 1828
rect 6778 1799 6891 1823
rect 6915 1804 7100 1823
rect 7124 1804 7137 1828
rect 6915 1799 7137 1804
rect 6778 1796 7137 1799
rect 7199 1796 7234 1833
rect 7302 1830 7402 1833
rect 7302 1826 7369 1830
rect 7302 1800 7314 1826
rect 7340 1804 7369 1826
rect 7395 1804 7402 1830
rect 7340 1800 7402 1804
rect 7302 1796 7402 1800
rect 5077 1786 5114 1795
rect 4789 1744 4826 1745
rect 4739 1735 4826 1744
rect 4739 1715 4797 1735
rect 4817 1715 4826 1735
rect 4739 1705 4826 1715
rect 4885 1735 4922 1745
rect 4885 1715 4893 1735
rect 4913 1715 4922 1735
rect 5422 1736 5459 1742
rect 5502 1736 5528 1795
rect 6035 1776 6056 1795
rect 5422 1733 5528 1736
rect 5080 1720 5117 1724
rect 4739 1704 4770 1705
rect 4885 1644 4922 1715
rect 4672 1620 4922 1644
rect 5078 1714 5117 1720
rect 5078 1696 5089 1714
rect 5107 1696 5117 1714
rect 5422 1715 5431 1733
rect 5449 1719 5528 1733
rect 5613 1751 5863 1775
rect 5449 1717 5525 1719
rect 5449 1715 5459 1717
rect 5422 1705 5459 1715
rect 5078 1687 5117 1696
rect 3828 1615 3865 1616
rect 3251 1594 3287 1615
rect 3677 1594 3708 1615
rect 4464 1596 4501 1619
rect 5078 1609 5113 1687
rect 5427 1640 5458 1705
rect 5613 1680 5650 1751
rect 5765 1690 5796 1691
rect 5613 1660 5622 1680
rect 5642 1660 5650 1680
rect 5613 1650 5650 1660
rect 5709 1680 5796 1690
rect 5709 1660 5718 1680
rect 5738 1660 5796 1680
rect 5709 1651 5796 1660
rect 5709 1650 5746 1651
rect 5075 1599 5113 1609
rect 5426 1631 5463 1640
rect 5426 1613 5436 1631
rect 5454 1613 5463 1631
rect 5426 1603 5463 1613
rect 4464 1595 4634 1596
rect 5075 1595 5085 1599
rect 3084 1590 3184 1594
rect 3084 1586 3146 1590
rect 3084 1560 3091 1586
rect 3117 1564 3146 1586
rect 3172 1564 3184 1590
rect 3117 1560 3184 1564
rect 3084 1557 3184 1560
rect 3252 1557 3287 1594
rect 3349 1591 3708 1594
rect 3349 1586 3571 1591
rect 3349 1562 3362 1586
rect 3386 1567 3571 1586
rect 3595 1567 3708 1591
rect 3386 1562 3708 1567
rect 3349 1558 3708 1562
rect 3775 1586 3924 1594
rect 3775 1566 3786 1586
rect 3806 1566 3924 1586
rect 4464 1581 5085 1595
rect 5103 1581 5113 1599
rect 5765 1598 5796 1651
rect 5826 1680 5863 1751
rect 6034 1756 6427 1776
rect 6447 1756 6450 1776
rect 6778 1775 6809 1796
rect 7199 1775 7235 1796
rect 6621 1774 6658 1775
rect 6034 1751 6450 1756
rect 6620 1765 6658 1774
rect 6034 1750 6375 1751
rect 5978 1690 6009 1691
rect 5826 1660 5835 1680
rect 5855 1660 5863 1680
rect 5826 1650 5863 1660
rect 5922 1683 6009 1690
rect 5922 1680 5983 1683
rect 5922 1660 5931 1680
rect 5951 1663 5983 1680
rect 6004 1663 6009 1683
rect 5951 1660 6009 1663
rect 5922 1653 6009 1660
rect 6034 1680 6071 1750
rect 6337 1749 6374 1750
rect 6620 1745 6629 1765
rect 6649 1745 6658 1765
rect 6620 1737 6658 1745
rect 6724 1769 6809 1775
rect 6834 1774 6871 1775
rect 6724 1749 6732 1769
rect 6752 1749 6809 1769
rect 6724 1741 6809 1749
rect 6833 1765 6871 1774
rect 6833 1745 6842 1765
rect 6862 1745 6871 1765
rect 6724 1740 6760 1741
rect 6833 1737 6871 1745
rect 6937 1769 7022 1775
rect 7042 1774 7079 1775
rect 6937 1749 6945 1769
rect 6965 1768 7022 1769
rect 6965 1749 6994 1768
rect 6937 1748 6994 1749
rect 7015 1748 7022 1768
rect 6937 1741 7022 1748
rect 7041 1765 7079 1774
rect 7041 1745 7050 1765
rect 7070 1745 7079 1765
rect 6937 1740 6973 1741
rect 7041 1737 7079 1745
rect 7145 1769 7289 1775
rect 7145 1749 7153 1769
rect 7173 1749 7205 1769
rect 7229 1749 7261 1769
rect 7281 1749 7289 1769
rect 7145 1741 7289 1749
rect 7145 1740 7181 1741
rect 7253 1740 7289 1741
rect 7355 1774 7392 1775
rect 7355 1773 7393 1774
rect 7355 1765 7419 1773
rect 7355 1745 7364 1765
rect 7384 1751 7419 1765
rect 7439 1751 7442 1771
rect 7384 1746 7442 1751
rect 7384 1745 7419 1746
rect 6621 1708 6658 1737
rect 6622 1706 6658 1708
rect 6834 1706 6871 1737
rect 6186 1690 6222 1691
rect 6034 1660 6043 1680
rect 6063 1660 6071 1680
rect 5922 1651 5978 1653
rect 5922 1650 5959 1651
rect 6034 1650 6071 1660
rect 6130 1680 6278 1690
rect 6378 1687 6474 1689
rect 6130 1660 6139 1680
rect 6159 1660 6249 1680
rect 6269 1660 6278 1680
rect 6130 1651 6278 1660
rect 6336 1680 6474 1687
rect 6622 1684 6871 1706
rect 7042 1705 7079 1737
rect 7355 1733 7419 1745
rect 7459 1707 7486 1885
rect 7318 1705 7486 1707
rect 7042 1701 7486 1705
rect 6336 1660 6345 1680
rect 6365 1660 6474 1680
rect 7042 1682 7091 1701
rect 7111 1682 7486 1701
rect 7042 1679 7486 1682
rect 7318 1678 7486 1679
rect 6336 1651 6474 1660
rect 6130 1650 6167 1651
rect 6186 1599 6222 1651
rect 6241 1650 6278 1651
rect 6337 1650 6374 1651
rect 5657 1597 5698 1598
rect 4464 1575 5113 1581
rect 5549 1590 5698 1597
rect 4464 1574 5112 1575
rect 5075 1572 5112 1574
rect 3775 1559 3924 1566
rect 5549 1570 5667 1590
rect 5687 1570 5698 1590
rect 5549 1562 5698 1570
rect 5765 1594 6124 1598
rect 5765 1589 6087 1594
rect 5765 1565 5878 1589
rect 5902 1570 6087 1589
rect 6111 1570 6124 1594
rect 5902 1565 6124 1570
rect 5765 1562 6124 1565
rect 6186 1562 6221 1599
rect 6289 1596 6389 1599
rect 6289 1592 6356 1596
rect 6289 1566 6301 1592
rect 6327 1570 6356 1592
rect 6382 1570 6389 1596
rect 6327 1566 6389 1570
rect 6289 1562 6389 1566
rect 3775 1558 3816 1559
rect 3099 1505 3136 1506
rect 3195 1505 3232 1506
rect 3251 1505 3287 1557
rect 3306 1505 3343 1506
rect 2999 1496 3137 1505
rect 2999 1476 3108 1496
rect 3128 1476 3137 1496
rect 2999 1469 3137 1476
rect 3195 1496 3343 1505
rect 3195 1476 3204 1496
rect 3224 1476 3314 1496
rect 3334 1476 3343 1496
rect 2999 1467 3095 1469
rect 3195 1466 3343 1476
rect 3402 1496 3439 1506
rect 3514 1505 3551 1506
rect 3495 1503 3551 1505
rect 3402 1476 3410 1496
rect 3430 1476 3439 1496
rect 3251 1465 3287 1466
rect 3099 1406 3136 1407
rect 3402 1406 3439 1476
rect 3464 1496 3551 1503
rect 3464 1493 3522 1496
rect 3464 1473 3469 1493
rect 3490 1476 3522 1493
rect 3542 1476 3551 1496
rect 3490 1473 3551 1476
rect 3464 1466 3551 1473
rect 3610 1496 3647 1506
rect 3610 1476 3618 1496
rect 3638 1476 3647 1496
rect 3464 1465 3495 1466
rect 3098 1405 3439 1406
rect 3023 1400 3439 1405
rect 3023 1380 3026 1400
rect 3046 1380 3439 1400
rect 3610 1405 3647 1476
rect 3677 1505 3708 1558
rect 5765 1541 5796 1562
rect 6186 1541 6222 1562
rect 5429 1532 5466 1541
rect 5608 1540 5645 1541
rect 5429 1514 5438 1532
rect 5456 1514 5466 1532
rect 3727 1505 3764 1506
rect 3677 1496 3764 1505
rect 3677 1476 3735 1496
rect 3755 1476 3764 1496
rect 3677 1466 3764 1476
rect 3823 1496 3860 1506
rect 3823 1476 3831 1496
rect 3851 1476 3860 1496
rect 3677 1465 3708 1466
rect 3823 1405 3860 1476
rect 5078 1500 5115 1510
rect 5429 1504 5466 1514
rect 5078 1482 5087 1500
rect 5105 1482 5115 1500
rect 5078 1473 5115 1482
rect 5078 1449 5113 1473
rect 5430 1469 5466 1504
rect 5607 1531 5645 1540
rect 5607 1511 5616 1531
rect 5636 1511 5645 1531
rect 5607 1503 5645 1511
rect 5711 1535 5796 1541
rect 5821 1540 5858 1541
rect 5711 1515 5719 1535
rect 5739 1515 5796 1535
rect 5711 1507 5796 1515
rect 5820 1531 5858 1540
rect 5820 1511 5829 1531
rect 5849 1511 5858 1531
rect 5711 1506 5747 1507
rect 5820 1503 5858 1511
rect 5924 1535 6009 1541
rect 6029 1540 6066 1541
rect 5924 1515 5932 1535
rect 5952 1534 6009 1535
rect 5952 1515 5981 1534
rect 5924 1514 5981 1515
rect 6002 1514 6009 1534
rect 5924 1507 6009 1514
rect 6028 1531 6066 1540
rect 6028 1511 6037 1531
rect 6057 1511 6066 1531
rect 5924 1506 5960 1507
rect 6028 1503 6066 1511
rect 6132 1535 6276 1541
rect 6132 1515 6140 1535
rect 6160 1534 6248 1535
rect 6160 1515 6188 1534
rect 6132 1513 6188 1515
rect 6210 1515 6248 1534
rect 6268 1515 6276 1535
rect 6210 1513 6276 1515
rect 6132 1507 6276 1513
rect 6132 1506 6168 1507
rect 6240 1506 6276 1507
rect 6342 1540 6379 1541
rect 6342 1539 6380 1540
rect 6342 1531 6406 1539
rect 6342 1511 6351 1531
rect 6371 1517 6406 1531
rect 6426 1517 6429 1537
rect 6371 1512 6429 1517
rect 6371 1511 6406 1512
rect 5608 1474 5645 1503
rect 5076 1425 5113 1449
rect 5075 1419 5113 1425
rect 3610 1381 3860 1405
rect 4486 1401 5113 1419
rect 4068 1384 4236 1385
rect 4487 1384 4511 1401
rect 4068 1358 4512 1384
rect 4068 1356 4236 1358
rect 4068 1178 4095 1356
rect 4135 1318 4199 1330
rect 4475 1326 4512 1358
rect 4683 1357 4932 1379
rect 4683 1326 4720 1357
rect 4896 1355 4932 1357
rect 5075 1360 5113 1401
rect 5428 1428 5466 1469
rect 5609 1472 5645 1474
rect 5821 1472 5858 1503
rect 5609 1450 5858 1472
rect 6029 1471 6066 1503
rect 6342 1499 6406 1511
rect 6446 1473 6473 1651
rect 6305 1471 6473 1473
rect 6029 1445 6473 1471
rect 6030 1428 6054 1445
rect 6305 1444 6473 1445
rect 5428 1410 6055 1428
rect 6681 1424 6931 1448
rect 5428 1404 5466 1410
rect 5428 1380 5465 1404
rect 4896 1326 4933 1355
rect 4135 1317 4170 1318
rect 4112 1312 4170 1317
rect 4112 1292 4115 1312
rect 4135 1298 4170 1312
rect 4190 1298 4199 1318
rect 4135 1290 4199 1298
rect 4161 1289 4199 1290
rect 4162 1288 4199 1289
rect 4265 1322 4301 1323
rect 4373 1322 4409 1323
rect 4265 1316 4409 1322
rect 4265 1314 4331 1316
rect 4265 1294 4273 1314
rect 4293 1295 4331 1314
rect 4353 1314 4409 1316
rect 4353 1295 4381 1314
rect 4293 1294 4381 1295
rect 4401 1294 4409 1314
rect 4265 1288 4409 1294
rect 4475 1318 4513 1326
rect 4581 1322 4617 1323
rect 4475 1298 4484 1318
rect 4504 1298 4513 1318
rect 4475 1289 4513 1298
rect 4532 1315 4617 1322
rect 4532 1295 4539 1315
rect 4560 1314 4617 1315
rect 4560 1295 4589 1314
rect 4532 1294 4589 1295
rect 4609 1294 4617 1314
rect 4475 1288 4512 1289
rect 4532 1288 4617 1294
rect 4683 1318 4721 1326
rect 4794 1322 4830 1323
rect 4683 1298 4692 1318
rect 4712 1298 4721 1318
rect 4683 1289 4721 1298
rect 4745 1314 4830 1322
rect 4745 1294 4802 1314
rect 4822 1294 4830 1314
rect 4683 1288 4720 1289
rect 4745 1288 4830 1294
rect 4896 1318 4934 1326
rect 4896 1298 4905 1318
rect 4925 1298 4934 1318
rect 4896 1289 4934 1298
rect 5075 1325 5111 1360
rect 5428 1356 5463 1380
rect 5426 1347 5463 1356
rect 5426 1329 5436 1347
rect 5454 1329 5463 1347
rect 5075 1315 5112 1325
rect 5426 1319 5463 1329
rect 6681 1353 6718 1424
rect 6833 1363 6864 1364
rect 6681 1333 6690 1353
rect 6710 1333 6718 1353
rect 6681 1323 6718 1333
rect 6777 1353 6864 1363
rect 6777 1333 6786 1353
rect 6806 1333 6864 1353
rect 6777 1324 6864 1333
rect 6777 1323 6814 1324
rect 5075 1297 5085 1315
rect 5103 1297 5112 1315
rect 4896 1288 4933 1289
rect 5075 1288 5112 1297
rect 4319 1267 4355 1288
rect 4745 1267 4776 1288
rect 6833 1271 6864 1324
rect 6894 1353 6931 1424
rect 7102 1429 7495 1449
rect 7515 1429 7518 1449
rect 7102 1424 7518 1429
rect 7102 1423 7443 1424
rect 7046 1363 7077 1364
rect 6894 1333 6903 1353
rect 6923 1333 6931 1353
rect 6894 1323 6931 1333
rect 6990 1356 7077 1363
rect 6990 1353 7051 1356
rect 6990 1333 6999 1353
rect 7019 1336 7051 1353
rect 7072 1336 7077 1356
rect 7019 1333 7077 1336
rect 6990 1326 7077 1333
rect 7102 1353 7139 1423
rect 7405 1422 7442 1423
rect 7254 1363 7290 1364
rect 7102 1333 7111 1353
rect 7131 1333 7139 1353
rect 6990 1324 7046 1326
rect 6990 1323 7027 1324
rect 7102 1323 7139 1333
rect 7198 1353 7346 1363
rect 7446 1360 7542 1362
rect 7198 1333 7207 1353
rect 7227 1333 7317 1353
rect 7337 1333 7346 1353
rect 7198 1324 7346 1333
rect 7404 1353 7542 1360
rect 7404 1333 7413 1353
rect 7433 1333 7542 1353
rect 7404 1324 7542 1333
rect 7198 1323 7235 1324
rect 7254 1272 7290 1324
rect 7309 1323 7346 1324
rect 7405 1323 7442 1324
rect 6725 1270 6766 1271
rect 4152 1263 4252 1267
rect 4152 1259 4214 1263
rect 4152 1233 4159 1259
rect 4185 1237 4214 1259
rect 4240 1237 4252 1263
rect 4185 1233 4252 1237
rect 4152 1230 4252 1233
rect 4320 1230 4355 1267
rect 4417 1264 4776 1267
rect 4417 1259 4639 1264
rect 4417 1235 4430 1259
rect 4454 1240 4639 1259
rect 4663 1240 4776 1264
rect 4454 1235 4776 1240
rect 4417 1231 4776 1235
rect 4843 1259 4992 1267
rect 4843 1239 4854 1259
rect 4874 1239 4992 1259
rect 6617 1263 6766 1270
rect 5429 1255 5466 1257
rect 5429 1254 6077 1255
rect 4843 1232 4992 1239
rect 5428 1248 6077 1254
rect 4843 1231 4884 1232
rect 4167 1178 4204 1179
rect 4263 1178 4300 1179
rect 4319 1178 4355 1230
rect 4374 1178 4411 1179
rect 4067 1169 4205 1178
rect 2323 1160 2355 1165
rect 1103 1142 1199 1144
rect 855 1115 864 1135
rect 884 1115 974 1135
rect 994 1115 1003 1135
rect 855 1106 1003 1115
rect 1061 1135 1199 1142
rect 1816 1139 2262 1154
rect 2092 1138 2262 1139
rect 1061 1115 1070 1135
rect 1090 1115 1199 1135
rect 1061 1106 1199 1115
rect 855 1105 892 1106
rect 911 1054 947 1106
rect 966 1105 1003 1106
rect 1062 1105 1099 1106
rect 382 1052 423 1053
rect 144 888 183 1037
rect 274 1045 423 1052
rect 274 1025 392 1045
rect 412 1025 423 1045
rect 274 1017 423 1025
rect 490 1049 849 1053
rect 490 1044 812 1049
rect 490 1020 603 1044
rect 627 1025 812 1044
rect 836 1025 849 1049
rect 627 1020 849 1025
rect 490 1017 849 1020
rect 911 1017 946 1054
rect 1014 1051 1114 1054
rect 1014 1047 1081 1051
rect 1014 1021 1026 1047
rect 1052 1025 1081 1047
rect 1107 1025 1114 1051
rect 1052 1021 1114 1025
rect 1014 1017 1114 1021
rect 490 996 521 1017
rect 911 996 947 1017
rect 333 995 370 996
rect 332 986 370 995
rect 332 966 341 986
rect 361 966 370 986
rect 332 958 370 966
rect 436 990 521 996
rect 546 995 583 996
rect 436 970 444 990
rect 464 970 521 990
rect 436 962 521 970
rect 545 986 583 995
rect 545 966 554 986
rect 574 966 583 986
rect 436 961 472 962
rect 545 958 583 966
rect 649 990 734 996
rect 754 995 791 996
rect 649 970 657 990
rect 677 989 734 990
rect 677 970 706 989
rect 649 969 706 970
rect 727 969 734 989
rect 649 962 734 969
rect 753 986 791 995
rect 753 966 762 986
rect 782 966 791 986
rect 649 961 685 962
rect 753 958 791 966
rect 857 991 1001 996
rect 857 990 922 991
rect 857 970 865 990
rect 885 970 922 990
rect 944 990 1001 991
rect 944 970 973 990
rect 993 970 1001 990
rect 857 962 1001 970
rect 857 961 893 962
rect 965 961 1001 962
rect 1067 995 1104 996
rect 1067 994 1105 995
rect 1067 986 1131 994
rect 1067 966 1076 986
rect 1096 972 1131 986
rect 1151 972 1154 992
rect 1096 967 1154 972
rect 1096 966 1131 967
rect 333 929 370 958
rect 334 927 370 929
rect 546 927 583 958
rect 334 905 583 927
rect 754 926 791 958
rect 1067 954 1131 966
rect 1171 928 1198 1106
rect 1030 926 1198 928
rect 754 900 1198 926
rect 1350 1025 1600 1049
rect 1350 954 1387 1025
rect 1502 964 1533 965
rect 1350 934 1359 954
rect 1379 934 1387 954
rect 1350 924 1387 934
rect 1446 954 1533 964
rect 1446 934 1455 954
rect 1475 934 1533 954
rect 1446 925 1533 934
rect 1446 924 1483 925
rect 754 890 776 900
rect 1030 899 1198 900
rect 714 888 776 890
rect 144 881 776 888
rect 143 872 776 881
rect 1502 872 1533 925
rect 1563 954 1600 1025
rect 1771 1030 2164 1050
rect 2184 1030 2187 1050
rect 1771 1025 2187 1030
rect 1771 1024 2112 1025
rect 1715 964 1746 965
rect 1563 934 1572 954
rect 1592 934 1600 954
rect 1563 924 1600 934
rect 1659 957 1746 964
rect 1659 954 1720 957
rect 1659 934 1668 954
rect 1688 937 1720 954
rect 1741 937 1746 957
rect 1688 934 1746 937
rect 1659 927 1746 934
rect 1771 954 1808 1024
rect 2074 1023 2111 1024
rect 1923 964 1959 965
rect 1771 934 1780 954
rect 1800 934 1808 954
rect 1659 925 1715 927
rect 1659 924 1696 925
rect 1771 924 1808 934
rect 1867 954 2015 964
rect 2115 961 2211 963
rect 1867 934 1876 954
rect 1896 934 1986 954
rect 2006 934 2015 954
rect 1867 925 2015 934
rect 2073 954 2211 961
rect 2073 934 2082 954
rect 2102 934 2211 954
rect 2073 925 2211 934
rect 1867 924 1904 925
rect 1923 873 1959 925
rect 1978 924 2015 925
rect 2074 924 2111 925
rect 143 854 153 872
rect 171 871 776 872
rect 1394 871 1435 872
rect 171 866 192 871
rect 171 854 183 866
rect 1286 864 1435 871
rect 143 846 183 854
rect 226 853 252 854
rect 143 844 180 846
rect 226 835 780 853
rect 1286 844 1404 864
rect 1424 844 1435 864
rect 1286 836 1435 844
rect 1502 868 1861 872
rect 1502 863 1824 868
rect 1502 839 1615 863
rect 1639 844 1824 863
rect 1848 844 1861 868
rect 1639 839 1861 844
rect 1502 836 1861 839
rect 1923 836 1958 873
rect 2026 870 2126 873
rect 2026 866 2093 870
rect 2026 840 2038 866
rect 2064 844 2093 866
rect 2119 844 2126 870
rect 2064 840 2126 844
rect 2026 836 2126 840
rect 146 776 183 782
rect 226 776 252 835
rect 759 816 780 835
rect 146 773 252 776
rect 146 755 155 773
rect 173 759 252 773
rect 337 791 587 815
rect 173 757 249 759
rect 173 755 183 757
rect 146 745 183 755
rect 151 680 182 745
rect 337 720 374 791
rect 489 730 520 731
rect 337 700 346 720
rect 366 700 374 720
rect 337 690 374 700
rect 433 720 520 730
rect 433 700 442 720
rect 462 700 520 720
rect 433 691 520 700
rect 433 690 470 691
rect 150 671 187 680
rect 150 653 160 671
rect 178 653 187 671
rect 150 643 187 653
rect 489 638 520 691
rect 550 720 587 791
rect 758 796 1151 816
rect 1171 796 1174 816
rect 1502 815 1533 836
rect 1923 815 1959 836
rect 1345 814 1382 815
rect 758 791 1174 796
rect 1344 805 1382 814
rect 758 790 1099 791
rect 702 730 733 731
rect 550 700 559 720
rect 579 700 587 720
rect 550 690 587 700
rect 646 723 733 730
rect 646 720 707 723
rect 646 700 655 720
rect 675 703 707 720
rect 728 703 733 723
rect 675 700 733 703
rect 646 693 733 700
rect 758 720 795 790
rect 1061 789 1098 790
rect 1344 785 1353 805
rect 1373 785 1382 805
rect 1344 777 1382 785
rect 1448 809 1533 815
rect 1558 814 1595 815
rect 1448 789 1456 809
rect 1476 789 1533 809
rect 1448 781 1533 789
rect 1557 805 1595 814
rect 1557 785 1566 805
rect 1586 785 1595 805
rect 1448 780 1484 781
rect 1557 777 1595 785
rect 1661 809 1746 815
rect 1766 814 1803 815
rect 1661 789 1669 809
rect 1689 808 1746 809
rect 1689 789 1718 808
rect 1661 788 1718 789
rect 1739 788 1746 808
rect 1661 781 1746 788
rect 1765 805 1803 814
rect 1765 785 1774 805
rect 1794 785 1803 805
rect 1661 780 1697 781
rect 1765 777 1803 785
rect 1869 810 2013 815
rect 1869 809 1928 810
rect 1869 789 1877 809
rect 1897 790 1928 809
rect 1952 809 2013 810
rect 1952 790 1985 809
rect 1897 789 1985 790
rect 2005 789 2013 809
rect 1869 781 2013 789
rect 1869 780 1905 781
rect 1977 780 2013 781
rect 2079 814 2116 815
rect 2079 813 2117 814
rect 2079 805 2143 813
rect 2079 785 2088 805
rect 2108 791 2143 805
rect 2163 791 2166 811
rect 2108 786 2166 791
rect 2108 785 2143 786
rect 1345 748 1382 777
rect 1346 746 1382 748
rect 1558 746 1595 777
rect 910 730 946 731
rect 758 700 767 720
rect 787 700 795 720
rect 646 691 702 693
rect 646 690 683 691
rect 758 690 795 700
rect 854 720 1002 730
rect 1102 727 1198 729
rect 854 700 863 720
rect 883 700 973 720
rect 993 700 1002 720
rect 854 691 1002 700
rect 1060 720 1198 727
rect 1346 724 1595 746
rect 1766 745 1803 777
rect 2079 773 2143 785
rect 2183 747 2210 925
rect 2042 745 2210 747
rect 1766 741 2210 745
rect 1060 700 1069 720
rect 1089 700 1198 720
rect 1766 722 1815 741
rect 1835 722 2210 741
rect 1766 719 2210 722
rect 2042 718 2210 719
rect 2231 744 2262 1138
rect 2323 1142 2328 1160
rect 2348 1142 2355 1160
rect 2323 1137 2355 1142
rect 2326 1135 2355 1137
rect 3055 1150 3223 1151
rect 3055 1147 3499 1150
rect 3055 1128 3430 1147
rect 3450 1128 3499 1147
rect 4067 1149 4176 1169
rect 4196 1149 4205 1169
rect 3055 1124 3499 1128
rect 3055 1122 3223 1124
rect 3055 944 3082 1122
rect 3122 1084 3186 1096
rect 3462 1092 3499 1124
rect 3670 1123 3919 1145
rect 4067 1142 4205 1149
rect 4263 1169 4411 1178
rect 4263 1149 4272 1169
rect 4292 1149 4382 1169
rect 4402 1149 4411 1169
rect 4067 1140 4163 1142
rect 4263 1139 4411 1149
rect 4470 1169 4507 1179
rect 4582 1178 4619 1179
rect 4563 1176 4619 1178
rect 4470 1149 4478 1169
rect 4498 1149 4507 1169
rect 4319 1138 4355 1139
rect 3670 1092 3707 1123
rect 3883 1121 3919 1123
rect 3883 1092 3920 1121
rect 3122 1083 3157 1084
rect 3099 1078 3157 1083
rect 3099 1058 3102 1078
rect 3122 1064 3157 1078
rect 3177 1064 3186 1084
rect 3122 1056 3186 1064
rect 3148 1055 3186 1056
rect 3149 1054 3186 1055
rect 3252 1088 3288 1089
rect 3360 1088 3396 1089
rect 3252 1080 3396 1088
rect 3252 1060 3260 1080
rect 3280 1060 3312 1080
rect 3336 1060 3368 1080
rect 3388 1060 3396 1080
rect 3252 1054 3396 1060
rect 3462 1084 3500 1092
rect 3568 1088 3604 1089
rect 3462 1064 3471 1084
rect 3491 1064 3500 1084
rect 3462 1055 3500 1064
rect 3519 1081 3604 1088
rect 3519 1061 3526 1081
rect 3547 1080 3604 1081
rect 3547 1061 3576 1080
rect 3519 1060 3576 1061
rect 3596 1060 3604 1080
rect 3462 1054 3499 1055
rect 3519 1054 3604 1060
rect 3670 1084 3708 1092
rect 3781 1088 3817 1089
rect 3670 1064 3679 1084
rect 3699 1064 3708 1084
rect 3670 1055 3708 1064
rect 3732 1080 3817 1088
rect 3732 1060 3789 1080
rect 3809 1060 3817 1080
rect 3670 1054 3707 1055
rect 3732 1054 3817 1060
rect 3883 1084 3921 1092
rect 3883 1064 3892 1084
rect 3912 1064 3921 1084
rect 4167 1079 4204 1080
rect 4470 1079 4507 1149
rect 4532 1169 4619 1176
rect 4532 1166 4590 1169
rect 4532 1146 4537 1166
rect 4558 1149 4590 1166
rect 4610 1149 4619 1169
rect 4558 1146 4619 1149
rect 4532 1139 4619 1146
rect 4678 1169 4715 1179
rect 4678 1149 4686 1169
rect 4706 1149 4715 1169
rect 4532 1138 4563 1139
rect 4166 1078 4507 1079
rect 3883 1055 3921 1064
rect 4091 1073 4507 1078
rect 3883 1054 3920 1055
rect 3306 1033 3342 1054
rect 3732 1033 3763 1054
rect 4091 1053 4094 1073
rect 4114 1053 4507 1073
rect 4678 1078 4715 1149
rect 4745 1178 4776 1231
rect 5428 1230 5438 1248
rect 5456 1234 6077 1248
rect 6617 1243 6735 1263
rect 6755 1243 6766 1263
rect 6617 1235 6766 1243
rect 6833 1267 7192 1271
rect 6833 1262 7155 1267
rect 6833 1238 6946 1262
rect 6970 1243 7155 1262
rect 7179 1243 7192 1267
rect 6970 1238 7192 1243
rect 6833 1235 7192 1238
rect 7254 1235 7289 1272
rect 7357 1269 7457 1272
rect 7357 1265 7424 1269
rect 7357 1239 7369 1265
rect 7395 1243 7424 1265
rect 7450 1243 7457 1269
rect 7395 1239 7457 1243
rect 7357 1235 7457 1239
rect 5456 1230 5466 1234
rect 5907 1233 6077 1234
rect 5078 1216 5115 1226
rect 5078 1198 5087 1216
rect 5105 1198 5115 1216
rect 5078 1189 5115 1198
rect 5428 1220 5466 1230
rect 4795 1178 4832 1179
rect 4745 1169 4832 1178
rect 4745 1149 4803 1169
rect 4823 1149 4832 1169
rect 4745 1139 4832 1149
rect 4891 1169 4928 1179
rect 4891 1149 4899 1169
rect 4919 1149 4928 1169
rect 4745 1138 4776 1139
rect 4891 1078 4928 1149
rect 5083 1124 5114 1189
rect 5428 1142 5463 1220
rect 6040 1210 6077 1233
rect 6833 1214 6864 1235
rect 7254 1214 7290 1235
rect 6676 1213 6713 1214
rect 5424 1133 5463 1142
rect 5082 1114 5119 1124
rect 5082 1112 5092 1114
rect 5016 1110 5092 1112
rect 4678 1054 4928 1078
rect 5013 1096 5092 1110
rect 5110 1096 5119 1114
rect 5424 1115 5434 1133
rect 5452 1115 5463 1133
rect 5424 1109 5463 1115
rect 5619 1185 5869 1209
rect 5619 1114 5656 1185
rect 5771 1124 5802 1125
rect 5424 1105 5461 1109
rect 5013 1093 5119 1096
rect 4485 1034 4506 1053
rect 5013 1034 5039 1093
rect 5082 1087 5119 1093
rect 5619 1094 5628 1114
rect 5648 1094 5656 1114
rect 5619 1084 5656 1094
rect 5715 1114 5802 1124
rect 5715 1094 5724 1114
rect 5744 1094 5802 1114
rect 5715 1085 5802 1094
rect 5715 1084 5752 1085
rect 5427 1034 5464 1043
rect 3139 1029 3239 1033
rect 3139 1025 3201 1029
rect 3139 999 3146 1025
rect 3172 1003 3201 1025
rect 3227 1003 3239 1029
rect 3172 999 3239 1003
rect 3139 996 3239 999
rect 3307 996 3342 1033
rect 3404 1030 3763 1033
rect 3404 1025 3626 1030
rect 3404 1001 3417 1025
rect 3441 1006 3626 1025
rect 3650 1006 3763 1030
rect 3441 1001 3763 1006
rect 3404 997 3763 1001
rect 3830 1025 3979 1033
rect 3830 1005 3841 1025
rect 3861 1005 3979 1025
rect 4485 1016 5039 1034
rect 5085 1023 5122 1025
rect 5013 1015 5039 1016
rect 5082 1015 5122 1023
rect 3830 998 3979 1005
rect 5082 1003 5094 1015
rect 5073 998 5094 1003
rect 3830 997 3871 998
rect 4489 997 5094 998
rect 5112 997 5122 1015
rect 3154 944 3191 945
rect 3250 944 3287 945
rect 3306 944 3342 996
rect 3361 944 3398 945
rect 3054 935 3192 944
rect 3054 915 3163 935
rect 3183 915 3192 935
rect 3054 908 3192 915
rect 3250 935 3398 944
rect 3250 915 3259 935
rect 3279 915 3369 935
rect 3389 915 3398 935
rect 3054 906 3150 908
rect 3250 905 3398 915
rect 3457 935 3494 945
rect 3569 944 3606 945
rect 3550 942 3606 944
rect 3457 915 3465 935
rect 3485 915 3494 935
rect 3306 904 3342 905
rect 3154 845 3191 846
rect 3457 845 3494 915
rect 3519 935 3606 942
rect 3519 932 3577 935
rect 3519 912 3524 932
rect 3545 915 3577 932
rect 3597 915 3606 935
rect 3545 912 3606 915
rect 3519 905 3606 912
rect 3665 935 3702 945
rect 3665 915 3673 935
rect 3693 915 3702 935
rect 3519 904 3550 905
rect 3153 844 3494 845
rect 3078 839 3494 844
rect 3078 819 3081 839
rect 3101 819 3494 839
rect 3665 844 3702 915
rect 3732 944 3763 997
rect 4489 988 5122 997
rect 5425 1016 5436 1034
rect 5454 1016 5464 1034
rect 5771 1032 5802 1085
rect 5832 1114 5869 1185
rect 6040 1190 6433 1210
rect 6453 1190 6456 1210
rect 6040 1185 6456 1190
rect 6675 1204 6713 1213
rect 6040 1184 6381 1185
rect 6675 1184 6684 1204
rect 6704 1184 6713 1204
rect 5984 1124 6015 1125
rect 5832 1094 5841 1114
rect 5861 1094 5869 1114
rect 5832 1084 5869 1094
rect 5928 1117 6015 1124
rect 5928 1114 5989 1117
rect 5928 1094 5937 1114
rect 5957 1097 5989 1114
rect 6010 1097 6015 1117
rect 5957 1094 6015 1097
rect 5928 1087 6015 1094
rect 6040 1114 6077 1184
rect 6343 1183 6380 1184
rect 6675 1176 6713 1184
rect 6779 1208 6864 1214
rect 6889 1213 6926 1214
rect 6779 1188 6787 1208
rect 6807 1188 6864 1208
rect 6779 1180 6864 1188
rect 6888 1204 6926 1213
rect 6888 1184 6897 1204
rect 6917 1184 6926 1204
rect 6779 1179 6815 1180
rect 6888 1176 6926 1184
rect 6992 1208 7077 1214
rect 7097 1213 7134 1214
rect 6992 1188 7000 1208
rect 7020 1207 7077 1208
rect 7020 1188 7049 1207
rect 6992 1187 7049 1188
rect 7070 1187 7077 1207
rect 6992 1180 7077 1187
rect 7096 1204 7134 1213
rect 7096 1184 7105 1204
rect 7125 1184 7134 1204
rect 6992 1179 7028 1180
rect 7096 1176 7134 1184
rect 7200 1208 7344 1214
rect 7200 1188 7208 1208
rect 7228 1207 7316 1208
rect 7228 1188 7261 1207
rect 7284 1188 7316 1207
rect 7336 1188 7344 1208
rect 7200 1180 7344 1188
rect 7200 1179 7236 1180
rect 7308 1179 7344 1180
rect 7410 1213 7447 1214
rect 7410 1212 7448 1213
rect 7410 1204 7474 1212
rect 7410 1184 7419 1204
rect 7439 1190 7474 1204
rect 7494 1190 7497 1210
rect 7439 1185 7497 1190
rect 7439 1184 7474 1185
rect 6676 1147 6713 1176
rect 6677 1145 6713 1147
rect 6889 1145 6926 1176
rect 6192 1124 6228 1125
rect 6040 1094 6049 1114
rect 6069 1094 6077 1114
rect 5928 1085 5984 1087
rect 5928 1084 5965 1085
rect 6040 1084 6077 1094
rect 6136 1114 6284 1124
rect 6677 1123 6926 1145
rect 7097 1144 7134 1176
rect 7410 1172 7474 1184
rect 7514 1146 7541 1324
rect 7373 1144 7541 1146
rect 7097 1133 7541 1144
rect 7604 1144 7634 2145
rect 7723 2138 7760 2149
rect 9344 2138 9371 2316
rect 9411 2278 9475 2290
rect 9751 2286 9788 2318
rect 9959 2317 10208 2339
rect 9959 2286 9996 2317
rect 10172 2315 10208 2317
rect 10351 2320 10389 2361
rect 10172 2286 10209 2315
rect 9411 2277 9446 2278
rect 9388 2272 9446 2277
rect 9388 2252 9391 2272
rect 9411 2258 9446 2272
rect 9466 2258 9475 2278
rect 9411 2250 9475 2258
rect 9437 2249 9475 2250
rect 9438 2248 9475 2249
rect 9541 2282 9577 2283
rect 9649 2282 9685 2283
rect 9541 2276 9685 2282
rect 9541 2274 9607 2276
rect 9541 2254 9549 2274
rect 9569 2255 9607 2274
rect 9629 2274 9685 2276
rect 9629 2255 9657 2274
rect 9569 2254 9657 2255
rect 9677 2254 9685 2274
rect 9541 2248 9685 2254
rect 9751 2278 9789 2286
rect 9857 2282 9893 2283
rect 9751 2258 9760 2278
rect 9780 2258 9789 2278
rect 9751 2249 9789 2258
rect 9808 2275 9893 2282
rect 9808 2255 9815 2275
rect 9836 2274 9893 2275
rect 9836 2255 9865 2274
rect 9808 2254 9865 2255
rect 9885 2254 9893 2274
rect 9751 2248 9788 2249
rect 9808 2248 9893 2254
rect 9959 2278 9997 2286
rect 10070 2282 10106 2283
rect 9959 2258 9968 2278
rect 9988 2258 9997 2278
rect 9959 2249 9997 2258
rect 10021 2274 10106 2282
rect 10021 2254 10078 2274
rect 10098 2254 10106 2274
rect 9959 2248 9996 2249
rect 10021 2248 10106 2254
rect 10172 2278 10210 2286
rect 10172 2258 10181 2278
rect 10201 2258 10210 2278
rect 10172 2249 10210 2258
rect 10351 2285 10387 2320
rect 10351 2275 10388 2285
rect 10351 2257 10361 2275
rect 10379 2257 10388 2275
rect 10172 2248 10209 2249
rect 10351 2248 10388 2257
rect 9595 2227 9631 2248
rect 10021 2227 10052 2248
rect 9428 2223 9528 2227
rect 9428 2219 9490 2223
rect 9428 2193 9435 2219
rect 9461 2197 9490 2219
rect 9516 2197 9528 2223
rect 9461 2193 9528 2197
rect 9428 2190 9528 2193
rect 9596 2190 9631 2227
rect 9693 2224 10052 2227
rect 9693 2219 9915 2224
rect 9693 2195 9706 2219
rect 9730 2200 9915 2219
rect 9939 2200 10052 2224
rect 9730 2195 10052 2200
rect 9693 2191 10052 2195
rect 10119 2219 10268 2227
rect 10119 2199 10130 2219
rect 10150 2199 10268 2219
rect 10119 2192 10268 2199
rect 10119 2191 10160 2192
rect 9443 2138 9480 2139
rect 9539 2138 9576 2139
rect 9595 2138 9631 2190
rect 9650 2138 9687 2139
rect 9343 2129 9481 2138
rect 8279 2111 8310 2114
rect 8279 2085 8286 2111
rect 8305 2085 8310 2111
rect 8279 1691 8310 2085
rect 8331 2110 8499 2111
rect 8331 2107 8775 2110
rect 8331 2088 8706 2107
rect 8726 2088 8775 2107
rect 9343 2109 9452 2129
rect 9472 2109 9481 2129
rect 8331 2084 8775 2088
rect 8331 2082 8499 2084
rect 8331 1904 8358 2082
rect 8398 2044 8462 2056
rect 8738 2052 8775 2084
rect 8946 2083 9195 2105
rect 9343 2102 9481 2109
rect 9539 2129 9687 2138
rect 9539 2109 9548 2129
rect 9568 2109 9658 2129
rect 9678 2109 9687 2129
rect 9343 2100 9439 2102
rect 9539 2099 9687 2109
rect 9746 2129 9783 2139
rect 9858 2138 9895 2139
rect 9839 2136 9895 2138
rect 9746 2109 9754 2129
rect 9774 2109 9783 2129
rect 9595 2098 9631 2099
rect 8946 2052 8983 2083
rect 9159 2081 9195 2083
rect 9159 2052 9196 2081
rect 8398 2043 8433 2044
rect 8375 2038 8433 2043
rect 8375 2018 8378 2038
rect 8398 2024 8433 2038
rect 8453 2024 8462 2044
rect 8398 2016 8462 2024
rect 8424 2015 8462 2016
rect 8425 2014 8462 2015
rect 8528 2048 8564 2049
rect 8636 2048 8672 2049
rect 8528 2040 8672 2048
rect 8528 2020 8536 2040
rect 8556 2039 8644 2040
rect 8556 2020 8589 2039
rect 8528 2019 8589 2020
rect 8613 2020 8644 2039
rect 8664 2020 8672 2040
rect 8613 2019 8672 2020
rect 8528 2014 8672 2019
rect 8738 2044 8776 2052
rect 8844 2048 8880 2049
rect 8738 2024 8747 2044
rect 8767 2024 8776 2044
rect 8738 2015 8776 2024
rect 8795 2041 8880 2048
rect 8795 2021 8802 2041
rect 8823 2040 8880 2041
rect 8823 2021 8852 2040
rect 8795 2020 8852 2021
rect 8872 2020 8880 2040
rect 8738 2014 8775 2015
rect 8795 2014 8880 2020
rect 8946 2044 8984 2052
rect 9057 2048 9093 2049
rect 8946 2024 8955 2044
rect 8975 2024 8984 2044
rect 8946 2015 8984 2024
rect 9008 2040 9093 2048
rect 9008 2020 9065 2040
rect 9085 2020 9093 2040
rect 8946 2014 8983 2015
rect 9008 2014 9093 2020
rect 9159 2044 9197 2052
rect 9159 2024 9168 2044
rect 9188 2024 9197 2044
rect 9443 2039 9480 2040
rect 9746 2039 9783 2109
rect 9808 2129 9895 2136
rect 9808 2126 9866 2129
rect 9808 2106 9813 2126
rect 9834 2109 9866 2126
rect 9886 2109 9895 2129
rect 9834 2106 9895 2109
rect 9808 2099 9895 2106
rect 9954 2129 9991 2139
rect 9954 2109 9962 2129
rect 9982 2109 9991 2129
rect 9808 2098 9839 2099
rect 9442 2038 9783 2039
rect 9159 2015 9197 2024
rect 9367 2033 9783 2038
rect 9159 2014 9196 2015
rect 8582 1993 8618 2014
rect 9008 1993 9039 2014
rect 9367 2013 9370 2033
rect 9390 2013 9783 2033
rect 9954 2038 9991 2109
rect 10021 2138 10052 2191
rect 10354 2176 10391 2186
rect 10354 2158 10363 2176
rect 10381 2158 10391 2176
rect 10354 2149 10391 2158
rect 10071 2138 10108 2139
rect 10021 2129 10108 2138
rect 10021 2109 10079 2129
rect 10099 2109 10108 2129
rect 10021 2099 10108 2109
rect 10167 2129 10204 2139
rect 10167 2109 10175 2129
rect 10195 2109 10204 2129
rect 10021 2098 10052 2099
rect 10167 2038 10204 2109
rect 10359 2084 10390 2149
rect 10358 2074 10395 2084
rect 10358 2072 10368 2074
rect 10292 2070 10368 2072
rect 9954 2014 10204 2038
rect 10289 2056 10368 2070
rect 10386 2056 10395 2074
rect 10289 2053 10395 2056
rect 9761 1994 9782 2013
rect 10289 1994 10315 2053
rect 10358 2047 10395 2053
rect 8415 1989 8515 1993
rect 8415 1985 8477 1989
rect 8415 1959 8422 1985
rect 8448 1963 8477 1985
rect 8503 1963 8515 1989
rect 8448 1959 8515 1963
rect 8415 1956 8515 1959
rect 8583 1956 8618 1993
rect 8680 1990 9039 1993
rect 8680 1985 8902 1990
rect 8680 1961 8693 1985
rect 8717 1966 8902 1985
rect 8926 1966 9039 1990
rect 8717 1961 9039 1966
rect 8680 1957 9039 1961
rect 9106 1985 9255 1993
rect 9106 1965 9117 1985
rect 9137 1965 9255 1985
rect 9761 1976 10315 1994
rect 10361 1983 10398 1985
rect 10289 1975 10315 1976
rect 10358 1975 10398 1983
rect 9106 1958 9255 1965
rect 10358 1963 10370 1975
rect 10349 1958 10370 1963
rect 9106 1957 9147 1958
rect 9765 1957 10370 1958
rect 10388 1957 10398 1975
rect 8430 1904 8467 1905
rect 8526 1904 8563 1905
rect 8582 1904 8618 1956
rect 8637 1904 8674 1905
rect 8330 1895 8468 1904
rect 8330 1875 8439 1895
rect 8459 1875 8468 1895
rect 8330 1868 8468 1875
rect 8526 1895 8674 1904
rect 8526 1875 8535 1895
rect 8555 1875 8645 1895
rect 8665 1875 8674 1895
rect 8330 1866 8426 1868
rect 8526 1865 8674 1875
rect 8733 1895 8770 1905
rect 8845 1904 8882 1905
rect 8826 1902 8882 1904
rect 8733 1875 8741 1895
rect 8761 1875 8770 1895
rect 8582 1864 8618 1865
rect 8430 1805 8467 1806
rect 8733 1805 8770 1875
rect 8795 1895 8882 1902
rect 8795 1892 8853 1895
rect 8795 1872 8800 1892
rect 8821 1875 8853 1892
rect 8873 1875 8882 1895
rect 8821 1872 8882 1875
rect 8795 1865 8882 1872
rect 8941 1895 8978 1905
rect 8941 1875 8949 1895
rect 8969 1875 8978 1895
rect 8795 1864 8826 1865
rect 8429 1804 8770 1805
rect 8354 1799 8770 1804
rect 8354 1779 8357 1799
rect 8377 1779 8770 1799
rect 8941 1804 8978 1875
rect 9008 1904 9039 1957
rect 9765 1948 10398 1957
rect 9765 1941 10397 1948
rect 9765 1939 9827 1941
rect 9343 1929 9511 1930
rect 9765 1929 9787 1939
rect 9058 1904 9095 1905
rect 9008 1895 9095 1904
rect 9008 1875 9066 1895
rect 9086 1875 9095 1895
rect 9008 1865 9095 1875
rect 9154 1895 9191 1905
rect 9154 1875 9162 1895
rect 9182 1875 9191 1895
rect 9008 1864 9039 1865
rect 9154 1804 9191 1875
rect 8941 1780 9191 1804
rect 9343 1903 9787 1929
rect 9343 1901 9511 1903
rect 9343 1723 9370 1901
rect 9410 1863 9474 1875
rect 9750 1871 9787 1903
rect 9958 1902 10207 1924
rect 9958 1871 9995 1902
rect 10171 1900 10207 1902
rect 10171 1871 10208 1900
rect 9410 1862 9445 1863
rect 9387 1857 9445 1862
rect 9387 1837 9390 1857
rect 9410 1843 9445 1857
rect 9465 1843 9474 1863
rect 9410 1835 9474 1843
rect 9436 1834 9474 1835
rect 9437 1833 9474 1834
rect 9540 1867 9576 1868
rect 9648 1867 9684 1868
rect 9540 1859 9684 1867
rect 9540 1839 9548 1859
rect 9568 1839 9597 1859
rect 9540 1838 9597 1839
rect 9619 1839 9656 1859
rect 9676 1839 9684 1859
rect 9619 1838 9684 1839
rect 9540 1833 9684 1838
rect 9750 1863 9788 1871
rect 9856 1867 9892 1868
rect 9750 1843 9759 1863
rect 9779 1843 9788 1863
rect 9750 1834 9788 1843
rect 9807 1860 9892 1867
rect 9807 1840 9814 1860
rect 9835 1859 9892 1860
rect 9835 1840 9864 1859
rect 9807 1839 9864 1840
rect 9884 1839 9892 1859
rect 9750 1833 9787 1834
rect 9807 1833 9892 1839
rect 9958 1863 9996 1871
rect 10069 1867 10105 1868
rect 9958 1843 9967 1863
rect 9987 1843 9996 1863
rect 9958 1834 9996 1843
rect 10020 1859 10105 1867
rect 10020 1839 10077 1859
rect 10097 1839 10105 1859
rect 9958 1833 9995 1834
rect 10020 1833 10105 1839
rect 10171 1863 10209 1871
rect 10171 1843 10180 1863
rect 10200 1843 10209 1863
rect 10171 1834 10209 1843
rect 10171 1833 10208 1834
rect 9594 1812 9630 1833
rect 10020 1812 10051 1833
rect 9427 1808 9527 1812
rect 9427 1804 9489 1808
rect 9427 1778 9434 1804
rect 9460 1782 9489 1804
rect 9515 1782 9527 1808
rect 9460 1778 9527 1782
rect 9427 1775 9527 1778
rect 9595 1775 9630 1812
rect 9692 1809 10051 1812
rect 9692 1804 9914 1809
rect 9692 1780 9705 1804
rect 9729 1785 9914 1804
rect 9938 1785 10051 1809
rect 9729 1780 10051 1785
rect 9692 1776 10051 1780
rect 10118 1804 10267 1812
rect 10118 1784 10129 1804
rect 10149 1784 10267 1804
rect 10118 1777 10267 1784
rect 10358 1792 10397 1941
rect 10118 1776 10159 1777
rect 9442 1723 9479 1724
rect 9538 1723 9575 1724
rect 9594 1723 9630 1775
rect 9649 1723 9686 1724
rect 9342 1714 9480 1723
rect 9342 1694 9451 1714
rect 9471 1694 9480 1714
rect 8279 1690 8449 1691
rect 8279 1675 8725 1690
rect 9342 1687 9480 1694
rect 9538 1714 9686 1723
rect 9538 1694 9547 1714
rect 9567 1694 9657 1714
rect 9677 1694 9686 1714
rect 9342 1685 9438 1687
rect 8281 1664 8725 1675
rect 8281 1662 8449 1664
rect 8281 1484 8308 1662
rect 8348 1624 8412 1636
rect 8688 1632 8725 1664
rect 8896 1663 9145 1685
rect 9538 1684 9686 1694
rect 9745 1714 9782 1724
rect 9857 1723 9894 1724
rect 9838 1721 9894 1723
rect 9745 1694 9753 1714
rect 9773 1694 9782 1714
rect 9594 1683 9630 1684
rect 8896 1632 8933 1663
rect 9109 1661 9145 1663
rect 9109 1632 9146 1661
rect 8348 1623 8383 1624
rect 8325 1618 8383 1623
rect 8325 1598 8328 1618
rect 8348 1604 8383 1618
rect 8403 1604 8412 1624
rect 8348 1596 8412 1604
rect 8374 1595 8412 1596
rect 8375 1594 8412 1595
rect 8478 1628 8514 1629
rect 8586 1628 8622 1629
rect 8478 1620 8622 1628
rect 8478 1600 8486 1620
rect 8506 1619 8594 1620
rect 8506 1602 8534 1619
rect 8558 1602 8594 1619
rect 8506 1600 8594 1602
rect 8614 1600 8622 1620
rect 8478 1594 8622 1600
rect 8688 1624 8726 1632
rect 8794 1628 8830 1629
rect 8688 1604 8697 1624
rect 8717 1604 8726 1624
rect 8688 1595 8726 1604
rect 8745 1621 8830 1628
rect 8745 1601 8752 1621
rect 8773 1620 8830 1621
rect 8773 1601 8802 1620
rect 8745 1600 8802 1601
rect 8822 1600 8830 1620
rect 8688 1594 8725 1595
rect 8745 1594 8830 1600
rect 8896 1624 8934 1632
rect 9007 1628 9043 1629
rect 8896 1604 8905 1624
rect 8925 1604 8934 1624
rect 8896 1595 8934 1604
rect 8958 1620 9043 1628
rect 8958 1600 9015 1620
rect 9035 1600 9043 1620
rect 8896 1594 8933 1595
rect 8958 1594 9043 1600
rect 9109 1624 9147 1632
rect 9442 1624 9479 1625
rect 9745 1624 9782 1694
rect 9807 1714 9894 1721
rect 9807 1711 9865 1714
rect 9807 1691 9812 1711
rect 9833 1694 9865 1711
rect 9885 1694 9894 1714
rect 9833 1691 9894 1694
rect 9807 1684 9894 1691
rect 9953 1714 9990 1724
rect 9953 1694 9961 1714
rect 9981 1694 9990 1714
rect 9807 1683 9838 1684
rect 9109 1604 9118 1624
rect 9138 1604 9147 1624
rect 9441 1623 9782 1624
rect 9109 1595 9147 1604
rect 9366 1618 9782 1623
rect 9366 1598 9369 1618
rect 9389 1598 9782 1618
rect 9953 1623 9990 1694
rect 10020 1723 10051 1776
rect 10358 1774 10368 1792
rect 10386 1774 10397 1792
rect 10358 1765 10395 1774
rect 10070 1723 10107 1724
rect 10020 1714 10107 1723
rect 10020 1694 10078 1714
rect 10098 1694 10107 1714
rect 10020 1684 10107 1694
rect 10166 1714 10203 1724
rect 10166 1694 10174 1714
rect 10194 1694 10203 1714
rect 10361 1699 10398 1703
rect 10020 1683 10051 1684
rect 10166 1623 10203 1694
rect 9953 1599 10203 1623
rect 10359 1693 10398 1699
rect 10359 1675 10370 1693
rect 10388 1675 10398 1693
rect 10359 1666 10398 1675
rect 9109 1594 9146 1595
rect 8532 1573 8568 1594
rect 8958 1573 8989 1594
rect 9745 1575 9782 1598
rect 10359 1588 10394 1666
rect 10356 1578 10394 1588
rect 9745 1574 9915 1575
rect 10356 1574 10366 1578
rect 8365 1569 8465 1573
rect 8365 1565 8427 1569
rect 8365 1539 8372 1565
rect 8398 1543 8427 1565
rect 8453 1543 8465 1569
rect 8398 1539 8465 1543
rect 8365 1536 8465 1539
rect 8533 1536 8568 1573
rect 8630 1570 8989 1573
rect 8630 1565 8852 1570
rect 8630 1541 8643 1565
rect 8667 1546 8852 1565
rect 8876 1546 8989 1570
rect 8667 1541 8989 1546
rect 8630 1537 8989 1541
rect 9056 1565 9205 1573
rect 9056 1545 9067 1565
rect 9087 1545 9205 1565
rect 9745 1560 10366 1574
rect 10384 1560 10394 1578
rect 9745 1554 10394 1560
rect 9745 1553 10393 1554
rect 10356 1551 10393 1553
rect 9056 1538 9205 1545
rect 9056 1537 9097 1538
rect 8380 1484 8417 1485
rect 8476 1484 8513 1485
rect 8532 1484 8568 1536
rect 8587 1484 8624 1485
rect 8280 1475 8418 1484
rect 8280 1455 8389 1475
rect 8409 1455 8418 1475
rect 8280 1448 8418 1455
rect 8476 1475 8624 1484
rect 8476 1455 8485 1475
rect 8505 1455 8595 1475
rect 8615 1455 8624 1475
rect 8280 1446 8376 1448
rect 8476 1445 8624 1455
rect 8683 1475 8720 1485
rect 8795 1484 8832 1485
rect 8776 1482 8832 1484
rect 8683 1455 8691 1475
rect 8711 1455 8720 1475
rect 8532 1444 8568 1445
rect 8380 1385 8417 1386
rect 8683 1385 8720 1455
rect 8745 1475 8832 1482
rect 8745 1472 8803 1475
rect 8745 1452 8750 1472
rect 8771 1455 8803 1472
rect 8823 1455 8832 1475
rect 8771 1452 8832 1455
rect 8745 1445 8832 1452
rect 8891 1475 8928 1485
rect 8891 1455 8899 1475
rect 8919 1455 8928 1475
rect 8745 1444 8776 1445
rect 8379 1384 8720 1385
rect 8304 1379 8720 1384
rect 8304 1359 8307 1379
rect 8327 1359 8720 1379
rect 8891 1384 8928 1455
rect 8958 1484 8989 1537
rect 9008 1484 9045 1485
rect 8958 1475 9045 1484
rect 8958 1455 9016 1475
rect 9036 1455 9045 1475
rect 8958 1445 9045 1455
rect 9104 1475 9141 1485
rect 9104 1455 9112 1475
rect 9132 1455 9141 1475
rect 8958 1444 8989 1445
rect 9104 1384 9141 1455
rect 10359 1479 10396 1489
rect 10359 1461 10368 1479
rect 10386 1461 10396 1479
rect 10359 1452 10396 1461
rect 10359 1428 10394 1452
rect 10357 1404 10394 1428
rect 10356 1398 10394 1404
rect 8891 1360 9141 1384
rect 9767 1380 10394 1398
rect 9349 1363 9517 1364
rect 9768 1363 9792 1380
rect 9349 1337 9793 1363
rect 9349 1335 9517 1337
rect 9349 1157 9376 1335
rect 9416 1297 9480 1309
rect 9756 1305 9793 1337
rect 9964 1336 10213 1358
rect 9964 1305 10001 1336
rect 10177 1334 10213 1336
rect 10356 1339 10394 1380
rect 10177 1305 10214 1334
rect 9416 1296 9451 1297
rect 9393 1291 9451 1296
rect 9393 1271 9396 1291
rect 9416 1277 9451 1291
rect 9471 1277 9480 1297
rect 9416 1269 9480 1277
rect 9442 1268 9480 1269
rect 9443 1267 9480 1268
rect 9546 1301 9582 1302
rect 9654 1301 9690 1302
rect 9546 1295 9690 1301
rect 9546 1293 9612 1295
rect 9546 1273 9554 1293
rect 9574 1274 9612 1293
rect 9634 1293 9690 1295
rect 9634 1274 9662 1293
rect 9574 1273 9662 1274
rect 9682 1273 9690 1293
rect 9546 1267 9690 1273
rect 9756 1297 9794 1305
rect 9862 1301 9898 1302
rect 9756 1277 9765 1297
rect 9785 1277 9794 1297
rect 9756 1268 9794 1277
rect 9813 1294 9898 1301
rect 9813 1274 9820 1294
rect 9841 1293 9898 1294
rect 9841 1274 9870 1293
rect 9813 1273 9870 1274
rect 9890 1273 9898 1293
rect 9756 1267 9793 1268
rect 9813 1267 9898 1273
rect 9964 1297 10002 1305
rect 10075 1301 10111 1302
rect 9964 1277 9973 1297
rect 9993 1277 10002 1297
rect 9964 1268 10002 1277
rect 10026 1293 10111 1301
rect 10026 1273 10083 1293
rect 10103 1273 10111 1293
rect 9964 1267 10001 1268
rect 10026 1267 10111 1273
rect 10177 1297 10215 1305
rect 10177 1277 10186 1297
rect 10206 1277 10215 1297
rect 10177 1268 10215 1277
rect 10356 1304 10392 1339
rect 10356 1294 10393 1304
rect 10356 1276 10366 1294
rect 10384 1276 10393 1294
rect 10177 1267 10214 1268
rect 10356 1267 10393 1276
rect 9600 1246 9636 1267
rect 10026 1246 10057 1267
rect 9433 1242 9533 1246
rect 9433 1238 9495 1242
rect 9433 1212 9440 1238
rect 9466 1216 9495 1238
rect 9521 1216 9533 1242
rect 9466 1212 9533 1216
rect 9433 1209 9533 1212
rect 9601 1209 9636 1246
rect 9698 1243 10057 1246
rect 9698 1238 9920 1243
rect 9698 1214 9711 1238
rect 9735 1219 9920 1238
rect 9944 1219 10057 1243
rect 9735 1214 10057 1219
rect 9698 1210 10057 1214
rect 10124 1238 10273 1246
rect 10124 1218 10135 1238
rect 10155 1218 10273 1238
rect 10124 1211 10273 1218
rect 10124 1210 10165 1211
rect 9448 1157 9485 1158
rect 9544 1157 9581 1158
rect 9600 1157 9636 1209
rect 9655 1157 9692 1158
rect 9348 1148 9486 1157
rect 7604 1139 7636 1144
rect 6384 1121 6480 1123
rect 6136 1094 6145 1114
rect 6165 1094 6255 1114
rect 6275 1094 6284 1114
rect 6136 1085 6284 1094
rect 6342 1114 6480 1121
rect 7097 1118 7543 1133
rect 7373 1117 7543 1118
rect 6342 1094 6351 1114
rect 6371 1094 6480 1114
rect 6342 1085 6480 1094
rect 6136 1084 6173 1085
rect 6192 1033 6228 1085
rect 6247 1084 6284 1085
rect 6343 1084 6380 1085
rect 5663 1031 5704 1032
rect 4489 981 5121 988
rect 4489 979 4551 981
rect 4067 969 4235 970
rect 4489 969 4511 979
rect 3782 944 3819 945
rect 3732 935 3819 944
rect 3732 915 3790 935
rect 3810 915 3819 935
rect 3732 905 3819 915
rect 3878 935 3915 945
rect 3878 915 3886 935
rect 3906 915 3915 935
rect 3732 904 3763 905
rect 3878 844 3915 915
rect 3665 820 3915 844
rect 4067 943 4511 969
rect 4067 941 4235 943
rect 4067 763 4094 941
rect 4134 903 4198 915
rect 4474 911 4511 943
rect 4682 942 4931 964
rect 4682 911 4719 942
rect 4895 940 4931 942
rect 4895 911 4932 940
rect 4134 902 4169 903
rect 4111 897 4169 902
rect 4111 877 4114 897
rect 4134 883 4169 897
rect 4189 883 4198 903
rect 4134 875 4198 883
rect 4160 874 4198 875
rect 4161 873 4198 874
rect 4264 907 4300 908
rect 4372 907 4408 908
rect 4264 899 4408 907
rect 4264 879 4272 899
rect 4292 879 4321 899
rect 4264 878 4321 879
rect 4343 879 4380 899
rect 4400 879 4408 899
rect 4343 878 4408 879
rect 4264 873 4408 878
rect 4474 903 4512 911
rect 4580 907 4616 908
rect 4474 883 4483 903
rect 4503 883 4512 903
rect 4474 874 4512 883
rect 4531 900 4616 907
rect 4531 880 4538 900
rect 4559 899 4616 900
rect 4559 880 4588 899
rect 4531 879 4588 880
rect 4608 879 4616 899
rect 4474 873 4511 874
rect 4531 873 4616 879
rect 4682 903 4720 911
rect 4793 907 4829 908
rect 4682 883 4691 903
rect 4711 883 4720 903
rect 4682 874 4720 883
rect 4744 899 4829 907
rect 4744 879 4801 899
rect 4821 879 4829 899
rect 4682 873 4719 874
rect 4744 873 4829 879
rect 4895 903 4933 911
rect 4895 883 4904 903
rect 4924 883 4933 903
rect 4895 874 4933 883
rect 4895 873 4932 874
rect 4318 852 4354 873
rect 4744 852 4775 873
rect 4151 848 4251 852
rect 4151 844 4213 848
rect 4151 818 4158 844
rect 4184 822 4213 844
rect 4239 822 4251 848
rect 4184 818 4251 822
rect 4151 815 4251 818
rect 4319 815 4354 852
rect 4416 849 4775 852
rect 4416 844 4638 849
rect 4416 820 4429 844
rect 4453 825 4638 844
rect 4662 825 4775 849
rect 4453 820 4775 825
rect 4416 816 4775 820
rect 4842 844 4991 852
rect 4842 824 4853 844
rect 4873 824 4991 844
rect 4842 817 4991 824
rect 5082 832 5121 981
rect 5425 867 5464 1016
rect 5555 1024 5704 1031
rect 5555 1004 5673 1024
rect 5693 1004 5704 1024
rect 5555 996 5704 1004
rect 5771 1028 6130 1032
rect 5771 1023 6093 1028
rect 5771 999 5884 1023
rect 5908 1004 6093 1023
rect 6117 1004 6130 1028
rect 5908 999 6130 1004
rect 5771 996 6130 999
rect 6192 996 6227 1033
rect 6295 1030 6395 1033
rect 6295 1026 6362 1030
rect 6295 1000 6307 1026
rect 6333 1004 6362 1026
rect 6388 1004 6395 1030
rect 6333 1000 6395 1004
rect 6295 996 6395 1000
rect 5771 975 5802 996
rect 6192 975 6228 996
rect 5614 974 5651 975
rect 5613 965 5651 974
rect 5613 945 5622 965
rect 5642 945 5651 965
rect 5613 937 5651 945
rect 5717 969 5802 975
rect 5827 974 5864 975
rect 5717 949 5725 969
rect 5745 949 5802 969
rect 5717 941 5802 949
rect 5826 965 5864 974
rect 5826 945 5835 965
rect 5855 945 5864 965
rect 5717 940 5753 941
rect 5826 937 5864 945
rect 5930 969 6015 975
rect 6035 974 6072 975
rect 5930 949 5938 969
rect 5958 968 6015 969
rect 5958 949 5987 968
rect 5930 948 5987 949
rect 6008 948 6015 968
rect 5930 941 6015 948
rect 6034 965 6072 974
rect 6034 945 6043 965
rect 6063 945 6072 965
rect 5930 940 5966 941
rect 6034 937 6072 945
rect 6138 970 6282 975
rect 6138 969 6203 970
rect 6138 949 6146 969
rect 6166 949 6203 969
rect 6225 969 6282 970
rect 6225 949 6254 969
rect 6274 949 6282 969
rect 6138 941 6282 949
rect 6138 940 6174 941
rect 6246 940 6282 941
rect 6348 974 6385 975
rect 6348 973 6386 974
rect 6348 965 6412 973
rect 6348 945 6357 965
rect 6377 951 6412 965
rect 6432 951 6435 971
rect 6377 946 6435 951
rect 6377 945 6412 946
rect 5614 908 5651 937
rect 5615 906 5651 908
rect 5827 906 5864 937
rect 5615 884 5864 906
rect 6035 905 6072 937
rect 6348 933 6412 945
rect 6452 907 6479 1085
rect 6311 905 6479 907
rect 6035 879 6479 905
rect 6631 1004 6881 1028
rect 6631 933 6668 1004
rect 6783 943 6814 944
rect 6631 913 6640 933
rect 6660 913 6668 933
rect 6631 903 6668 913
rect 6727 933 6814 943
rect 6727 913 6736 933
rect 6756 913 6814 933
rect 6727 904 6814 913
rect 6727 903 6764 904
rect 6035 869 6057 879
rect 6311 878 6479 879
rect 5995 867 6057 869
rect 5425 860 6057 867
rect 4842 816 4883 817
rect 4166 763 4203 764
rect 4262 763 4299 764
rect 4318 763 4354 815
rect 4373 763 4410 764
rect 2231 718 2236 744
rect 2255 718 2262 744
rect 4066 754 4204 763
rect 4066 734 4175 754
rect 4195 734 4204 754
rect 4066 727 4204 734
rect 4262 754 4410 763
rect 4262 734 4271 754
rect 4291 734 4381 754
rect 4401 734 4410 754
rect 4066 725 4162 727
rect 4262 724 4410 734
rect 4469 754 4506 764
rect 4581 763 4618 764
rect 4562 761 4618 763
rect 4469 734 4477 754
rect 4497 734 4506 754
rect 4318 723 4354 724
rect 2231 715 2262 718
rect 1060 691 1198 700
rect 854 690 891 691
rect 910 639 946 691
rect 965 690 1002 691
rect 1061 690 1098 691
rect 381 637 422 638
rect 273 630 422 637
rect 273 610 391 630
rect 411 610 422 630
rect 273 602 422 610
rect 489 634 848 638
rect 489 629 811 634
rect 489 605 602 629
rect 626 610 811 629
rect 835 610 848 634
rect 626 605 848 610
rect 489 602 848 605
rect 910 602 945 639
rect 1013 636 1113 639
rect 1013 632 1080 636
rect 1013 606 1025 632
rect 1051 610 1080 632
rect 1106 610 1113 636
rect 1051 606 1113 610
rect 1013 602 1113 606
rect 489 581 520 602
rect 910 581 946 602
rect 153 572 190 581
rect 332 580 369 581
rect 153 554 162 572
rect 180 554 190 572
rect 153 544 190 554
rect 154 509 190 544
rect 331 571 369 580
rect 331 551 340 571
rect 360 551 369 571
rect 331 543 369 551
rect 435 575 520 581
rect 545 580 582 581
rect 435 555 443 575
rect 463 555 520 575
rect 435 547 520 555
rect 544 571 582 580
rect 544 551 553 571
rect 573 551 582 571
rect 435 546 471 547
rect 544 543 582 551
rect 648 575 733 581
rect 753 580 790 581
rect 648 555 656 575
rect 676 574 733 575
rect 676 555 705 574
rect 648 554 705 555
rect 726 554 733 574
rect 648 547 733 554
rect 752 571 790 580
rect 752 551 761 571
rect 781 551 790 571
rect 648 546 684 547
rect 752 543 790 551
rect 856 575 1000 581
rect 856 555 864 575
rect 884 574 972 575
rect 884 555 912 574
rect 856 553 912 555
rect 934 555 972 574
rect 992 555 1000 575
rect 934 553 1000 555
rect 856 547 1000 553
rect 856 546 892 547
rect 964 546 1000 547
rect 1066 580 1103 581
rect 1066 579 1104 580
rect 1066 571 1130 579
rect 1066 551 1075 571
rect 1095 557 1130 571
rect 1150 557 1153 577
rect 1095 552 1153 557
rect 1095 551 1130 552
rect 332 514 369 543
rect 152 444 190 509
rect 333 512 369 514
rect 545 512 582 543
rect 333 490 582 512
rect 753 511 790 543
rect 1066 539 1130 551
rect 1170 513 1197 691
rect 4166 664 4203 665
rect 4469 664 4506 734
rect 4531 754 4618 761
rect 4531 751 4589 754
rect 4531 731 4536 751
rect 4557 734 4589 751
rect 4609 734 4618 754
rect 4557 731 4618 734
rect 4531 724 4618 731
rect 4677 754 4714 764
rect 4677 734 4685 754
rect 4705 734 4714 754
rect 4531 723 4562 724
rect 4165 663 4506 664
rect 4090 658 4506 663
rect 4090 638 4093 658
rect 4113 638 4506 658
rect 4677 663 4714 734
rect 4744 763 4775 816
rect 5082 814 5092 832
rect 5110 814 5121 832
rect 5424 851 6057 860
rect 6783 851 6814 904
rect 6844 933 6881 1004
rect 7052 1009 7445 1029
rect 7465 1009 7468 1029
rect 7052 1004 7468 1009
rect 7052 1003 7393 1004
rect 6996 943 7027 944
rect 6844 913 6853 933
rect 6873 913 6881 933
rect 6844 903 6881 913
rect 6940 936 7027 943
rect 6940 933 7001 936
rect 6940 913 6949 933
rect 6969 916 7001 933
rect 7022 916 7027 936
rect 6969 913 7027 916
rect 6940 906 7027 913
rect 7052 933 7089 1003
rect 7355 1002 7392 1003
rect 7204 943 7240 944
rect 7052 913 7061 933
rect 7081 913 7089 933
rect 6940 904 6996 906
rect 6940 903 6977 904
rect 7052 903 7089 913
rect 7148 933 7296 943
rect 7396 940 7492 942
rect 7148 913 7157 933
rect 7177 913 7267 933
rect 7287 913 7296 933
rect 7148 904 7296 913
rect 7354 933 7492 940
rect 7354 913 7363 933
rect 7383 913 7492 933
rect 7354 904 7492 913
rect 7148 903 7185 904
rect 7204 852 7240 904
rect 7259 903 7296 904
rect 7355 903 7392 904
rect 5424 833 5434 851
rect 5452 850 6057 851
rect 6675 850 6716 851
rect 5452 845 5473 850
rect 5452 833 5464 845
rect 6567 843 6716 850
rect 5424 825 5464 833
rect 5507 832 5533 833
rect 5424 823 5461 825
rect 5507 814 6061 832
rect 6567 823 6685 843
rect 6705 823 6716 843
rect 6567 815 6716 823
rect 6783 847 7142 851
rect 6783 842 7105 847
rect 6783 818 6896 842
rect 6920 823 7105 842
rect 7129 823 7142 847
rect 6920 818 7142 823
rect 6783 815 7142 818
rect 7204 815 7239 852
rect 7307 849 7407 852
rect 7307 845 7374 849
rect 7307 819 7319 845
rect 7345 823 7374 845
rect 7400 823 7407 849
rect 7345 819 7407 823
rect 7307 815 7407 819
rect 5082 805 5119 814
rect 4794 763 4831 764
rect 4744 754 4831 763
rect 4744 734 4802 754
rect 4822 734 4831 754
rect 4744 724 4831 734
rect 4890 754 4927 764
rect 4890 734 4898 754
rect 4918 734 4927 754
rect 5427 755 5464 761
rect 5507 755 5533 814
rect 6040 795 6061 814
rect 5427 752 5533 755
rect 5085 739 5122 743
rect 4744 723 4775 724
rect 4890 663 4927 734
rect 4677 639 4927 663
rect 5083 733 5122 739
rect 5083 715 5094 733
rect 5112 715 5122 733
rect 5427 734 5436 752
rect 5454 738 5533 752
rect 5618 770 5868 794
rect 5454 736 5530 738
rect 5454 734 5464 736
rect 5427 724 5464 734
rect 5083 706 5122 715
rect 4469 615 4506 638
rect 5083 628 5118 706
rect 5432 659 5463 724
rect 5618 699 5655 770
rect 5770 709 5801 710
rect 5618 679 5627 699
rect 5647 679 5655 699
rect 5618 669 5655 679
rect 5714 699 5801 709
rect 5714 679 5723 699
rect 5743 679 5801 699
rect 5714 670 5801 679
rect 5714 669 5751 670
rect 5080 618 5118 628
rect 5431 650 5468 659
rect 5431 632 5441 650
rect 5459 632 5468 650
rect 5431 622 5468 632
rect 4469 614 4639 615
rect 5080 614 5090 618
rect 4469 600 5090 614
rect 5108 600 5118 618
rect 5770 617 5801 670
rect 5831 699 5868 770
rect 6039 775 6432 795
rect 6452 775 6455 795
rect 6783 794 6814 815
rect 7204 794 7240 815
rect 6626 793 6663 794
rect 6039 770 6455 775
rect 6625 784 6663 793
rect 6039 769 6380 770
rect 5983 709 6014 710
rect 5831 679 5840 699
rect 5860 679 5868 699
rect 5831 669 5868 679
rect 5927 702 6014 709
rect 5927 699 5988 702
rect 5927 679 5936 699
rect 5956 682 5988 699
rect 6009 682 6014 702
rect 5956 679 6014 682
rect 5927 672 6014 679
rect 6039 699 6076 769
rect 6342 768 6379 769
rect 6625 764 6634 784
rect 6654 764 6663 784
rect 6625 756 6663 764
rect 6729 788 6814 794
rect 6839 793 6876 794
rect 6729 768 6737 788
rect 6757 768 6814 788
rect 6729 760 6814 768
rect 6838 784 6876 793
rect 6838 764 6847 784
rect 6867 764 6876 784
rect 6729 759 6765 760
rect 6838 756 6876 764
rect 6942 788 7027 794
rect 7047 793 7084 794
rect 6942 768 6950 788
rect 6970 787 7027 788
rect 6970 768 6999 787
rect 6942 767 6999 768
rect 7020 767 7027 787
rect 6942 760 7027 767
rect 7046 784 7084 793
rect 7046 764 7055 784
rect 7075 764 7084 784
rect 6942 759 6978 760
rect 7046 756 7084 764
rect 7150 789 7294 794
rect 7150 788 7209 789
rect 7150 768 7158 788
rect 7178 769 7209 788
rect 7233 788 7294 789
rect 7233 769 7266 788
rect 7178 768 7266 769
rect 7286 768 7294 788
rect 7150 760 7294 768
rect 7150 759 7186 760
rect 7258 759 7294 760
rect 7360 793 7397 794
rect 7360 792 7398 793
rect 7360 784 7424 792
rect 7360 764 7369 784
rect 7389 770 7424 784
rect 7444 770 7447 790
rect 7389 765 7447 770
rect 7389 764 7424 765
rect 6626 727 6663 756
rect 6627 725 6663 727
rect 6839 725 6876 756
rect 6191 709 6227 710
rect 6039 679 6048 699
rect 6068 679 6076 699
rect 5927 670 5983 672
rect 5927 669 5964 670
rect 6039 669 6076 679
rect 6135 699 6283 709
rect 6383 706 6479 708
rect 6135 679 6144 699
rect 6164 679 6254 699
rect 6274 679 6283 699
rect 6135 670 6283 679
rect 6341 699 6479 706
rect 6627 703 6876 725
rect 7047 724 7084 756
rect 7360 752 7424 764
rect 7464 726 7491 904
rect 7323 724 7491 726
rect 7047 720 7491 724
rect 6341 679 6350 699
rect 6370 679 6479 699
rect 7047 701 7096 720
rect 7116 701 7491 720
rect 7047 698 7491 701
rect 7323 697 7491 698
rect 7512 723 7543 1117
rect 7604 1121 7609 1139
rect 7629 1121 7636 1139
rect 7604 1116 7636 1121
rect 7607 1114 7636 1116
rect 8336 1129 8504 1130
rect 8336 1126 8780 1129
rect 8336 1107 8711 1126
rect 8731 1107 8780 1126
rect 9348 1128 9457 1148
rect 9477 1128 9486 1148
rect 8336 1103 8780 1107
rect 8336 1101 8504 1103
rect 8336 923 8363 1101
rect 8403 1063 8467 1075
rect 8743 1071 8780 1103
rect 8951 1102 9200 1124
rect 9348 1121 9486 1128
rect 9544 1148 9692 1157
rect 9544 1128 9553 1148
rect 9573 1128 9663 1148
rect 9683 1128 9692 1148
rect 9348 1119 9444 1121
rect 9544 1118 9692 1128
rect 9751 1148 9788 1158
rect 9863 1157 9900 1158
rect 9844 1155 9900 1157
rect 9751 1128 9759 1148
rect 9779 1128 9788 1148
rect 9600 1117 9636 1118
rect 8951 1071 8988 1102
rect 9164 1100 9200 1102
rect 9164 1071 9201 1100
rect 8403 1062 8438 1063
rect 8380 1057 8438 1062
rect 8380 1037 8383 1057
rect 8403 1043 8438 1057
rect 8458 1043 8467 1063
rect 8403 1035 8467 1043
rect 8429 1034 8467 1035
rect 8430 1033 8467 1034
rect 8533 1067 8569 1068
rect 8641 1067 8677 1068
rect 8533 1059 8677 1067
rect 8533 1039 8541 1059
rect 8561 1039 8593 1059
rect 8617 1039 8649 1059
rect 8669 1039 8677 1059
rect 8533 1033 8677 1039
rect 8743 1063 8781 1071
rect 8849 1067 8885 1068
rect 8743 1043 8752 1063
rect 8772 1043 8781 1063
rect 8743 1034 8781 1043
rect 8800 1060 8885 1067
rect 8800 1040 8807 1060
rect 8828 1059 8885 1060
rect 8828 1040 8857 1059
rect 8800 1039 8857 1040
rect 8877 1039 8885 1059
rect 8743 1033 8780 1034
rect 8800 1033 8885 1039
rect 8951 1063 8989 1071
rect 9062 1067 9098 1068
rect 8951 1043 8960 1063
rect 8980 1043 8989 1063
rect 8951 1034 8989 1043
rect 9013 1059 9098 1067
rect 9013 1039 9070 1059
rect 9090 1039 9098 1059
rect 8951 1033 8988 1034
rect 9013 1033 9098 1039
rect 9164 1063 9202 1071
rect 9164 1043 9173 1063
rect 9193 1043 9202 1063
rect 9448 1058 9485 1059
rect 9751 1058 9788 1128
rect 9813 1148 9900 1155
rect 9813 1145 9871 1148
rect 9813 1125 9818 1145
rect 9839 1128 9871 1145
rect 9891 1128 9900 1148
rect 9839 1125 9900 1128
rect 9813 1118 9900 1125
rect 9959 1148 9996 1158
rect 9959 1128 9967 1148
rect 9987 1128 9996 1148
rect 9813 1117 9844 1118
rect 9447 1057 9788 1058
rect 9164 1034 9202 1043
rect 9372 1052 9788 1057
rect 9164 1033 9201 1034
rect 8587 1012 8623 1033
rect 9013 1012 9044 1033
rect 9372 1032 9375 1052
rect 9395 1032 9788 1052
rect 9959 1057 9996 1128
rect 10026 1157 10057 1210
rect 10359 1195 10396 1205
rect 10359 1177 10368 1195
rect 10386 1177 10396 1195
rect 10359 1168 10396 1177
rect 10076 1157 10113 1158
rect 10026 1148 10113 1157
rect 10026 1128 10084 1148
rect 10104 1128 10113 1148
rect 10026 1118 10113 1128
rect 10172 1148 10209 1158
rect 10172 1128 10180 1148
rect 10200 1128 10209 1148
rect 10026 1117 10057 1118
rect 10172 1057 10209 1128
rect 10364 1103 10395 1168
rect 10363 1093 10400 1103
rect 10363 1091 10373 1093
rect 10297 1089 10373 1091
rect 9959 1033 10209 1057
rect 10294 1075 10373 1089
rect 10391 1075 10400 1093
rect 10294 1072 10400 1075
rect 9766 1013 9787 1032
rect 10294 1013 10320 1072
rect 10363 1066 10400 1072
rect 8420 1008 8520 1012
rect 8420 1004 8482 1008
rect 8420 978 8427 1004
rect 8453 982 8482 1004
rect 8508 982 8520 1008
rect 8453 978 8520 982
rect 8420 975 8520 978
rect 8588 975 8623 1012
rect 8685 1009 9044 1012
rect 8685 1004 8907 1009
rect 8685 980 8698 1004
rect 8722 985 8907 1004
rect 8931 985 9044 1009
rect 8722 980 9044 985
rect 8685 976 9044 980
rect 9111 1004 9260 1012
rect 9111 984 9122 1004
rect 9142 984 9260 1004
rect 9766 995 10320 1013
rect 10366 1002 10403 1004
rect 10294 994 10320 995
rect 10363 994 10403 1002
rect 9111 977 9260 984
rect 10363 982 10375 994
rect 10354 977 10375 982
rect 9111 976 9152 977
rect 9770 976 10375 977
rect 10393 976 10403 994
rect 8435 923 8472 924
rect 8531 923 8568 924
rect 8587 923 8623 975
rect 8642 923 8679 924
rect 8335 914 8473 923
rect 8335 894 8444 914
rect 8464 894 8473 914
rect 8335 887 8473 894
rect 8531 914 8679 923
rect 8531 894 8540 914
rect 8560 894 8650 914
rect 8670 894 8679 914
rect 8335 885 8431 887
rect 8531 884 8679 894
rect 8738 914 8775 924
rect 8850 923 8887 924
rect 8831 921 8887 923
rect 8738 894 8746 914
rect 8766 894 8775 914
rect 8587 883 8623 884
rect 8435 824 8472 825
rect 8738 824 8775 894
rect 8800 914 8887 921
rect 8800 911 8858 914
rect 8800 891 8805 911
rect 8826 894 8858 911
rect 8878 894 8887 914
rect 8826 891 8887 894
rect 8800 884 8887 891
rect 8946 914 8983 924
rect 8946 894 8954 914
rect 8974 894 8983 914
rect 8800 883 8831 884
rect 8434 823 8775 824
rect 8359 818 8775 823
rect 8359 798 8362 818
rect 8382 798 8775 818
rect 8946 823 8983 894
rect 9013 923 9044 976
rect 9770 967 10403 976
rect 9770 960 10402 967
rect 9770 958 9832 960
rect 9348 948 9516 949
rect 9770 948 9792 958
rect 9063 923 9100 924
rect 9013 914 9100 923
rect 9013 894 9071 914
rect 9091 894 9100 914
rect 9013 884 9100 894
rect 9159 914 9196 924
rect 9159 894 9167 914
rect 9187 894 9196 914
rect 9013 883 9044 884
rect 9159 823 9196 894
rect 8946 799 9196 823
rect 9348 922 9792 948
rect 9348 920 9516 922
rect 9348 742 9375 920
rect 9415 882 9479 894
rect 9755 890 9792 922
rect 9963 921 10212 943
rect 9963 890 10000 921
rect 10176 919 10212 921
rect 10176 890 10213 919
rect 9415 881 9450 882
rect 9392 876 9450 881
rect 9392 856 9395 876
rect 9415 862 9450 876
rect 9470 862 9479 882
rect 9415 854 9479 862
rect 9441 853 9479 854
rect 9442 852 9479 853
rect 9545 886 9581 887
rect 9653 886 9689 887
rect 9545 878 9689 886
rect 9545 858 9553 878
rect 9573 858 9602 878
rect 9545 857 9602 858
rect 9624 858 9661 878
rect 9681 858 9689 878
rect 9624 857 9689 858
rect 9545 852 9689 857
rect 9755 882 9793 890
rect 9861 886 9897 887
rect 9755 862 9764 882
rect 9784 862 9793 882
rect 9755 853 9793 862
rect 9812 879 9897 886
rect 9812 859 9819 879
rect 9840 878 9897 879
rect 9840 859 9869 878
rect 9812 858 9869 859
rect 9889 858 9897 878
rect 9755 852 9792 853
rect 9812 852 9897 858
rect 9963 882 10001 890
rect 10074 886 10110 887
rect 9963 862 9972 882
rect 9992 862 10001 882
rect 9963 853 10001 862
rect 10025 878 10110 886
rect 10025 858 10082 878
rect 10102 858 10110 878
rect 9963 852 10000 853
rect 10025 852 10110 858
rect 10176 882 10214 890
rect 10176 862 10185 882
rect 10205 862 10214 882
rect 10176 853 10214 862
rect 10176 852 10213 853
rect 9599 831 9635 852
rect 10025 831 10056 852
rect 9432 827 9532 831
rect 9432 823 9494 827
rect 9432 797 9439 823
rect 9465 801 9494 823
rect 9520 801 9532 827
rect 9465 797 9532 801
rect 9432 794 9532 797
rect 9600 794 9635 831
rect 9697 828 10056 831
rect 9697 823 9919 828
rect 9697 799 9710 823
rect 9734 804 9919 823
rect 9943 804 10056 828
rect 9734 799 10056 804
rect 9697 795 10056 799
rect 10123 823 10272 831
rect 10123 803 10134 823
rect 10154 803 10272 823
rect 10123 796 10272 803
rect 10363 811 10402 960
rect 10123 795 10164 796
rect 9447 742 9484 743
rect 9543 742 9580 743
rect 9599 742 9635 794
rect 9654 742 9691 743
rect 7512 697 7517 723
rect 7536 697 7543 723
rect 9347 733 9485 742
rect 9347 713 9456 733
rect 9476 713 9485 733
rect 9347 706 9485 713
rect 9543 733 9691 742
rect 9543 713 9552 733
rect 9572 713 9662 733
rect 9682 713 9691 733
rect 9347 704 9443 706
rect 9543 703 9691 713
rect 9750 733 9787 743
rect 9862 742 9899 743
rect 9843 740 9899 742
rect 9750 713 9758 733
rect 9778 713 9787 733
rect 9599 702 9635 703
rect 7512 694 7543 697
rect 6341 670 6479 679
rect 6135 669 6172 670
rect 6191 618 6227 670
rect 6246 669 6283 670
rect 6342 669 6379 670
rect 5662 616 5703 617
rect 4469 594 5118 600
rect 5554 609 5703 616
rect 4469 593 5117 594
rect 5080 591 5117 593
rect 5554 589 5672 609
rect 5692 589 5703 609
rect 5554 581 5703 589
rect 5770 613 6129 617
rect 5770 608 6092 613
rect 5770 584 5883 608
rect 5907 589 6092 608
rect 6116 589 6129 613
rect 5907 584 6129 589
rect 5770 581 6129 584
rect 6191 581 6226 618
rect 6294 615 6394 618
rect 6294 611 6361 615
rect 6294 585 6306 611
rect 6332 589 6361 611
rect 6387 589 6394 615
rect 6332 585 6394 589
rect 6294 581 6394 585
rect 5770 560 5801 581
rect 6191 560 6227 581
rect 5434 551 5471 560
rect 5613 559 5650 560
rect 5434 533 5443 551
rect 5461 533 5471 551
rect 5083 527 5120 529
rect 1029 511 1197 513
rect 753 485 1197 511
rect 754 459 778 485
rect 1029 484 1197 485
rect 5078 519 5120 527
rect 5434 523 5471 533
rect 5078 501 5092 519
rect 5110 501 5120 519
rect 5078 492 5120 501
rect 747 451 787 459
rect 747 444 756 451
rect 152 429 756 444
rect 779 429 787 451
rect 152 426 787 429
rect 152 420 190 426
rect 747 414 787 426
rect 5078 451 5119 492
rect 5435 488 5471 523
rect 5612 550 5650 559
rect 5612 530 5621 550
rect 5641 530 5650 550
rect 5612 522 5650 530
rect 5716 554 5801 560
rect 5826 559 5863 560
rect 5716 534 5724 554
rect 5744 534 5801 554
rect 5716 526 5801 534
rect 5825 550 5863 559
rect 5825 530 5834 550
rect 5854 530 5863 550
rect 5716 525 5752 526
rect 5825 522 5863 530
rect 5929 554 6014 560
rect 6034 559 6071 560
rect 5929 534 5937 554
rect 5957 553 6014 554
rect 5957 534 5986 553
rect 5929 533 5986 534
rect 6007 533 6014 553
rect 5929 526 6014 533
rect 6033 550 6071 559
rect 6033 530 6042 550
rect 6062 530 6071 550
rect 5929 525 5965 526
rect 6033 522 6071 530
rect 6137 554 6281 560
rect 6137 534 6145 554
rect 6165 553 6253 554
rect 6165 534 6193 553
rect 6137 532 6193 534
rect 6215 534 6253 553
rect 6273 534 6281 554
rect 6215 532 6281 534
rect 6137 526 6281 532
rect 6137 525 6173 526
rect 6245 525 6281 526
rect 6347 559 6384 560
rect 6347 558 6385 559
rect 6347 550 6411 558
rect 6347 530 6356 550
rect 6376 536 6411 550
rect 6431 536 6434 556
rect 6376 531 6434 536
rect 6376 530 6411 531
rect 5613 493 5650 522
rect 5078 429 5089 451
rect 5112 429 5119 451
rect 5078 424 5119 429
rect 5433 423 5471 488
rect 5614 491 5650 493
rect 5826 491 5863 522
rect 5614 469 5863 491
rect 6034 490 6071 522
rect 6347 518 6411 530
rect 6451 492 6478 670
rect 9447 643 9484 644
rect 9750 643 9787 713
rect 9812 733 9899 740
rect 9812 730 9870 733
rect 9812 710 9817 730
rect 9838 713 9870 730
rect 9890 713 9899 733
rect 9838 710 9899 713
rect 9812 703 9899 710
rect 9958 733 9995 743
rect 9958 713 9966 733
rect 9986 713 9995 733
rect 9812 702 9843 703
rect 9446 642 9787 643
rect 9371 637 9787 642
rect 9371 617 9374 637
rect 9394 617 9787 637
rect 9958 642 9995 713
rect 10025 742 10056 795
rect 10363 793 10373 811
rect 10391 793 10402 811
rect 10363 784 10400 793
rect 10075 742 10112 743
rect 10025 733 10112 742
rect 10025 713 10083 733
rect 10103 713 10112 733
rect 10025 703 10112 713
rect 10171 733 10208 743
rect 10171 713 10179 733
rect 10199 713 10208 733
rect 10366 718 10403 722
rect 10025 702 10056 703
rect 10171 642 10208 713
rect 9958 618 10208 642
rect 10364 712 10403 718
rect 10364 694 10375 712
rect 10393 694 10403 712
rect 10364 685 10403 694
rect 9750 594 9787 617
rect 10364 607 10399 685
rect 10361 597 10399 607
rect 9750 593 9920 594
rect 10361 593 10371 597
rect 9750 579 10371 593
rect 10389 579 10399 597
rect 9750 573 10399 579
rect 9750 572 10398 573
rect 10361 570 10398 572
rect 10364 506 10401 508
rect 6310 490 6478 492
rect 6034 464 6478 490
rect 6035 438 6059 464
rect 6310 463 6478 464
rect 10359 498 10401 506
rect 10359 480 10373 498
rect 10391 480 10401 498
rect 10359 471 10401 480
rect 6028 430 6068 438
rect 6028 423 6037 430
rect 5433 408 6037 423
rect 6060 408 6068 430
rect 5433 405 6068 408
rect 5433 399 5471 405
rect 6028 393 6068 405
rect 10359 430 10400 471
rect 10359 408 10370 430
rect 10393 408 10400 430
rect 10359 403 10400 408
rect 1740 310 1990 334
rect 1740 239 1777 310
rect 1892 249 1923 250
rect 1740 219 1749 239
rect 1769 219 1777 239
rect 1740 209 1777 219
rect 1836 239 1923 249
rect 1836 219 1845 239
rect 1865 219 1923 239
rect 1836 210 1923 219
rect 1836 209 1873 210
rect 1892 157 1923 210
rect 1953 239 1990 310
rect 2161 315 2554 335
rect 2574 315 2577 335
rect 2161 310 2577 315
rect 2161 309 2502 310
rect 2105 249 2136 250
rect 1953 219 1962 239
rect 1982 219 1990 239
rect 1953 209 1990 219
rect 2049 242 2136 249
rect 2049 239 2110 242
rect 2049 219 2058 239
rect 2078 222 2110 239
rect 2131 222 2136 242
rect 2078 219 2136 222
rect 2049 212 2136 219
rect 2161 239 2198 309
rect 2464 308 2501 309
rect 7021 289 7271 313
rect 2313 249 2349 250
rect 2161 219 2170 239
rect 2190 219 2198 239
rect 2049 210 2105 212
rect 2049 209 2086 210
rect 2161 209 2198 219
rect 2257 239 2405 249
rect 2505 246 2601 248
rect 2257 219 2266 239
rect 2286 219 2376 239
rect 2396 219 2405 239
rect 2257 210 2405 219
rect 2463 245 2601 246
rect 2463 240 2687 245
rect 2463 239 2651 240
rect 2463 219 2472 239
rect 2492 220 2651 239
rect 2679 220 2687 240
rect 2492 219 2687 220
rect 2463 212 2687 219
rect 4830 222 5080 246
rect 2463 210 2601 212
rect 2257 209 2294 210
rect 2313 158 2349 210
rect 2368 209 2405 210
rect 2464 209 2501 210
rect 1784 156 1825 157
rect 1676 149 1825 156
rect 1676 129 1794 149
rect 1814 129 1825 149
rect 1676 121 1825 129
rect 1892 153 2251 157
rect 1892 148 2214 153
rect 1892 124 2005 148
rect 2029 129 2214 148
rect 2238 129 2251 153
rect 2029 124 2251 129
rect 1892 121 2251 124
rect 2313 121 2348 158
rect 2416 155 2516 158
rect 2416 151 2483 155
rect 2416 125 2428 151
rect 2454 129 2483 151
rect 2509 129 2516 155
rect 2454 125 2516 129
rect 2416 121 2516 125
rect 1892 100 1923 121
rect 2313 100 2349 121
rect 1735 99 1772 100
rect 1734 90 1772 99
rect 1734 70 1743 90
rect 1763 70 1772 90
rect 1734 62 1772 70
rect 1838 94 1923 100
rect 1948 99 1985 100
rect 1838 74 1846 94
rect 1866 74 1923 94
rect 1838 66 1923 74
rect 1947 90 1985 99
rect 1947 70 1956 90
rect 1976 70 1985 90
rect 1838 65 1874 66
rect 1947 62 1985 70
rect 2051 94 2136 100
rect 2156 99 2193 100
rect 2051 74 2059 94
rect 2079 93 2136 94
rect 2079 74 2108 93
rect 2051 73 2108 74
rect 2129 73 2136 93
rect 2051 66 2136 73
rect 2155 90 2193 99
rect 2155 70 2164 90
rect 2184 70 2193 90
rect 2051 65 2087 66
rect 2155 62 2193 70
rect 2259 94 2403 100
rect 2259 74 2267 94
rect 2287 93 2375 94
rect 2287 74 2322 93
rect 2259 71 2322 74
rect 2347 74 2375 93
rect 2395 74 2403 94
rect 2347 71 2403 74
rect 2259 66 2403 71
rect 2259 65 2295 66
rect 2367 65 2403 66
rect 2469 99 2506 100
rect 2469 98 2507 99
rect 2469 90 2533 98
rect 2469 70 2478 90
rect 2498 76 2533 90
rect 2553 76 2556 96
rect 2498 71 2556 76
rect 2498 70 2533 71
rect 1735 33 1772 62
rect 1736 31 1772 33
rect 1948 31 1985 62
rect 1736 9 1985 31
rect 2156 30 2193 62
rect 2469 58 2533 70
rect 2573 32 2600 210
rect 4830 151 4867 222
rect 4982 161 5013 162
rect 4830 131 4839 151
rect 4859 131 4867 151
rect 4830 121 4867 131
rect 4926 151 5013 161
rect 4926 131 4935 151
rect 4955 131 5013 151
rect 4926 122 5013 131
rect 4926 121 4963 122
rect 4982 69 5013 122
rect 5043 151 5080 222
rect 5251 227 5644 247
rect 5664 227 5667 247
rect 5251 222 5667 227
rect 5251 221 5592 222
rect 5195 161 5226 162
rect 5043 131 5052 151
rect 5072 131 5080 151
rect 5043 121 5080 131
rect 5139 154 5226 161
rect 5139 151 5200 154
rect 5139 131 5148 151
rect 5168 134 5200 151
rect 5221 134 5226 154
rect 5168 131 5226 134
rect 5139 124 5226 131
rect 5251 151 5288 221
rect 5554 220 5591 221
rect 7021 218 7058 289
rect 7173 228 7204 229
rect 7021 198 7030 218
rect 7050 198 7058 218
rect 7021 188 7058 198
rect 7117 218 7204 228
rect 7117 198 7126 218
rect 7146 198 7204 218
rect 7117 189 7204 198
rect 7117 188 7154 189
rect 5403 161 5439 162
rect 5251 131 5260 151
rect 5280 131 5288 151
rect 5139 122 5195 124
rect 5139 121 5176 122
rect 5251 121 5288 131
rect 5347 151 5495 161
rect 5595 158 5691 160
rect 5347 131 5356 151
rect 5376 131 5466 151
rect 5486 131 5495 151
rect 5347 122 5495 131
rect 5553 151 5691 158
rect 5553 131 5562 151
rect 5582 131 5691 151
rect 7173 136 7204 189
rect 7234 218 7271 289
rect 7442 294 7835 314
rect 7855 294 7858 314
rect 7442 289 7858 294
rect 7442 288 7783 289
rect 7386 228 7417 229
rect 7234 198 7243 218
rect 7263 198 7271 218
rect 7234 188 7271 198
rect 7330 221 7417 228
rect 7330 218 7391 221
rect 7330 198 7339 218
rect 7359 201 7391 218
rect 7412 201 7417 221
rect 7359 198 7417 201
rect 7330 191 7417 198
rect 7442 218 7479 288
rect 7745 287 7782 288
rect 7594 228 7630 229
rect 7442 198 7451 218
rect 7471 198 7479 218
rect 7330 189 7386 191
rect 7330 188 7367 189
rect 7442 188 7479 198
rect 7538 218 7686 228
rect 7786 225 7882 227
rect 7538 198 7547 218
rect 7567 198 7657 218
rect 7677 198 7686 218
rect 7538 189 7686 198
rect 7744 224 7882 225
rect 7744 219 7968 224
rect 7744 218 7932 219
rect 7744 198 7753 218
rect 7773 199 7932 218
rect 7960 199 7968 219
rect 7773 198 7968 199
rect 7744 191 7968 198
rect 7744 189 7882 191
rect 7538 188 7575 189
rect 7594 137 7630 189
rect 7649 188 7686 189
rect 7745 188 7782 189
rect 7065 135 7106 136
rect 5553 122 5691 131
rect 6957 128 7106 135
rect 5347 121 5384 122
rect 5403 70 5439 122
rect 5458 121 5495 122
rect 5554 121 5591 122
rect 4874 68 4915 69
rect 4766 61 4915 68
rect 4766 41 4884 61
rect 4904 41 4915 61
rect 4766 33 4915 41
rect 4982 65 5341 69
rect 4982 60 5304 65
rect 4982 36 5095 60
rect 5119 41 5304 60
rect 5328 41 5341 65
rect 5119 36 5341 41
rect 4982 33 5341 36
rect 5403 33 5438 70
rect 5506 67 5606 70
rect 5506 63 5573 67
rect 5506 37 5518 63
rect 5544 41 5573 63
rect 5599 41 5606 67
rect 5544 37 5606 41
rect 5506 33 5606 37
rect 2432 30 2600 32
rect 2156 4 2600 30
rect 4982 12 5013 33
rect 5403 12 5439 33
rect 4825 11 4862 12
rect 2432 3 2600 4
rect 4824 2 4862 11
rect 4824 -18 4833 2
rect 4853 -18 4862 2
rect 4824 -26 4862 -18
rect 4928 6 5013 12
rect 5038 11 5075 12
rect 4928 -14 4936 6
rect 4956 -14 5013 6
rect 4928 -22 5013 -14
rect 5037 2 5075 11
rect 5037 -18 5046 2
rect 5066 -18 5075 2
rect 4928 -23 4964 -22
rect 5037 -26 5075 -18
rect 5141 6 5226 12
rect 5246 11 5283 12
rect 5141 -14 5149 6
rect 5169 5 5226 6
rect 5169 -14 5198 5
rect 5141 -15 5198 -14
rect 5219 -15 5226 5
rect 5141 -22 5226 -15
rect 5245 2 5283 11
rect 5245 -18 5254 2
rect 5274 -18 5283 2
rect 5141 -23 5177 -22
rect 5245 -26 5283 -18
rect 5349 6 5493 12
rect 5349 -14 5357 6
rect 5377 2 5465 6
rect 5377 -14 5409 2
rect 5349 -15 5409 -14
rect 5430 -14 5465 2
rect 5485 -14 5493 6
rect 5430 -15 5493 -14
rect 5349 -22 5493 -15
rect 5349 -23 5385 -22
rect 5457 -23 5493 -22
rect 5559 11 5596 12
rect 5559 10 5597 11
rect 5559 2 5623 10
rect 5559 -18 5568 2
rect 5588 -12 5623 2
rect 5643 -12 5646 8
rect 5588 -17 5646 -12
rect 5588 -18 5623 -17
rect 4825 -55 4862 -26
rect 4826 -57 4862 -55
rect 5038 -57 5075 -26
rect 4826 -79 5075 -57
rect 5246 -58 5283 -26
rect 5559 -30 5623 -18
rect 5663 -56 5690 122
rect 6957 108 7075 128
rect 7095 108 7106 128
rect 6957 100 7106 108
rect 7173 132 7532 136
rect 7173 127 7495 132
rect 7173 103 7286 127
rect 7310 108 7495 127
rect 7519 108 7532 132
rect 7310 103 7532 108
rect 7173 100 7532 103
rect 7594 100 7629 137
rect 7697 134 7797 137
rect 7697 130 7764 134
rect 7697 104 7709 130
rect 7735 108 7764 130
rect 7790 108 7797 134
rect 7735 104 7797 108
rect 7697 100 7797 104
rect 7173 79 7204 100
rect 7594 79 7630 100
rect 7016 78 7053 79
rect 7015 69 7053 78
rect 7015 49 7024 69
rect 7044 49 7053 69
rect 7015 41 7053 49
rect 7119 73 7204 79
rect 7229 78 7266 79
rect 7119 53 7127 73
rect 7147 53 7204 73
rect 7119 45 7204 53
rect 7228 69 7266 78
rect 7228 49 7237 69
rect 7257 49 7266 69
rect 7119 44 7155 45
rect 7228 41 7266 49
rect 7332 73 7417 79
rect 7437 78 7474 79
rect 7332 53 7340 73
rect 7360 72 7417 73
rect 7360 53 7389 72
rect 7332 52 7389 53
rect 7410 52 7417 72
rect 7332 45 7417 52
rect 7436 69 7474 78
rect 7436 49 7445 69
rect 7465 49 7474 69
rect 7332 44 7368 45
rect 7436 41 7474 49
rect 7540 73 7684 79
rect 7540 53 7548 73
rect 7568 72 7656 73
rect 7568 53 7603 72
rect 7540 50 7603 53
rect 7628 53 7656 72
rect 7676 53 7684 73
rect 7628 50 7684 53
rect 7540 45 7684 50
rect 7540 44 7576 45
rect 7648 44 7684 45
rect 7750 78 7787 79
rect 7750 77 7788 78
rect 7750 69 7814 77
rect 7750 49 7759 69
rect 7779 55 7814 69
rect 7834 55 7837 75
rect 7779 50 7837 55
rect 7779 49 7814 50
rect 7016 12 7053 41
rect 7017 10 7053 12
rect 7229 10 7266 41
rect 7017 -12 7266 10
rect 7437 9 7474 41
rect 7750 37 7814 49
rect 7854 33 7881 189
rect 7851 10 7882 33
rect 7579 9 7882 10
rect 7437 -16 7882 9
rect 7437 -17 7622 -16
rect 5522 -58 5690 -56
rect 5246 -65 5690 -58
rect 5246 -82 5659 -65
rect 5683 -82 5690 -65
rect 5246 -84 5690 -82
rect 5522 -85 5690 -84
<< viali >>
rect 1115 8069 1135 8089
rect 671 7976 692 7996
rect 4078 8150 4098 8170
rect 4294 8153 4316 8174
rect 4502 8153 4523 8173
rect 4122 8091 4148 8117
rect 2973 7983 2992 8009
rect 1044 7883 1070 7909
rect 669 7827 690 7847
rect 885 7828 907 7849
rect 1094 7830 1114 7850
rect 2127 7888 2147 7908
rect 1683 7795 1704 7815
rect 2056 7702 2082 7728
rect 1114 7654 1134 7674
rect 670 7561 691 7581
rect 1681 7646 1702 7666
rect 1892 7647 1916 7667
rect 2106 7649 2126 7669
rect 1778 7580 1798 7599
rect 2880 7567 2900 7585
rect 3393 7986 3413 8005
rect 3065 7916 3085 7936
rect 3276 7917 3300 7937
rect 3489 7919 3510 7939
rect 4500 8004 4521 8024
rect 4057 7911 4077 7931
rect 3109 7857 3135 7883
rect 3487 7770 3508 7790
rect 3044 7677 3064 7697
rect 6396 8048 6416 8068
rect 5952 7955 5973 7975
rect 9359 8129 9379 8149
rect 9575 8132 9597 8153
rect 9783 8132 9804 8152
rect 9403 8070 9429 8096
rect 8254 7962 8273 7988
rect 4077 7735 4097 7755
rect 4284 7736 4306 7757
rect 4501 7738 4522 7758
rect 4121 7676 4147 7702
rect 6325 7862 6351 7888
rect 5950 7806 5971 7826
rect 6166 7807 6188 7828
rect 6375 7809 6395 7829
rect 1043 7468 1069 7494
rect 668 7412 689 7432
rect 875 7411 897 7432
rect 1093 7415 1113 7435
rect 2182 7327 2202 7347
rect 1738 7234 1759 7254
rect 2111 7141 2137 7167
rect 1120 7088 1140 7108
rect 676 6995 697 7015
rect 1736 7085 1757 7105
rect 1951 7087 1975 7104
rect 2161 7088 2181 7108
rect 1049 6902 1075 6928
rect 674 6846 695 6866
rect 890 6847 912 6868
rect 1099 6849 1119 6869
rect 2132 6907 2152 6927
rect 1688 6814 1709 6834
rect 2061 6721 2087 6747
rect 1119 6673 1139 6693
rect 675 6580 696 6600
rect 1686 6665 1707 6685
rect 1896 6667 1920 6687
rect 2111 6668 2131 6688
rect 1783 6599 1803 6618
rect 2204 6595 2223 6621
rect 1048 6487 1074 6513
rect 673 6431 694 6451
rect 880 6430 902 6451
rect 1098 6434 1118 6454
rect 3015 7496 3035 7516
rect 3225 7499 3248 7518
rect 3439 7499 3460 7519
rect 4499 7589 4520 7609
rect 4056 7496 4076 7516
rect 7408 7867 7428 7887
rect 6964 7774 6985 7794
rect 7337 7681 7363 7707
rect 3059 7437 3085 7463
rect 6395 7633 6415 7653
rect 5951 7540 5972 7560
rect 6962 7625 6983 7645
rect 7173 7626 7197 7646
rect 7387 7628 7407 7648
rect 7059 7559 7079 7578
rect 8161 7546 8181 7564
rect 8674 7965 8694 7984
rect 8346 7895 8366 7915
rect 8557 7896 8581 7916
rect 8770 7898 8791 7918
rect 9781 7983 9802 8003
rect 9338 7890 9358 7910
rect 8390 7836 8416 7862
rect 8768 7749 8789 7769
rect 8325 7656 8345 7676
rect 9358 7714 9378 7734
rect 9565 7715 9587 7736
rect 9782 7717 9803 7737
rect 9402 7655 9428 7681
rect 6324 7447 6350 7473
rect 3437 7350 3458 7370
rect 2994 7257 3014 7277
rect 5949 7391 5970 7411
rect 6156 7390 6178 7411
rect 6374 7394 6394 7414
rect 4083 7169 4103 7189
rect 4299 7172 4321 7193
rect 4507 7172 4528 7192
rect 7463 7306 7483 7326
rect 7019 7213 7040 7233
rect 4127 7110 4153 7136
rect 3398 7005 3418 7024
rect 3070 6935 3090 6955
rect 3280 6937 3304 6957
rect 3494 6938 3515 6958
rect 4505 7023 4526 7043
rect 4062 6930 4082 6950
rect 7392 7120 7418 7146
rect 3114 6876 3140 6902
rect 3492 6789 3513 6809
rect 3049 6696 3069 6716
rect 6401 7067 6421 7087
rect 5957 6974 5978 6994
rect 7017 7064 7038 7084
rect 7232 7066 7256 7083
rect 7442 7067 7462 7087
rect 4082 6754 4102 6774
rect 4289 6755 4311 6776
rect 4506 6757 4527 6777
rect 4126 6695 4152 6721
rect 6330 6881 6356 6907
rect 5955 6825 5976 6845
rect 6171 6826 6193 6847
rect 6380 6828 6400 6848
rect 2757 6538 2780 6557
rect 2347 6395 2367 6415
rect 1903 6302 1924 6322
rect 2276 6209 2302 6235
rect 1901 6153 1922 6173
rect 2110 6152 2135 6178
rect 2326 6156 2346 6176
rect 1127 6109 1147 6129
rect 683 6016 704 6036
rect 1056 5923 1082 5949
rect 681 5867 702 5887
rect 897 5868 919 5889
rect 1106 5870 1126 5890
rect 2139 5928 2159 5948
rect 1695 5835 1716 5855
rect 2068 5742 2094 5768
rect 1126 5694 1146 5714
rect 682 5601 703 5621
rect 1693 5686 1714 5706
rect 1904 5687 1928 5707
rect 2118 5689 2138 5709
rect 1790 5620 1810 5639
rect 1055 5508 1081 5534
rect 680 5452 701 5472
rect 887 5451 909 5472
rect 1105 5455 1125 5475
rect 2194 5367 2214 5387
rect 1750 5274 1771 5294
rect 2123 5181 2149 5207
rect 1132 5128 1152 5148
rect 688 5035 709 5055
rect 1748 5125 1769 5145
rect 1960 5126 1983 5145
rect 2173 5128 2193 5148
rect 1061 4942 1087 4968
rect 686 4886 707 4906
rect 902 4887 924 4908
rect 1111 4889 1131 4909
rect 2144 4947 2164 4967
rect 1700 4854 1721 4874
rect 2073 4761 2099 4787
rect 1131 4713 1151 4733
rect 687 4620 708 4640
rect 1698 4705 1719 4725
rect 1908 4707 1932 4727
rect 2123 4708 2143 4728
rect 1795 4639 1815 4658
rect 2308 5059 2328 5077
rect 2216 4635 2235 4661
rect 4504 6608 4525 6628
rect 4061 6515 4081 6535
rect 7413 6886 7433 6906
rect 6969 6793 6990 6813
rect 7342 6700 7368 6726
rect 2862 6468 2882 6488
rect 3069 6470 3092 6489
rect 3286 6471 3307 6491
rect 6400 6652 6420 6672
rect 5956 6559 5977 6579
rect 6967 6644 6988 6664
rect 7177 6646 7201 6666
rect 7392 6647 7412 6667
rect 7064 6578 7084 6597
rect 7485 6574 7504 6600
rect 6329 6466 6355 6492
rect 2906 6409 2932 6435
rect 3284 6322 3305 6342
rect 2841 6229 2861 6249
rect 5954 6410 5975 6430
rect 6161 6409 6183 6430
rect 6379 6413 6399 6433
rect 8296 7475 8316 7495
rect 8506 7478 8529 7497
rect 8720 7478 8741 7498
rect 9780 7568 9801 7588
rect 9337 7475 9357 7495
rect 8340 7416 8366 7442
rect 8718 7329 8739 7349
rect 8275 7236 8295 7256
rect 9364 7148 9384 7168
rect 9580 7151 9602 7172
rect 9788 7151 9809 7171
rect 9408 7089 9434 7115
rect 8679 6984 8699 7003
rect 8351 6914 8371 6934
rect 8561 6916 8585 6936
rect 8775 6917 8796 6937
rect 9786 7002 9807 7022
rect 9343 6909 9363 6929
rect 8395 6855 8421 6881
rect 8773 6768 8794 6788
rect 8330 6675 8350 6695
rect 9363 6733 9383 6753
rect 9570 6734 9592 6755
rect 9787 6736 9808 6756
rect 9407 6674 9433 6700
rect 8038 6517 8061 6536
rect 4090 6190 4110 6210
rect 4306 6193 4328 6214
rect 4514 6193 4535 6213
rect 7628 6374 7648 6394
rect 7184 6281 7205 6301
rect 7557 6188 7583 6214
rect 4134 6131 4160 6157
rect 2985 6023 3004 6049
rect 3405 6026 3425 6045
rect 3077 5956 3097 5976
rect 3288 5957 3312 5977
rect 3501 5959 3522 5979
rect 4512 6044 4533 6064
rect 4069 5951 4089 5971
rect 7182 6132 7203 6152
rect 7391 6131 7416 6157
rect 7607 6135 7627 6155
rect 3121 5897 3147 5923
rect 3499 5810 3520 5830
rect 3056 5717 3076 5737
rect 6408 6088 6428 6108
rect 5964 5995 5985 6015
rect 4089 5775 4109 5795
rect 4296 5776 4318 5797
rect 4513 5778 4534 5798
rect 4133 5716 4159 5742
rect 6337 5902 6363 5928
rect 5962 5846 5983 5866
rect 6178 5847 6200 5868
rect 6387 5849 6407 5869
rect 3027 5536 3047 5556
rect 3233 5540 3257 5557
rect 3451 5539 3472 5559
rect 4511 5629 4532 5649
rect 4068 5536 4088 5556
rect 7420 5907 7440 5927
rect 6976 5814 6997 5834
rect 7349 5721 7375 5747
rect 3071 5477 3097 5503
rect 6407 5673 6427 5693
rect 5963 5580 5984 5600
rect 6974 5665 6995 5685
rect 7185 5666 7209 5686
rect 7399 5668 7419 5688
rect 7071 5599 7091 5618
rect 6336 5487 6362 5513
rect 3449 5390 3470 5410
rect 3006 5297 3026 5317
rect 5961 5431 5982 5451
rect 6168 5430 6190 5451
rect 6386 5434 6406 5454
rect 4095 5209 4115 5229
rect 4311 5212 4333 5233
rect 4519 5212 4540 5232
rect 7475 5346 7495 5366
rect 7031 5253 7052 5273
rect 4139 5150 4165 5176
rect 3410 5045 3430 5064
rect 3082 4975 3102 4995
rect 3292 4977 3316 4997
rect 3506 4978 3527 4998
rect 4517 5063 4538 5083
rect 4074 4970 4094 4990
rect 7404 5160 7430 5186
rect 3126 4916 3152 4942
rect 3504 4829 3525 4849
rect 3061 4736 3081 4756
rect 6413 5107 6433 5127
rect 5969 5014 5990 5034
rect 7029 5104 7050 5124
rect 7241 5105 7264 5124
rect 7454 5107 7474 5127
rect 4094 4794 4114 4814
rect 4301 4795 4323 4816
rect 4518 4797 4539 4817
rect 4138 4735 4164 4761
rect 6342 4921 6368 4947
rect 5967 4865 5988 4885
rect 6183 4866 6205 4887
rect 6392 4868 6412 4888
rect 1060 4527 1086 4553
rect 685 4471 706 4491
rect 892 4470 914 4491
rect 1110 4474 1130 4494
rect 4516 4648 4537 4668
rect 2787 4543 2807 4563
rect 2991 4544 3017 4563
rect 3211 4546 3232 4566
rect 4073 4555 4093 4575
rect 7425 4926 7445 4946
rect 6981 4833 7002 4853
rect 7354 4740 7380 4766
rect 2831 4484 2857 4510
rect 6412 4692 6432 4712
rect 5968 4599 5989 4619
rect 6979 4684 7000 4704
rect 7189 4686 7213 4706
rect 7404 4687 7424 4707
rect 7076 4618 7096 4637
rect 7589 5038 7609 5056
rect 7497 4614 7516 4640
rect 9785 6587 9806 6607
rect 9342 6494 9362 6514
rect 8143 6447 8163 6467
rect 8350 6449 8373 6468
rect 8567 6450 8588 6470
rect 8187 6388 8213 6414
rect 8565 6301 8586 6321
rect 8122 6208 8142 6228
rect 9371 6169 9391 6189
rect 9587 6172 9609 6193
rect 9795 6172 9816 6192
rect 9415 6110 9441 6136
rect 8266 6002 8285 6028
rect 8686 6005 8706 6024
rect 8358 5935 8378 5955
rect 8569 5936 8593 5956
rect 8782 5938 8803 5958
rect 9793 6023 9814 6043
rect 9350 5930 9370 5950
rect 8402 5876 8428 5902
rect 8780 5789 8801 5809
rect 8337 5696 8357 5716
rect 9370 5754 9390 5774
rect 9577 5755 9599 5776
rect 9794 5757 9815 5777
rect 9414 5695 9440 5721
rect 8308 5515 8328 5535
rect 8514 5519 8538 5536
rect 8732 5518 8753 5538
rect 9792 5608 9813 5628
rect 9349 5515 9369 5535
rect 8352 5456 8378 5482
rect 8730 5369 8751 5389
rect 8287 5276 8307 5296
rect 9376 5188 9396 5208
rect 9592 5191 9614 5212
rect 9800 5191 9821 5211
rect 9420 5129 9446 5155
rect 8691 5024 8711 5043
rect 8363 4954 8383 4974
rect 8573 4956 8597 4976
rect 8787 4957 8808 4977
rect 9798 5042 9819 5062
rect 9355 4949 9375 4969
rect 8407 4895 8433 4921
rect 8785 4808 8806 4828
rect 8342 4715 8362 4735
rect 9375 4773 9395 4793
rect 9582 4774 9604 4795
rect 9799 4776 9820 4796
rect 9419 4714 9445 4740
rect 6341 4506 6367 4532
rect 2442 4403 2462 4423
rect 1998 4310 2019 4330
rect 3209 4397 3230 4417
rect 2766 4304 2786 4324
rect 5966 4450 5987 4470
rect 6173 4449 6195 4470
rect 6391 4453 6411 4473
rect 9797 4627 9818 4647
rect 8068 4522 8088 4542
rect 8272 4523 8298 4542
rect 8492 4525 8513 4545
rect 9354 4534 9374 4554
rect 8112 4463 8138 4489
rect 2371 4217 2397 4243
rect 1135 4152 1155 4172
rect 1996 4161 2017 4181
rect 2211 4164 2237 4183
rect 2421 4164 2441 4184
rect 691 4059 712 4079
rect 4098 4233 4118 4253
rect 4314 4236 4336 4257
rect 4522 4236 4543 4256
rect 7723 4382 7743 4402
rect 7279 4289 7300 4309
rect 8490 4376 8511 4396
rect 8047 4283 8067 4303
rect 4142 4174 4168 4200
rect 1064 3966 1090 3992
rect 689 3910 710 3930
rect 905 3911 927 3932
rect 1114 3913 1134 3933
rect 2147 3971 2167 3991
rect 1703 3878 1724 3898
rect 2076 3785 2102 3811
rect 1134 3737 1154 3757
rect 690 3644 711 3664
rect 1701 3729 1722 3749
rect 1912 3730 1936 3750
rect 2126 3732 2146 3752
rect 1798 3663 1818 3682
rect 1063 3551 1089 3577
rect 688 3495 709 3515
rect 895 3494 917 3515
rect 1113 3498 1133 3518
rect 2202 3410 2222 3430
rect 1758 3317 1779 3337
rect 2131 3224 2157 3250
rect 1140 3171 1160 3191
rect 696 3078 717 3098
rect 1756 3168 1777 3188
rect 1971 3170 1995 3187
rect 2181 3171 2201 3191
rect 1069 2985 1095 3011
rect 694 2929 715 2949
rect 910 2930 932 2951
rect 1119 2932 1139 2952
rect 2152 2990 2172 3010
rect 1708 2897 1729 2917
rect 2081 2804 2107 2830
rect 1139 2756 1159 2776
rect 695 2663 716 2683
rect 1706 2748 1727 2768
rect 1916 2750 1940 2770
rect 2131 2751 2151 2771
rect 1803 2682 1823 2701
rect 2224 2678 2243 2704
rect 1068 2570 1094 2596
rect 693 2514 714 2534
rect 900 2513 922 2534
rect 1118 2517 1138 2537
rect 2367 2478 2387 2498
rect 1923 2385 1944 2405
rect 2296 2292 2322 2318
rect 1921 2236 1942 2256
rect 2136 2238 2159 2257
rect 2346 2239 2366 2259
rect 1147 2192 1167 2212
rect 703 2099 724 2119
rect 2993 4066 3012 4092
rect 2900 3650 2920 3668
rect 3413 4069 3433 4088
rect 3085 3999 3105 4019
rect 3296 4000 3320 4020
rect 3509 4002 3530 4022
rect 4520 4087 4541 4107
rect 4077 3994 4097 4014
rect 7652 4196 7678 4222
rect 3129 3940 3155 3966
rect 3507 3853 3528 3873
rect 3064 3760 3084 3780
rect 6416 4131 6436 4151
rect 7277 4140 7298 4160
rect 7492 4143 7518 4162
rect 7702 4143 7722 4163
rect 5972 4038 5993 4058
rect 9379 4212 9399 4232
rect 9595 4215 9617 4236
rect 9803 4215 9824 4235
rect 9423 4153 9449 4179
rect 4097 3818 4117 3838
rect 4304 3819 4326 3840
rect 4521 3821 4542 3841
rect 4141 3759 4167 3785
rect 6345 3945 6371 3971
rect 5970 3889 5991 3909
rect 6186 3890 6208 3911
rect 6395 3892 6415 3912
rect 3035 3579 3055 3599
rect 3245 3582 3268 3601
rect 3459 3582 3480 3602
rect 4519 3672 4540 3692
rect 4076 3579 4096 3599
rect 7428 3950 7448 3970
rect 6984 3857 7005 3877
rect 7357 3764 7383 3790
rect 3079 3520 3105 3546
rect 6415 3716 6435 3736
rect 5971 3623 5992 3643
rect 6982 3708 7003 3728
rect 7193 3709 7217 3729
rect 7407 3711 7427 3731
rect 7079 3642 7099 3661
rect 6344 3530 6370 3556
rect 3457 3433 3478 3453
rect 3014 3340 3034 3360
rect 5969 3474 5990 3494
rect 6176 3473 6198 3494
rect 6394 3477 6414 3497
rect 4103 3252 4123 3272
rect 4319 3255 4341 3276
rect 4527 3255 4548 3275
rect 7483 3389 7503 3409
rect 7039 3296 7060 3316
rect 4147 3193 4173 3219
rect 3418 3088 3438 3107
rect 3090 3018 3110 3038
rect 3300 3020 3324 3040
rect 3514 3021 3535 3041
rect 4525 3106 4546 3126
rect 4082 3013 4102 3033
rect 7412 3203 7438 3229
rect 3134 2959 3160 2985
rect 3512 2872 3533 2892
rect 3069 2779 3089 2799
rect 6421 3150 6441 3170
rect 5977 3057 5998 3077
rect 7037 3147 7058 3167
rect 7252 3149 7276 3166
rect 7462 3150 7482 3170
rect 4102 2837 4122 2857
rect 4309 2838 4331 2859
rect 4526 2840 4547 2860
rect 4146 2778 4172 2804
rect 6350 2964 6376 2990
rect 5975 2908 5996 2928
rect 6191 2909 6213 2930
rect 6400 2911 6420 2931
rect 4524 2691 4545 2711
rect 4081 2598 4101 2618
rect 7433 2969 7453 2989
rect 6989 2876 7010 2896
rect 7362 2783 7388 2809
rect 2882 2551 2902 2571
rect 3093 2549 3118 2575
rect 3306 2554 3327 2574
rect 6420 2735 6440 2755
rect 5976 2642 5997 2662
rect 6987 2727 7008 2747
rect 7197 2729 7221 2749
rect 7412 2730 7432 2750
rect 7084 2661 7104 2680
rect 7505 2657 7524 2683
rect 6349 2549 6375 2575
rect 2926 2492 2952 2518
rect 3304 2405 3325 2425
rect 2861 2312 2881 2332
rect 5974 2493 5995 2513
rect 6181 2492 6203 2513
rect 6399 2496 6419 2516
rect 2448 2170 2471 2189
rect 1076 2006 1102 2032
rect 701 1950 722 1970
rect 917 1951 939 1972
rect 1126 1953 1146 1973
rect 2159 2011 2179 2031
rect 1715 1918 1736 1938
rect 2088 1825 2114 1851
rect 1146 1777 1166 1797
rect 702 1684 723 1704
rect 1713 1769 1734 1789
rect 1924 1770 1948 1790
rect 2138 1772 2158 1792
rect 1810 1703 1830 1722
rect 1075 1591 1101 1617
rect 700 1535 721 1555
rect 907 1534 929 1555
rect 1125 1538 1145 1558
rect 2214 1450 2234 1470
rect 1770 1357 1791 1377
rect 2143 1264 2169 1290
rect 1152 1211 1172 1231
rect 708 1118 729 1138
rect 1768 1208 1789 1228
rect 1980 1209 2003 1228
rect 2193 1211 2213 1231
rect 4110 2273 4130 2293
rect 4326 2276 4348 2297
rect 4534 2276 4555 2296
rect 7648 2457 7668 2477
rect 7204 2364 7225 2384
rect 7577 2271 7603 2297
rect 4154 2214 4180 2240
rect 3005 2106 3024 2132
rect 3425 2109 3445 2128
rect 3097 2039 3117 2059
rect 3308 2040 3332 2060
rect 3521 2042 3542 2062
rect 4532 2127 4553 2147
rect 4089 2034 4109 2054
rect 7202 2215 7223 2235
rect 7417 2217 7440 2236
rect 7627 2218 7647 2238
rect 3141 1980 3167 2006
rect 3519 1893 3540 1913
rect 3076 1800 3096 1820
rect 6428 2171 6448 2191
rect 5984 2078 6005 2098
rect 8274 4045 8293 4071
rect 8181 3629 8201 3647
rect 8694 4048 8714 4067
rect 8366 3978 8386 3998
rect 8577 3979 8601 3999
rect 8790 3981 8811 4001
rect 9801 4066 9822 4086
rect 9358 3973 9378 3993
rect 8410 3919 8436 3945
rect 8788 3832 8809 3852
rect 8345 3739 8365 3759
rect 9378 3797 9398 3817
rect 9585 3798 9607 3819
rect 9802 3800 9823 3820
rect 9422 3738 9448 3764
rect 8316 3558 8336 3578
rect 8526 3561 8549 3580
rect 8740 3561 8761 3581
rect 9800 3651 9821 3671
rect 9357 3558 9377 3578
rect 8360 3499 8386 3525
rect 8738 3412 8759 3432
rect 8295 3319 8315 3339
rect 9384 3231 9404 3251
rect 9600 3234 9622 3255
rect 9808 3234 9829 3254
rect 9428 3172 9454 3198
rect 8699 3067 8719 3086
rect 8371 2997 8391 3017
rect 8581 2999 8605 3019
rect 8795 3000 8816 3020
rect 9806 3085 9827 3105
rect 9363 2992 9383 3012
rect 8415 2938 8441 2964
rect 8793 2851 8814 2871
rect 8350 2758 8370 2778
rect 9383 2816 9403 2836
rect 9590 2817 9612 2838
rect 9807 2819 9828 2839
rect 9427 2757 9453 2783
rect 9805 2670 9826 2690
rect 9362 2577 9382 2597
rect 8163 2530 8183 2550
rect 8374 2528 8399 2554
rect 8587 2533 8608 2553
rect 8207 2471 8233 2497
rect 8585 2384 8606 2404
rect 8142 2291 8162 2311
rect 7729 2149 7752 2168
rect 4109 1858 4129 1878
rect 4316 1859 4338 1880
rect 4533 1861 4554 1881
rect 4153 1799 4179 1825
rect 6357 1985 6383 2011
rect 5982 1929 6003 1949
rect 6198 1930 6220 1951
rect 6407 1932 6427 1952
rect 3047 1619 3067 1639
rect 3253 1623 3277 1640
rect 3471 1622 3492 1642
rect 4531 1712 4552 1732
rect 4088 1619 4108 1639
rect 7440 1990 7460 2010
rect 6996 1897 7017 1917
rect 7369 1804 7395 1830
rect 3091 1560 3117 1586
rect 6427 1756 6447 1776
rect 5983 1663 6004 1683
rect 6994 1748 7015 1768
rect 7205 1749 7229 1769
rect 7419 1751 7439 1771
rect 7091 1682 7111 1701
rect 6356 1570 6382 1596
rect 3469 1473 3490 1493
rect 3026 1380 3046 1400
rect 5981 1514 6002 1534
rect 6188 1513 6210 1534
rect 6406 1517 6426 1537
rect 4115 1292 4135 1312
rect 4331 1295 4353 1316
rect 4539 1295 4560 1315
rect 7495 1429 7515 1449
rect 7051 1336 7072 1356
rect 4159 1233 4185 1259
rect 1081 1025 1107 1051
rect 706 969 727 989
rect 922 970 944 991
rect 1131 972 1151 992
rect 2164 1030 2184 1050
rect 1720 937 1741 957
rect 2093 844 2119 870
rect 1151 796 1171 816
rect 707 703 728 723
rect 1718 788 1739 808
rect 1928 790 1952 810
rect 2143 791 2163 811
rect 1815 722 1835 741
rect 2328 1142 2348 1160
rect 3430 1128 3450 1147
rect 3102 1058 3122 1078
rect 3312 1060 3336 1080
rect 3526 1061 3547 1081
rect 4537 1146 4558 1166
rect 4094 1053 4114 1073
rect 7424 1243 7450 1269
rect 3146 999 3172 1025
rect 3524 912 3545 932
rect 3081 819 3101 839
rect 6433 1190 6453 1210
rect 5989 1097 6010 1117
rect 7049 1187 7070 1207
rect 7261 1188 7284 1207
rect 7474 1190 7494 1210
rect 9391 2252 9411 2272
rect 9607 2255 9629 2276
rect 9815 2255 9836 2275
rect 9435 2193 9461 2219
rect 8286 2085 8305 2111
rect 8706 2088 8726 2107
rect 8378 2018 8398 2038
rect 8589 2019 8613 2039
rect 8802 2021 8823 2041
rect 9813 2106 9834 2126
rect 9370 2013 9390 2033
rect 8422 1959 8448 1985
rect 8800 1872 8821 1892
rect 8357 1779 8377 1799
rect 9390 1837 9410 1857
rect 9597 1838 9619 1859
rect 9814 1840 9835 1860
rect 9434 1778 9460 1804
rect 8328 1598 8348 1618
rect 8534 1602 8558 1619
rect 8752 1601 8773 1621
rect 9812 1691 9833 1711
rect 9369 1598 9389 1618
rect 8372 1539 8398 1565
rect 8750 1452 8771 1472
rect 8307 1359 8327 1379
rect 9396 1271 9416 1291
rect 9612 1274 9634 1295
rect 9820 1274 9841 1294
rect 9440 1212 9466 1238
rect 4114 877 4134 897
rect 4321 878 4343 899
rect 4538 880 4559 900
rect 4158 818 4184 844
rect 6362 1004 6388 1030
rect 5987 948 6008 968
rect 6203 949 6225 970
rect 6412 951 6432 971
rect 2236 718 2255 744
rect 1080 610 1106 636
rect 705 554 726 574
rect 912 553 934 574
rect 1130 557 1150 577
rect 4536 731 4557 751
rect 4093 638 4113 658
rect 7445 1009 7465 1029
rect 7001 916 7022 936
rect 7374 823 7400 849
rect 6432 775 6452 795
rect 5988 682 6009 702
rect 6999 767 7020 787
rect 7209 769 7233 789
rect 7424 770 7444 790
rect 7096 701 7116 720
rect 7609 1121 7629 1139
rect 8711 1107 8731 1126
rect 8383 1037 8403 1057
rect 8593 1039 8617 1059
rect 8807 1040 8828 1060
rect 9818 1125 9839 1145
rect 9375 1032 9395 1052
rect 8427 978 8453 1004
rect 8805 891 8826 911
rect 8362 798 8382 818
rect 9395 856 9415 876
rect 9602 857 9624 878
rect 9819 859 9840 879
rect 9439 797 9465 823
rect 7517 697 7536 723
rect 6361 589 6387 615
rect 756 429 779 451
rect 5986 533 6007 553
rect 6193 532 6215 553
rect 6411 536 6431 556
rect 5089 429 5112 451
rect 9817 710 9838 730
rect 9374 617 9394 637
rect 6037 408 6060 430
rect 10370 408 10393 430
rect 2554 315 2574 335
rect 2110 222 2131 242
rect 2651 220 2679 240
rect 2483 129 2509 155
rect 2108 73 2129 93
rect 2322 71 2347 93
rect 2533 76 2553 96
rect 5644 227 5664 247
rect 5200 134 5221 154
rect 7835 294 7855 314
rect 7391 201 7412 221
rect 7932 199 7960 219
rect 5573 41 5599 67
rect 5198 -15 5219 5
rect 5409 -15 5430 2
rect 5623 -12 5643 8
rect 7764 108 7790 134
rect 7389 52 7410 72
rect 7603 50 7628 72
rect 7814 55 7834 75
rect 5659 -82 5683 -65
<< metal1 >>
rect 3914 8244 4323 8245
rect 3908 8215 4323 8244
rect 9195 8223 9604 8224
rect 1111 8094 1143 8095
rect 1108 8089 1143 8094
rect 1108 8069 1115 8089
rect 1135 8069 1143 8089
rect 1108 8061 1143 8069
rect 3908 8064 3948 8215
rect 4282 8182 4323 8215
rect 9189 8194 9604 8223
rect 4070 8177 4105 8178
rect 664 7996 696 8003
rect 664 7976 671 7996
rect 692 7976 696 7996
rect 664 7911 696 7976
rect 1034 7911 1074 7912
rect 664 7909 1076 7911
rect 664 7883 1044 7909
rect 1070 7883 1076 7909
rect 664 7875 1076 7883
rect 664 7847 696 7875
rect 1109 7855 1143 8061
rect 3385 8036 3948 8064
rect 4049 8170 4105 8177
rect 4049 8150 4078 8170
rect 4098 8150 4105 8170
rect 4049 8145 4105 8150
rect 4278 8174 4328 8182
rect 4278 8153 4294 8174
rect 4316 8153 4328 8174
rect 2964 8009 3311 8013
rect 2964 7983 2973 8009
rect 2992 7983 3311 8009
rect 3386 8008 3420 8036
rect 2964 7978 3311 7983
rect 3385 8005 3421 8008
rect 3385 7986 3393 8005
rect 3413 7986 3421 8005
rect 3385 7982 3421 7986
rect 3271 7948 3311 7978
rect 3057 7943 3092 7944
rect 664 7827 669 7847
rect 690 7827 696 7847
rect 664 7820 696 7827
rect 873 7849 913 7854
rect 873 7828 885 7849
rect 907 7828 913 7849
rect 873 7816 913 7828
rect 1087 7850 1143 7855
rect 1087 7830 1094 7850
rect 1114 7830 1143 7850
rect 1087 7823 1143 7830
rect 1200 7924 2157 7943
rect 3036 7936 3092 7943
rect 1087 7822 1122 7823
rect 879 7784 907 7816
rect 1200 7784 1231 7924
rect 2120 7908 2155 7924
rect 2120 7888 2127 7908
rect 2147 7888 2155 7908
rect 2120 7880 2155 7888
rect 879 7753 1231 7784
rect 1676 7815 1708 7822
rect 1676 7795 1683 7815
rect 1704 7795 1708 7815
rect 1676 7730 1708 7795
rect 2046 7730 2086 7731
rect 1676 7728 2088 7730
rect 1676 7702 2056 7728
rect 2082 7702 2088 7728
rect 1676 7694 2088 7702
rect 1110 7679 1142 7680
rect 1107 7674 1142 7679
rect 1107 7654 1114 7674
rect 1134 7654 1142 7674
rect 1107 7646 1142 7654
rect 663 7581 695 7588
rect 663 7561 670 7581
rect 691 7561 695 7581
rect 663 7496 695 7561
rect 1033 7496 1073 7497
rect 663 7494 1075 7496
rect 663 7468 1043 7494
rect 1069 7468 1075 7494
rect 663 7460 1075 7468
rect 663 7432 695 7460
rect 663 7412 668 7432
rect 689 7412 695 7432
rect 663 7405 695 7412
rect 863 7432 913 7441
rect 1108 7440 1142 7646
rect 1676 7666 1708 7694
rect 1676 7646 1681 7666
rect 1702 7646 1708 7666
rect 1676 7639 1708 7646
rect 1883 7667 1925 7675
rect 2121 7674 2155 7880
rect 1883 7647 1892 7667
rect 1916 7647 1925 7667
rect 1883 7635 1925 7647
rect 2099 7669 2155 7674
rect 2099 7649 2106 7669
rect 2126 7649 2155 7669
rect 3036 7916 3065 7936
rect 3085 7916 3092 7936
rect 3036 7911 3092 7916
rect 3268 7937 3311 7948
rect 3268 7917 3276 7937
rect 3300 7931 3311 7937
rect 3483 7939 3515 7946
rect 3300 7917 3310 7931
rect 3036 7705 3070 7911
rect 3268 7908 3310 7917
rect 3483 7919 3489 7939
rect 3510 7919 3515 7939
rect 3483 7891 3515 7919
rect 4049 7939 4083 8145
rect 4278 8144 4328 8153
rect 4496 8173 4528 8180
rect 4496 8153 4502 8173
rect 4523 8153 4528 8173
rect 4496 8125 4528 8153
rect 4116 8117 4528 8125
rect 4116 8091 4122 8117
rect 4148 8091 4528 8117
rect 4116 8089 4528 8091
rect 4118 8088 4158 8089
rect 4496 8024 4528 8089
rect 6392 8073 6424 8074
rect 6389 8068 6424 8073
rect 6389 8048 6396 8068
rect 6416 8048 6424 8068
rect 6389 8040 6424 8048
rect 9189 8043 9229 8194
rect 9563 8161 9604 8194
rect 9351 8156 9386 8157
rect 4496 8004 4500 8024
rect 4521 8004 4528 8024
rect 4496 7997 4528 8004
rect 5945 7975 5977 7982
rect 5945 7955 5952 7975
rect 5973 7955 5977 7975
rect 4049 7931 4084 7939
rect 4049 7911 4057 7931
rect 4077 7911 4084 7931
rect 4049 7906 4084 7911
rect 4049 7905 4081 7906
rect 3103 7883 3515 7891
rect 3103 7857 3109 7883
rect 3135 7857 3515 7883
rect 3103 7855 3515 7857
rect 3105 7854 3145 7855
rect 3483 7790 3515 7855
rect 5945 7890 5977 7955
rect 6315 7890 6355 7891
rect 5945 7888 6357 7890
rect 5945 7862 6325 7888
rect 6351 7862 6357 7888
rect 5945 7854 6357 7862
rect 3483 7770 3487 7790
rect 3508 7770 3515 7790
rect 3483 7763 3515 7770
rect 3960 7801 4312 7832
rect 3036 7697 3071 7705
rect 3036 7677 3044 7697
rect 3064 7677 3071 7697
rect 3036 7661 3071 7677
rect 3960 7661 3991 7801
rect 4284 7769 4312 7801
rect 5945 7826 5977 7854
rect 6390 7834 6424 8040
rect 8666 8015 9229 8043
rect 9330 8149 9386 8156
rect 9330 8129 9359 8149
rect 9379 8129 9386 8149
rect 9330 8124 9386 8129
rect 9559 8153 9609 8161
rect 9559 8132 9575 8153
rect 9597 8132 9609 8153
rect 8245 7988 8592 7992
rect 8245 7962 8254 7988
rect 8273 7962 8592 7988
rect 8667 7987 8701 8015
rect 8245 7957 8592 7962
rect 8666 7984 8702 7987
rect 8666 7965 8674 7984
rect 8694 7965 8702 7984
rect 8666 7961 8702 7965
rect 8552 7927 8592 7957
rect 8338 7922 8373 7923
rect 5945 7806 5950 7826
rect 5971 7806 5977 7826
rect 5945 7799 5977 7806
rect 6154 7828 6194 7833
rect 6154 7807 6166 7828
rect 6188 7807 6194 7828
rect 6154 7795 6194 7807
rect 6368 7829 6424 7834
rect 6368 7809 6375 7829
rect 6395 7809 6424 7829
rect 6368 7802 6424 7809
rect 6481 7903 7438 7922
rect 8317 7915 8373 7922
rect 6368 7801 6403 7802
rect 4069 7762 4104 7763
rect 2099 7642 2155 7649
rect 3034 7642 3991 7661
rect 4048 7755 4104 7762
rect 4048 7735 4077 7755
rect 4097 7735 4104 7755
rect 4048 7730 4104 7735
rect 4278 7757 4318 7769
rect 4278 7736 4284 7757
rect 4306 7736 4318 7757
rect 4278 7731 4318 7736
rect 4495 7758 4527 7765
rect 4495 7738 4501 7758
rect 4522 7738 4527 7758
rect 2099 7641 2134 7642
rect 1885 7606 1920 7635
rect 1885 7605 2195 7606
rect 1770 7599 1806 7603
rect 1770 7580 1778 7599
rect 1798 7580 1806 7599
rect 1770 7577 1806 7580
rect 1771 7549 1805 7577
rect 1885 7571 2212 7605
rect 863 7411 875 7432
rect 897 7411 913 7432
rect 863 7403 913 7411
rect 1086 7435 1142 7440
rect 1086 7415 1093 7435
rect 1113 7415 1142 7435
rect 1086 7408 1142 7415
rect 1243 7521 1806 7549
rect 1086 7407 1121 7408
rect 868 7370 909 7403
rect 1243 7370 1283 7521
rect 868 7341 1283 7370
rect 2172 7347 2212 7571
rect 2873 7590 2902 7592
rect 2873 7585 3246 7590
rect 2873 7567 2880 7585
rect 2900 7567 3246 7585
rect 2873 7562 3246 7567
rect 2878 7560 3246 7562
rect 3007 7523 3042 7524
rect 3222 7523 3246 7560
rect 868 7340 1277 7341
rect 2172 7327 2182 7347
rect 2202 7327 2212 7347
rect 2172 7317 2212 7327
rect 2986 7516 3042 7523
rect 2986 7496 3015 7516
rect 3035 7496 3042 7516
rect 2986 7491 3042 7496
rect 3217 7518 3254 7523
rect 3217 7499 3225 7518
rect 3248 7499 3254 7518
rect 3217 7493 3254 7499
rect 3433 7519 3465 7526
rect 3433 7499 3439 7519
rect 3460 7499 3465 7519
rect 1731 7254 1763 7261
rect 1731 7234 1738 7254
rect 1759 7234 1763 7254
rect 1731 7169 1763 7234
rect 2101 7169 2141 7170
rect 1731 7167 2143 7169
rect 1731 7141 2111 7167
rect 2137 7141 2143 7167
rect 1731 7133 2143 7141
rect 1116 7113 1148 7114
rect 1113 7108 1148 7113
rect 1113 7088 1120 7108
rect 1140 7088 1148 7108
rect 1113 7080 1148 7088
rect 669 7015 701 7022
rect 669 6995 676 7015
rect 697 6995 701 7015
rect 669 6930 701 6995
rect 1039 6930 1079 6931
rect 669 6928 1081 6930
rect 669 6902 1049 6928
rect 1075 6902 1081 6928
rect 669 6894 1081 6902
rect 669 6866 701 6894
rect 1114 6874 1148 7080
rect 1731 7105 1763 7133
rect 1731 7085 1736 7105
rect 1757 7085 1763 7105
rect 1731 7078 1763 7085
rect 1942 7104 1980 7116
rect 2176 7113 2210 7317
rect 2986 7287 3020 7491
rect 3433 7471 3465 7499
rect 4048 7524 4082 7730
rect 4495 7710 4527 7738
rect 6160 7763 6188 7795
rect 6481 7763 6512 7903
rect 7401 7887 7436 7903
rect 7401 7867 7408 7887
rect 7428 7867 7436 7887
rect 7401 7859 7436 7867
rect 6160 7732 6512 7763
rect 6957 7794 6989 7801
rect 6957 7774 6964 7794
rect 6985 7774 6989 7794
rect 4115 7702 4527 7710
rect 4115 7676 4121 7702
rect 4147 7676 4527 7702
rect 4115 7674 4527 7676
rect 4117 7673 4157 7674
rect 4495 7609 4527 7674
rect 6957 7709 6989 7774
rect 7327 7709 7367 7710
rect 6957 7707 7369 7709
rect 6957 7681 7337 7707
rect 7363 7681 7369 7707
rect 6957 7673 7369 7681
rect 6391 7658 6423 7659
rect 6388 7653 6423 7658
rect 6388 7633 6395 7653
rect 6415 7633 6423 7653
rect 6388 7625 6423 7633
rect 4495 7589 4499 7609
rect 4520 7589 4527 7609
rect 4495 7582 4527 7589
rect 5944 7560 5976 7567
rect 5944 7540 5951 7560
rect 5972 7540 5976 7560
rect 4048 7516 4083 7524
rect 4048 7496 4056 7516
rect 4076 7496 4083 7516
rect 4048 7491 4083 7496
rect 4048 7490 4080 7491
rect 3053 7463 3465 7471
rect 3053 7437 3059 7463
rect 3085 7437 3465 7463
rect 3053 7435 3465 7437
rect 3055 7434 3095 7435
rect 3433 7370 3465 7435
rect 5944 7475 5976 7540
rect 6314 7475 6354 7476
rect 5944 7473 6356 7475
rect 5944 7447 6324 7473
rect 6350 7447 6356 7473
rect 5944 7439 6356 7447
rect 5944 7411 5976 7439
rect 5944 7391 5949 7411
rect 5970 7391 5976 7411
rect 5944 7384 5976 7391
rect 6144 7411 6194 7420
rect 6389 7419 6423 7625
rect 6957 7645 6989 7673
rect 6957 7625 6962 7645
rect 6983 7625 6989 7645
rect 6957 7618 6989 7625
rect 7164 7646 7206 7654
rect 7402 7653 7436 7859
rect 7164 7626 7173 7646
rect 7197 7626 7206 7646
rect 7164 7614 7206 7626
rect 7380 7648 7436 7653
rect 7380 7628 7387 7648
rect 7407 7628 7436 7648
rect 8317 7895 8346 7915
rect 8366 7895 8373 7915
rect 8317 7890 8373 7895
rect 8549 7916 8592 7927
rect 8549 7896 8557 7916
rect 8581 7910 8592 7916
rect 8764 7918 8796 7925
rect 8581 7896 8591 7910
rect 8317 7684 8351 7890
rect 8549 7887 8591 7896
rect 8764 7898 8770 7918
rect 8791 7898 8796 7918
rect 8764 7870 8796 7898
rect 9330 7918 9364 8124
rect 9559 8123 9609 8132
rect 9777 8152 9809 8159
rect 9777 8132 9783 8152
rect 9804 8132 9809 8152
rect 9777 8104 9809 8132
rect 9397 8096 9809 8104
rect 9397 8070 9403 8096
rect 9429 8070 9809 8096
rect 9397 8068 9809 8070
rect 9399 8067 9439 8068
rect 9777 8003 9809 8068
rect 9777 7983 9781 8003
rect 9802 7983 9809 8003
rect 9777 7976 9809 7983
rect 9330 7910 9365 7918
rect 9330 7890 9338 7910
rect 9358 7890 9365 7910
rect 9330 7885 9365 7890
rect 9330 7884 9362 7885
rect 8384 7862 8796 7870
rect 8384 7836 8390 7862
rect 8416 7836 8796 7862
rect 8384 7834 8796 7836
rect 8386 7833 8426 7834
rect 8764 7769 8796 7834
rect 8764 7749 8768 7769
rect 8789 7749 8796 7769
rect 8764 7742 8796 7749
rect 9241 7780 9593 7811
rect 8317 7676 8352 7684
rect 8317 7656 8325 7676
rect 8345 7656 8352 7676
rect 8317 7640 8352 7656
rect 9241 7640 9272 7780
rect 9565 7748 9593 7780
rect 9350 7741 9385 7742
rect 7380 7621 7436 7628
rect 8315 7621 9272 7640
rect 9329 7734 9385 7741
rect 9329 7714 9358 7734
rect 9378 7714 9385 7734
rect 9329 7709 9385 7714
rect 9559 7736 9599 7748
rect 9559 7715 9565 7736
rect 9587 7715 9599 7736
rect 9559 7710 9599 7715
rect 9776 7737 9808 7744
rect 9776 7717 9782 7737
rect 9803 7717 9808 7737
rect 7380 7620 7415 7621
rect 7166 7585 7201 7614
rect 7166 7584 7476 7585
rect 7051 7578 7087 7582
rect 7051 7559 7059 7578
rect 7079 7559 7087 7578
rect 7051 7556 7087 7559
rect 7052 7528 7086 7556
rect 7166 7550 7493 7584
rect 6144 7390 6156 7411
rect 6178 7390 6194 7411
rect 6144 7382 6194 7390
rect 6367 7414 6423 7419
rect 6367 7394 6374 7414
rect 6394 7394 6423 7414
rect 6367 7387 6423 7394
rect 6524 7500 7087 7528
rect 6367 7386 6402 7387
rect 3433 7350 3437 7370
rect 3458 7350 3465 7370
rect 3433 7343 3465 7350
rect 6149 7349 6190 7382
rect 6524 7349 6564 7500
rect 6149 7320 6564 7349
rect 7453 7326 7493 7550
rect 8154 7569 8183 7571
rect 8154 7564 8527 7569
rect 8154 7546 8161 7564
rect 8181 7546 8527 7564
rect 8154 7541 8527 7546
rect 8159 7539 8527 7541
rect 8288 7502 8323 7503
rect 8503 7502 8527 7539
rect 6149 7319 6558 7320
rect 7453 7306 7463 7326
rect 7483 7306 7493 7326
rect 7453 7296 7493 7306
rect 8267 7495 8323 7502
rect 8267 7475 8296 7495
rect 8316 7475 8323 7495
rect 8267 7470 8323 7475
rect 8498 7497 8535 7502
rect 8498 7478 8506 7497
rect 8529 7478 8535 7497
rect 8498 7472 8535 7478
rect 8714 7498 8746 7505
rect 8714 7478 8720 7498
rect 8741 7478 8746 7498
rect 1942 7087 1951 7104
rect 1975 7087 1980 7104
rect 1942 7044 1980 7087
rect 2154 7108 2210 7113
rect 2154 7088 2161 7108
rect 2181 7088 2210 7108
rect 2154 7081 2210 7088
rect 2984 7277 3024 7287
rect 2984 7257 2994 7277
rect 3014 7257 3024 7277
rect 3919 7263 4328 7264
rect 2154 7080 2189 7081
rect 2288 7044 2372 7049
rect 1942 7015 2372 7044
rect 669 6846 674 6866
rect 695 6846 701 6866
rect 669 6839 701 6846
rect 878 6868 918 6873
rect 878 6847 890 6868
rect 912 6847 918 6868
rect 878 6835 918 6847
rect 1092 6869 1148 6874
rect 1092 6849 1099 6869
rect 1119 6849 1148 6869
rect 1092 6842 1148 6849
rect 1205 6943 2162 6962
rect 1092 6841 1127 6842
rect 884 6803 912 6835
rect 1205 6803 1236 6943
rect 2125 6927 2160 6943
rect 2125 6907 2132 6927
rect 2152 6907 2160 6927
rect 2125 6899 2160 6907
rect 884 6772 1236 6803
rect 1681 6834 1713 6841
rect 1681 6814 1688 6834
rect 1709 6814 1713 6834
rect 1681 6749 1713 6814
rect 2051 6749 2091 6750
rect 1681 6747 2093 6749
rect 1681 6721 2061 6747
rect 2087 6721 2093 6747
rect 1681 6713 2093 6721
rect 1115 6698 1147 6699
rect 1112 6693 1147 6698
rect 1112 6673 1119 6693
rect 1139 6673 1147 6693
rect 1112 6665 1147 6673
rect 668 6600 700 6607
rect 668 6580 675 6600
rect 696 6580 700 6600
rect 668 6515 700 6580
rect 1038 6515 1078 6516
rect 668 6513 1080 6515
rect 668 6487 1048 6513
rect 1074 6487 1080 6513
rect 668 6479 1080 6487
rect 668 6451 700 6479
rect 668 6431 673 6451
rect 694 6431 700 6451
rect 668 6424 700 6431
rect 868 6451 918 6460
rect 1113 6459 1147 6665
rect 1681 6685 1713 6713
rect 1681 6665 1686 6685
rect 1707 6665 1713 6685
rect 1886 6687 1928 6696
rect 2126 6693 2160 6899
rect 1886 6673 1896 6687
rect 1681 6658 1713 6665
rect 1885 6667 1896 6673
rect 1920 6667 1928 6687
rect 1885 6656 1928 6667
rect 2104 6688 2160 6693
rect 2104 6668 2111 6688
rect 2131 6668 2160 6688
rect 2104 6661 2160 6668
rect 2104 6660 2139 6661
rect 1885 6626 1925 6656
rect 1775 6618 1811 6622
rect 1775 6599 1783 6618
rect 1803 6599 1811 6618
rect 1775 6596 1811 6599
rect 1885 6621 2232 6626
rect 1776 6568 1810 6596
rect 1885 6595 2204 6621
rect 2223 6595 2232 6621
rect 1885 6591 2232 6595
rect 868 6430 880 6451
rect 902 6430 918 6451
rect 868 6422 918 6430
rect 1091 6454 1147 6459
rect 1091 6434 1098 6454
rect 1118 6434 1147 6454
rect 1091 6427 1147 6434
rect 1248 6540 1811 6568
rect 1091 6426 1126 6427
rect 873 6389 914 6422
rect 1248 6389 1288 6540
rect 2337 6421 2372 7015
rect 2984 7033 3024 7257
rect 3913 7234 4328 7263
rect 3913 7083 3953 7234
rect 4287 7201 4328 7234
rect 7012 7233 7044 7240
rect 7012 7213 7019 7233
rect 7040 7213 7044 7233
rect 4075 7196 4110 7197
rect 3390 7055 3953 7083
rect 4054 7189 4110 7196
rect 4054 7169 4083 7189
rect 4103 7169 4110 7189
rect 4054 7164 4110 7169
rect 4283 7193 4333 7201
rect 4283 7172 4299 7193
rect 4321 7172 4333 7193
rect 2984 6999 3311 7033
rect 3391 7027 3425 7055
rect 3390 7024 3426 7027
rect 3390 7005 3398 7024
rect 3418 7005 3426 7024
rect 3390 7001 3426 7005
rect 3001 6998 3311 6999
rect 3276 6969 3311 6998
rect 3062 6962 3097 6963
rect 3041 6955 3097 6962
rect 3041 6935 3070 6955
rect 3090 6935 3097 6955
rect 3041 6930 3097 6935
rect 3271 6957 3313 6969
rect 3271 6937 3280 6957
rect 3304 6937 3313 6957
rect 3041 6724 3075 6930
rect 3271 6929 3313 6937
rect 3488 6958 3520 6965
rect 3488 6938 3494 6958
rect 3515 6938 3520 6958
rect 3488 6910 3520 6938
rect 4054 6958 4088 7164
rect 4283 7163 4333 7172
rect 4501 7192 4533 7199
rect 4501 7172 4507 7192
rect 4528 7172 4533 7192
rect 4501 7144 4533 7172
rect 4121 7136 4533 7144
rect 4121 7110 4127 7136
rect 4153 7110 4533 7136
rect 4121 7108 4533 7110
rect 4123 7107 4163 7108
rect 4501 7043 4533 7108
rect 7012 7148 7044 7213
rect 7382 7148 7422 7149
rect 7012 7146 7424 7148
rect 7012 7120 7392 7146
rect 7418 7120 7424 7146
rect 7012 7112 7424 7120
rect 6397 7092 6429 7093
rect 6394 7087 6429 7092
rect 6394 7067 6401 7087
rect 6421 7067 6429 7087
rect 6394 7059 6429 7067
rect 4501 7023 4505 7043
rect 4526 7023 4533 7043
rect 4501 7016 4533 7023
rect 5950 6994 5982 7001
rect 5950 6974 5957 6994
rect 5978 6974 5982 6994
rect 4054 6950 4089 6958
rect 4054 6930 4062 6950
rect 4082 6930 4089 6950
rect 4054 6925 4089 6930
rect 4054 6924 4086 6925
rect 3108 6902 3520 6910
rect 3108 6876 3114 6902
rect 3140 6876 3520 6902
rect 3108 6874 3520 6876
rect 3110 6873 3150 6874
rect 3488 6809 3520 6874
rect 5950 6909 5982 6974
rect 6320 6909 6360 6910
rect 5950 6907 6362 6909
rect 5950 6881 6330 6907
rect 6356 6881 6362 6907
rect 5950 6873 6362 6881
rect 3488 6789 3492 6809
rect 3513 6789 3520 6809
rect 3488 6782 3520 6789
rect 3965 6820 4317 6851
rect 3041 6716 3076 6724
rect 3041 6696 3049 6716
rect 3069 6696 3076 6716
rect 3041 6680 3076 6696
rect 3965 6680 3996 6820
rect 4289 6788 4317 6820
rect 5950 6845 5982 6873
rect 6395 6853 6429 7059
rect 7012 7084 7044 7112
rect 7012 7064 7017 7084
rect 7038 7064 7044 7084
rect 7012 7057 7044 7064
rect 7223 7083 7261 7095
rect 7457 7092 7491 7296
rect 8267 7266 8301 7470
rect 8714 7450 8746 7478
rect 9329 7503 9363 7709
rect 9776 7689 9808 7717
rect 9396 7681 9808 7689
rect 9396 7655 9402 7681
rect 9428 7655 9808 7681
rect 9396 7653 9808 7655
rect 9398 7652 9438 7653
rect 9776 7588 9808 7653
rect 9776 7568 9780 7588
rect 9801 7568 9808 7588
rect 9776 7561 9808 7568
rect 9329 7495 9364 7503
rect 9329 7475 9337 7495
rect 9357 7475 9364 7495
rect 9329 7470 9364 7475
rect 9329 7469 9361 7470
rect 8334 7442 8746 7450
rect 8334 7416 8340 7442
rect 8366 7416 8746 7442
rect 8334 7414 8746 7416
rect 8336 7413 8376 7414
rect 8714 7349 8746 7414
rect 8714 7329 8718 7349
rect 8739 7329 8746 7349
rect 8714 7322 8746 7329
rect 7223 7066 7232 7083
rect 7256 7066 7261 7083
rect 7223 7023 7261 7066
rect 7435 7087 7491 7092
rect 7435 7067 7442 7087
rect 7462 7067 7491 7087
rect 7435 7060 7491 7067
rect 8265 7256 8305 7266
rect 8265 7236 8275 7256
rect 8295 7236 8305 7256
rect 9200 7242 9609 7243
rect 7435 7059 7470 7060
rect 7569 7023 7653 7028
rect 7223 6994 7653 7023
rect 5950 6825 5955 6845
rect 5976 6825 5982 6845
rect 5950 6818 5982 6825
rect 6159 6847 6199 6852
rect 6159 6826 6171 6847
rect 6193 6826 6199 6847
rect 6159 6814 6199 6826
rect 6373 6848 6429 6853
rect 6373 6828 6380 6848
rect 6400 6828 6429 6848
rect 6373 6821 6429 6828
rect 6486 6922 7443 6941
rect 6373 6820 6408 6821
rect 4074 6781 4109 6782
rect 3039 6661 3996 6680
rect 4053 6774 4109 6781
rect 4053 6754 4082 6774
rect 4102 6754 4109 6774
rect 4053 6749 4109 6754
rect 4283 6776 4323 6788
rect 4283 6755 4289 6776
rect 4311 6755 4323 6776
rect 4283 6750 4323 6755
rect 4500 6777 4532 6784
rect 4500 6757 4506 6777
rect 4527 6757 4532 6777
rect 2749 6563 2786 6568
rect 2749 6557 3096 6563
rect 2749 6538 2757 6557
rect 2780 6538 3096 6557
rect 2749 6533 3096 6538
rect 2749 6527 2786 6533
rect 3066 6502 3096 6533
rect 4053 6543 4087 6749
rect 4500 6729 4532 6757
rect 6165 6782 6193 6814
rect 6486 6782 6517 6922
rect 7406 6906 7441 6922
rect 7406 6886 7413 6906
rect 7433 6886 7441 6906
rect 7406 6878 7441 6886
rect 6165 6751 6517 6782
rect 6962 6813 6994 6820
rect 6962 6793 6969 6813
rect 6990 6793 6994 6813
rect 4120 6721 4532 6729
rect 4120 6695 4126 6721
rect 4152 6695 4532 6721
rect 4120 6693 4532 6695
rect 4122 6692 4162 6693
rect 4500 6628 4532 6693
rect 6962 6728 6994 6793
rect 7332 6728 7372 6729
rect 6962 6726 7374 6728
rect 6962 6700 7342 6726
rect 7368 6700 7374 6726
rect 6962 6692 7374 6700
rect 6396 6677 6428 6678
rect 6393 6672 6428 6677
rect 6393 6652 6400 6672
rect 6420 6652 6428 6672
rect 6393 6644 6428 6652
rect 4500 6608 4504 6628
rect 4525 6608 4532 6628
rect 4500 6601 4532 6608
rect 5949 6579 5981 6586
rect 5949 6559 5956 6579
rect 5977 6559 5981 6579
rect 4053 6535 4088 6543
rect 4053 6515 4061 6535
rect 4081 6515 4088 6535
rect 4053 6510 4088 6515
rect 4053 6509 4085 6510
rect 2854 6495 2889 6496
rect 2833 6488 2889 6495
rect 2833 6468 2862 6488
rect 2882 6468 2889 6488
rect 2833 6463 2889 6468
rect 3064 6489 3103 6502
rect 3064 6470 3069 6489
rect 3092 6470 3103 6489
rect 3064 6464 3103 6470
rect 3280 6491 3312 6498
rect 3280 6471 3286 6491
rect 3307 6471 3312 6491
rect 2337 6415 2375 6421
rect 2337 6395 2347 6415
rect 2367 6395 2375 6415
rect 2337 6393 2375 6395
rect 873 6360 1288 6389
rect 2340 6387 2375 6393
rect 873 6359 1282 6360
rect 1896 6322 1928 6329
rect 1896 6302 1903 6322
rect 1924 6302 1928 6322
rect 1896 6237 1928 6302
rect 2266 6237 2306 6238
rect 1896 6235 2308 6237
rect 1896 6209 2276 6235
rect 2302 6209 2308 6235
rect 1896 6201 2308 6209
rect 1896 6173 1928 6201
rect 1896 6153 1901 6173
rect 1922 6153 1928 6173
rect 1896 6146 1928 6153
rect 2100 6178 2147 6184
rect 2341 6181 2375 6387
rect 2833 6257 2867 6463
rect 3280 6443 3312 6471
rect 2900 6435 3312 6443
rect 2900 6409 2906 6435
rect 2932 6409 3312 6435
rect 2900 6407 3312 6409
rect 2902 6406 2942 6407
rect 3280 6342 3312 6407
rect 5949 6494 5981 6559
rect 6319 6494 6359 6495
rect 5949 6492 6361 6494
rect 5949 6466 6329 6492
rect 6355 6466 6361 6492
rect 5949 6458 6361 6466
rect 5949 6430 5981 6458
rect 5949 6410 5954 6430
rect 5975 6410 5981 6430
rect 5949 6403 5981 6410
rect 6149 6430 6199 6439
rect 6394 6438 6428 6644
rect 6962 6664 6994 6692
rect 6962 6644 6967 6664
rect 6988 6644 6994 6664
rect 7167 6666 7209 6675
rect 7407 6672 7441 6878
rect 7167 6652 7177 6666
rect 6962 6637 6994 6644
rect 7166 6646 7177 6652
rect 7201 6646 7209 6666
rect 7166 6635 7209 6646
rect 7385 6667 7441 6672
rect 7385 6647 7392 6667
rect 7412 6647 7441 6667
rect 7385 6640 7441 6647
rect 7385 6639 7420 6640
rect 7166 6605 7206 6635
rect 7056 6597 7092 6601
rect 7056 6578 7064 6597
rect 7084 6578 7092 6597
rect 7056 6575 7092 6578
rect 7166 6600 7513 6605
rect 7057 6547 7091 6575
rect 7166 6574 7485 6600
rect 7504 6574 7513 6600
rect 7166 6570 7513 6574
rect 6149 6409 6161 6430
rect 6183 6409 6199 6430
rect 6149 6401 6199 6409
rect 6372 6433 6428 6438
rect 6372 6413 6379 6433
rect 6399 6413 6428 6433
rect 6372 6406 6428 6413
rect 6529 6519 7092 6547
rect 6372 6405 6407 6406
rect 3280 6322 3284 6342
rect 3305 6322 3312 6342
rect 6154 6368 6195 6401
rect 6529 6368 6569 6519
rect 7618 6400 7653 6994
rect 8265 7012 8305 7236
rect 9194 7213 9609 7242
rect 9194 7062 9234 7213
rect 9568 7180 9609 7213
rect 9356 7175 9391 7176
rect 8671 7034 9234 7062
rect 9335 7168 9391 7175
rect 9335 7148 9364 7168
rect 9384 7148 9391 7168
rect 9335 7143 9391 7148
rect 9564 7172 9614 7180
rect 9564 7151 9580 7172
rect 9602 7151 9614 7172
rect 8265 6978 8592 7012
rect 8672 7006 8706 7034
rect 8671 7003 8707 7006
rect 8671 6984 8679 7003
rect 8699 6984 8707 7003
rect 8671 6980 8707 6984
rect 8282 6977 8592 6978
rect 8557 6948 8592 6977
rect 8343 6941 8378 6942
rect 8322 6934 8378 6941
rect 8322 6914 8351 6934
rect 8371 6914 8378 6934
rect 8322 6909 8378 6914
rect 8552 6936 8594 6948
rect 8552 6916 8561 6936
rect 8585 6916 8594 6936
rect 8322 6703 8356 6909
rect 8552 6908 8594 6916
rect 8769 6937 8801 6944
rect 8769 6917 8775 6937
rect 8796 6917 8801 6937
rect 8769 6889 8801 6917
rect 9335 6937 9369 7143
rect 9564 7142 9614 7151
rect 9782 7171 9814 7178
rect 9782 7151 9788 7171
rect 9809 7151 9814 7171
rect 9782 7123 9814 7151
rect 9402 7115 9814 7123
rect 9402 7089 9408 7115
rect 9434 7089 9814 7115
rect 9402 7087 9814 7089
rect 9404 7086 9444 7087
rect 9782 7022 9814 7087
rect 9782 7002 9786 7022
rect 9807 7002 9814 7022
rect 9782 6995 9814 7002
rect 9335 6929 9370 6937
rect 9335 6909 9343 6929
rect 9363 6909 9370 6929
rect 9335 6904 9370 6909
rect 9335 6903 9367 6904
rect 8389 6881 8801 6889
rect 8389 6855 8395 6881
rect 8421 6855 8801 6881
rect 8389 6853 8801 6855
rect 8391 6852 8431 6853
rect 8769 6788 8801 6853
rect 8769 6768 8773 6788
rect 8794 6768 8801 6788
rect 8769 6761 8801 6768
rect 9246 6799 9598 6830
rect 8322 6695 8357 6703
rect 8322 6675 8330 6695
rect 8350 6675 8357 6695
rect 8322 6659 8357 6675
rect 9246 6659 9277 6799
rect 9570 6767 9598 6799
rect 9355 6760 9390 6761
rect 8320 6640 9277 6659
rect 9334 6753 9390 6760
rect 9334 6733 9363 6753
rect 9383 6733 9390 6753
rect 9334 6728 9390 6733
rect 9564 6755 9604 6767
rect 9564 6734 9570 6755
rect 9592 6734 9604 6755
rect 9564 6729 9604 6734
rect 9781 6756 9813 6763
rect 9781 6736 9787 6756
rect 9808 6736 9813 6756
rect 8030 6542 8067 6547
rect 8030 6536 8377 6542
rect 8030 6517 8038 6536
rect 8061 6517 8377 6536
rect 8030 6512 8377 6517
rect 8030 6506 8067 6512
rect 8347 6481 8377 6512
rect 9334 6522 9368 6728
rect 9781 6708 9813 6736
rect 9401 6700 9813 6708
rect 9401 6674 9407 6700
rect 9433 6674 9813 6700
rect 9401 6672 9813 6674
rect 9403 6671 9443 6672
rect 9781 6607 9813 6672
rect 9781 6587 9785 6607
rect 9806 6587 9813 6607
rect 9781 6580 9813 6587
rect 9334 6514 9369 6522
rect 9334 6494 9342 6514
rect 9362 6494 9369 6514
rect 9334 6489 9369 6494
rect 9334 6488 9366 6489
rect 8135 6474 8170 6475
rect 8114 6467 8170 6474
rect 8114 6447 8143 6467
rect 8163 6447 8170 6467
rect 8114 6442 8170 6447
rect 8345 6468 8384 6481
rect 8345 6449 8350 6468
rect 8373 6449 8384 6468
rect 8345 6443 8384 6449
rect 8561 6470 8593 6477
rect 8561 6450 8567 6470
rect 8588 6450 8593 6470
rect 7618 6394 7656 6400
rect 7618 6374 7628 6394
rect 7648 6374 7656 6394
rect 7618 6372 7656 6374
rect 6154 6339 6569 6368
rect 7621 6366 7656 6372
rect 6154 6338 6563 6339
rect 3280 6315 3312 6322
rect 7177 6301 7209 6308
rect 3926 6284 4335 6285
rect 2833 6251 2868 6257
rect 3920 6255 4335 6284
rect 2833 6249 2871 6251
rect 2833 6229 2841 6249
rect 2861 6229 2871 6249
rect 2833 6223 2871 6229
rect 2100 6152 2110 6178
rect 2135 6152 2147 6178
rect 2100 6150 2147 6152
rect 2319 6176 2375 6181
rect 2319 6156 2326 6176
rect 2346 6156 2375 6176
rect 1123 6134 1155 6135
rect 1120 6129 1155 6134
rect 1120 6109 1127 6129
rect 1147 6109 1155 6129
rect 1120 6101 1155 6109
rect 676 6036 708 6043
rect 676 6016 683 6036
rect 704 6016 708 6036
rect 676 5951 708 6016
rect 1046 5951 1086 5952
rect 676 5949 1088 5951
rect 676 5923 1056 5949
rect 1082 5923 1088 5949
rect 676 5915 1088 5923
rect 676 5887 708 5915
rect 1121 5895 1155 6101
rect 2105 6115 2142 6150
rect 2319 6149 2375 6156
rect 2319 6148 2354 6149
rect 2439 6115 2471 6117
rect 2105 6082 2475 6115
rect 676 5867 681 5887
rect 702 5867 708 5887
rect 676 5860 708 5867
rect 885 5889 925 5894
rect 885 5868 897 5889
rect 919 5868 925 5889
rect 885 5856 925 5868
rect 1099 5890 1155 5895
rect 1099 5870 1106 5890
rect 1126 5870 1155 5890
rect 1099 5863 1155 5870
rect 1212 5964 2169 5983
rect 1099 5862 1134 5863
rect 891 5824 919 5856
rect 1212 5824 1243 5964
rect 2132 5948 2167 5964
rect 2132 5928 2139 5948
rect 2159 5928 2167 5948
rect 2132 5920 2167 5928
rect 891 5793 1243 5824
rect 1688 5855 1720 5862
rect 1688 5835 1695 5855
rect 1716 5835 1720 5855
rect 1688 5770 1720 5835
rect 2058 5770 2098 5771
rect 1688 5768 2100 5770
rect 1688 5742 2068 5768
rect 2094 5742 2100 5768
rect 1688 5734 2100 5742
rect 1122 5719 1154 5720
rect 1119 5714 1154 5719
rect 1119 5694 1126 5714
rect 1146 5694 1154 5714
rect 1119 5686 1154 5694
rect 675 5621 707 5628
rect 675 5601 682 5621
rect 703 5601 707 5621
rect 675 5536 707 5601
rect 1045 5536 1085 5537
rect 675 5534 1087 5536
rect 675 5508 1055 5534
rect 1081 5508 1087 5534
rect 675 5500 1087 5508
rect 675 5472 707 5500
rect 675 5452 680 5472
rect 701 5452 707 5472
rect 675 5445 707 5452
rect 875 5472 925 5481
rect 1120 5480 1154 5686
rect 1688 5706 1720 5734
rect 1688 5686 1693 5706
rect 1714 5686 1720 5706
rect 1688 5679 1720 5686
rect 1895 5707 1937 5715
rect 2133 5714 2167 5920
rect 1895 5687 1904 5707
rect 1928 5687 1937 5707
rect 1895 5675 1937 5687
rect 2111 5709 2167 5714
rect 2111 5689 2118 5709
rect 2138 5689 2167 5709
rect 2111 5682 2167 5689
rect 2111 5681 2146 5682
rect 1897 5646 1932 5675
rect 1897 5645 2207 5646
rect 1782 5639 1818 5643
rect 1782 5620 1790 5639
rect 1810 5620 1818 5639
rect 1782 5617 1818 5620
rect 1783 5589 1817 5617
rect 1897 5611 2224 5645
rect 875 5451 887 5472
rect 909 5451 925 5472
rect 875 5443 925 5451
rect 1098 5475 1154 5480
rect 1098 5455 1105 5475
rect 1125 5455 1154 5475
rect 1098 5448 1154 5455
rect 1255 5561 1818 5589
rect 1098 5447 1133 5448
rect 880 5410 921 5443
rect 1255 5410 1295 5561
rect 880 5381 1295 5410
rect 2184 5387 2224 5611
rect 880 5380 1289 5381
rect 2184 5367 2194 5387
rect 2214 5367 2224 5387
rect 2184 5357 2224 5367
rect 1743 5294 1775 5301
rect 1743 5274 1750 5294
rect 1771 5274 1775 5294
rect 1743 5209 1775 5274
rect 2113 5209 2153 5210
rect 1743 5207 2155 5209
rect 1743 5181 2123 5207
rect 2149 5181 2155 5207
rect 1743 5173 2155 5181
rect 1128 5153 1160 5154
rect 1125 5148 1160 5153
rect 1125 5128 1132 5148
rect 1152 5128 1160 5148
rect 1125 5120 1160 5128
rect 681 5055 713 5062
rect 681 5035 688 5055
rect 709 5035 713 5055
rect 681 4970 713 5035
rect 1051 4970 1091 4971
rect 681 4968 1093 4970
rect 681 4942 1061 4968
rect 1087 4942 1093 4968
rect 681 4934 1093 4942
rect 681 4906 713 4934
rect 1126 4914 1160 5120
rect 1743 5145 1775 5173
rect 2188 5153 2222 5357
rect 1743 5125 1748 5145
rect 1769 5125 1775 5145
rect 1743 5118 1775 5125
rect 1954 5145 1991 5151
rect 1954 5126 1960 5145
rect 1983 5126 1991 5145
rect 1954 5121 1991 5126
rect 2166 5148 2222 5153
rect 2166 5128 2173 5148
rect 2193 5128 2222 5148
rect 2166 5121 2222 5128
rect 1962 5084 1986 5121
rect 2166 5120 2201 5121
rect 1962 5082 2330 5084
rect 1962 5077 2335 5082
rect 1962 5059 2308 5077
rect 2328 5059 2335 5077
rect 1962 5054 2335 5059
rect 2306 5052 2335 5054
rect 681 4886 686 4906
rect 707 4886 713 4906
rect 681 4879 713 4886
rect 890 4908 930 4913
rect 890 4887 902 4908
rect 924 4887 930 4908
rect 890 4875 930 4887
rect 1104 4909 1160 4914
rect 1104 4889 1111 4909
rect 1131 4889 1160 4909
rect 1104 4882 1160 4889
rect 1217 4983 2174 5002
rect 1104 4881 1139 4882
rect 896 4843 924 4875
rect 1217 4843 1248 4983
rect 2137 4967 2172 4983
rect 2137 4947 2144 4967
rect 2164 4947 2172 4967
rect 2137 4939 2172 4947
rect 896 4812 1248 4843
rect 1693 4874 1725 4881
rect 1693 4854 1700 4874
rect 1721 4854 1725 4874
rect 1693 4789 1725 4854
rect 2063 4789 2103 4790
rect 1693 4787 2105 4789
rect 1693 4761 2073 4787
rect 2099 4761 2105 4787
rect 1693 4753 2105 4761
rect 1127 4738 1159 4739
rect 1124 4733 1159 4738
rect 1124 4713 1131 4733
rect 1151 4713 1159 4733
rect 1124 4705 1159 4713
rect 680 4640 712 4647
rect 680 4620 687 4640
rect 708 4620 712 4640
rect 680 4555 712 4620
rect 1050 4555 1090 4556
rect 680 4553 1092 4555
rect 680 4527 1060 4553
rect 1086 4527 1092 4553
rect 680 4519 1092 4527
rect 680 4491 712 4519
rect 680 4471 685 4491
rect 706 4471 712 4491
rect 680 4464 712 4471
rect 880 4491 930 4500
rect 1125 4499 1159 4705
rect 1693 4725 1725 4753
rect 1693 4705 1698 4725
rect 1719 4705 1725 4725
rect 1898 4727 1940 4736
rect 2138 4733 2172 4939
rect 1898 4713 1908 4727
rect 1693 4698 1725 4705
rect 1897 4707 1908 4713
rect 1932 4707 1940 4727
rect 1897 4696 1940 4707
rect 2116 4728 2172 4733
rect 2116 4708 2123 4728
rect 2143 4708 2172 4728
rect 2116 4701 2172 4708
rect 2116 4700 2151 4701
rect 1897 4666 1937 4696
rect 1787 4658 1823 4662
rect 1787 4639 1795 4658
rect 1815 4639 1823 4658
rect 1787 4636 1823 4639
rect 1897 4661 2244 4666
rect 1788 4608 1822 4636
rect 1897 4635 2216 4661
rect 2235 4635 2244 4661
rect 1897 4631 2244 4635
rect 880 4470 892 4491
rect 914 4470 930 4491
rect 880 4462 930 4470
rect 1103 4494 1159 4499
rect 1103 4474 1110 4494
rect 1130 4474 1159 4494
rect 1103 4467 1159 4474
rect 1260 4580 1823 4608
rect 1103 4466 1138 4467
rect 885 4429 926 4462
rect 1260 4429 1300 4580
rect 2439 4429 2471 6082
rect 2836 5629 2871 6223
rect 3920 6104 3960 6255
rect 4294 6222 4335 6255
rect 7177 6281 7184 6301
rect 7205 6281 7209 6301
rect 4082 6217 4117 6218
rect 3397 6076 3960 6104
rect 4061 6210 4117 6217
rect 4061 6190 4090 6210
rect 4110 6190 4117 6210
rect 4061 6185 4117 6190
rect 4290 6214 4340 6222
rect 4290 6193 4306 6214
rect 4328 6193 4340 6214
rect 2976 6049 3323 6053
rect 2976 6023 2985 6049
rect 3004 6023 3323 6049
rect 3398 6048 3432 6076
rect 2976 6018 3323 6023
rect 3397 6045 3433 6048
rect 3397 6026 3405 6045
rect 3425 6026 3433 6045
rect 3397 6022 3433 6026
rect 3283 5988 3323 6018
rect 3069 5983 3104 5984
rect 3048 5976 3104 5983
rect 3048 5956 3077 5976
rect 3097 5956 3104 5976
rect 3048 5951 3104 5956
rect 3280 5977 3323 5988
rect 3280 5957 3288 5977
rect 3312 5971 3323 5977
rect 3495 5979 3527 5986
rect 3312 5957 3322 5971
rect 3048 5745 3082 5951
rect 3280 5948 3322 5957
rect 3495 5959 3501 5979
rect 3522 5959 3527 5979
rect 3495 5931 3527 5959
rect 4061 5979 4095 6185
rect 4290 6184 4340 6193
rect 4508 6213 4540 6220
rect 4508 6193 4514 6213
rect 4535 6193 4540 6213
rect 4508 6165 4540 6193
rect 4128 6157 4540 6165
rect 4128 6131 4134 6157
rect 4160 6131 4540 6157
rect 4128 6129 4540 6131
rect 4130 6128 4170 6129
rect 4508 6064 4540 6129
rect 7177 6216 7209 6281
rect 7547 6216 7587 6217
rect 7177 6214 7589 6216
rect 7177 6188 7557 6214
rect 7583 6188 7589 6214
rect 7177 6180 7589 6188
rect 7177 6152 7209 6180
rect 7177 6132 7182 6152
rect 7203 6132 7209 6152
rect 7177 6125 7209 6132
rect 7381 6157 7428 6163
rect 7622 6160 7656 6366
rect 8114 6236 8148 6442
rect 8561 6422 8593 6450
rect 8181 6414 8593 6422
rect 8181 6388 8187 6414
rect 8213 6388 8593 6414
rect 8181 6386 8593 6388
rect 8183 6385 8223 6386
rect 8561 6321 8593 6386
rect 8561 6301 8565 6321
rect 8586 6301 8593 6321
rect 8561 6294 8593 6301
rect 9207 6263 9616 6264
rect 8114 6230 8149 6236
rect 9201 6234 9616 6263
rect 8114 6228 8152 6230
rect 8114 6208 8122 6228
rect 8142 6208 8152 6228
rect 8114 6202 8152 6208
rect 7381 6131 7391 6157
rect 7416 6131 7428 6157
rect 7381 6129 7428 6131
rect 7600 6155 7656 6160
rect 7600 6135 7607 6155
rect 7627 6135 7656 6155
rect 6404 6113 6436 6114
rect 6401 6108 6436 6113
rect 6401 6088 6408 6108
rect 6428 6088 6436 6108
rect 6401 6080 6436 6088
rect 4508 6044 4512 6064
rect 4533 6044 4540 6064
rect 4508 6037 4540 6044
rect 5957 6015 5989 6022
rect 5957 5995 5964 6015
rect 5985 5995 5989 6015
rect 4061 5971 4096 5979
rect 4061 5951 4069 5971
rect 4089 5951 4096 5971
rect 4061 5946 4096 5951
rect 4061 5945 4093 5946
rect 3115 5923 3527 5931
rect 3115 5897 3121 5923
rect 3147 5897 3527 5923
rect 3115 5895 3527 5897
rect 3117 5894 3157 5895
rect 3495 5830 3527 5895
rect 5957 5930 5989 5995
rect 6327 5930 6367 5931
rect 5957 5928 6369 5930
rect 5957 5902 6337 5928
rect 6363 5902 6369 5928
rect 5957 5894 6369 5902
rect 3495 5810 3499 5830
rect 3520 5810 3527 5830
rect 3495 5803 3527 5810
rect 3972 5841 4324 5872
rect 3048 5737 3083 5745
rect 3048 5717 3056 5737
rect 3076 5717 3083 5737
rect 3048 5701 3083 5717
rect 3972 5701 4003 5841
rect 4296 5809 4324 5841
rect 5957 5866 5989 5894
rect 6402 5874 6436 6080
rect 7386 6094 7423 6129
rect 7600 6128 7656 6135
rect 7600 6127 7635 6128
rect 7720 6094 7752 6096
rect 7386 6061 7756 6094
rect 5957 5846 5962 5866
rect 5983 5846 5989 5866
rect 5957 5839 5989 5846
rect 6166 5868 6206 5873
rect 6166 5847 6178 5868
rect 6200 5847 6206 5868
rect 6166 5835 6206 5847
rect 6380 5869 6436 5874
rect 6380 5849 6387 5869
rect 6407 5849 6436 5869
rect 6380 5842 6436 5849
rect 6493 5943 7450 5962
rect 6380 5841 6415 5842
rect 4081 5802 4116 5803
rect 3046 5682 4003 5701
rect 4060 5795 4116 5802
rect 4060 5775 4089 5795
rect 4109 5775 4116 5795
rect 4060 5770 4116 5775
rect 4290 5797 4330 5809
rect 4290 5776 4296 5797
rect 4318 5776 4330 5797
rect 4290 5771 4330 5776
rect 4507 5798 4539 5805
rect 4507 5778 4513 5798
rect 4534 5778 4539 5798
rect 2836 5600 3266 5629
rect 2836 5595 2920 5600
rect 3019 5563 3054 5564
rect 2998 5556 3054 5563
rect 2998 5536 3027 5556
rect 3047 5536 3054 5556
rect 2998 5531 3054 5536
rect 3228 5557 3266 5600
rect 3228 5540 3233 5557
rect 3257 5540 3266 5557
rect 2998 5327 3032 5531
rect 3228 5528 3266 5540
rect 3445 5559 3477 5566
rect 3445 5539 3451 5559
rect 3472 5539 3477 5559
rect 3445 5511 3477 5539
rect 4060 5564 4094 5770
rect 4507 5750 4539 5778
rect 6172 5803 6200 5835
rect 6493 5803 6524 5943
rect 7413 5927 7448 5943
rect 7413 5907 7420 5927
rect 7440 5907 7448 5927
rect 7413 5899 7448 5907
rect 6172 5772 6524 5803
rect 6969 5834 7001 5841
rect 6969 5814 6976 5834
rect 6997 5814 7001 5834
rect 4127 5742 4539 5750
rect 4127 5716 4133 5742
rect 4159 5716 4539 5742
rect 4127 5714 4539 5716
rect 4129 5713 4169 5714
rect 4507 5649 4539 5714
rect 6969 5749 7001 5814
rect 7339 5749 7379 5750
rect 6969 5747 7381 5749
rect 6969 5721 7349 5747
rect 7375 5721 7381 5747
rect 6969 5713 7381 5721
rect 6403 5698 6435 5699
rect 6400 5693 6435 5698
rect 6400 5673 6407 5693
rect 6427 5673 6435 5693
rect 6400 5665 6435 5673
rect 4507 5629 4511 5649
rect 4532 5629 4539 5649
rect 4507 5622 4539 5629
rect 5956 5600 5988 5607
rect 5956 5580 5963 5600
rect 5984 5580 5988 5600
rect 4060 5556 4095 5564
rect 4060 5536 4068 5556
rect 4088 5536 4095 5556
rect 4060 5531 4095 5536
rect 4060 5530 4092 5531
rect 3065 5503 3477 5511
rect 3065 5477 3071 5503
rect 3097 5477 3477 5503
rect 3065 5475 3477 5477
rect 3067 5474 3107 5475
rect 3445 5410 3477 5475
rect 5956 5515 5988 5580
rect 6326 5515 6366 5516
rect 5956 5513 6368 5515
rect 5956 5487 6336 5513
rect 6362 5487 6368 5513
rect 5956 5479 6368 5487
rect 5956 5451 5988 5479
rect 5956 5431 5961 5451
rect 5982 5431 5988 5451
rect 5956 5424 5988 5431
rect 6156 5451 6206 5460
rect 6401 5459 6435 5665
rect 6969 5685 7001 5713
rect 6969 5665 6974 5685
rect 6995 5665 7001 5685
rect 6969 5658 7001 5665
rect 7176 5686 7218 5694
rect 7414 5693 7448 5899
rect 7176 5666 7185 5686
rect 7209 5666 7218 5686
rect 7176 5654 7218 5666
rect 7392 5688 7448 5693
rect 7392 5668 7399 5688
rect 7419 5668 7448 5688
rect 7392 5661 7448 5668
rect 7392 5660 7427 5661
rect 7178 5625 7213 5654
rect 7178 5624 7488 5625
rect 7063 5618 7099 5622
rect 7063 5599 7071 5618
rect 7091 5599 7099 5618
rect 7063 5596 7099 5599
rect 7064 5568 7098 5596
rect 7178 5590 7505 5624
rect 6156 5430 6168 5451
rect 6190 5430 6206 5451
rect 6156 5422 6206 5430
rect 6379 5454 6435 5459
rect 6379 5434 6386 5454
rect 6406 5434 6435 5454
rect 6379 5427 6435 5434
rect 6536 5540 7099 5568
rect 6379 5426 6414 5427
rect 3445 5390 3449 5410
rect 3470 5390 3477 5410
rect 3445 5383 3477 5390
rect 6161 5389 6202 5422
rect 6536 5389 6576 5540
rect 6161 5360 6576 5389
rect 7465 5366 7505 5590
rect 6161 5359 6570 5360
rect 7465 5346 7475 5366
rect 7495 5346 7505 5366
rect 7465 5336 7505 5346
rect 2996 5317 3036 5327
rect 2996 5297 3006 5317
rect 3026 5297 3036 5317
rect 3931 5303 4340 5304
rect 2996 5073 3036 5297
rect 3925 5274 4340 5303
rect 3925 5123 3965 5274
rect 4299 5241 4340 5274
rect 7024 5273 7056 5280
rect 7024 5253 7031 5273
rect 7052 5253 7056 5273
rect 4087 5236 4122 5237
rect 3402 5095 3965 5123
rect 4066 5229 4122 5236
rect 4066 5209 4095 5229
rect 4115 5209 4122 5229
rect 4066 5204 4122 5209
rect 4295 5233 4345 5241
rect 4295 5212 4311 5233
rect 4333 5212 4345 5233
rect 2996 5039 3323 5073
rect 3403 5067 3437 5095
rect 3402 5064 3438 5067
rect 3402 5045 3410 5064
rect 3430 5045 3438 5064
rect 3402 5041 3438 5045
rect 3013 5038 3323 5039
rect 3288 5009 3323 5038
rect 3074 5002 3109 5003
rect 3053 4995 3109 5002
rect 3053 4975 3082 4995
rect 3102 4975 3109 4995
rect 3053 4970 3109 4975
rect 3283 4997 3325 5009
rect 3283 4977 3292 4997
rect 3316 4977 3325 4997
rect 3053 4764 3087 4970
rect 3283 4969 3325 4977
rect 3500 4998 3532 5005
rect 3500 4978 3506 4998
rect 3527 4978 3532 4998
rect 3500 4950 3532 4978
rect 4066 4998 4100 5204
rect 4295 5203 4345 5212
rect 4513 5232 4545 5239
rect 4513 5212 4519 5232
rect 4540 5212 4545 5232
rect 4513 5184 4545 5212
rect 4133 5176 4545 5184
rect 4133 5150 4139 5176
rect 4165 5150 4545 5176
rect 4133 5148 4545 5150
rect 4135 5147 4175 5148
rect 4513 5083 4545 5148
rect 7024 5188 7056 5253
rect 7394 5188 7434 5189
rect 7024 5186 7436 5188
rect 7024 5160 7404 5186
rect 7430 5160 7436 5186
rect 7024 5152 7436 5160
rect 6409 5132 6441 5133
rect 6406 5127 6441 5132
rect 6406 5107 6413 5127
rect 6433 5107 6441 5127
rect 6406 5099 6441 5107
rect 4513 5063 4517 5083
rect 4538 5063 4545 5083
rect 4513 5056 4545 5063
rect 5962 5034 5994 5041
rect 5962 5014 5969 5034
rect 5990 5014 5994 5034
rect 4066 4990 4101 4998
rect 4066 4970 4074 4990
rect 4094 4970 4101 4990
rect 4066 4965 4101 4970
rect 4066 4964 4098 4965
rect 3120 4942 3532 4950
rect 3120 4916 3126 4942
rect 3152 4916 3532 4942
rect 3120 4914 3532 4916
rect 3122 4913 3162 4914
rect 3500 4849 3532 4914
rect 5962 4949 5994 5014
rect 6332 4949 6372 4950
rect 5962 4947 6374 4949
rect 5962 4921 6342 4947
rect 6368 4921 6374 4947
rect 5962 4913 6374 4921
rect 3500 4829 3504 4849
rect 3525 4829 3532 4849
rect 3500 4822 3532 4829
rect 3977 4860 4329 4891
rect 3053 4756 3088 4764
rect 3053 4736 3061 4756
rect 3081 4736 3088 4756
rect 3053 4720 3088 4736
rect 3977 4720 4008 4860
rect 4301 4828 4329 4860
rect 5962 4885 5994 4913
rect 6407 4893 6441 5099
rect 7024 5124 7056 5152
rect 7469 5132 7503 5336
rect 7024 5104 7029 5124
rect 7050 5104 7056 5124
rect 7024 5097 7056 5104
rect 7235 5124 7272 5130
rect 7235 5105 7241 5124
rect 7264 5105 7272 5124
rect 7235 5100 7272 5105
rect 7447 5127 7503 5132
rect 7447 5107 7454 5127
rect 7474 5107 7503 5127
rect 7447 5100 7503 5107
rect 7243 5063 7267 5100
rect 7447 5099 7482 5100
rect 7243 5061 7611 5063
rect 7243 5056 7616 5061
rect 7243 5038 7589 5056
rect 7609 5038 7616 5056
rect 7243 5033 7616 5038
rect 7587 5031 7616 5033
rect 5962 4865 5967 4885
rect 5988 4865 5994 4885
rect 5962 4858 5994 4865
rect 6171 4887 6211 4892
rect 6171 4866 6183 4887
rect 6205 4866 6211 4887
rect 6171 4854 6211 4866
rect 6385 4888 6441 4893
rect 6385 4868 6392 4888
rect 6412 4868 6441 4888
rect 6385 4861 6441 4868
rect 6498 4962 7455 4981
rect 6385 4860 6420 4861
rect 4086 4821 4121 4822
rect 3051 4701 4008 4720
rect 4065 4814 4121 4821
rect 4065 4794 4094 4814
rect 4114 4794 4121 4814
rect 4065 4789 4121 4794
rect 4295 4816 4335 4828
rect 4295 4795 4301 4816
rect 4323 4795 4335 4816
rect 4295 4790 4335 4795
rect 4512 4817 4544 4824
rect 4512 4797 4518 4817
rect 4539 4797 4544 4817
rect 2649 4644 2734 4647
rect 2642 4640 2734 4644
rect 2642 4639 3023 4640
rect 2642 4609 2649 4639
rect 2686 4610 3023 4639
rect 2686 4609 2734 4610
rect 2642 4607 2734 4609
rect 2642 4604 2727 4607
rect 2988 4572 3023 4610
rect 4065 4583 4099 4789
rect 4512 4769 4544 4797
rect 6177 4822 6205 4854
rect 6498 4822 6529 4962
rect 7418 4946 7453 4962
rect 7418 4926 7425 4946
rect 7445 4926 7453 4946
rect 7418 4918 7453 4926
rect 6177 4791 6529 4822
rect 6974 4853 7006 4860
rect 6974 4833 6981 4853
rect 7002 4833 7006 4853
rect 4132 4761 4544 4769
rect 4132 4735 4138 4761
rect 4164 4735 4544 4761
rect 4132 4733 4544 4735
rect 4134 4732 4174 4733
rect 4512 4668 4544 4733
rect 6974 4768 7006 4833
rect 7344 4768 7384 4769
rect 6974 4766 7386 4768
rect 6974 4740 7354 4766
rect 7380 4740 7386 4766
rect 6974 4732 7386 4740
rect 6408 4717 6440 4718
rect 6405 4712 6440 4717
rect 6405 4692 6412 4712
rect 6432 4692 6440 4712
rect 6405 4684 6440 4692
rect 4512 4648 4516 4668
rect 4537 4648 4544 4668
rect 4512 4641 4544 4648
rect 5961 4619 5993 4626
rect 5961 4599 5968 4619
rect 5989 4599 5993 4619
rect 4065 4575 4100 4583
rect 2779 4570 2814 4571
rect 885 4400 1300 4429
rect 2438 4428 2471 4429
rect 2435 4423 2471 4428
rect 2435 4403 2442 4423
rect 2462 4403 2471 4423
rect 885 4399 1294 4400
rect 2435 4398 2471 4403
rect 2758 4563 2814 4570
rect 2758 4543 2787 4563
rect 2807 4543 2814 4563
rect 2758 4538 2814 4543
rect 2983 4563 3032 4572
rect 2983 4544 2991 4563
rect 3017 4544 3032 4563
rect 2435 4395 2470 4398
rect 1991 4330 2023 4337
rect 1991 4310 1998 4330
rect 2019 4310 2023 4330
rect 1991 4245 2023 4310
rect 2361 4245 2401 4246
rect 1991 4243 2403 4245
rect 1991 4217 2371 4243
rect 2397 4217 2403 4243
rect 1991 4209 2403 4217
rect 1991 4181 2023 4209
rect 1131 4177 1163 4178
rect 1128 4172 1163 4177
rect 1128 4152 1135 4172
rect 1155 4152 1163 4172
rect 1991 4161 1996 4181
rect 2017 4161 2023 4181
rect 1991 4154 2023 4161
rect 2196 4183 2245 4193
rect 2436 4189 2470 4395
rect 2758 4332 2792 4538
rect 2983 4534 3032 4544
rect 3205 4566 3237 4573
rect 3205 4546 3211 4566
rect 3232 4546 3237 4566
rect 4065 4555 4073 4575
rect 4093 4555 4100 4575
rect 4065 4550 4100 4555
rect 4065 4549 4097 4550
rect 3205 4518 3237 4546
rect 2825 4510 3237 4518
rect 2825 4484 2831 4510
rect 2857 4484 3237 4510
rect 2825 4482 3237 4484
rect 2827 4481 2867 4482
rect 3205 4417 3237 4482
rect 5961 4534 5993 4599
rect 6331 4534 6371 4535
rect 5961 4532 6373 4534
rect 5961 4506 6341 4532
rect 6367 4506 6373 4532
rect 5961 4498 6373 4506
rect 5961 4470 5993 4498
rect 5961 4450 5966 4470
rect 5987 4450 5993 4470
rect 5961 4443 5993 4450
rect 6161 4470 6211 4479
rect 6406 4478 6440 4684
rect 6974 4704 7006 4732
rect 6974 4684 6979 4704
rect 7000 4684 7006 4704
rect 7179 4706 7221 4715
rect 7419 4712 7453 4918
rect 7179 4692 7189 4706
rect 6974 4677 7006 4684
rect 7178 4686 7189 4692
rect 7213 4686 7221 4706
rect 7178 4675 7221 4686
rect 7397 4707 7453 4712
rect 7397 4687 7404 4707
rect 7424 4687 7453 4707
rect 7397 4680 7453 4687
rect 7397 4679 7432 4680
rect 7178 4645 7218 4675
rect 7068 4637 7104 4641
rect 7068 4618 7076 4637
rect 7096 4618 7104 4637
rect 7068 4615 7104 4618
rect 7178 4640 7525 4645
rect 7069 4587 7103 4615
rect 7178 4614 7497 4640
rect 7516 4614 7525 4640
rect 7178 4610 7525 4614
rect 6161 4449 6173 4470
rect 6195 4449 6211 4470
rect 6161 4441 6211 4449
rect 6384 4473 6440 4478
rect 6384 4453 6391 4473
rect 6411 4453 6440 4473
rect 6384 4446 6440 4453
rect 6541 4559 7104 4587
rect 6384 4445 6419 4446
rect 3205 4397 3209 4417
rect 3230 4397 3237 4417
rect 3205 4390 3237 4397
rect 6166 4408 6207 4441
rect 6541 4408 6581 4559
rect 7720 4408 7752 6061
rect 8117 5608 8152 6202
rect 9201 6083 9241 6234
rect 9575 6201 9616 6234
rect 9363 6196 9398 6197
rect 8678 6055 9241 6083
rect 9342 6189 9398 6196
rect 9342 6169 9371 6189
rect 9391 6169 9398 6189
rect 9342 6164 9398 6169
rect 9571 6193 9621 6201
rect 9571 6172 9587 6193
rect 9609 6172 9621 6193
rect 8257 6028 8604 6032
rect 8257 6002 8266 6028
rect 8285 6002 8604 6028
rect 8679 6027 8713 6055
rect 8257 5997 8604 6002
rect 8678 6024 8714 6027
rect 8678 6005 8686 6024
rect 8706 6005 8714 6024
rect 8678 6001 8714 6005
rect 8564 5967 8604 5997
rect 8350 5962 8385 5963
rect 8329 5955 8385 5962
rect 8329 5935 8358 5955
rect 8378 5935 8385 5955
rect 8329 5930 8385 5935
rect 8561 5956 8604 5967
rect 8561 5936 8569 5956
rect 8593 5950 8604 5956
rect 8776 5958 8808 5965
rect 8593 5936 8603 5950
rect 8329 5724 8363 5930
rect 8561 5927 8603 5936
rect 8776 5938 8782 5958
rect 8803 5938 8808 5958
rect 8776 5910 8808 5938
rect 9342 5958 9376 6164
rect 9571 6163 9621 6172
rect 9789 6192 9821 6199
rect 9789 6172 9795 6192
rect 9816 6172 9821 6192
rect 9789 6144 9821 6172
rect 9409 6136 9821 6144
rect 9409 6110 9415 6136
rect 9441 6110 9821 6136
rect 9409 6108 9821 6110
rect 9411 6107 9451 6108
rect 9789 6043 9821 6108
rect 9789 6023 9793 6043
rect 9814 6023 9821 6043
rect 9789 6016 9821 6023
rect 9342 5950 9377 5958
rect 9342 5930 9350 5950
rect 9370 5930 9377 5950
rect 9342 5925 9377 5930
rect 9342 5924 9374 5925
rect 8396 5902 8808 5910
rect 8396 5876 8402 5902
rect 8428 5876 8808 5902
rect 8396 5874 8808 5876
rect 8398 5873 8438 5874
rect 8776 5809 8808 5874
rect 8776 5789 8780 5809
rect 8801 5789 8808 5809
rect 8776 5782 8808 5789
rect 9253 5820 9605 5851
rect 8329 5716 8364 5724
rect 8329 5696 8337 5716
rect 8357 5696 8364 5716
rect 8329 5680 8364 5696
rect 9253 5680 9284 5820
rect 9577 5788 9605 5820
rect 9362 5781 9397 5782
rect 8327 5661 9284 5680
rect 9341 5774 9397 5781
rect 9341 5754 9370 5774
rect 9390 5754 9397 5774
rect 9341 5749 9397 5754
rect 9571 5776 9611 5788
rect 9571 5755 9577 5776
rect 9599 5755 9611 5776
rect 9571 5750 9611 5755
rect 9788 5777 9820 5784
rect 9788 5757 9794 5777
rect 9815 5757 9820 5777
rect 8117 5579 8547 5608
rect 8117 5574 8201 5579
rect 8300 5542 8335 5543
rect 8279 5535 8335 5542
rect 8279 5515 8308 5535
rect 8328 5515 8335 5535
rect 8279 5510 8335 5515
rect 8509 5536 8547 5579
rect 8509 5519 8514 5536
rect 8538 5519 8547 5536
rect 8279 5306 8313 5510
rect 8509 5507 8547 5519
rect 8726 5538 8758 5545
rect 8726 5518 8732 5538
rect 8753 5518 8758 5538
rect 8726 5490 8758 5518
rect 9341 5543 9375 5749
rect 9788 5729 9820 5757
rect 9408 5721 9820 5729
rect 9408 5695 9414 5721
rect 9440 5695 9820 5721
rect 9408 5693 9820 5695
rect 9410 5692 9450 5693
rect 9788 5628 9820 5693
rect 9788 5608 9792 5628
rect 9813 5608 9820 5628
rect 9788 5601 9820 5608
rect 9341 5535 9376 5543
rect 9341 5515 9349 5535
rect 9369 5515 9376 5535
rect 9341 5510 9376 5515
rect 9341 5509 9373 5510
rect 8346 5482 8758 5490
rect 8346 5456 8352 5482
rect 8378 5456 8758 5482
rect 8346 5454 8758 5456
rect 8348 5453 8388 5454
rect 8726 5389 8758 5454
rect 8726 5369 8730 5389
rect 8751 5369 8758 5389
rect 8726 5362 8758 5369
rect 8277 5296 8317 5306
rect 8277 5276 8287 5296
rect 8307 5276 8317 5296
rect 9212 5282 9621 5283
rect 8277 5052 8317 5276
rect 9206 5253 9621 5282
rect 9206 5102 9246 5253
rect 9580 5220 9621 5253
rect 9368 5215 9403 5216
rect 8683 5074 9246 5102
rect 9347 5208 9403 5215
rect 9347 5188 9376 5208
rect 9396 5188 9403 5208
rect 9347 5183 9403 5188
rect 9576 5212 9626 5220
rect 9576 5191 9592 5212
rect 9614 5191 9626 5212
rect 8277 5018 8604 5052
rect 8684 5046 8718 5074
rect 8683 5043 8719 5046
rect 8683 5024 8691 5043
rect 8711 5024 8719 5043
rect 8683 5020 8719 5024
rect 8294 5017 8604 5018
rect 8569 4988 8604 5017
rect 8355 4981 8390 4982
rect 8334 4974 8390 4981
rect 8334 4954 8363 4974
rect 8383 4954 8390 4974
rect 8334 4949 8390 4954
rect 8564 4976 8606 4988
rect 8564 4956 8573 4976
rect 8597 4956 8606 4976
rect 8334 4743 8368 4949
rect 8564 4948 8606 4956
rect 8781 4977 8813 4984
rect 8781 4957 8787 4977
rect 8808 4957 8813 4977
rect 8781 4929 8813 4957
rect 9347 4977 9381 5183
rect 9576 5182 9626 5191
rect 9794 5211 9826 5218
rect 9794 5191 9800 5211
rect 9821 5191 9826 5211
rect 9794 5163 9826 5191
rect 9414 5155 9826 5163
rect 9414 5129 9420 5155
rect 9446 5129 9826 5155
rect 9414 5127 9826 5129
rect 9416 5126 9456 5127
rect 9794 5062 9826 5127
rect 9794 5042 9798 5062
rect 9819 5042 9826 5062
rect 9794 5035 9826 5042
rect 9347 4969 9382 4977
rect 9347 4949 9355 4969
rect 9375 4949 9382 4969
rect 9347 4944 9382 4949
rect 9347 4943 9379 4944
rect 8401 4921 8813 4929
rect 8401 4895 8407 4921
rect 8433 4895 8813 4921
rect 8401 4893 8813 4895
rect 8403 4892 8443 4893
rect 8781 4828 8813 4893
rect 8781 4808 8785 4828
rect 8806 4808 8813 4828
rect 8781 4801 8813 4808
rect 9258 4839 9610 4870
rect 8334 4735 8369 4743
rect 8334 4715 8342 4735
rect 8362 4715 8369 4735
rect 8334 4699 8369 4715
rect 9258 4699 9289 4839
rect 9582 4807 9610 4839
rect 9367 4800 9402 4801
rect 8332 4680 9289 4699
rect 9346 4793 9402 4800
rect 9346 4773 9375 4793
rect 9395 4773 9402 4793
rect 9346 4768 9402 4773
rect 9576 4795 9616 4807
rect 9576 4774 9582 4795
rect 9604 4774 9616 4795
rect 9576 4769 9616 4774
rect 9793 4796 9825 4803
rect 9793 4776 9799 4796
rect 9820 4776 9825 4796
rect 7930 4623 8015 4626
rect 7923 4619 8015 4623
rect 7923 4618 8304 4619
rect 7923 4588 7930 4618
rect 7967 4589 8304 4618
rect 7967 4588 8015 4589
rect 7923 4586 8015 4588
rect 7923 4583 8008 4586
rect 8269 4551 8304 4589
rect 9346 4562 9380 4768
rect 9793 4748 9825 4776
rect 9413 4740 9825 4748
rect 9413 4714 9419 4740
rect 9445 4714 9825 4740
rect 9413 4712 9825 4714
rect 9415 4711 9455 4712
rect 9793 4647 9825 4712
rect 9793 4627 9797 4647
rect 9818 4627 9825 4647
rect 9793 4620 9825 4627
rect 9346 4554 9381 4562
rect 8060 4549 8095 4550
rect 6166 4379 6581 4408
rect 7719 4407 7752 4408
rect 7716 4402 7752 4407
rect 7716 4382 7723 4402
rect 7743 4382 7752 4402
rect 6166 4378 6575 4379
rect 7716 4377 7752 4382
rect 8039 4542 8095 4549
rect 8039 4522 8068 4542
rect 8088 4522 8095 4542
rect 8039 4517 8095 4522
rect 8264 4542 8313 4551
rect 8264 4523 8272 4542
rect 8298 4523 8313 4542
rect 7716 4374 7751 4377
rect 2758 4329 2793 4332
rect 2196 4164 2211 4183
rect 2237 4164 2245 4183
rect 2196 4155 2245 4164
rect 2414 4184 2470 4189
rect 2414 4164 2421 4184
rect 2441 4164 2470 4184
rect 2414 4157 2470 4164
rect 2757 4324 2793 4329
rect 3934 4327 4343 4328
rect 2757 4304 2766 4324
rect 2786 4304 2793 4324
rect 2757 4299 2793 4304
rect 2757 4298 2790 4299
rect 3928 4298 4343 4327
rect 2414 4156 2449 4157
rect 1128 4144 1163 4152
rect 684 4079 716 4086
rect 684 4059 691 4079
rect 712 4059 716 4079
rect 684 3994 716 4059
rect 1054 3994 1094 3995
rect 684 3992 1096 3994
rect 684 3966 1064 3992
rect 1090 3966 1096 3992
rect 684 3958 1096 3966
rect 684 3930 716 3958
rect 1129 3938 1163 4144
rect 2205 4117 2240 4155
rect 2463 4117 2586 4122
rect 2205 4116 2586 4117
rect 2205 4088 2548 4116
rect 2582 4115 2586 4116
rect 2582 4088 2587 4115
rect 2205 4087 2587 4088
rect 2463 4082 2587 4087
rect 684 3910 689 3930
rect 710 3910 716 3930
rect 684 3903 716 3910
rect 893 3932 933 3937
rect 893 3911 905 3932
rect 927 3911 933 3932
rect 893 3899 933 3911
rect 1107 3933 1163 3938
rect 1107 3913 1114 3933
rect 1134 3913 1163 3933
rect 1107 3906 1163 3913
rect 1220 4007 2177 4026
rect 1107 3905 1142 3906
rect 899 3867 927 3899
rect 1220 3867 1251 4007
rect 2140 3991 2175 4007
rect 2140 3971 2147 3991
rect 2167 3971 2175 3991
rect 2140 3963 2175 3971
rect 899 3836 1251 3867
rect 1696 3898 1728 3905
rect 1696 3878 1703 3898
rect 1724 3878 1728 3898
rect 1696 3813 1728 3878
rect 2066 3813 2106 3814
rect 1696 3811 2108 3813
rect 1696 3785 2076 3811
rect 2102 3785 2108 3811
rect 1696 3777 2108 3785
rect 1130 3762 1162 3763
rect 1127 3757 1162 3762
rect 1127 3737 1134 3757
rect 1154 3737 1162 3757
rect 1127 3729 1162 3737
rect 683 3664 715 3671
rect 683 3644 690 3664
rect 711 3644 715 3664
rect 683 3579 715 3644
rect 1053 3579 1093 3580
rect 683 3577 1095 3579
rect 683 3551 1063 3577
rect 1089 3551 1095 3577
rect 683 3543 1095 3551
rect 683 3515 715 3543
rect 683 3495 688 3515
rect 709 3495 715 3515
rect 683 3488 715 3495
rect 883 3515 933 3524
rect 1128 3523 1162 3729
rect 1696 3749 1728 3777
rect 1696 3729 1701 3749
rect 1722 3729 1728 3749
rect 1696 3722 1728 3729
rect 1903 3750 1945 3758
rect 2141 3757 2175 3963
rect 1903 3730 1912 3750
rect 1936 3730 1945 3750
rect 1903 3718 1945 3730
rect 2119 3752 2175 3757
rect 2119 3732 2126 3752
rect 2146 3732 2175 3752
rect 2119 3725 2175 3732
rect 2119 3724 2154 3725
rect 1905 3689 1940 3718
rect 1905 3688 2215 3689
rect 1790 3682 1826 3686
rect 1790 3663 1798 3682
rect 1818 3663 1826 3682
rect 1790 3660 1826 3663
rect 1791 3632 1825 3660
rect 1905 3654 2232 3688
rect 883 3494 895 3515
rect 917 3494 933 3515
rect 883 3486 933 3494
rect 1106 3518 1162 3523
rect 1106 3498 1113 3518
rect 1133 3498 1162 3518
rect 1106 3491 1162 3498
rect 1263 3604 1826 3632
rect 1106 3490 1141 3491
rect 888 3453 929 3486
rect 1263 3453 1303 3604
rect 888 3424 1303 3453
rect 2192 3430 2232 3654
rect 888 3423 1297 3424
rect 2192 3410 2202 3430
rect 2222 3410 2232 3430
rect 2192 3400 2232 3410
rect 1751 3337 1783 3344
rect 1751 3317 1758 3337
rect 1779 3317 1783 3337
rect 1751 3252 1783 3317
rect 2121 3252 2161 3253
rect 1751 3250 2163 3252
rect 1751 3224 2131 3250
rect 2157 3224 2163 3250
rect 1751 3216 2163 3224
rect 1136 3196 1168 3197
rect 1133 3191 1168 3196
rect 1133 3171 1140 3191
rect 1160 3171 1168 3191
rect 1133 3163 1168 3171
rect 689 3098 721 3105
rect 689 3078 696 3098
rect 717 3078 721 3098
rect 689 3013 721 3078
rect 1059 3013 1099 3014
rect 689 3011 1101 3013
rect 689 2985 1069 3011
rect 1095 2985 1101 3011
rect 689 2977 1101 2985
rect 689 2949 721 2977
rect 1134 2957 1168 3163
rect 1751 3188 1783 3216
rect 1751 3168 1756 3188
rect 1777 3168 1783 3188
rect 1751 3161 1783 3168
rect 1962 3187 2000 3199
rect 2196 3196 2230 3400
rect 1962 3170 1971 3187
rect 1995 3170 2000 3187
rect 1962 3127 2000 3170
rect 2174 3191 2230 3196
rect 2174 3171 2181 3191
rect 2201 3171 2230 3191
rect 2174 3164 2230 3171
rect 2174 3163 2209 3164
rect 2308 3127 2392 3132
rect 1962 3098 2392 3127
rect 689 2929 694 2949
rect 715 2929 721 2949
rect 689 2922 721 2929
rect 898 2951 938 2956
rect 898 2930 910 2951
rect 932 2930 938 2951
rect 898 2918 938 2930
rect 1112 2952 1168 2957
rect 1112 2932 1119 2952
rect 1139 2932 1168 2952
rect 1112 2925 1168 2932
rect 1225 3026 2182 3045
rect 1112 2924 1147 2925
rect 904 2886 932 2918
rect 1225 2886 1256 3026
rect 2145 3010 2180 3026
rect 2145 2990 2152 3010
rect 2172 2990 2180 3010
rect 2145 2982 2180 2990
rect 904 2855 1256 2886
rect 1701 2917 1733 2924
rect 1701 2897 1708 2917
rect 1729 2897 1733 2917
rect 1701 2832 1733 2897
rect 2071 2832 2111 2833
rect 1701 2830 2113 2832
rect 1701 2804 2081 2830
rect 2107 2804 2113 2830
rect 1701 2796 2113 2804
rect 1135 2781 1167 2782
rect 1132 2776 1167 2781
rect 1132 2756 1139 2776
rect 1159 2756 1167 2776
rect 1132 2748 1167 2756
rect 688 2683 720 2690
rect 688 2663 695 2683
rect 716 2663 720 2683
rect 688 2598 720 2663
rect 1058 2598 1098 2599
rect 688 2596 1100 2598
rect 688 2570 1068 2596
rect 1094 2570 1100 2596
rect 688 2562 1100 2570
rect 688 2534 720 2562
rect 688 2514 693 2534
rect 714 2514 720 2534
rect 688 2507 720 2514
rect 888 2534 938 2543
rect 1133 2542 1167 2748
rect 1701 2768 1733 2796
rect 1701 2748 1706 2768
rect 1727 2748 1733 2768
rect 1906 2770 1948 2779
rect 2146 2776 2180 2982
rect 1906 2756 1916 2770
rect 1701 2741 1733 2748
rect 1905 2750 1916 2756
rect 1940 2750 1948 2770
rect 1905 2739 1948 2750
rect 2124 2771 2180 2776
rect 2124 2751 2131 2771
rect 2151 2751 2180 2771
rect 2124 2744 2180 2751
rect 2124 2743 2159 2744
rect 1905 2709 1945 2739
rect 1795 2701 1831 2705
rect 1795 2682 1803 2701
rect 1823 2682 1831 2701
rect 1795 2679 1831 2682
rect 1905 2704 2252 2709
rect 1796 2651 1830 2679
rect 1905 2678 2224 2704
rect 2243 2678 2252 2704
rect 1905 2674 2252 2678
rect 888 2513 900 2534
rect 922 2513 938 2534
rect 888 2505 938 2513
rect 1111 2537 1167 2542
rect 1111 2517 1118 2537
rect 1138 2517 1167 2537
rect 1111 2510 1167 2517
rect 1268 2623 1831 2651
rect 1111 2509 1146 2510
rect 893 2472 934 2505
rect 1268 2472 1308 2623
rect 2357 2504 2392 3098
rect 2757 2645 2789 4298
rect 3928 4147 3968 4298
rect 4302 4265 4343 4298
rect 7272 4309 7304 4316
rect 7272 4289 7279 4309
rect 7300 4289 7304 4309
rect 4090 4260 4125 4261
rect 3405 4119 3968 4147
rect 4069 4253 4125 4260
rect 4069 4233 4098 4253
rect 4118 4233 4125 4253
rect 4069 4228 4125 4233
rect 4298 4257 4348 4265
rect 4298 4236 4314 4257
rect 4336 4236 4348 4257
rect 2984 4092 3331 4096
rect 2984 4066 2993 4092
rect 3012 4066 3331 4092
rect 3406 4091 3440 4119
rect 2984 4061 3331 4066
rect 3405 4088 3441 4091
rect 3405 4069 3413 4088
rect 3433 4069 3441 4088
rect 3405 4065 3441 4069
rect 3291 4031 3331 4061
rect 3077 4026 3112 4027
rect 3056 4019 3112 4026
rect 3056 3999 3085 4019
rect 3105 3999 3112 4019
rect 3056 3994 3112 3999
rect 3288 4020 3331 4031
rect 3288 4000 3296 4020
rect 3320 4014 3331 4020
rect 3503 4022 3535 4029
rect 3320 4000 3330 4014
rect 3056 3788 3090 3994
rect 3288 3991 3330 4000
rect 3503 4002 3509 4022
rect 3530 4002 3535 4022
rect 3503 3974 3535 4002
rect 4069 4022 4103 4228
rect 4298 4227 4348 4236
rect 4516 4256 4548 4263
rect 4516 4236 4522 4256
rect 4543 4236 4548 4256
rect 4516 4208 4548 4236
rect 4136 4200 4548 4208
rect 4136 4174 4142 4200
rect 4168 4174 4548 4200
rect 4136 4172 4548 4174
rect 4138 4171 4178 4172
rect 4516 4107 4548 4172
rect 7272 4224 7304 4289
rect 7642 4224 7682 4225
rect 7272 4222 7684 4224
rect 7272 4196 7652 4222
rect 7678 4196 7684 4222
rect 7272 4188 7684 4196
rect 7272 4160 7304 4188
rect 6412 4156 6444 4157
rect 6409 4151 6444 4156
rect 6409 4131 6416 4151
rect 6436 4131 6444 4151
rect 7272 4140 7277 4160
rect 7298 4140 7304 4160
rect 7272 4133 7304 4140
rect 7477 4162 7526 4172
rect 7717 4168 7751 4374
rect 8039 4311 8073 4517
rect 8264 4513 8313 4523
rect 8486 4545 8518 4552
rect 8486 4525 8492 4545
rect 8513 4525 8518 4545
rect 9346 4534 9354 4554
rect 9374 4534 9381 4554
rect 9346 4529 9381 4534
rect 9346 4528 9378 4529
rect 8486 4497 8518 4525
rect 8106 4489 8518 4497
rect 8106 4463 8112 4489
rect 8138 4463 8518 4489
rect 8106 4461 8518 4463
rect 8108 4460 8148 4461
rect 8486 4396 8518 4461
rect 8486 4376 8490 4396
rect 8511 4376 8518 4396
rect 8486 4369 8518 4376
rect 8039 4308 8074 4311
rect 7477 4143 7492 4162
rect 7518 4143 7526 4162
rect 7477 4134 7526 4143
rect 7695 4163 7751 4168
rect 7695 4143 7702 4163
rect 7722 4143 7751 4163
rect 7695 4136 7751 4143
rect 8038 4303 8074 4308
rect 9215 4306 9624 4307
rect 8038 4283 8047 4303
rect 8067 4283 8074 4303
rect 8038 4278 8074 4283
rect 8038 4277 8071 4278
rect 9209 4277 9624 4306
rect 7695 4135 7730 4136
rect 6409 4123 6444 4131
rect 4516 4087 4520 4107
rect 4541 4087 4548 4107
rect 4516 4080 4548 4087
rect 5965 4058 5997 4065
rect 5965 4038 5972 4058
rect 5993 4038 5997 4058
rect 4069 4014 4104 4022
rect 4069 3994 4077 4014
rect 4097 3994 4104 4014
rect 4069 3989 4104 3994
rect 4069 3988 4101 3989
rect 3123 3966 3535 3974
rect 3123 3940 3129 3966
rect 3155 3940 3535 3966
rect 3123 3938 3535 3940
rect 3125 3937 3165 3938
rect 3503 3873 3535 3938
rect 5965 3973 5997 4038
rect 6335 3973 6375 3974
rect 5965 3971 6377 3973
rect 5965 3945 6345 3971
rect 6371 3945 6377 3971
rect 5965 3937 6377 3945
rect 3503 3853 3507 3873
rect 3528 3853 3535 3873
rect 3503 3846 3535 3853
rect 3980 3884 4332 3915
rect 3056 3780 3091 3788
rect 3056 3760 3064 3780
rect 3084 3760 3091 3780
rect 3056 3744 3091 3760
rect 3980 3744 4011 3884
rect 4304 3852 4332 3884
rect 5965 3909 5997 3937
rect 6410 3917 6444 4123
rect 7486 4096 7521 4134
rect 7744 4096 7867 4101
rect 7486 4095 7867 4096
rect 7486 4067 7829 4095
rect 7863 4094 7867 4095
rect 7863 4067 7868 4094
rect 7486 4066 7868 4067
rect 7744 4061 7868 4066
rect 5965 3889 5970 3909
rect 5991 3889 5997 3909
rect 5965 3882 5997 3889
rect 6174 3911 6214 3916
rect 6174 3890 6186 3911
rect 6208 3890 6214 3911
rect 6174 3878 6214 3890
rect 6388 3912 6444 3917
rect 6388 3892 6395 3912
rect 6415 3892 6444 3912
rect 6388 3885 6444 3892
rect 6501 3986 7458 4005
rect 6388 3884 6423 3885
rect 4089 3845 4124 3846
rect 3054 3725 4011 3744
rect 4068 3838 4124 3845
rect 4068 3818 4097 3838
rect 4117 3818 4124 3838
rect 4068 3813 4124 3818
rect 4298 3840 4338 3852
rect 4298 3819 4304 3840
rect 4326 3819 4338 3840
rect 4298 3814 4338 3819
rect 4515 3841 4547 3848
rect 4515 3821 4521 3841
rect 4542 3821 4547 3841
rect 2893 3673 2922 3675
rect 2893 3668 3266 3673
rect 2893 3650 2900 3668
rect 2920 3650 3266 3668
rect 2893 3645 3266 3650
rect 2898 3643 3266 3645
rect 3027 3606 3062 3607
rect 3242 3606 3266 3643
rect 3006 3599 3062 3606
rect 3006 3579 3035 3599
rect 3055 3579 3062 3599
rect 3006 3574 3062 3579
rect 3237 3601 3274 3606
rect 3237 3582 3245 3601
rect 3268 3582 3274 3601
rect 3237 3576 3274 3582
rect 3453 3602 3485 3609
rect 3453 3582 3459 3602
rect 3480 3582 3485 3602
rect 3006 3370 3040 3574
rect 3453 3554 3485 3582
rect 4068 3607 4102 3813
rect 4515 3793 4547 3821
rect 6180 3846 6208 3878
rect 6501 3846 6532 3986
rect 7421 3970 7456 3986
rect 7421 3950 7428 3970
rect 7448 3950 7456 3970
rect 7421 3942 7456 3950
rect 6180 3815 6532 3846
rect 6977 3877 7009 3884
rect 6977 3857 6984 3877
rect 7005 3857 7009 3877
rect 4135 3785 4547 3793
rect 4135 3759 4141 3785
rect 4167 3759 4547 3785
rect 4135 3757 4547 3759
rect 4137 3756 4177 3757
rect 4515 3692 4547 3757
rect 6977 3792 7009 3857
rect 7347 3792 7387 3793
rect 6977 3790 7389 3792
rect 6977 3764 7357 3790
rect 7383 3764 7389 3790
rect 6977 3756 7389 3764
rect 6411 3741 6443 3742
rect 6408 3736 6443 3741
rect 6408 3716 6415 3736
rect 6435 3716 6443 3736
rect 6408 3708 6443 3716
rect 4515 3672 4519 3692
rect 4540 3672 4547 3692
rect 4515 3665 4547 3672
rect 5964 3643 5996 3650
rect 5964 3623 5971 3643
rect 5992 3623 5996 3643
rect 4068 3599 4103 3607
rect 4068 3579 4076 3599
rect 4096 3579 4103 3599
rect 4068 3574 4103 3579
rect 4068 3573 4100 3574
rect 3073 3546 3485 3554
rect 3073 3520 3079 3546
rect 3105 3520 3485 3546
rect 3073 3518 3485 3520
rect 3075 3517 3115 3518
rect 3453 3453 3485 3518
rect 5964 3558 5996 3623
rect 6334 3558 6374 3559
rect 5964 3556 6376 3558
rect 5964 3530 6344 3556
rect 6370 3530 6376 3556
rect 5964 3522 6376 3530
rect 5964 3494 5996 3522
rect 5964 3474 5969 3494
rect 5990 3474 5996 3494
rect 5964 3467 5996 3474
rect 6164 3494 6214 3503
rect 6409 3502 6443 3708
rect 6977 3728 7009 3756
rect 6977 3708 6982 3728
rect 7003 3708 7009 3728
rect 6977 3701 7009 3708
rect 7184 3729 7226 3737
rect 7422 3736 7456 3942
rect 7184 3709 7193 3729
rect 7217 3709 7226 3729
rect 7184 3697 7226 3709
rect 7400 3731 7456 3736
rect 7400 3711 7407 3731
rect 7427 3711 7456 3731
rect 7400 3704 7456 3711
rect 7400 3703 7435 3704
rect 7186 3668 7221 3697
rect 7186 3667 7496 3668
rect 7071 3661 7107 3665
rect 7071 3642 7079 3661
rect 7099 3642 7107 3661
rect 7071 3639 7107 3642
rect 7072 3611 7106 3639
rect 7186 3633 7513 3667
rect 6164 3473 6176 3494
rect 6198 3473 6214 3494
rect 6164 3465 6214 3473
rect 6387 3497 6443 3502
rect 6387 3477 6394 3497
rect 6414 3477 6443 3497
rect 6387 3470 6443 3477
rect 6544 3583 7107 3611
rect 6387 3469 6422 3470
rect 3453 3433 3457 3453
rect 3478 3433 3485 3453
rect 3453 3426 3485 3433
rect 6169 3432 6210 3465
rect 6544 3432 6584 3583
rect 6169 3403 6584 3432
rect 7473 3409 7513 3633
rect 6169 3402 6578 3403
rect 7473 3389 7483 3409
rect 7503 3389 7513 3409
rect 7473 3379 7513 3389
rect 3004 3360 3044 3370
rect 3004 3340 3014 3360
rect 3034 3340 3044 3360
rect 3939 3346 4348 3347
rect 3004 3116 3044 3340
rect 3933 3317 4348 3346
rect 3933 3166 3973 3317
rect 4307 3284 4348 3317
rect 7032 3316 7064 3323
rect 7032 3296 7039 3316
rect 7060 3296 7064 3316
rect 4095 3279 4130 3280
rect 3410 3138 3973 3166
rect 4074 3272 4130 3279
rect 4074 3252 4103 3272
rect 4123 3252 4130 3272
rect 4074 3247 4130 3252
rect 4303 3276 4353 3284
rect 4303 3255 4319 3276
rect 4341 3255 4353 3276
rect 3004 3082 3331 3116
rect 3411 3110 3445 3138
rect 3410 3107 3446 3110
rect 3410 3088 3418 3107
rect 3438 3088 3446 3107
rect 3410 3084 3446 3088
rect 3021 3081 3331 3082
rect 3296 3052 3331 3081
rect 3082 3045 3117 3046
rect 3061 3038 3117 3045
rect 3061 3018 3090 3038
rect 3110 3018 3117 3038
rect 3061 3013 3117 3018
rect 3291 3040 3333 3052
rect 3291 3020 3300 3040
rect 3324 3020 3333 3040
rect 3061 2807 3095 3013
rect 3291 3012 3333 3020
rect 3508 3041 3540 3048
rect 3508 3021 3514 3041
rect 3535 3021 3540 3041
rect 3508 2993 3540 3021
rect 4074 3041 4108 3247
rect 4303 3246 4353 3255
rect 4521 3275 4553 3282
rect 4521 3255 4527 3275
rect 4548 3255 4553 3275
rect 4521 3227 4553 3255
rect 4141 3219 4553 3227
rect 4141 3193 4147 3219
rect 4173 3193 4553 3219
rect 4141 3191 4553 3193
rect 4143 3190 4183 3191
rect 4521 3126 4553 3191
rect 7032 3231 7064 3296
rect 7402 3231 7442 3232
rect 7032 3229 7444 3231
rect 7032 3203 7412 3229
rect 7438 3203 7444 3229
rect 7032 3195 7444 3203
rect 6417 3175 6449 3176
rect 6414 3170 6449 3175
rect 6414 3150 6421 3170
rect 6441 3150 6449 3170
rect 6414 3142 6449 3150
rect 4521 3106 4525 3126
rect 4546 3106 4553 3126
rect 4521 3099 4553 3106
rect 5970 3077 6002 3084
rect 5970 3057 5977 3077
rect 5998 3057 6002 3077
rect 4074 3033 4109 3041
rect 4074 3013 4082 3033
rect 4102 3013 4109 3033
rect 4074 3008 4109 3013
rect 4074 3007 4106 3008
rect 3128 2985 3540 2993
rect 3128 2959 3134 2985
rect 3160 2959 3540 2985
rect 3128 2957 3540 2959
rect 3130 2956 3170 2957
rect 3508 2892 3540 2957
rect 5970 2992 6002 3057
rect 6340 2992 6380 2993
rect 5970 2990 6382 2992
rect 5970 2964 6350 2990
rect 6376 2964 6382 2990
rect 5970 2956 6382 2964
rect 3508 2872 3512 2892
rect 3533 2872 3540 2892
rect 3508 2865 3540 2872
rect 3985 2903 4337 2934
rect 3061 2799 3096 2807
rect 3061 2779 3069 2799
rect 3089 2779 3096 2799
rect 3061 2763 3096 2779
rect 3985 2763 4016 2903
rect 4309 2871 4337 2903
rect 5970 2928 6002 2956
rect 6415 2936 6449 3142
rect 7032 3167 7064 3195
rect 7032 3147 7037 3167
rect 7058 3147 7064 3167
rect 7032 3140 7064 3147
rect 7243 3166 7281 3178
rect 7477 3175 7511 3379
rect 7243 3149 7252 3166
rect 7276 3149 7281 3166
rect 7243 3106 7281 3149
rect 7455 3170 7511 3175
rect 7455 3150 7462 3170
rect 7482 3150 7511 3170
rect 7455 3143 7511 3150
rect 7455 3142 7490 3143
rect 7589 3106 7673 3111
rect 7243 3077 7673 3106
rect 5970 2908 5975 2928
rect 5996 2908 6002 2928
rect 5970 2901 6002 2908
rect 6179 2930 6219 2935
rect 6179 2909 6191 2930
rect 6213 2909 6219 2930
rect 6179 2897 6219 2909
rect 6393 2931 6449 2936
rect 6393 2911 6400 2931
rect 6420 2911 6449 2931
rect 6393 2904 6449 2911
rect 6506 3005 7463 3024
rect 6393 2903 6428 2904
rect 4094 2864 4129 2865
rect 3059 2744 4016 2763
rect 4073 2857 4129 2864
rect 4073 2837 4102 2857
rect 4122 2837 4129 2857
rect 4073 2832 4129 2837
rect 4303 2859 4343 2871
rect 4303 2838 4309 2859
rect 4331 2838 4343 2859
rect 4303 2833 4343 2838
rect 4520 2860 4552 2867
rect 4520 2840 4526 2860
rect 4547 2840 4552 2860
rect 2753 2612 3123 2645
rect 2757 2610 2789 2612
rect 2874 2578 2909 2579
rect 2853 2571 2909 2578
rect 3086 2577 3123 2612
rect 4073 2626 4107 2832
rect 4520 2812 4552 2840
rect 6185 2865 6213 2897
rect 6506 2865 6537 3005
rect 7426 2989 7461 3005
rect 7426 2969 7433 2989
rect 7453 2969 7461 2989
rect 7426 2961 7461 2969
rect 6185 2834 6537 2865
rect 6982 2896 7014 2903
rect 6982 2876 6989 2896
rect 7010 2876 7014 2896
rect 4140 2804 4552 2812
rect 4140 2778 4146 2804
rect 4172 2778 4552 2804
rect 4140 2776 4552 2778
rect 4142 2775 4182 2776
rect 4520 2711 4552 2776
rect 6982 2811 7014 2876
rect 7352 2811 7392 2812
rect 6982 2809 7394 2811
rect 6982 2783 7362 2809
rect 7388 2783 7394 2809
rect 6982 2775 7394 2783
rect 6416 2760 6448 2761
rect 6413 2755 6448 2760
rect 6413 2735 6420 2755
rect 6440 2735 6448 2755
rect 6413 2727 6448 2735
rect 4520 2691 4524 2711
rect 4545 2691 4552 2711
rect 4520 2684 4552 2691
rect 5969 2662 6001 2669
rect 5969 2642 5976 2662
rect 5997 2642 6001 2662
rect 4073 2618 4108 2626
rect 4073 2598 4081 2618
rect 4101 2598 4108 2618
rect 4073 2593 4108 2598
rect 4073 2592 4105 2593
rect 2853 2551 2882 2571
rect 2902 2551 2909 2571
rect 2853 2546 2909 2551
rect 3081 2575 3128 2577
rect 3081 2549 3093 2575
rect 3118 2549 3128 2575
rect 2357 2498 2395 2504
rect 2357 2478 2367 2498
rect 2387 2478 2395 2498
rect 2357 2476 2395 2478
rect 893 2443 1308 2472
rect 2360 2470 2395 2476
rect 893 2442 1302 2443
rect 1916 2405 1948 2412
rect 1916 2385 1923 2405
rect 1944 2385 1948 2405
rect 1916 2320 1948 2385
rect 2286 2320 2326 2321
rect 1916 2318 2328 2320
rect 1916 2292 2296 2318
rect 2322 2292 2328 2318
rect 1916 2284 2328 2292
rect 1916 2256 1948 2284
rect 2361 2264 2395 2470
rect 2853 2340 2887 2546
rect 3081 2543 3128 2549
rect 3300 2574 3332 2581
rect 3300 2554 3306 2574
rect 3327 2554 3332 2574
rect 3300 2526 3332 2554
rect 2920 2518 3332 2526
rect 2920 2492 2926 2518
rect 2952 2492 3332 2518
rect 2920 2490 3332 2492
rect 2922 2489 2962 2490
rect 3300 2425 3332 2490
rect 5969 2577 6001 2642
rect 6339 2577 6379 2578
rect 5969 2575 6381 2577
rect 5969 2549 6349 2575
rect 6375 2549 6381 2575
rect 5969 2541 6381 2549
rect 5969 2513 6001 2541
rect 5969 2493 5974 2513
rect 5995 2493 6001 2513
rect 5969 2486 6001 2493
rect 6169 2513 6219 2522
rect 6414 2521 6448 2727
rect 6982 2747 7014 2775
rect 6982 2727 6987 2747
rect 7008 2727 7014 2747
rect 7187 2749 7229 2758
rect 7427 2755 7461 2961
rect 7187 2735 7197 2749
rect 6982 2720 7014 2727
rect 7186 2729 7197 2735
rect 7221 2729 7229 2749
rect 7186 2718 7229 2729
rect 7405 2750 7461 2755
rect 7405 2730 7412 2750
rect 7432 2730 7461 2750
rect 7405 2723 7461 2730
rect 7405 2722 7440 2723
rect 7186 2688 7226 2718
rect 7076 2680 7112 2684
rect 7076 2661 7084 2680
rect 7104 2661 7112 2680
rect 7076 2658 7112 2661
rect 7186 2683 7533 2688
rect 7077 2630 7111 2658
rect 7186 2657 7505 2683
rect 7524 2657 7533 2683
rect 7186 2653 7533 2657
rect 6169 2492 6181 2513
rect 6203 2492 6219 2513
rect 6169 2484 6219 2492
rect 6392 2516 6448 2521
rect 6392 2496 6399 2516
rect 6419 2496 6448 2516
rect 6392 2489 6448 2496
rect 6549 2602 7112 2630
rect 6392 2488 6427 2489
rect 3300 2405 3304 2425
rect 3325 2405 3332 2425
rect 6174 2451 6215 2484
rect 6549 2451 6589 2602
rect 7638 2483 7673 3077
rect 8038 2624 8070 4277
rect 9209 4126 9249 4277
rect 9583 4244 9624 4277
rect 9371 4239 9406 4240
rect 8686 4098 9249 4126
rect 9350 4232 9406 4239
rect 9350 4212 9379 4232
rect 9399 4212 9406 4232
rect 9350 4207 9406 4212
rect 9579 4236 9629 4244
rect 9579 4215 9595 4236
rect 9617 4215 9629 4236
rect 8265 4071 8612 4075
rect 8265 4045 8274 4071
rect 8293 4045 8612 4071
rect 8687 4070 8721 4098
rect 8265 4040 8612 4045
rect 8686 4067 8722 4070
rect 8686 4048 8694 4067
rect 8714 4048 8722 4067
rect 8686 4044 8722 4048
rect 8572 4010 8612 4040
rect 8358 4005 8393 4006
rect 8337 3998 8393 4005
rect 8337 3978 8366 3998
rect 8386 3978 8393 3998
rect 8337 3973 8393 3978
rect 8569 3999 8612 4010
rect 8569 3979 8577 3999
rect 8601 3993 8612 3999
rect 8784 4001 8816 4008
rect 8601 3979 8611 3993
rect 8337 3767 8371 3973
rect 8569 3970 8611 3979
rect 8784 3981 8790 4001
rect 8811 3981 8816 4001
rect 8784 3953 8816 3981
rect 9350 4001 9384 4207
rect 9579 4206 9629 4215
rect 9797 4235 9829 4242
rect 9797 4215 9803 4235
rect 9824 4215 9829 4235
rect 9797 4187 9829 4215
rect 9417 4179 9829 4187
rect 9417 4153 9423 4179
rect 9449 4153 9829 4179
rect 9417 4151 9829 4153
rect 9419 4150 9459 4151
rect 9797 4086 9829 4151
rect 9797 4066 9801 4086
rect 9822 4066 9829 4086
rect 9797 4059 9829 4066
rect 9350 3993 9385 4001
rect 9350 3973 9358 3993
rect 9378 3973 9385 3993
rect 9350 3968 9385 3973
rect 9350 3967 9382 3968
rect 8404 3945 8816 3953
rect 8404 3919 8410 3945
rect 8436 3919 8816 3945
rect 8404 3917 8816 3919
rect 8406 3916 8446 3917
rect 8784 3852 8816 3917
rect 8784 3832 8788 3852
rect 8809 3832 8816 3852
rect 8784 3825 8816 3832
rect 9261 3863 9613 3894
rect 8337 3759 8372 3767
rect 8337 3739 8345 3759
rect 8365 3739 8372 3759
rect 8337 3723 8372 3739
rect 9261 3723 9292 3863
rect 9585 3831 9613 3863
rect 9370 3824 9405 3825
rect 8335 3704 9292 3723
rect 9349 3817 9405 3824
rect 9349 3797 9378 3817
rect 9398 3797 9405 3817
rect 9349 3792 9405 3797
rect 9579 3819 9619 3831
rect 9579 3798 9585 3819
rect 9607 3798 9619 3819
rect 9579 3793 9619 3798
rect 9796 3820 9828 3827
rect 9796 3800 9802 3820
rect 9823 3800 9828 3820
rect 8174 3652 8203 3654
rect 8174 3647 8547 3652
rect 8174 3629 8181 3647
rect 8201 3629 8547 3647
rect 8174 3624 8547 3629
rect 8179 3622 8547 3624
rect 8308 3585 8343 3586
rect 8523 3585 8547 3622
rect 8287 3578 8343 3585
rect 8287 3558 8316 3578
rect 8336 3558 8343 3578
rect 8287 3553 8343 3558
rect 8518 3580 8555 3585
rect 8518 3561 8526 3580
rect 8549 3561 8555 3580
rect 8518 3555 8555 3561
rect 8734 3581 8766 3588
rect 8734 3561 8740 3581
rect 8761 3561 8766 3581
rect 8287 3349 8321 3553
rect 8734 3533 8766 3561
rect 9349 3586 9383 3792
rect 9796 3772 9828 3800
rect 9416 3764 9828 3772
rect 9416 3738 9422 3764
rect 9448 3738 9828 3764
rect 9416 3736 9828 3738
rect 9418 3735 9458 3736
rect 9796 3671 9828 3736
rect 9796 3651 9800 3671
rect 9821 3651 9828 3671
rect 9796 3644 9828 3651
rect 9349 3578 9384 3586
rect 9349 3558 9357 3578
rect 9377 3558 9384 3578
rect 9349 3553 9384 3558
rect 9349 3552 9381 3553
rect 8354 3525 8766 3533
rect 8354 3499 8360 3525
rect 8386 3499 8766 3525
rect 8354 3497 8766 3499
rect 8356 3496 8396 3497
rect 8734 3432 8766 3497
rect 8734 3412 8738 3432
rect 8759 3412 8766 3432
rect 8734 3405 8766 3412
rect 8285 3339 8325 3349
rect 8285 3319 8295 3339
rect 8315 3319 8325 3339
rect 9220 3325 9629 3326
rect 8285 3095 8325 3319
rect 9214 3296 9629 3325
rect 9214 3145 9254 3296
rect 9588 3263 9629 3296
rect 9376 3258 9411 3259
rect 8691 3117 9254 3145
rect 9355 3251 9411 3258
rect 9355 3231 9384 3251
rect 9404 3231 9411 3251
rect 9355 3226 9411 3231
rect 9584 3255 9634 3263
rect 9584 3234 9600 3255
rect 9622 3234 9634 3255
rect 8285 3061 8612 3095
rect 8692 3089 8726 3117
rect 8691 3086 8727 3089
rect 8691 3067 8699 3086
rect 8719 3067 8727 3086
rect 8691 3063 8727 3067
rect 8302 3060 8612 3061
rect 8577 3031 8612 3060
rect 8363 3024 8398 3025
rect 8342 3017 8398 3024
rect 8342 2997 8371 3017
rect 8391 2997 8398 3017
rect 8342 2992 8398 2997
rect 8572 3019 8614 3031
rect 8572 2999 8581 3019
rect 8605 2999 8614 3019
rect 8342 2786 8376 2992
rect 8572 2991 8614 2999
rect 8789 3020 8821 3027
rect 8789 3000 8795 3020
rect 8816 3000 8821 3020
rect 8789 2972 8821 3000
rect 9355 3020 9389 3226
rect 9584 3225 9634 3234
rect 9802 3254 9834 3261
rect 9802 3234 9808 3254
rect 9829 3234 9834 3254
rect 9802 3206 9834 3234
rect 9422 3198 9834 3206
rect 9422 3172 9428 3198
rect 9454 3172 9834 3198
rect 9422 3170 9834 3172
rect 9424 3169 9464 3170
rect 9802 3105 9834 3170
rect 9802 3085 9806 3105
rect 9827 3085 9834 3105
rect 9802 3078 9834 3085
rect 9355 3012 9390 3020
rect 9355 2992 9363 3012
rect 9383 2992 9390 3012
rect 9355 2987 9390 2992
rect 9355 2986 9387 2987
rect 8409 2964 8821 2972
rect 8409 2938 8415 2964
rect 8441 2938 8821 2964
rect 8409 2936 8821 2938
rect 8411 2935 8451 2936
rect 8789 2871 8821 2936
rect 8789 2851 8793 2871
rect 8814 2851 8821 2871
rect 8789 2844 8821 2851
rect 9266 2882 9618 2913
rect 8342 2778 8377 2786
rect 8342 2758 8350 2778
rect 8370 2758 8377 2778
rect 8342 2742 8377 2758
rect 9266 2742 9297 2882
rect 9590 2850 9618 2882
rect 9375 2843 9410 2844
rect 8340 2723 9297 2742
rect 9354 2836 9410 2843
rect 9354 2816 9383 2836
rect 9403 2816 9410 2836
rect 9354 2811 9410 2816
rect 9584 2838 9624 2850
rect 9584 2817 9590 2838
rect 9612 2817 9624 2838
rect 9584 2812 9624 2817
rect 9801 2839 9833 2846
rect 9801 2819 9807 2839
rect 9828 2819 9833 2839
rect 8034 2591 8404 2624
rect 8038 2589 8070 2591
rect 8155 2557 8190 2558
rect 8134 2550 8190 2557
rect 8367 2556 8404 2591
rect 9354 2605 9388 2811
rect 9801 2791 9833 2819
rect 9421 2783 9833 2791
rect 9421 2757 9427 2783
rect 9453 2757 9833 2783
rect 9421 2755 9833 2757
rect 9423 2754 9463 2755
rect 9801 2690 9833 2755
rect 9801 2670 9805 2690
rect 9826 2670 9833 2690
rect 9801 2663 9833 2670
rect 9354 2597 9389 2605
rect 9354 2577 9362 2597
rect 9382 2577 9389 2597
rect 9354 2572 9389 2577
rect 9354 2571 9386 2572
rect 8134 2530 8163 2550
rect 8183 2530 8190 2550
rect 8134 2525 8190 2530
rect 8362 2554 8409 2556
rect 8362 2528 8374 2554
rect 8399 2528 8409 2554
rect 7638 2477 7676 2483
rect 7638 2457 7648 2477
rect 7668 2457 7676 2477
rect 7638 2455 7676 2457
rect 6174 2422 6589 2451
rect 7641 2449 7676 2455
rect 6174 2421 6583 2422
rect 3300 2398 3332 2405
rect 7197 2384 7229 2391
rect 3946 2367 4355 2368
rect 2853 2334 2888 2340
rect 3940 2338 4355 2367
rect 2853 2332 2891 2334
rect 2853 2312 2861 2332
rect 2881 2312 2891 2332
rect 2853 2306 2891 2312
rect 1916 2236 1921 2256
rect 1942 2236 1948 2256
rect 1916 2229 1948 2236
rect 2125 2257 2164 2263
rect 2125 2238 2136 2257
rect 2159 2238 2164 2257
rect 2125 2225 2164 2238
rect 2339 2259 2395 2264
rect 2339 2239 2346 2259
rect 2366 2239 2395 2259
rect 2339 2232 2395 2239
rect 2339 2231 2374 2232
rect 1143 2217 1175 2218
rect 1140 2212 1175 2217
rect 1140 2192 1147 2212
rect 1167 2192 1175 2212
rect 1140 2184 1175 2192
rect 696 2119 728 2126
rect 696 2099 703 2119
rect 724 2099 728 2119
rect 696 2034 728 2099
rect 1066 2034 1106 2035
rect 696 2032 1108 2034
rect 696 2006 1076 2032
rect 1102 2006 1108 2032
rect 696 1998 1108 2006
rect 696 1970 728 1998
rect 1141 1978 1175 2184
rect 2132 2194 2162 2225
rect 2442 2194 2479 2200
rect 2132 2189 2479 2194
rect 2132 2170 2448 2189
rect 2471 2170 2479 2189
rect 2132 2164 2479 2170
rect 2442 2159 2479 2164
rect 696 1950 701 1970
rect 722 1950 728 1970
rect 696 1943 728 1950
rect 905 1972 945 1977
rect 905 1951 917 1972
rect 939 1951 945 1972
rect 905 1939 945 1951
rect 1119 1973 1175 1978
rect 1119 1953 1126 1973
rect 1146 1953 1175 1973
rect 1119 1946 1175 1953
rect 1232 2047 2189 2066
rect 1119 1945 1154 1946
rect 911 1907 939 1939
rect 1232 1907 1263 2047
rect 2152 2031 2187 2047
rect 2152 2011 2159 2031
rect 2179 2011 2187 2031
rect 2152 2003 2187 2011
rect 911 1876 1263 1907
rect 1708 1938 1740 1945
rect 1708 1918 1715 1938
rect 1736 1918 1740 1938
rect 1708 1853 1740 1918
rect 2078 1853 2118 1854
rect 1708 1851 2120 1853
rect 1708 1825 2088 1851
rect 2114 1825 2120 1851
rect 1708 1817 2120 1825
rect 1142 1802 1174 1803
rect 1139 1797 1174 1802
rect 1139 1777 1146 1797
rect 1166 1777 1174 1797
rect 1139 1769 1174 1777
rect 695 1704 727 1711
rect 695 1684 702 1704
rect 723 1684 727 1704
rect 695 1619 727 1684
rect 1065 1619 1105 1620
rect 695 1617 1107 1619
rect 695 1591 1075 1617
rect 1101 1591 1107 1617
rect 695 1583 1107 1591
rect 695 1555 727 1583
rect 695 1535 700 1555
rect 721 1535 727 1555
rect 695 1528 727 1535
rect 895 1555 945 1564
rect 1140 1563 1174 1769
rect 1708 1789 1740 1817
rect 1708 1769 1713 1789
rect 1734 1769 1740 1789
rect 1708 1762 1740 1769
rect 1915 1790 1957 1798
rect 2153 1797 2187 2003
rect 1915 1770 1924 1790
rect 1948 1770 1957 1790
rect 1915 1758 1957 1770
rect 2131 1792 2187 1797
rect 2131 1772 2138 1792
rect 2158 1772 2187 1792
rect 2131 1765 2187 1772
rect 2131 1764 2166 1765
rect 1917 1729 1952 1758
rect 1917 1728 2227 1729
rect 1802 1722 1838 1726
rect 1802 1703 1810 1722
rect 1830 1703 1838 1722
rect 1802 1700 1838 1703
rect 1803 1672 1837 1700
rect 1917 1694 2244 1728
rect 895 1534 907 1555
rect 929 1534 945 1555
rect 895 1526 945 1534
rect 1118 1558 1174 1563
rect 1118 1538 1125 1558
rect 1145 1538 1174 1558
rect 1118 1531 1174 1538
rect 1275 1644 1838 1672
rect 1118 1530 1153 1531
rect 900 1493 941 1526
rect 1275 1493 1315 1644
rect 900 1464 1315 1493
rect 2204 1470 2244 1694
rect 2856 1712 2891 2306
rect 3940 2187 3980 2338
rect 4314 2305 4355 2338
rect 7197 2364 7204 2384
rect 7225 2364 7229 2384
rect 4102 2300 4137 2301
rect 3417 2159 3980 2187
rect 4081 2293 4137 2300
rect 4081 2273 4110 2293
rect 4130 2273 4137 2293
rect 4081 2268 4137 2273
rect 4310 2297 4360 2305
rect 4310 2276 4326 2297
rect 4348 2276 4360 2297
rect 2996 2132 3343 2136
rect 2996 2106 3005 2132
rect 3024 2106 3343 2132
rect 3418 2131 3452 2159
rect 2996 2101 3343 2106
rect 3417 2128 3453 2131
rect 3417 2109 3425 2128
rect 3445 2109 3453 2128
rect 3417 2105 3453 2109
rect 3303 2071 3343 2101
rect 3089 2066 3124 2067
rect 3068 2059 3124 2066
rect 3068 2039 3097 2059
rect 3117 2039 3124 2059
rect 3068 2034 3124 2039
rect 3300 2060 3343 2071
rect 3300 2040 3308 2060
rect 3332 2054 3343 2060
rect 3515 2062 3547 2069
rect 3332 2040 3342 2054
rect 3068 1828 3102 2034
rect 3300 2031 3342 2040
rect 3515 2042 3521 2062
rect 3542 2042 3547 2062
rect 3515 2014 3547 2042
rect 4081 2062 4115 2268
rect 4310 2267 4360 2276
rect 4528 2296 4560 2303
rect 4528 2276 4534 2296
rect 4555 2276 4560 2296
rect 4528 2248 4560 2276
rect 4148 2240 4560 2248
rect 4148 2214 4154 2240
rect 4180 2214 4560 2240
rect 4148 2212 4560 2214
rect 4150 2211 4190 2212
rect 4528 2147 4560 2212
rect 7197 2299 7229 2364
rect 7567 2299 7607 2300
rect 7197 2297 7609 2299
rect 7197 2271 7577 2297
rect 7603 2271 7609 2297
rect 7197 2263 7609 2271
rect 7197 2235 7229 2263
rect 7642 2243 7676 2449
rect 8134 2319 8168 2525
rect 8362 2522 8409 2528
rect 8581 2553 8613 2560
rect 8581 2533 8587 2553
rect 8608 2533 8613 2553
rect 8581 2505 8613 2533
rect 8201 2497 8613 2505
rect 8201 2471 8207 2497
rect 8233 2471 8613 2497
rect 8201 2469 8613 2471
rect 8203 2468 8243 2469
rect 8581 2404 8613 2469
rect 8581 2384 8585 2404
rect 8606 2384 8613 2404
rect 8581 2377 8613 2384
rect 9227 2346 9636 2347
rect 8134 2313 8169 2319
rect 9221 2317 9636 2346
rect 8134 2311 8172 2313
rect 8134 2291 8142 2311
rect 8162 2291 8172 2311
rect 8134 2285 8172 2291
rect 7197 2215 7202 2235
rect 7223 2215 7229 2235
rect 7197 2208 7229 2215
rect 7406 2236 7445 2242
rect 7406 2217 7417 2236
rect 7440 2217 7445 2236
rect 7406 2204 7445 2217
rect 7620 2238 7676 2243
rect 7620 2218 7627 2238
rect 7647 2218 7676 2238
rect 7620 2211 7676 2218
rect 7620 2210 7655 2211
rect 6424 2196 6456 2197
rect 6421 2191 6456 2196
rect 6421 2171 6428 2191
rect 6448 2171 6456 2191
rect 6421 2163 6456 2171
rect 4528 2127 4532 2147
rect 4553 2127 4560 2147
rect 4528 2120 4560 2127
rect 5977 2098 6009 2105
rect 5977 2078 5984 2098
rect 6005 2078 6009 2098
rect 4081 2054 4116 2062
rect 4081 2034 4089 2054
rect 4109 2034 4116 2054
rect 4081 2029 4116 2034
rect 4081 2028 4113 2029
rect 3135 2006 3547 2014
rect 3135 1980 3141 2006
rect 3167 1980 3547 2006
rect 3135 1978 3547 1980
rect 3137 1977 3177 1978
rect 3515 1913 3547 1978
rect 5977 2013 6009 2078
rect 6347 2013 6387 2014
rect 5977 2011 6389 2013
rect 5977 1985 6357 2011
rect 6383 1985 6389 2011
rect 5977 1977 6389 1985
rect 3515 1893 3519 1913
rect 3540 1893 3547 1913
rect 3515 1886 3547 1893
rect 3992 1924 4344 1955
rect 3068 1820 3103 1828
rect 3068 1800 3076 1820
rect 3096 1800 3103 1820
rect 3068 1784 3103 1800
rect 3992 1784 4023 1924
rect 4316 1892 4344 1924
rect 5977 1949 6009 1977
rect 6422 1957 6456 2163
rect 7413 2173 7443 2204
rect 7723 2173 7760 2179
rect 7413 2168 7760 2173
rect 7413 2149 7729 2168
rect 7752 2149 7760 2168
rect 7413 2143 7760 2149
rect 7723 2138 7760 2143
rect 5977 1929 5982 1949
rect 6003 1929 6009 1949
rect 5977 1922 6009 1929
rect 6186 1951 6226 1956
rect 6186 1930 6198 1951
rect 6220 1930 6226 1951
rect 6186 1918 6226 1930
rect 6400 1952 6456 1957
rect 6400 1932 6407 1952
rect 6427 1932 6456 1952
rect 6400 1925 6456 1932
rect 6513 2026 7470 2045
rect 6400 1924 6435 1925
rect 4101 1885 4136 1886
rect 3066 1765 4023 1784
rect 4080 1878 4136 1885
rect 4080 1858 4109 1878
rect 4129 1858 4136 1878
rect 4080 1853 4136 1858
rect 4310 1880 4350 1892
rect 4310 1859 4316 1880
rect 4338 1859 4350 1880
rect 4310 1854 4350 1859
rect 4527 1881 4559 1888
rect 4527 1861 4533 1881
rect 4554 1861 4559 1881
rect 2856 1683 3286 1712
rect 2856 1678 2940 1683
rect 3039 1646 3074 1647
rect 900 1463 1309 1464
rect 2204 1450 2214 1470
rect 2234 1450 2244 1470
rect 2204 1440 2244 1450
rect 3018 1639 3074 1646
rect 3018 1619 3047 1639
rect 3067 1619 3074 1639
rect 3018 1614 3074 1619
rect 3248 1640 3286 1683
rect 3248 1623 3253 1640
rect 3277 1623 3286 1640
rect 1763 1377 1795 1384
rect 1763 1357 1770 1377
rect 1791 1357 1795 1377
rect 1763 1292 1795 1357
rect 2133 1292 2173 1293
rect 1763 1290 2175 1292
rect 1763 1264 2143 1290
rect 2169 1264 2175 1290
rect 1763 1256 2175 1264
rect 1148 1236 1180 1237
rect 1145 1231 1180 1236
rect 1145 1211 1152 1231
rect 1172 1211 1180 1231
rect 1145 1203 1180 1211
rect 701 1138 733 1145
rect 701 1118 708 1138
rect 729 1118 733 1138
rect 701 1053 733 1118
rect 1071 1053 1111 1054
rect 701 1051 1113 1053
rect 701 1025 1081 1051
rect 1107 1025 1113 1051
rect 701 1017 1113 1025
rect 701 989 733 1017
rect 1146 997 1180 1203
rect 1763 1228 1795 1256
rect 2208 1236 2242 1440
rect 3018 1410 3052 1614
rect 3248 1611 3286 1623
rect 3465 1642 3497 1649
rect 3465 1622 3471 1642
rect 3492 1622 3497 1642
rect 3465 1594 3497 1622
rect 4080 1647 4114 1853
rect 4527 1833 4559 1861
rect 6192 1886 6220 1918
rect 6513 1886 6544 2026
rect 7433 2010 7468 2026
rect 7433 1990 7440 2010
rect 7460 1990 7468 2010
rect 7433 1982 7468 1990
rect 6192 1855 6544 1886
rect 6989 1917 7021 1924
rect 6989 1897 6996 1917
rect 7017 1897 7021 1917
rect 4147 1825 4559 1833
rect 4147 1799 4153 1825
rect 4179 1799 4559 1825
rect 4147 1797 4559 1799
rect 4149 1796 4189 1797
rect 4527 1732 4559 1797
rect 6989 1832 7021 1897
rect 7359 1832 7399 1833
rect 6989 1830 7401 1832
rect 6989 1804 7369 1830
rect 7395 1804 7401 1830
rect 6989 1796 7401 1804
rect 6423 1781 6455 1782
rect 6420 1776 6455 1781
rect 6420 1756 6427 1776
rect 6447 1756 6455 1776
rect 6420 1748 6455 1756
rect 4527 1712 4531 1732
rect 4552 1712 4559 1732
rect 4527 1705 4559 1712
rect 5976 1683 6008 1690
rect 5976 1663 5983 1683
rect 6004 1663 6008 1683
rect 4080 1639 4115 1647
rect 4080 1619 4088 1639
rect 4108 1619 4115 1639
rect 4080 1614 4115 1619
rect 4080 1613 4112 1614
rect 3085 1586 3497 1594
rect 3085 1560 3091 1586
rect 3117 1560 3497 1586
rect 3085 1558 3497 1560
rect 3087 1557 3127 1558
rect 3465 1493 3497 1558
rect 5976 1598 6008 1663
rect 6346 1598 6386 1599
rect 5976 1596 6388 1598
rect 5976 1570 6356 1596
rect 6382 1570 6388 1596
rect 5976 1562 6388 1570
rect 5976 1534 6008 1562
rect 5976 1514 5981 1534
rect 6002 1514 6008 1534
rect 5976 1507 6008 1514
rect 6176 1534 6226 1543
rect 6421 1542 6455 1748
rect 6989 1768 7021 1796
rect 6989 1748 6994 1768
rect 7015 1748 7021 1768
rect 6989 1741 7021 1748
rect 7196 1769 7238 1777
rect 7434 1776 7468 1982
rect 7196 1749 7205 1769
rect 7229 1749 7238 1769
rect 7196 1737 7238 1749
rect 7412 1771 7468 1776
rect 7412 1751 7419 1771
rect 7439 1751 7468 1771
rect 7412 1744 7468 1751
rect 7412 1743 7447 1744
rect 7198 1708 7233 1737
rect 7198 1707 7508 1708
rect 7083 1701 7119 1705
rect 7083 1682 7091 1701
rect 7111 1682 7119 1701
rect 7083 1679 7119 1682
rect 7084 1651 7118 1679
rect 7198 1673 7525 1707
rect 6176 1513 6188 1534
rect 6210 1513 6226 1534
rect 6176 1505 6226 1513
rect 6399 1537 6455 1542
rect 6399 1517 6406 1537
rect 6426 1517 6455 1537
rect 6399 1510 6455 1517
rect 6556 1623 7119 1651
rect 6399 1509 6434 1510
rect 3465 1473 3469 1493
rect 3490 1473 3497 1493
rect 3465 1466 3497 1473
rect 6181 1472 6222 1505
rect 6556 1472 6596 1623
rect 6181 1443 6596 1472
rect 7485 1449 7525 1673
rect 8137 1691 8172 2285
rect 9221 2166 9261 2317
rect 9595 2284 9636 2317
rect 9383 2279 9418 2280
rect 8698 2138 9261 2166
rect 9362 2272 9418 2279
rect 9362 2252 9391 2272
rect 9411 2252 9418 2272
rect 9362 2247 9418 2252
rect 9591 2276 9641 2284
rect 9591 2255 9607 2276
rect 9629 2255 9641 2276
rect 8277 2111 8624 2115
rect 8277 2085 8286 2111
rect 8305 2085 8624 2111
rect 8699 2110 8733 2138
rect 8277 2080 8624 2085
rect 8698 2107 8734 2110
rect 8698 2088 8706 2107
rect 8726 2088 8734 2107
rect 8698 2084 8734 2088
rect 8584 2050 8624 2080
rect 8370 2045 8405 2046
rect 8349 2038 8405 2045
rect 8349 2018 8378 2038
rect 8398 2018 8405 2038
rect 8349 2013 8405 2018
rect 8581 2039 8624 2050
rect 8581 2019 8589 2039
rect 8613 2033 8624 2039
rect 8796 2041 8828 2048
rect 8613 2019 8623 2033
rect 8349 1807 8383 2013
rect 8581 2010 8623 2019
rect 8796 2021 8802 2041
rect 8823 2021 8828 2041
rect 8796 1993 8828 2021
rect 9362 2041 9396 2247
rect 9591 2246 9641 2255
rect 9809 2275 9841 2282
rect 9809 2255 9815 2275
rect 9836 2255 9841 2275
rect 9809 2227 9841 2255
rect 9429 2219 9841 2227
rect 9429 2193 9435 2219
rect 9461 2193 9841 2219
rect 9429 2191 9841 2193
rect 9431 2190 9471 2191
rect 9809 2126 9841 2191
rect 9809 2106 9813 2126
rect 9834 2106 9841 2126
rect 9809 2099 9841 2106
rect 9362 2033 9397 2041
rect 9362 2013 9370 2033
rect 9390 2013 9397 2033
rect 9362 2008 9397 2013
rect 9362 2007 9394 2008
rect 8416 1985 8828 1993
rect 8416 1959 8422 1985
rect 8448 1959 8828 1985
rect 8416 1957 8828 1959
rect 8418 1956 8458 1957
rect 8796 1892 8828 1957
rect 8796 1872 8800 1892
rect 8821 1872 8828 1892
rect 8796 1865 8828 1872
rect 9273 1903 9625 1934
rect 8349 1799 8384 1807
rect 8349 1779 8357 1799
rect 8377 1779 8384 1799
rect 8349 1763 8384 1779
rect 9273 1763 9304 1903
rect 9597 1871 9625 1903
rect 9382 1864 9417 1865
rect 8347 1744 9304 1763
rect 9361 1857 9417 1864
rect 9361 1837 9390 1857
rect 9410 1837 9417 1857
rect 9361 1832 9417 1837
rect 9591 1859 9631 1871
rect 9591 1838 9597 1859
rect 9619 1838 9631 1859
rect 9591 1833 9631 1838
rect 9808 1860 9840 1867
rect 9808 1840 9814 1860
rect 9835 1840 9840 1860
rect 8137 1662 8567 1691
rect 8137 1657 8221 1662
rect 8320 1625 8355 1626
rect 6181 1442 6590 1443
rect 7485 1429 7495 1449
rect 7515 1429 7525 1449
rect 7485 1419 7525 1429
rect 8299 1618 8355 1625
rect 8299 1598 8328 1618
rect 8348 1598 8355 1618
rect 8299 1593 8355 1598
rect 8529 1619 8567 1662
rect 8529 1602 8534 1619
rect 8558 1602 8567 1619
rect 1763 1208 1768 1228
rect 1789 1208 1795 1228
rect 1763 1201 1795 1208
rect 1974 1228 2011 1234
rect 1974 1209 1980 1228
rect 2003 1209 2011 1228
rect 1974 1204 2011 1209
rect 2186 1231 2242 1236
rect 2186 1211 2193 1231
rect 2213 1211 2242 1231
rect 2186 1204 2242 1211
rect 3016 1400 3056 1410
rect 3016 1380 3026 1400
rect 3046 1380 3056 1400
rect 3951 1386 4360 1387
rect 1982 1167 2006 1204
rect 2186 1203 2221 1204
rect 1982 1165 2350 1167
rect 1982 1160 2355 1165
rect 1982 1142 2328 1160
rect 2348 1142 2355 1160
rect 1982 1137 2355 1142
rect 2326 1135 2355 1137
rect 3016 1156 3056 1380
rect 3945 1357 4360 1386
rect 3945 1206 3985 1357
rect 4319 1324 4360 1357
rect 7044 1356 7076 1363
rect 7044 1336 7051 1356
rect 7072 1336 7076 1356
rect 4107 1319 4142 1320
rect 3422 1178 3985 1206
rect 4086 1312 4142 1319
rect 4086 1292 4115 1312
rect 4135 1292 4142 1312
rect 4086 1287 4142 1292
rect 4315 1316 4365 1324
rect 4315 1295 4331 1316
rect 4353 1295 4365 1316
rect 3016 1122 3343 1156
rect 3423 1150 3457 1178
rect 3422 1147 3458 1150
rect 3422 1128 3430 1147
rect 3450 1128 3458 1147
rect 3422 1124 3458 1128
rect 3033 1121 3343 1122
rect 3308 1092 3343 1121
rect 3094 1085 3129 1086
rect 701 969 706 989
rect 727 969 733 989
rect 701 962 733 969
rect 910 991 950 996
rect 910 970 922 991
rect 944 970 950 991
rect 910 958 950 970
rect 1124 992 1180 997
rect 1124 972 1131 992
rect 1151 972 1180 992
rect 1124 965 1180 972
rect 1237 1066 2194 1085
rect 3073 1078 3129 1085
rect 1124 964 1159 965
rect 916 926 944 958
rect 1237 926 1268 1066
rect 2157 1050 2192 1066
rect 2157 1030 2164 1050
rect 2184 1030 2192 1050
rect 2157 1022 2192 1030
rect 916 895 1268 926
rect 1713 957 1745 964
rect 1713 937 1720 957
rect 1741 937 1745 957
rect 1713 872 1745 937
rect 2083 872 2123 873
rect 1713 870 2125 872
rect 1713 844 2093 870
rect 2119 844 2125 870
rect 1713 836 2125 844
rect 1147 821 1179 822
rect 1144 816 1179 821
rect 1144 796 1151 816
rect 1171 796 1179 816
rect 1144 788 1179 796
rect 700 723 732 730
rect 700 703 707 723
rect 728 703 732 723
rect 700 638 732 703
rect 1070 638 1110 639
rect 700 636 1112 638
rect 700 610 1080 636
rect 1106 610 1112 636
rect 700 602 1112 610
rect 700 574 732 602
rect 700 554 705 574
rect 726 554 732 574
rect 700 547 732 554
rect 900 574 950 583
rect 1145 582 1179 788
rect 1713 808 1745 836
rect 1713 788 1718 808
rect 1739 788 1745 808
rect 1918 810 1960 819
rect 2158 816 2192 1022
rect 1918 796 1928 810
rect 1713 781 1745 788
rect 1917 790 1928 796
rect 1952 790 1960 810
rect 1917 779 1960 790
rect 2136 811 2192 816
rect 2136 791 2143 811
rect 2163 791 2192 811
rect 3073 1058 3102 1078
rect 3122 1058 3129 1078
rect 3073 1053 3129 1058
rect 3303 1080 3345 1092
rect 3303 1060 3312 1080
rect 3336 1060 3345 1080
rect 3073 847 3107 1053
rect 3303 1052 3345 1060
rect 3520 1081 3552 1088
rect 3520 1061 3526 1081
rect 3547 1061 3552 1081
rect 3520 1033 3552 1061
rect 4086 1081 4120 1287
rect 4315 1286 4365 1295
rect 4533 1315 4565 1322
rect 4533 1295 4539 1315
rect 4560 1295 4565 1315
rect 4533 1267 4565 1295
rect 4153 1259 4565 1267
rect 4153 1233 4159 1259
rect 4185 1233 4565 1259
rect 4153 1231 4565 1233
rect 4155 1230 4195 1231
rect 4533 1166 4565 1231
rect 7044 1271 7076 1336
rect 7414 1271 7454 1272
rect 7044 1269 7456 1271
rect 7044 1243 7424 1269
rect 7450 1243 7456 1269
rect 7044 1235 7456 1243
rect 6429 1215 6461 1216
rect 6426 1210 6461 1215
rect 6426 1190 6433 1210
rect 6453 1190 6461 1210
rect 6426 1182 6461 1190
rect 4533 1146 4537 1166
rect 4558 1146 4565 1166
rect 4533 1139 4565 1146
rect 5982 1117 6014 1124
rect 5982 1097 5989 1117
rect 6010 1097 6014 1117
rect 4086 1073 4121 1081
rect 4086 1053 4094 1073
rect 4114 1053 4121 1073
rect 4086 1048 4121 1053
rect 4086 1047 4118 1048
rect 3140 1025 3552 1033
rect 3140 999 3146 1025
rect 3172 999 3552 1025
rect 3140 997 3552 999
rect 3142 996 3182 997
rect 3520 932 3552 997
rect 5982 1032 6014 1097
rect 6352 1032 6392 1033
rect 5982 1030 6394 1032
rect 5982 1004 6362 1030
rect 6388 1004 6394 1030
rect 5982 996 6394 1004
rect 3520 912 3524 932
rect 3545 912 3552 932
rect 3520 905 3552 912
rect 3997 943 4349 974
rect 3073 839 3108 847
rect 3073 819 3081 839
rect 3101 819 3108 839
rect 3073 803 3108 819
rect 3997 803 4028 943
rect 4321 911 4349 943
rect 5982 968 6014 996
rect 6427 976 6461 1182
rect 7044 1207 7076 1235
rect 7489 1215 7523 1419
rect 8299 1389 8333 1593
rect 8529 1590 8567 1602
rect 8746 1621 8778 1628
rect 8746 1601 8752 1621
rect 8773 1601 8778 1621
rect 8746 1573 8778 1601
rect 9361 1626 9395 1832
rect 9808 1812 9840 1840
rect 9428 1804 9840 1812
rect 9428 1778 9434 1804
rect 9460 1778 9840 1804
rect 9428 1776 9840 1778
rect 9430 1775 9470 1776
rect 9808 1711 9840 1776
rect 9808 1691 9812 1711
rect 9833 1691 9840 1711
rect 9808 1684 9840 1691
rect 9361 1618 9396 1626
rect 9361 1598 9369 1618
rect 9389 1598 9396 1618
rect 9361 1593 9396 1598
rect 9361 1592 9393 1593
rect 8366 1565 8778 1573
rect 8366 1539 8372 1565
rect 8398 1539 8778 1565
rect 8366 1537 8778 1539
rect 8368 1536 8408 1537
rect 8746 1472 8778 1537
rect 8746 1452 8750 1472
rect 8771 1452 8778 1472
rect 8746 1445 8778 1452
rect 7044 1187 7049 1207
rect 7070 1187 7076 1207
rect 7044 1180 7076 1187
rect 7255 1207 7292 1213
rect 7255 1188 7261 1207
rect 7284 1188 7292 1207
rect 7255 1183 7292 1188
rect 7467 1210 7523 1215
rect 7467 1190 7474 1210
rect 7494 1190 7523 1210
rect 7467 1183 7523 1190
rect 8297 1379 8337 1389
rect 8297 1359 8307 1379
rect 8327 1359 8337 1379
rect 9232 1365 9641 1366
rect 7263 1146 7287 1183
rect 7467 1182 7502 1183
rect 7263 1144 7631 1146
rect 7263 1139 7636 1144
rect 7263 1121 7609 1139
rect 7629 1121 7636 1139
rect 7263 1116 7636 1121
rect 7607 1114 7636 1116
rect 8297 1135 8337 1359
rect 9226 1336 9641 1365
rect 9226 1185 9266 1336
rect 9600 1303 9641 1336
rect 9388 1298 9423 1299
rect 8703 1157 9266 1185
rect 9367 1291 9423 1298
rect 9367 1271 9396 1291
rect 9416 1271 9423 1291
rect 9367 1266 9423 1271
rect 9596 1295 9646 1303
rect 9596 1274 9612 1295
rect 9634 1274 9646 1295
rect 8297 1101 8624 1135
rect 8704 1129 8738 1157
rect 8703 1126 8739 1129
rect 8703 1107 8711 1126
rect 8731 1107 8739 1126
rect 8703 1103 8739 1107
rect 8314 1100 8624 1101
rect 8589 1071 8624 1100
rect 8375 1064 8410 1065
rect 5982 948 5987 968
rect 6008 948 6014 968
rect 5982 941 6014 948
rect 6191 970 6231 975
rect 6191 949 6203 970
rect 6225 949 6231 970
rect 6191 937 6231 949
rect 6405 971 6461 976
rect 6405 951 6412 971
rect 6432 951 6461 971
rect 6405 944 6461 951
rect 6518 1045 7475 1064
rect 8354 1057 8410 1064
rect 6405 943 6440 944
rect 4106 904 4141 905
rect 2136 784 2192 791
rect 3071 784 4028 803
rect 4085 897 4141 904
rect 4085 877 4114 897
rect 4134 877 4141 897
rect 4085 872 4141 877
rect 4315 899 4355 911
rect 4315 878 4321 899
rect 4343 878 4355 899
rect 4315 873 4355 878
rect 4532 900 4564 907
rect 4532 880 4538 900
rect 4559 880 4564 900
rect 2136 783 2171 784
rect 1917 749 1957 779
rect 1807 741 1843 745
rect 1807 722 1815 741
rect 1835 722 1843 741
rect 1807 719 1843 722
rect 1917 744 2264 749
rect 1808 691 1842 719
rect 1917 718 2236 744
rect 2255 718 2264 744
rect 1917 714 2264 718
rect 900 553 912 574
rect 934 553 950 574
rect 900 545 950 553
rect 1123 577 1179 582
rect 1123 557 1130 577
rect 1150 557 1179 577
rect 1123 550 1179 557
rect 1280 663 1843 691
rect 4085 666 4119 872
rect 4532 852 4564 880
rect 6197 905 6225 937
rect 6518 905 6549 1045
rect 7438 1029 7473 1045
rect 7438 1009 7445 1029
rect 7465 1009 7473 1029
rect 7438 1001 7473 1009
rect 6197 874 6549 905
rect 6994 936 7026 943
rect 6994 916 7001 936
rect 7022 916 7026 936
rect 4152 844 4564 852
rect 4152 818 4158 844
rect 4184 818 4564 844
rect 4152 816 4564 818
rect 4154 815 4194 816
rect 4532 751 4564 816
rect 6994 851 7026 916
rect 7364 851 7404 852
rect 6994 849 7406 851
rect 6994 823 7374 849
rect 7400 823 7406 849
rect 6994 815 7406 823
rect 6428 800 6460 801
rect 6425 795 6460 800
rect 6425 775 6432 795
rect 6452 775 6460 795
rect 6425 767 6460 775
rect 4532 731 4536 751
rect 4557 731 4564 751
rect 4532 724 4564 731
rect 5981 702 6013 709
rect 5981 682 5988 702
rect 6009 682 6013 702
rect 1123 549 1158 550
rect 905 512 946 545
rect 1280 512 1320 663
rect 4085 658 4120 666
rect 4085 638 4093 658
rect 4113 638 4120 658
rect 4085 633 4120 638
rect 4085 632 4117 633
rect 5981 617 6013 682
rect 6351 617 6391 618
rect 5981 615 6393 617
rect 5981 589 6361 615
rect 6387 589 6393 615
rect 5981 581 6393 589
rect 5981 553 6013 581
rect 5981 533 5986 553
rect 6007 533 6013 553
rect 5981 526 6013 533
rect 6181 553 6231 562
rect 6426 561 6460 767
rect 6994 787 7026 815
rect 6994 767 6999 787
rect 7020 767 7026 787
rect 7199 789 7241 798
rect 7439 795 7473 1001
rect 7199 775 7209 789
rect 6994 760 7026 767
rect 7198 769 7209 775
rect 7233 769 7241 789
rect 7198 758 7241 769
rect 7417 790 7473 795
rect 7417 770 7424 790
rect 7444 770 7473 790
rect 8354 1037 8383 1057
rect 8403 1037 8410 1057
rect 8354 1032 8410 1037
rect 8584 1059 8626 1071
rect 8584 1039 8593 1059
rect 8617 1039 8626 1059
rect 8354 826 8388 1032
rect 8584 1031 8626 1039
rect 8801 1060 8833 1067
rect 8801 1040 8807 1060
rect 8828 1040 8833 1060
rect 8801 1012 8833 1040
rect 9367 1060 9401 1266
rect 9596 1265 9646 1274
rect 9814 1294 9846 1301
rect 9814 1274 9820 1294
rect 9841 1274 9846 1294
rect 9814 1246 9846 1274
rect 9434 1238 9846 1246
rect 9434 1212 9440 1238
rect 9466 1212 9846 1238
rect 9434 1210 9846 1212
rect 9436 1209 9476 1210
rect 9814 1145 9846 1210
rect 9814 1125 9818 1145
rect 9839 1125 9846 1145
rect 9814 1118 9846 1125
rect 9367 1052 9402 1060
rect 9367 1032 9375 1052
rect 9395 1032 9402 1052
rect 9367 1027 9402 1032
rect 9367 1026 9399 1027
rect 8421 1004 8833 1012
rect 8421 978 8427 1004
rect 8453 978 8833 1004
rect 8421 976 8833 978
rect 8423 975 8463 976
rect 8801 911 8833 976
rect 8801 891 8805 911
rect 8826 891 8833 911
rect 8801 884 8833 891
rect 9278 922 9630 953
rect 8354 818 8389 826
rect 8354 798 8362 818
rect 8382 798 8389 818
rect 8354 782 8389 798
rect 9278 782 9309 922
rect 9602 890 9630 922
rect 9387 883 9422 884
rect 7417 763 7473 770
rect 8352 763 9309 782
rect 9366 876 9422 883
rect 9366 856 9395 876
rect 9415 856 9422 876
rect 9366 851 9422 856
rect 9596 878 9636 890
rect 9596 857 9602 878
rect 9624 857 9636 878
rect 9596 852 9636 857
rect 9813 879 9845 886
rect 9813 859 9819 879
rect 9840 859 9845 879
rect 7417 762 7452 763
rect 7198 728 7238 758
rect 7088 720 7124 724
rect 7088 701 7096 720
rect 7116 701 7124 720
rect 7088 698 7124 701
rect 7198 723 7545 728
rect 7089 670 7123 698
rect 7198 697 7517 723
rect 7536 697 7545 723
rect 7198 693 7545 697
rect 6181 532 6193 553
rect 6215 532 6231 553
rect 6181 524 6231 532
rect 6404 556 6460 561
rect 6404 536 6411 556
rect 6431 536 6460 556
rect 6404 529 6460 536
rect 6561 642 7124 670
rect 9366 645 9400 851
rect 9813 831 9845 859
rect 9433 823 9845 831
rect 9433 797 9439 823
rect 9465 797 9845 823
rect 9433 795 9845 797
rect 9435 794 9475 795
rect 9813 730 9845 795
rect 9813 710 9817 730
rect 9838 710 9845 730
rect 9813 703 9845 710
rect 6404 528 6439 529
rect 905 483 1320 512
rect 6186 491 6227 524
rect 6561 491 6601 642
rect 9366 637 9401 645
rect 9366 617 9374 637
rect 9394 617 9401 637
rect 9366 612 9401 617
rect 9366 611 9398 612
rect 905 482 1314 483
rect 6186 462 6601 491
rect 6186 461 6595 462
rect 747 454 787 459
rect 694 451 5119 454
rect 694 429 756 451
rect 779 429 5089 451
rect 5112 429 5119 451
rect 6028 433 6068 438
rect 694 424 5119 429
rect 5975 430 10400 433
rect 747 414 787 424
rect 5975 408 6037 430
rect 6060 408 10370 430
rect 10393 408 10400 430
rect 5975 403 10400 408
rect 6028 393 6068 403
rect 2543 382 2592 386
rect 2543 381 2553 382
rect 2543 352 2552 381
rect 2584 352 2592 382
rect 2543 351 2592 352
rect 2542 343 2592 351
rect 2542 335 2591 343
rect 2542 315 2554 335
rect 2574 315 2591 335
rect 2542 308 2591 315
rect 2646 334 2694 337
rect 2547 307 2582 308
rect 2103 242 2135 249
rect 2103 222 2110 242
rect 2131 222 2135 242
rect 2103 157 2135 222
rect 2473 157 2513 158
rect 2103 155 2515 157
rect 2103 129 2483 155
rect 2509 129 2515 155
rect 2103 121 2515 129
rect 2103 93 2135 121
rect 2548 101 2582 307
rect 2646 307 2649 334
rect 2684 307 2694 334
rect 2646 240 2694 307
rect 2646 220 2651 240
rect 2679 220 2694 240
rect 2646 210 2694 220
rect 2775 327 2811 372
rect 7824 361 7873 365
rect 7824 360 7834 361
rect 5636 327 5672 333
rect 7824 331 7833 360
rect 7865 331 7873 361
rect 7824 330 7873 331
rect 2775 299 5672 327
rect 2103 73 2108 93
rect 2129 73 2135 93
rect 2103 66 2135 73
rect 2311 93 2355 100
rect 2311 71 2322 93
rect 2347 71 2355 93
rect 2311 63 2355 71
rect 2526 96 2582 101
rect 2526 76 2533 96
rect 2553 76 2582 96
rect 2526 69 2582 76
rect 2526 68 2561 69
rect 2317 33 2342 63
rect 2775 35 2813 299
rect 5636 247 5672 299
rect 7823 322 7873 330
rect 7823 314 7872 322
rect 7823 294 7835 314
rect 7855 294 7872 314
rect 7823 287 7872 294
rect 7927 313 7975 316
rect 7828 286 7863 287
rect 5636 227 5644 247
rect 5664 227 5672 247
rect 5636 224 5672 227
rect 5637 219 5672 224
rect 5193 154 5225 161
rect 5193 134 5200 154
rect 5221 134 5225 154
rect 5193 69 5225 134
rect 5563 69 5603 70
rect 5193 67 5605 69
rect 5193 41 5573 67
rect 5599 41 5605 67
rect 2725 33 2814 35
rect 2317 0 2814 33
rect 2725 -4 2814 0
rect 5193 33 5605 41
rect 5193 5 5225 33
rect 5638 13 5672 219
rect 7384 221 7416 228
rect 7384 201 7391 221
rect 7412 201 7416 221
rect 7384 136 7416 201
rect 7754 136 7794 137
rect 7384 134 7796 136
rect 7384 108 7764 134
rect 7790 108 7796 134
rect 7384 100 7796 108
rect 7384 72 7416 100
rect 7829 80 7863 286
rect 7927 286 7930 313
rect 7965 286 7975 313
rect 7927 219 7975 286
rect 7927 199 7932 219
rect 7960 199 7975 219
rect 7927 189 7975 199
rect 7384 52 7389 72
rect 7410 52 7416 72
rect 7384 45 7416 52
rect 7592 72 7636 79
rect 7592 50 7603 72
rect 7628 50 7636 72
rect 7592 42 7636 50
rect 7807 75 7863 80
rect 7807 55 7814 75
rect 7834 55 7863 75
rect 7807 48 7863 55
rect 7807 47 7842 48
rect 5193 -15 5198 5
rect 5219 -15 5225 5
rect 5193 -22 5225 -15
rect 5399 2 5444 11
rect 5399 -15 5409 2
rect 5430 -15 5444 2
rect 5399 -86 5444 -15
rect 5616 8 5672 13
rect 5616 -12 5623 8
rect 5643 -12 5672 8
rect 5616 -19 5672 -12
rect 7598 13 7623 42
rect 7598 -18 7622 13
rect 6914 -19 7622 -18
rect 5616 -20 5651 -19
rect 5796 -20 7622 -19
rect 5787 -21 7622 -20
rect 5787 -40 7621 -21
rect 5787 -51 6959 -40
rect 5787 -57 5834 -51
rect 5650 -65 5834 -57
rect 5650 -82 5659 -65
rect 5683 -82 5834 -65
rect 5650 -90 5834 -82
rect 5650 -91 5833 -90
<< via1 >>
rect 2649 4609 2686 4639
rect 7930 4588 7967 4618
rect 2548 4088 2582 4116
rect 7829 4067 7863 4095
rect 2553 381 2584 382
rect 2552 352 2584 381
rect 2649 307 2684 334
rect 7834 360 7865 361
rect 7833 331 7865 360
rect 7930 286 7965 313
<< metal2 >>
rect 2644 4639 2693 4645
rect 2644 4609 2649 4639
rect 2686 4609 2693 4639
rect 2542 4116 2587 4122
rect 2542 4088 2548 4116
rect 2582 4088 2587 4116
rect 2542 478 2587 4088
rect 2644 509 2693 4609
rect 7925 4618 7974 4624
rect 7925 4588 7930 4618
rect 7967 4588 7974 4618
rect 7823 4095 7868 4101
rect 7823 4067 7829 4095
rect 7863 4067 7868 4095
rect 2548 386 2586 478
rect 2543 382 2592 386
rect 2543 381 2553 382
rect 2543 352 2552 381
rect 2584 352 2592 382
rect 2543 343 2592 352
rect 2646 334 2692 509
rect 7823 457 7868 4067
rect 7925 488 7974 4588
rect 7829 365 7867 457
rect 2646 307 2649 334
rect 2684 307 2692 334
rect 7824 361 7873 365
rect 7824 360 7834 361
rect 7824 331 7833 360
rect 7865 331 7873 361
rect 7824 322 7873 331
rect 2646 292 2692 307
rect 7927 313 7973 488
rect 7927 286 7930 313
rect 7965 286 7973 313
rect 7927 271 7973 286
<< labels >>
rlabel locali 304 8073 333 8079 1 vdd
rlabel locali 517 8070 546 8076 1 vdd
rlabel locali 250 7885 272 7900 1 d0
rlabel nwell 671 8040 694 8043 1 vdd
rlabel locali 301 7774 330 7780 1 gnd
rlabel locali 514 7774 543 7780 1 gnd
rlabel space 611 7769 640 7778 1 gnd
rlabel locali 303 7658 332 7664 1 vdd
rlabel locali 516 7655 545 7661 1 vdd
rlabel locali 249 7470 271 7485 1 d0
rlabel nwell 670 7625 693 7628 1 vdd
rlabel locali 300 7359 329 7365 1 gnd
rlabel locali 513 7359 542 7365 1 gnd
rlabel space 610 7354 639 7363 1 gnd
rlabel locali 1316 7892 1345 7898 1 vdd
rlabel locali 1529 7889 1558 7895 1 vdd
rlabel nwell 1683 7859 1706 7862 1 vdd
rlabel locali 1313 7593 1342 7599 1 gnd
rlabel locali 1526 7593 1555 7599 1 gnd
rlabel space 1623 7588 1652 7597 1 gnd
rlabel locali 1254 7703 1301 7724 1 d1
rlabel locali 116 8265 141 8274 1 vref
rlabel locali 309 7092 338 7098 1 vdd
rlabel locali 522 7089 551 7095 1 vdd
rlabel locali 255 6904 277 6919 1 d0
rlabel nwell 676 7059 699 7062 1 vdd
rlabel locali 306 6793 335 6799 1 gnd
rlabel locali 519 6793 548 6799 1 gnd
rlabel space 616 6788 645 6797 1 gnd
rlabel locali 308 6677 337 6683 1 vdd
rlabel locali 521 6674 550 6680 1 vdd
rlabel locali 254 6489 276 6504 1 d0
rlabel nwell 675 6644 698 6647 1 vdd
rlabel locali 305 6378 334 6384 1 gnd
rlabel locali 518 6378 547 6384 1 gnd
rlabel locali 1321 6911 1350 6917 1 vdd
rlabel locali 1534 6908 1563 6914 1 vdd
rlabel nwell 1688 6878 1711 6881 1 vdd
rlabel locali 1318 6612 1347 6618 1 gnd
rlabel locali 1531 6612 1560 6618 1 gnd
rlabel space 1628 6607 1657 6616 1 gnd
rlabel locali 1259 6722 1306 6743 1 d1
rlabel locali 1371 7331 1400 7337 1 vdd
rlabel locali 1584 7328 1613 7334 1 vdd
rlabel nwell 1738 7298 1761 7301 1 vdd
rlabel locali 1368 7032 1397 7038 1 gnd
rlabel locali 1581 7032 1610 7038 1 gnd
rlabel space 1678 7027 1707 7036 1 gnd
rlabel locali 1314 7143 1337 7158 1 d2
rlabel space 615 6373 644 6382 1 gnd
rlabel locali 1326 5183 1349 5198 1 d2
rlabel space 1690 5067 1719 5076 1 gnd
rlabel locali 1593 5072 1622 5078 1 gnd
rlabel locali 1380 5072 1409 5078 1 gnd
rlabel nwell 1750 5338 1773 5341 1 vdd
rlabel locali 1596 5368 1625 5374 1 vdd
rlabel locali 1383 5371 1412 5377 1 vdd
rlabel locali 1271 4762 1318 4783 1 d1
rlabel space 1640 4647 1669 4656 1 gnd
rlabel locali 1543 4652 1572 4658 1 gnd
rlabel locali 1330 4652 1359 4658 1 gnd
rlabel nwell 1700 4918 1723 4921 1 vdd
rlabel locali 1546 4948 1575 4954 1 vdd
rlabel locali 1333 4951 1362 4957 1 vdd
rlabel space 627 4413 656 4422 1 gnd
rlabel locali 530 4418 559 4424 1 gnd
rlabel locali 317 4418 346 4424 1 gnd
rlabel nwell 687 4684 710 4687 1 vdd
rlabel locali 266 4529 288 4544 1 d0
rlabel locali 533 4714 562 4720 1 vdd
rlabel locali 320 4717 349 4723 1 vdd
rlabel space 628 4828 657 4837 1 gnd
rlabel locali 531 4833 560 4839 1 gnd
rlabel locali 318 4833 347 4839 1 gnd
rlabel nwell 688 5099 711 5102 1 vdd
rlabel locali 267 4944 289 4959 1 d0
rlabel locali 534 5129 563 5135 1 vdd
rlabel locali 321 5132 350 5138 1 vdd
rlabel locali 1266 5743 1313 5764 1 d1
rlabel space 1635 5628 1664 5637 1 gnd
rlabel locali 1538 5633 1567 5639 1 gnd
rlabel locali 1325 5633 1354 5639 1 gnd
rlabel nwell 1695 5899 1718 5902 1 vdd
rlabel locali 1541 5929 1570 5935 1 vdd
rlabel locali 1328 5932 1357 5938 1 vdd
rlabel space 622 5394 651 5403 1 gnd
rlabel locali 525 5399 554 5405 1 gnd
rlabel locali 312 5399 341 5405 1 gnd
rlabel nwell 682 5665 705 5668 1 vdd
rlabel locali 261 5510 283 5525 1 d0
rlabel locali 528 5695 557 5701 1 vdd
rlabel locali 315 5698 344 5704 1 vdd
rlabel space 623 5809 652 5818 1 gnd
rlabel locali 526 5814 555 5820 1 gnd
rlabel locali 313 5814 342 5820 1 gnd
rlabel nwell 683 6080 706 6083 1 vdd
rlabel locali 262 5925 284 5940 1 d0
rlabel locali 529 6110 558 6116 1 vdd
rlabel locali 316 6113 345 6119 1 vdd
rlabel locali 1536 6399 1565 6405 1 vdd
rlabel locali 1749 6396 1778 6402 1 vdd
rlabel nwell 1903 6366 1926 6369 1 vdd
rlabel locali 1533 6100 1562 6106 1 gnd
rlabel locali 1746 6100 1775 6106 1 gnd
rlabel space 1843 6095 1872 6104 1 gnd
rlabel locali 1474 6209 1506 6228 1 d3
rlabel locali 1494 2292 1526 2311 1 d3
rlabel space 1863 2178 1892 2187 1 gnd
rlabel locali 1766 2183 1795 2189 1 gnd
rlabel locali 1553 2183 1582 2189 1 gnd
rlabel nwell 1923 2449 1946 2452 1 vdd
rlabel locali 1769 2479 1798 2485 1 vdd
rlabel locali 1556 2482 1585 2488 1 vdd
rlabel locali 336 2196 365 2202 1 vdd
rlabel locali 549 2193 578 2199 1 vdd
rlabel locali 282 2008 304 2023 1 d0
rlabel nwell 703 2163 726 2166 1 vdd
rlabel locali 333 1897 362 1903 1 gnd
rlabel locali 546 1897 575 1903 1 gnd
rlabel space 643 1892 672 1901 1 gnd
rlabel locali 335 1781 364 1787 1 vdd
rlabel locali 548 1778 577 1784 1 vdd
rlabel locali 281 1593 303 1608 1 d0
rlabel nwell 702 1748 725 1751 1 vdd
rlabel locali 332 1482 361 1488 1 gnd
rlabel locali 545 1482 574 1488 1 gnd
rlabel space 642 1477 671 1486 1 gnd
rlabel locali 1348 2015 1377 2021 1 vdd
rlabel locali 1561 2012 1590 2018 1 vdd
rlabel nwell 1715 1982 1738 1985 1 vdd
rlabel locali 1345 1716 1374 1722 1 gnd
rlabel locali 1558 1716 1587 1722 1 gnd
rlabel space 1655 1711 1684 1720 1 gnd
rlabel locali 1286 1826 1333 1847 1 d1
rlabel locali 341 1215 370 1221 1 vdd
rlabel locali 554 1212 583 1218 1 vdd
rlabel locali 287 1027 309 1042 1 d0
rlabel nwell 708 1182 731 1185 1 vdd
rlabel locali 338 916 367 922 1 gnd
rlabel locali 551 916 580 922 1 gnd
rlabel space 648 911 677 920 1 gnd
rlabel locali 340 800 369 806 1 vdd
rlabel locali 553 797 582 803 1 vdd
rlabel locali 286 612 308 627 1 d0
rlabel nwell 707 767 730 770 1 vdd
rlabel locali 337 501 366 507 1 gnd
rlabel locali 550 501 579 507 1 gnd
rlabel space 647 496 676 505 1 gnd
rlabel locali 1353 1034 1382 1040 1 vdd
rlabel locali 1566 1031 1595 1037 1 vdd
rlabel nwell 1720 1001 1743 1004 1 vdd
rlabel locali 1350 735 1379 741 1 gnd
rlabel locali 1563 735 1592 741 1 gnd
rlabel space 1660 730 1689 739 1 gnd
rlabel locali 1291 845 1338 866 1 d1
rlabel locali 1403 1454 1432 1460 1 vdd
rlabel locali 1616 1451 1645 1457 1 vdd
rlabel nwell 1770 1421 1793 1424 1 vdd
rlabel locali 1400 1155 1429 1161 1 gnd
rlabel locali 1613 1155 1642 1161 1 gnd
rlabel space 1710 1150 1739 1159 1 gnd
rlabel locali 1346 1266 1369 1281 1 d2
rlabel space 635 2456 664 2465 1 gnd
rlabel locali 1334 3226 1357 3241 1 d2
rlabel space 1698 3110 1727 3119 1 gnd
rlabel locali 1601 3115 1630 3121 1 gnd
rlabel locali 1388 3115 1417 3121 1 gnd
rlabel nwell 1758 3381 1781 3384 1 vdd
rlabel locali 1604 3411 1633 3417 1 vdd
rlabel locali 1391 3414 1420 3420 1 vdd
rlabel locali 1279 2805 1326 2826 1 d1
rlabel space 1648 2690 1677 2699 1 gnd
rlabel locali 1551 2695 1580 2701 1 gnd
rlabel locali 1338 2695 1367 2701 1 gnd
rlabel nwell 1708 2961 1731 2964 1 vdd
rlabel locali 1554 2991 1583 2997 1 vdd
rlabel locali 1341 2994 1370 3000 1 vdd
rlabel locali 538 2461 567 2467 1 gnd
rlabel locali 325 2461 354 2467 1 gnd
rlabel nwell 695 2727 718 2730 1 vdd
rlabel locali 274 2572 296 2587 1 d0
rlabel locali 541 2757 570 2763 1 vdd
rlabel locali 328 2760 357 2766 1 vdd
rlabel space 636 2871 665 2880 1 gnd
rlabel locali 539 2876 568 2882 1 gnd
rlabel locali 326 2876 355 2882 1 gnd
rlabel nwell 696 3142 719 3145 1 vdd
rlabel locali 275 2987 297 3002 1 d0
rlabel locali 542 3172 571 3178 1 vdd
rlabel locali 329 3175 358 3181 1 vdd
rlabel locali 1274 3786 1321 3807 1 d1
rlabel space 1643 3671 1672 3680 1 gnd
rlabel locali 1546 3676 1575 3682 1 gnd
rlabel locali 1333 3676 1362 3682 1 gnd
rlabel nwell 1703 3942 1726 3945 1 vdd
rlabel locali 1549 3972 1578 3978 1 vdd
rlabel locali 1336 3975 1365 3981 1 vdd
rlabel space 630 3437 659 3446 1 gnd
rlabel locali 533 3442 562 3448 1 gnd
rlabel locali 320 3442 349 3448 1 gnd
rlabel nwell 690 3708 713 3711 1 vdd
rlabel locali 269 3553 291 3568 1 d0
rlabel locali 536 3738 565 3744 1 vdd
rlabel locali 323 3741 352 3747 1 vdd
rlabel space 631 3852 660 3861 1 gnd
rlabel locali 534 3857 563 3863 1 gnd
rlabel locali 321 3857 350 3863 1 gnd
rlabel nwell 691 4123 714 4126 1 vdd
rlabel locali 270 3968 292 3983 1 d0
rlabel locali 537 4153 566 4159 1 vdd
rlabel locali 324 4156 353 4162 1 vdd
rlabel locali 1631 4407 1660 4413 1 vdd
rlabel locali 1844 4404 1873 4410 1 vdd
rlabel nwell 1998 4374 2021 4377 1 vdd
rlabel locali 1628 4108 1657 4114 1 gnd
rlabel locali 1841 4108 1870 4114 1 gnd
rlabel space 1938 4103 1967 4112 1 gnd
rlabel locali 1573 4213 1595 4237 1 d4
rlabel locali 4895 648 4924 654 5 vdd
rlabel locali 4682 651 4711 657 5 vdd
rlabel locali 4956 827 4978 842 5 d0
rlabel nwell 4534 684 4557 687 5 vdd
rlabel locali 4898 947 4927 953 5 gnd
rlabel locali 4685 947 4714 953 5 gnd
rlabel space 4588 949 4617 958 5 gnd
rlabel locali 4896 1063 4925 1069 5 vdd
rlabel locali 4683 1066 4712 1072 5 vdd
rlabel locali 4957 1242 4979 1257 5 d0
rlabel nwell 4535 1099 4558 1102 5 vdd
rlabel locali 4899 1362 4928 1368 5 gnd
rlabel locali 4686 1362 4715 1368 5 gnd
rlabel space 4589 1364 4618 1373 5 gnd
rlabel locali 3883 829 3912 835 5 vdd
rlabel locali 3670 832 3699 838 5 vdd
rlabel nwell 3522 865 3545 868 5 vdd
rlabel locali 3886 1128 3915 1134 5 gnd
rlabel locali 3673 1128 3702 1134 5 gnd
rlabel space 3576 1130 3605 1139 5 gnd
rlabel locali 3927 1003 3974 1024 5 d1
rlabel locali 4890 1629 4919 1635 5 vdd
rlabel locali 4677 1632 4706 1638 5 vdd
rlabel locali 4951 1808 4973 1823 5 d0
rlabel nwell 4529 1665 4552 1668 5 vdd
rlabel locali 4893 1928 4922 1934 5 gnd
rlabel locali 4680 1928 4709 1934 5 gnd
rlabel space 4583 1930 4612 1939 5 gnd
rlabel locali 4891 2044 4920 2050 5 vdd
rlabel locali 4678 2047 4707 2053 5 vdd
rlabel locali 4952 2223 4974 2238 5 d0
rlabel nwell 4530 2080 4553 2083 5 vdd
rlabel locali 4894 2343 4923 2349 5 gnd
rlabel locali 4681 2343 4710 2349 5 gnd
rlabel locali 3878 1810 3907 1816 5 vdd
rlabel locali 3665 1813 3694 1819 5 vdd
rlabel nwell 3517 1846 3540 1849 5 vdd
rlabel locali 3881 2109 3910 2115 5 gnd
rlabel locali 3668 2109 3697 2115 5 gnd
rlabel space 3571 2111 3600 2120 5 gnd
rlabel locali 3922 1984 3969 2005 5 d1
rlabel locali 3828 1390 3857 1396 5 vdd
rlabel locali 3615 1393 3644 1399 5 vdd
rlabel nwell 3467 1426 3490 1429 5 vdd
rlabel locali 3831 1689 3860 1695 5 gnd
rlabel locali 3618 1689 3647 1695 5 gnd
rlabel space 3521 1691 3550 1700 5 gnd
rlabel locali 3891 1569 3914 1584 5 d2
rlabel space 4584 2345 4613 2354 5 gnd
rlabel locali 3879 3529 3902 3544 5 d2
rlabel space 3509 3651 3538 3660 5 gnd
rlabel locali 3606 3649 3635 3655 5 gnd
rlabel locali 3819 3649 3848 3655 5 gnd
rlabel nwell 3455 3386 3478 3389 5 vdd
rlabel locali 3603 3353 3632 3359 5 vdd
rlabel locali 3816 3350 3845 3356 5 vdd
rlabel locali 3910 3944 3957 3965 5 d1
rlabel space 3559 4071 3588 4080 5 gnd
rlabel locali 3656 4069 3685 4075 5 gnd
rlabel locali 3869 4069 3898 4075 5 gnd
rlabel nwell 3505 3806 3528 3809 5 vdd
rlabel locali 3653 3773 3682 3779 5 vdd
rlabel locali 3866 3770 3895 3776 5 vdd
rlabel space 4572 4305 4601 4314 5 gnd
rlabel locali 4669 4303 4698 4309 5 gnd
rlabel locali 4882 4303 4911 4309 5 gnd
rlabel nwell 4518 4040 4541 4043 5 vdd
rlabel locali 4940 4183 4962 4198 5 d0
rlabel locali 4666 4007 4695 4013 5 vdd
rlabel locali 4879 4004 4908 4010 5 vdd
rlabel space 4571 3890 4600 3899 5 gnd
rlabel locali 4668 3888 4697 3894 5 gnd
rlabel locali 4881 3888 4910 3894 5 gnd
rlabel nwell 4517 3625 4540 3628 5 vdd
rlabel locali 4939 3768 4961 3783 5 d0
rlabel locali 4665 3592 4694 3598 5 vdd
rlabel locali 4878 3589 4907 3595 5 vdd
rlabel locali 3915 2963 3962 2984 5 d1
rlabel space 3564 3090 3593 3099 5 gnd
rlabel locali 3661 3088 3690 3094 5 gnd
rlabel locali 3874 3088 3903 3094 5 gnd
rlabel nwell 3510 2825 3533 2828 5 vdd
rlabel locali 3658 2792 3687 2798 5 vdd
rlabel locali 3871 2789 3900 2795 5 vdd
rlabel space 4577 3324 4606 3333 5 gnd
rlabel locali 4674 3322 4703 3328 5 gnd
rlabel locali 4887 3322 4916 3328 5 gnd
rlabel nwell 4523 3059 4546 3062 5 vdd
rlabel locali 4945 3202 4967 3217 5 d0
rlabel locali 4671 3026 4700 3032 5 vdd
rlabel locali 4884 3023 4913 3029 5 vdd
rlabel space 4576 2909 4605 2918 5 gnd
rlabel locali 4673 2907 4702 2913 5 gnd
rlabel locali 4886 2907 4915 2913 5 gnd
rlabel nwell 4522 2644 4545 2647 5 vdd
rlabel locali 4944 2787 4966 2802 5 d0
rlabel locali 4670 2611 4699 2617 5 vdd
rlabel locali 4883 2608 4912 2614 5 vdd
rlabel locali 3663 2322 3692 2328 5 vdd
rlabel locali 3450 2325 3479 2331 5 vdd
rlabel nwell 3302 2358 3325 2361 5 vdd
rlabel locali 3666 2621 3695 2627 5 gnd
rlabel locali 3453 2621 3482 2627 5 gnd
rlabel space 3356 2623 3385 2632 5 gnd
rlabel locali 3722 2499 3754 2518 5 d3
rlabel locali 3702 6416 3734 6435 5 d3
rlabel space 3336 6540 3365 6549 5 gnd
rlabel locali 3433 6538 3462 6544 5 gnd
rlabel locali 3646 6538 3675 6544 5 gnd
rlabel nwell 3282 6275 3305 6278 5 vdd
rlabel locali 3430 6242 3459 6248 5 vdd
rlabel locali 3643 6239 3672 6245 5 vdd
rlabel locali 4863 6525 4892 6531 5 vdd
rlabel locali 4650 6528 4679 6534 5 vdd
rlabel locali 4924 6704 4946 6719 5 d0
rlabel nwell 4502 6561 4525 6564 5 vdd
rlabel locali 4866 6824 4895 6830 5 gnd
rlabel locali 4653 6824 4682 6830 5 gnd
rlabel space 4556 6826 4585 6835 5 gnd
rlabel locali 4864 6940 4893 6946 5 vdd
rlabel locali 4651 6943 4680 6949 5 vdd
rlabel locali 4925 7119 4947 7134 5 d0
rlabel nwell 4503 6976 4526 6979 5 vdd
rlabel locali 4867 7239 4896 7245 5 gnd
rlabel locali 4654 7239 4683 7245 5 gnd
rlabel space 4557 7241 4586 7250 5 gnd
rlabel locali 3851 6706 3880 6712 5 vdd
rlabel locali 3638 6709 3667 6715 5 vdd
rlabel nwell 3490 6742 3513 6745 5 vdd
rlabel locali 3854 7005 3883 7011 5 gnd
rlabel locali 3641 7005 3670 7011 5 gnd
rlabel space 3544 7007 3573 7016 5 gnd
rlabel locali 3895 6880 3942 6901 5 d1
rlabel locali 4858 7506 4887 7512 5 vdd
rlabel locali 4645 7509 4674 7515 5 vdd
rlabel locali 4919 7685 4941 7700 5 d0
rlabel nwell 4497 7542 4520 7545 5 vdd
rlabel locali 4861 7805 4890 7811 5 gnd
rlabel locali 4648 7805 4677 7811 5 gnd
rlabel space 4551 7807 4580 7816 5 gnd
rlabel locali 4859 7921 4888 7927 5 vdd
rlabel locali 4646 7924 4675 7930 5 vdd
rlabel locali 4920 8100 4942 8115 5 d0
rlabel nwell 4498 7957 4521 7960 5 vdd
rlabel locali 4862 8220 4891 8226 5 gnd
rlabel locali 4649 8220 4678 8226 5 gnd
rlabel space 4552 8222 4581 8231 5 gnd
rlabel locali 3846 7687 3875 7693 5 vdd
rlabel locali 3633 7690 3662 7696 5 vdd
rlabel nwell 3485 7723 3508 7726 5 vdd
rlabel locali 3849 7986 3878 7992 5 gnd
rlabel locali 3636 7986 3665 7992 5 gnd
rlabel space 3539 7988 3568 7997 5 gnd
rlabel locali 3890 7861 3937 7882 5 d1
rlabel locali 3796 7267 3825 7273 5 vdd
rlabel locali 3583 7270 3612 7276 5 vdd
rlabel nwell 3435 7303 3458 7306 5 vdd
rlabel locali 3799 7566 3828 7572 5 gnd
rlabel locali 3586 7566 3615 7572 5 gnd
rlabel space 3489 7568 3518 7577 5 gnd
rlabel locali 3859 7446 3882 7461 5 d2
rlabel space 4564 6262 4593 6271 5 gnd
rlabel locali 3871 5486 3894 5501 5 d2
rlabel space 3501 5608 3530 5617 5 gnd
rlabel locali 3598 5606 3627 5612 5 gnd
rlabel locali 3811 5606 3840 5612 5 gnd
rlabel nwell 3447 5343 3470 5346 5 vdd
rlabel locali 3595 5310 3624 5316 5 vdd
rlabel locali 3808 5307 3837 5313 5 vdd
rlabel locali 3902 5901 3949 5922 5 d1
rlabel space 3551 6028 3580 6037 5 gnd
rlabel locali 3648 6026 3677 6032 5 gnd
rlabel locali 3861 6026 3890 6032 5 gnd
rlabel nwell 3497 5763 3520 5766 5 vdd
rlabel locali 3645 5730 3674 5736 5 vdd
rlabel locali 3858 5727 3887 5733 5 vdd
rlabel locali 4661 6260 4690 6266 5 gnd
rlabel locali 4874 6260 4903 6266 5 gnd
rlabel nwell 4510 5997 4533 6000 5 vdd
rlabel locali 4932 6140 4954 6155 5 d0
rlabel locali 4658 5964 4687 5970 5 vdd
rlabel locali 4871 5961 4900 5967 5 vdd
rlabel space 4563 5847 4592 5856 5 gnd
rlabel locali 4660 5845 4689 5851 5 gnd
rlabel locali 4873 5845 4902 5851 5 gnd
rlabel nwell 4509 5582 4532 5585 5 vdd
rlabel locali 4931 5725 4953 5740 5 d0
rlabel locali 4657 5549 4686 5555 5 vdd
rlabel locali 4870 5546 4899 5552 5 vdd
rlabel locali 3907 4920 3954 4941 5 d1
rlabel space 3556 5047 3585 5056 5 gnd
rlabel locali 3653 5045 3682 5051 5 gnd
rlabel locali 3866 5045 3895 5051 5 gnd
rlabel nwell 3502 4782 3525 4785 5 vdd
rlabel locali 3650 4749 3679 4755 5 vdd
rlabel locali 3863 4746 3892 4752 5 vdd
rlabel space 4569 5281 4598 5290 5 gnd
rlabel locali 4666 5279 4695 5285 5 gnd
rlabel locali 4879 5279 4908 5285 5 gnd
rlabel nwell 4515 5016 4538 5019 5 vdd
rlabel locali 4937 5159 4959 5174 5 d0
rlabel locali 4663 4983 4692 4989 5 vdd
rlabel locali 4876 4980 4905 4986 5 vdd
rlabel space 4568 4866 4597 4875 5 gnd
rlabel locali 4665 4864 4694 4870 5 gnd
rlabel locali 4878 4864 4907 4870 5 gnd
rlabel nwell 4514 4601 4537 4604 5 vdd
rlabel locali 4936 4744 4958 4759 5 d0
rlabel locali 4662 4568 4691 4574 5 vdd
rlabel locali 4875 4565 4904 4571 5 vdd
rlabel locali 3568 4314 3597 4320 5 vdd
rlabel locali 3355 4317 3384 4323 5 vdd
rlabel nwell 3207 4350 3230 4353 5 vdd
rlabel locali 3571 4613 3600 4619 5 gnd
rlabel locali 3358 4613 3387 4619 5 gnd
rlabel space 3261 4615 3290 4624 5 gnd
rlabel locali 3633 4490 3655 4514 5 d4
rlabel locali 1743 319 1772 325 1 vdd
rlabel locali 1956 316 1985 322 1 vdd
rlabel nwell 2110 286 2133 289 1 vdd
rlabel locali 1740 20 1769 26 1 gnd
rlabel locali 1953 20 1982 26 1 gnd
rlabel space 2050 15 2079 24 1 gnd
rlabel locali 1685 128 1709 145 1 d5
rlabel locali 5585 8052 5614 8058 1 vdd
rlabel locali 5798 8049 5827 8055 1 vdd
rlabel locali 5531 7864 5553 7879 1 d0
rlabel nwell 5952 8019 5975 8022 1 vdd
rlabel locali 5582 7753 5611 7759 1 gnd
rlabel locali 5795 7753 5824 7759 1 gnd
rlabel space 5892 7748 5921 7757 1 gnd
rlabel locali 5584 7637 5613 7643 1 vdd
rlabel locali 5797 7634 5826 7640 1 vdd
rlabel locali 5530 7449 5552 7464 1 d0
rlabel nwell 5951 7604 5974 7607 1 vdd
rlabel locali 5581 7338 5610 7344 1 gnd
rlabel locali 5794 7338 5823 7344 1 gnd
rlabel space 5891 7333 5920 7342 1 gnd
rlabel locali 6597 7871 6626 7877 1 vdd
rlabel locali 6810 7868 6839 7874 1 vdd
rlabel nwell 6964 7838 6987 7841 1 vdd
rlabel locali 6594 7572 6623 7578 1 gnd
rlabel locali 6807 7572 6836 7578 1 gnd
rlabel space 6904 7567 6933 7576 1 gnd
rlabel locali 6535 7682 6582 7703 1 d1
rlabel locali 5590 7071 5619 7077 1 vdd
rlabel locali 5803 7068 5832 7074 1 vdd
rlabel locali 5536 6883 5558 6898 1 d0
rlabel nwell 5957 7038 5980 7041 1 vdd
rlabel locali 5587 6772 5616 6778 1 gnd
rlabel locali 5800 6772 5829 6778 1 gnd
rlabel space 5897 6767 5926 6776 1 gnd
rlabel locali 5589 6656 5618 6662 1 vdd
rlabel locali 5802 6653 5831 6659 1 vdd
rlabel locali 5535 6468 5557 6483 1 d0
rlabel nwell 5956 6623 5979 6626 1 vdd
rlabel locali 5586 6357 5615 6363 1 gnd
rlabel locali 5799 6357 5828 6363 1 gnd
rlabel locali 6602 6890 6631 6896 1 vdd
rlabel locali 6815 6887 6844 6893 1 vdd
rlabel nwell 6969 6857 6992 6860 1 vdd
rlabel locali 6599 6591 6628 6597 1 gnd
rlabel locali 6812 6591 6841 6597 1 gnd
rlabel space 6909 6586 6938 6595 1 gnd
rlabel locali 6540 6701 6587 6722 1 d1
rlabel locali 6652 7310 6681 7316 1 vdd
rlabel locali 6865 7307 6894 7313 1 vdd
rlabel nwell 7019 7277 7042 7280 1 vdd
rlabel locali 6649 7011 6678 7017 1 gnd
rlabel locali 6862 7011 6891 7017 1 gnd
rlabel space 6959 7006 6988 7015 1 gnd
rlabel locali 6595 7122 6618 7137 1 d2
rlabel space 5896 6352 5925 6361 1 gnd
rlabel locali 6607 5162 6630 5177 1 d2
rlabel space 6971 5046 7000 5055 1 gnd
rlabel locali 6874 5051 6903 5057 1 gnd
rlabel locali 6661 5051 6690 5057 1 gnd
rlabel nwell 7031 5317 7054 5320 1 vdd
rlabel locali 6877 5347 6906 5353 1 vdd
rlabel locali 6664 5350 6693 5356 1 vdd
rlabel locali 6552 4741 6599 4762 1 d1
rlabel space 6921 4626 6950 4635 1 gnd
rlabel locali 6824 4631 6853 4637 1 gnd
rlabel locali 6611 4631 6640 4637 1 gnd
rlabel nwell 6981 4897 7004 4900 1 vdd
rlabel locali 6827 4927 6856 4933 1 vdd
rlabel locali 6614 4930 6643 4936 1 vdd
rlabel space 5908 4392 5937 4401 1 gnd
rlabel locali 5811 4397 5840 4403 1 gnd
rlabel locali 5598 4397 5627 4403 1 gnd
rlabel nwell 5968 4663 5991 4666 1 vdd
rlabel locali 5547 4508 5569 4523 1 d0
rlabel locali 5814 4693 5843 4699 1 vdd
rlabel locali 5601 4696 5630 4702 1 vdd
rlabel space 5909 4807 5938 4816 1 gnd
rlabel locali 5812 4812 5841 4818 1 gnd
rlabel locali 5599 4812 5628 4818 1 gnd
rlabel nwell 5969 5078 5992 5081 1 vdd
rlabel locali 5548 4923 5570 4938 1 d0
rlabel locali 5815 5108 5844 5114 1 vdd
rlabel locali 5602 5111 5631 5117 1 vdd
rlabel locali 6547 5722 6594 5743 1 d1
rlabel space 6916 5607 6945 5616 1 gnd
rlabel locali 6819 5612 6848 5618 1 gnd
rlabel locali 6606 5612 6635 5618 1 gnd
rlabel nwell 6976 5878 6999 5881 1 vdd
rlabel locali 6822 5908 6851 5914 1 vdd
rlabel locali 6609 5911 6638 5917 1 vdd
rlabel space 5903 5373 5932 5382 1 gnd
rlabel locali 5806 5378 5835 5384 1 gnd
rlabel locali 5593 5378 5622 5384 1 gnd
rlabel nwell 5963 5644 5986 5647 1 vdd
rlabel locali 5542 5489 5564 5504 1 d0
rlabel locali 5809 5674 5838 5680 1 vdd
rlabel locali 5596 5677 5625 5683 1 vdd
rlabel space 5904 5788 5933 5797 1 gnd
rlabel locali 5807 5793 5836 5799 1 gnd
rlabel locali 5594 5793 5623 5799 1 gnd
rlabel nwell 5964 6059 5987 6062 1 vdd
rlabel locali 5543 5904 5565 5919 1 d0
rlabel locali 5810 6089 5839 6095 1 vdd
rlabel locali 5597 6092 5626 6098 1 vdd
rlabel locali 6817 6378 6846 6384 1 vdd
rlabel locali 7030 6375 7059 6381 1 vdd
rlabel nwell 7184 6345 7207 6348 1 vdd
rlabel locali 6814 6079 6843 6085 1 gnd
rlabel locali 7027 6079 7056 6085 1 gnd
rlabel space 7124 6074 7153 6083 1 gnd
rlabel locali 6755 6188 6787 6207 1 d3
rlabel locali 6775 2271 6807 2290 1 d3
rlabel space 7144 2157 7173 2166 1 gnd
rlabel locali 7047 2162 7076 2168 1 gnd
rlabel locali 6834 2162 6863 2168 1 gnd
rlabel nwell 7204 2428 7227 2431 1 vdd
rlabel locali 7050 2458 7079 2464 1 vdd
rlabel locali 6837 2461 6866 2467 1 vdd
rlabel locali 5617 2175 5646 2181 1 vdd
rlabel locali 5830 2172 5859 2178 1 vdd
rlabel locali 5563 1987 5585 2002 1 d0
rlabel nwell 5984 2142 6007 2145 1 vdd
rlabel locali 5614 1876 5643 1882 1 gnd
rlabel locali 5827 1876 5856 1882 1 gnd
rlabel space 5924 1871 5953 1880 1 gnd
rlabel locali 5616 1760 5645 1766 1 vdd
rlabel locali 5829 1757 5858 1763 1 vdd
rlabel locali 5562 1572 5584 1587 1 d0
rlabel nwell 5983 1727 6006 1730 1 vdd
rlabel locali 5613 1461 5642 1467 1 gnd
rlabel locali 5826 1461 5855 1467 1 gnd
rlabel space 5923 1456 5952 1465 1 gnd
rlabel locali 6629 1994 6658 2000 1 vdd
rlabel locali 6842 1991 6871 1997 1 vdd
rlabel nwell 6996 1961 7019 1964 1 vdd
rlabel locali 6626 1695 6655 1701 1 gnd
rlabel locali 6839 1695 6868 1701 1 gnd
rlabel space 6936 1690 6965 1699 1 gnd
rlabel locali 6567 1805 6614 1826 1 d1
rlabel locali 5622 1194 5651 1200 1 vdd
rlabel locali 5835 1191 5864 1197 1 vdd
rlabel locali 5568 1006 5590 1021 1 d0
rlabel nwell 5989 1161 6012 1164 1 vdd
rlabel locali 5619 895 5648 901 1 gnd
rlabel locali 5832 895 5861 901 1 gnd
rlabel space 5929 890 5958 899 1 gnd
rlabel locali 5621 779 5650 785 1 vdd
rlabel locali 5834 776 5863 782 1 vdd
rlabel locali 5567 591 5589 606 1 d0
rlabel nwell 5988 746 6011 749 1 vdd
rlabel locali 5618 480 5647 486 1 gnd
rlabel locali 5831 480 5860 486 1 gnd
rlabel space 5928 475 5957 484 1 gnd
rlabel locali 6634 1013 6663 1019 1 vdd
rlabel locali 6847 1010 6876 1016 1 vdd
rlabel nwell 7001 980 7024 983 1 vdd
rlabel locali 6631 714 6660 720 1 gnd
rlabel locali 6844 714 6873 720 1 gnd
rlabel space 6941 709 6970 718 1 gnd
rlabel locali 6572 824 6619 845 1 d1
rlabel locali 6684 1433 6713 1439 1 vdd
rlabel locali 6897 1430 6926 1436 1 vdd
rlabel nwell 7051 1400 7074 1403 1 vdd
rlabel locali 6681 1134 6710 1140 1 gnd
rlabel locali 6894 1134 6923 1140 1 gnd
rlabel space 6991 1129 7020 1138 1 gnd
rlabel locali 6627 1245 6650 1260 1 d2
rlabel space 5916 2435 5945 2444 1 gnd
rlabel locali 6615 3205 6638 3220 1 d2
rlabel space 6979 3089 7008 3098 1 gnd
rlabel locali 6882 3094 6911 3100 1 gnd
rlabel locali 6669 3094 6698 3100 1 gnd
rlabel nwell 7039 3360 7062 3363 1 vdd
rlabel locali 6885 3390 6914 3396 1 vdd
rlabel locali 6672 3393 6701 3399 1 vdd
rlabel locali 6560 2784 6607 2805 1 d1
rlabel space 6929 2669 6958 2678 1 gnd
rlabel locali 6832 2674 6861 2680 1 gnd
rlabel locali 6619 2674 6648 2680 1 gnd
rlabel nwell 6989 2940 7012 2943 1 vdd
rlabel locali 6835 2970 6864 2976 1 vdd
rlabel locali 6622 2973 6651 2979 1 vdd
rlabel locali 5819 2440 5848 2446 1 gnd
rlabel locali 5606 2440 5635 2446 1 gnd
rlabel nwell 5976 2706 5999 2709 1 vdd
rlabel locali 5555 2551 5577 2566 1 d0
rlabel locali 5822 2736 5851 2742 1 vdd
rlabel locali 5609 2739 5638 2745 1 vdd
rlabel space 5917 2850 5946 2859 1 gnd
rlabel locali 5820 2855 5849 2861 1 gnd
rlabel locali 5607 2855 5636 2861 1 gnd
rlabel nwell 5977 3121 6000 3124 1 vdd
rlabel locali 5556 2966 5578 2981 1 d0
rlabel locali 5823 3151 5852 3157 1 vdd
rlabel locali 5610 3154 5639 3160 1 vdd
rlabel locali 6555 3765 6602 3786 1 d1
rlabel space 6924 3650 6953 3659 1 gnd
rlabel locali 6827 3655 6856 3661 1 gnd
rlabel locali 6614 3655 6643 3661 1 gnd
rlabel nwell 6984 3921 7007 3924 1 vdd
rlabel locali 6830 3951 6859 3957 1 vdd
rlabel locali 6617 3954 6646 3960 1 vdd
rlabel space 5911 3416 5940 3425 1 gnd
rlabel locali 5814 3421 5843 3427 1 gnd
rlabel locali 5601 3421 5630 3427 1 gnd
rlabel nwell 5971 3687 5994 3690 1 vdd
rlabel locali 5550 3532 5572 3547 1 d0
rlabel locali 5817 3717 5846 3723 1 vdd
rlabel locali 5604 3720 5633 3726 1 vdd
rlabel space 5912 3831 5941 3840 1 gnd
rlabel locali 5815 3836 5844 3842 1 gnd
rlabel locali 5602 3836 5631 3842 1 gnd
rlabel nwell 5972 4102 5995 4105 1 vdd
rlabel locali 5551 3947 5573 3962 1 d0
rlabel locali 5818 4132 5847 4138 1 vdd
rlabel locali 5605 4135 5634 4141 1 vdd
rlabel locali 6912 4386 6941 4392 1 vdd
rlabel locali 7125 4383 7154 4389 1 vdd
rlabel nwell 7279 4353 7302 4356 1 vdd
rlabel locali 6909 4087 6938 4093 1 gnd
rlabel locali 7122 4087 7151 4093 1 gnd
rlabel space 7219 4082 7248 4091 1 gnd
rlabel locali 6854 4192 6876 4216 1 d4
rlabel locali 10176 627 10205 633 5 vdd
rlabel locali 9963 630 9992 636 5 vdd
rlabel locali 10237 806 10259 821 5 d0
rlabel nwell 9815 663 9838 666 5 vdd
rlabel locali 10179 926 10208 932 5 gnd
rlabel locali 9966 926 9995 932 5 gnd
rlabel space 9869 928 9898 937 5 gnd
rlabel locali 10177 1042 10206 1048 5 vdd
rlabel locali 9964 1045 9993 1051 5 vdd
rlabel locali 10238 1221 10260 1236 5 d0
rlabel nwell 9816 1078 9839 1081 5 vdd
rlabel locali 10180 1341 10209 1347 5 gnd
rlabel locali 9967 1341 9996 1347 5 gnd
rlabel space 9870 1343 9899 1352 5 gnd
rlabel locali 9164 808 9193 814 5 vdd
rlabel locali 8951 811 8980 817 5 vdd
rlabel nwell 8803 844 8826 847 5 vdd
rlabel locali 9167 1107 9196 1113 5 gnd
rlabel locali 8954 1107 8983 1113 5 gnd
rlabel space 8857 1109 8886 1118 5 gnd
rlabel locali 9208 982 9255 1003 5 d1
rlabel locali 10171 1608 10200 1614 5 vdd
rlabel locali 9958 1611 9987 1617 5 vdd
rlabel locali 10232 1787 10254 1802 5 d0
rlabel nwell 9810 1644 9833 1647 5 vdd
rlabel locali 10174 1907 10203 1913 5 gnd
rlabel locali 9961 1907 9990 1913 5 gnd
rlabel space 9864 1909 9893 1918 5 gnd
rlabel locali 10172 2023 10201 2029 5 vdd
rlabel locali 9959 2026 9988 2032 5 vdd
rlabel locali 10233 2202 10255 2217 5 d0
rlabel nwell 9811 2059 9834 2062 5 vdd
rlabel locali 10175 2322 10204 2328 5 gnd
rlabel locali 9962 2322 9991 2328 5 gnd
rlabel locali 9159 1789 9188 1795 5 vdd
rlabel locali 8946 1792 8975 1798 5 vdd
rlabel nwell 8798 1825 8821 1828 5 vdd
rlabel locali 9162 2088 9191 2094 5 gnd
rlabel locali 8949 2088 8978 2094 5 gnd
rlabel space 8852 2090 8881 2099 5 gnd
rlabel locali 9203 1963 9250 1984 5 d1
rlabel locali 9109 1369 9138 1375 5 vdd
rlabel locali 8896 1372 8925 1378 5 vdd
rlabel nwell 8748 1405 8771 1408 5 vdd
rlabel locali 9112 1668 9141 1674 5 gnd
rlabel locali 8899 1668 8928 1674 5 gnd
rlabel space 8802 1670 8831 1679 5 gnd
rlabel locali 9172 1548 9195 1563 5 d2
rlabel space 9865 2324 9894 2333 5 gnd
rlabel locali 9160 3508 9183 3523 5 d2
rlabel space 8790 3630 8819 3639 5 gnd
rlabel locali 8887 3628 8916 3634 5 gnd
rlabel locali 9100 3628 9129 3634 5 gnd
rlabel nwell 8736 3365 8759 3368 5 vdd
rlabel locali 8884 3332 8913 3338 5 vdd
rlabel locali 9097 3329 9126 3335 5 vdd
rlabel locali 9191 3923 9238 3944 5 d1
rlabel space 8840 4050 8869 4059 5 gnd
rlabel locali 8937 4048 8966 4054 5 gnd
rlabel locali 9150 4048 9179 4054 5 gnd
rlabel nwell 8786 3785 8809 3788 5 vdd
rlabel locali 8934 3752 8963 3758 5 vdd
rlabel locali 9147 3749 9176 3755 5 vdd
rlabel space 9853 4284 9882 4293 5 gnd
rlabel locali 9950 4282 9979 4288 5 gnd
rlabel locali 10163 4282 10192 4288 5 gnd
rlabel nwell 9799 4019 9822 4022 5 vdd
rlabel locali 10221 4162 10243 4177 5 d0
rlabel locali 9947 3986 9976 3992 5 vdd
rlabel locali 10160 3983 10189 3989 5 vdd
rlabel space 9852 3869 9881 3878 5 gnd
rlabel locali 9949 3867 9978 3873 5 gnd
rlabel locali 10162 3867 10191 3873 5 gnd
rlabel nwell 9798 3604 9821 3607 5 vdd
rlabel locali 10220 3747 10242 3762 5 d0
rlabel locali 9946 3571 9975 3577 5 vdd
rlabel locali 10159 3568 10188 3574 5 vdd
rlabel locali 9196 2942 9243 2963 5 d1
rlabel space 8845 3069 8874 3078 5 gnd
rlabel locali 8942 3067 8971 3073 5 gnd
rlabel locali 9155 3067 9184 3073 5 gnd
rlabel nwell 8791 2804 8814 2807 5 vdd
rlabel locali 8939 2771 8968 2777 5 vdd
rlabel locali 9152 2768 9181 2774 5 vdd
rlabel space 9858 3303 9887 3312 5 gnd
rlabel locali 9955 3301 9984 3307 5 gnd
rlabel locali 10168 3301 10197 3307 5 gnd
rlabel nwell 9804 3038 9827 3041 5 vdd
rlabel locali 10226 3181 10248 3196 5 d0
rlabel locali 9952 3005 9981 3011 5 vdd
rlabel locali 10165 3002 10194 3008 5 vdd
rlabel space 9857 2888 9886 2897 5 gnd
rlabel locali 9954 2886 9983 2892 5 gnd
rlabel locali 10167 2886 10196 2892 5 gnd
rlabel nwell 9803 2623 9826 2626 5 vdd
rlabel locali 10225 2766 10247 2781 5 d0
rlabel locali 9951 2590 9980 2596 5 vdd
rlabel locali 10164 2587 10193 2593 5 vdd
rlabel locali 8944 2301 8973 2307 5 vdd
rlabel locali 8731 2304 8760 2310 5 vdd
rlabel nwell 8583 2337 8606 2340 5 vdd
rlabel locali 8947 2600 8976 2606 5 gnd
rlabel locali 8734 2600 8763 2606 5 gnd
rlabel space 8637 2602 8666 2611 5 gnd
rlabel locali 9003 2478 9035 2497 5 d3
rlabel locali 8983 6395 9015 6414 5 d3
rlabel space 8617 6519 8646 6528 5 gnd
rlabel locali 8714 6517 8743 6523 5 gnd
rlabel locali 8927 6517 8956 6523 5 gnd
rlabel nwell 8563 6254 8586 6257 5 vdd
rlabel locali 8711 6221 8740 6227 5 vdd
rlabel locali 8924 6218 8953 6224 5 vdd
rlabel locali 10144 6504 10173 6510 5 vdd
rlabel locali 9931 6507 9960 6513 5 vdd
rlabel locali 10205 6683 10227 6698 5 d0
rlabel nwell 9783 6540 9806 6543 5 vdd
rlabel locali 10147 6803 10176 6809 5 gnd
rlabel locali 9934 6803 9963 6809 5 gnd
rlabel space 9837 6805 9866 6814 5 gnd
rlabel locali 10145 6919 10174 6925 5 vdd
rlabel locali 9932 6922 9961 6928 5 vdd
rlabel locali 10206 7098 10228 7113 5 d0
rlabel nwell 9784 6955 9807 6958 5 vdd
rlabel locali 10148 7218 10177 7224 5 gnd
rlabel locali 9935 7218 9964 7224 5 gnd
rlabel space 9838 7220 9867 7229 5 gnd
rlabel locali 9132 6685 9161 6691 5 vdd
rlabel locali 8919 6688 8948 6694 5 vdd
rlabel nwell 8771 6721 8794 6724 5 vdd
rlabel locali 9135 6984 9164 6990 5 gnd
rlabel locali 8922 6984 8951 6990 5 gnd
rlabel space 8825 6986 8854 6995 5 gnd
rlabel locali 9176 6859 9223 6880 5 d1
rlabel locali 10139 7485 10168 7491 5 vdd
rlabel locali 9926 7488 9955 7494 5 vdd
rlabel locali 10200 7664 10222 7679 5 d0
rlabel nwell 9778 7521 9801 7524 5 vdd
rlabel locali 10142 7784 10171 7790 5 gnd
rlabel locali 9929 7784 9958 7790 5 gnd
rlabel space 9832 7786 9861 7795 5 gnd
rlabel locali 10140 7900 10169 7906 5 vdd
rlabel locali 9927 7903 9956 7909 5 vdd
rlabel locali 10201 8079 10223 8094 5 d0
rlabel nwell 9779 7936 9802 7939 5 vdd
rlabel locali 10143 8199 10172 8205 5 gnd
rlabel locali 9930 8199 9959 8205 5 gnd
rlabel space 9833 8201 9862 8210 5 gnd
rlabel locali 9127 7666 9156 7672 5 vdd
rlabel locali 8914 7669 8943 7675 5 vdd
rlabel nwell 8766 7702 8789 7705 5 vdd
rlabel locali 9130 7965 9159 7971 5 gnd
rlabel locali 8917 7965 8946 7971 5 gnd
rlabel space 8820 7967 8849 7976 5 gnd
rlabel locali 9171 7840 9218 7861 5 d1
rlabel locali 10324 8241 10351 8254 5 gnd
rlabel locali 9077 7246 9106 7252 5 vdd
rlabel locali 8864 7249 8893 7255 5 vdd
rlabel nwell 8716 7282 8739 7285 5 vdd
rlabel locali 9080 7545 9109 7551 5 gnd
rlabel locali 8867 7545 8896 7551 5 gnd
rlabel space 8770 7547 8799 7556 5 gnd
rlabel locali 9140 7425 9163 7440 5 d2
rlabel space 9845 6241 9874 6250 5 gnd
rlabel locali 9152 5465 9175 5480 5 d2
rlabel space 8782 5587 8811 5596 5 gnd
rlabel locali 8879 5585 8908 5591 5 gnd
rlabel locali 9092 5585 9121 5591 5 gnd
rlabel nwell 8728 5322 8751 5325 5 vdd
rlabel locali 8876 5289 8905 5295 5 vdd
rlabel locali 9089 5286 9118 5292 5 vdd
rlabel locali 9183 5880 9230 5901 5 d1
rlabel space 8832 6007 8861 6016 5 gnd
rlabel locali 8929 6005 8958 6011 5 gnd
rlabel locali 9142 6005 9171 6011 5 gnd
rlabel nwell 8778 5742 8801 5745 5 vdd
rlabel locali 8926 5709 8955 5715 5 vdd
rlabel locali 9139 5706 9168 5712 5 vdd
rlabel locali 9942 6239 9971 6245 5 gnd
rlabel locali 10155 6239 10184 6245 5 gnd
rlabel nwell 9791 5976 9814 5979 5 vdd
rlabel locali 10213 6119 10235 6134 5 d0
rlabel locali 9939 5943 9968 5949 5 vdd
rlabel locali 10152 5940 10181 5946 5 vdd
rlabel space 9844 5826 9873 5835 5 gnd
rlabel locali 9941 5824 9970 5830 5 gnd
rlabel locali 10154 5824 10183 5830 5 gnd
rlabel nwell 9790 5561 9813 5564 5 vdd
rlabel locali 10212 5704 10234 5719 5 d0
rlabel locali 9938 5528 9967 5534 5 vdd
rlabel locali 10151 5525 10180 5531 5 vdd
rlabel locali 9188 4899 9235 4920 5 d1
rlabel space 8837 5026 8866 5035 5 gnd
rlabel locali 8934 5024 8963 5030 5 gnd
rlabel locali 9147 5024 9176 5030 5 gnd
rlabel nwell 8783 4761 8806 4764 5 vdd
rlabel locali 8931 4728 8960 4734 5 vdd
rlabel locali 9144 4725 9173 4731 5 vdd
rlabel space 9850 5260 9879 5269 5 gnd
rlabel locali 9947 5258 9976 5264 5 gnd
rlabel locali 10160 5258 10189 5264 5 gnd
rlabel nwell 9796 4995 9819 4998 5 vdd
rlabel locali 10218 5138 10240 5153 5 d0
rlabel locali 9944 4962 9973 4968 5 vdd
rlabel locali 10157 4959 10186 4965 5 vdd
rlabel space 9849 4845 9878 4854 5 gnd
rlabel locali 9946 4843 9975 4849 5 gnd
rlabel locali 10159 4843 10188 4849 5 gnd
rlabel nwell 9795 4580 9818 4583 5 vdd
rlabel locali 10217 4723 10239 4738 5 d0
rlabel locali 9943 4547 9972 4553 5 vdd
rlabel locali 10156 4544 10185 4550 5 vdd
rlabel locali 8849 4293 8878 4299 5 vdd
rlabel locali 8636 4296 8665 4302 5 vdd
rlabel nwell 8488 4329 8511 4332 5 vdd
rlabel locali 8852 4592 8881 4598 5 gnd
rlabel locali 8639 4592 8668 4598 5 gnd
rlabel space 8542 4594 8571 4603 5 gnd
rlabel locali 8914 4469 8936 4493 5 d4
rlabel locali 7024 298 7053 304 1 vdd
rlabel locali 7237 295 7266 301 1 vdd
rlabel nwell 7391 265 7414 268 1 vdd
rlabel locali 7021 -1 7050 5 1 gnd
rlabel locali 7234 -1 7263 5 1 gnd
rlabel space 7331 -6 7360 3 1 gnd
rlabel locali 6966 107 6990 124 1 d5
rlabel locali 4833 231 4862 237 1 vdd
rlabel locali 5046 228 5075 234 1 vdd
rlabel locali 5409 78 5431 93 1 vout
rlabel nwell 5200 198 5223 201 1 vdd
rlabel locali 4830 -68 4859 -62 1 gnd
rlabel locali 5043 -68 5072 -62 1 gnd
rlabel space 5140 -73 5169 -64 1 gnd
rlabel locali 4777 38 4796 58 1 d6
<< end >>
