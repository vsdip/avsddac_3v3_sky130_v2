magic
tech sky130A
timestamp 1620567848
<< nwell >>
rect 318 9221 645 9295
rect 5374 9262 5701 9336
rect 318 9071 1129 9221
rect 1256 8977 1583 9051
rect 3801 9001 4612 9151
rect 5374 9112 6185 9262
rect 1256 8827 2067 8977
rect 4285 8927 4612 9001
rect 6312 9018 6639 9092
rect 8857 9042 9668 9192
rect 6312 8868 7123 9018
rect 9341 8968 9668 9042
rect 317 8667 644 8741
rect 2862 8691 3673 8841
rect 317 8517 1128 8667
rect 3346 8617 3673 8691
rect 5373 8708 5700 8782
rect 7918 8732 8729 8882
rect 1397 8385 1724 8459
rect 3800 8447 4611 8597
rect 5373 8558 6184 8708
rect 8402 8658 8729 8732
rect 1397 8235 2208 8385
rect 4284 8373 4611 8447
rect 6453 8426 6780 8500
rect 8856 8488 9667 8638
rect 319 8118 646 8192
rect 2722 8180 3533 8330
rect 6453 8276 7264 8426
rect 9340 8414 9667 8488
rect 319 7968 1130 8118
rect 3206 8106 3533 8180
rect 5375 8159 5702 8233
rect 7778 8221 8589 8371
rect 1257 7874 1584 7948
rect 3802 7898 4613 8048
rect 5375 8009 6186 8159
rect 8262 8147 8589 8221
rect 1257 7724 2068 7874
rect 4286 7824 4613 7898
rect 6313 7915 6640 7989
rect 8858 7939 9669 8089
rect 6313 7765 7124 7915
rect 9342 7865 9669 7939
rect 318 7564 645 7638
rect 2863 7588 3674 7738
rect 318 7414 1129 7564
rect 3347 7514 3674 7588
rect 5374 7605 5701 7679
rect 7919 7629 8730 7779
rect 1367 7295 1694 7369
rect 3801 7344 4612 7494
rect 5374 7455 6185 7605
rect 8403 7555 8730 7629
rect 1367 7145 2178 7295
rect 4285 7270 4612 7344
rect 6423 7336 6750 7410
rect 8857 7385 9668 7535
rect 319 7015 646 7089
rect 2753 7064 3564 7214
rect 6423 7186 7234 7336
rect 9341 7311 9668 7385
rect 319 6865 1130 7015
rect 3237 6990 3564 7064
rect 5375 7056 5702 7130
rect 7809 7105 8620 7255
rect 1257 6771 1584 6845
rect 3802 6795 4613 6945
rect 5375 6906 6186 7056
rect 8293 7031 8620 7105
rect 1257 6621 2068 6771
rect 4286 6721 4613 6795
rect 6313 6812 6640 6886
rect 8858 6836 9669 6986
rect 6313 6662 7124 6812
rect 9342 6762 9669 6836
rect 318 6461 645 6535
rect 2863 6485 3674 6635
rect 318 6311 1129 6461
rect 3347 6411 3674 6485
rect 5374 6502 5701 6576
rect 7919 6526 8730 6676
rect 1398 6179 1725 6253
rect 3801 6241 4612 6391
rect 5374 6352 6185 6502
rect 8403 6452 8730 6526
rect 1398 6029 2209 6179
rect 4285 6167 4612 6241
rect 6454 6220 6781 6294
rect 8857 6282 9668 6432
rect 320 5912 647 5986
rect 2723 5974 3534 6124
rect 6454 6070 7265 6220
rect 9341 6208 9668 6282
rect 320 5762 1131 5912
rect 3207 5900 3534 5974
rect 5376 5953 5703 6027
rect 7779 6015 8590 6165
rect 1258 5668 1585 5742
rect 3803 5692 4614 5842
rect 5376 5803 6187 5953
rect 8263 5941 8590 6015
rect 1258 5518 2069 5668
rect 4287 5618 4614 5692
rect 6314 5709 6641 5783
rect 8859 5733 9670 5883
rect 6314 5559 7125 5709
rect 9343 5659 9670 5733
rect 319 5358 646 5432
rect 2864 5382 3675 5532
rect 319 5208 1130 5358
rect 3348 5308 3675 5382
rect 5375 5399 5702 5473
rect 7920 5423 8731 5573
rect 1367 5095 1694 5169
rect 3802 5138 4613 5288
rect 5375 5249 6186 5399
rect 8404 5349 8731 5423
rect 1367 4945 2178 5095
rect 4286 5064 4613 5138
rect 6423 5136 6750 5210
rect 8858 5179 9669 5329
rect 320 4809 647 4883
rect 2755 4852 3566 5002
rect 6423 4986 7234 5136
rect 9342 5105 9669 5179
rect 320 4659 1131 4809
rect 3239 4778 3566 4852
rect 5376 4850 5703 4924
rect 7811 4893 8622 5043
rect 1258 4565 1585 4639
rect 3803 4589 4614 4739
rect 5376 4700 6187 4850
rect 8295 4819 8622 4893
rect 1258 4415 2069 4565
rect 4287 4515 4614 4589
rect 6314 4606 6641 4680
rect 8859 4630 9670 4780
rect 6314 4456 7125 4606
rect 9343 4556 9670 4630
rect 319 4255 646 4329
rect 2864 4279 3675 4429
rect 319 4105 1130 4255
rect 3348 4205 3675 4279
rect 5375 4296 5702 4370
rect 7920 4320 8731 4470
rect 1399 3973 1726 4047
rect 3802 4035 4613 4185
rect 5375 4146 6186 4296
rect 8404 4246 8731 4320
rect 1399 3823 2210 3973
rect 4286 3961 4613 4035
rect 6455 4014 6782 4088
rect 8858 4076 9669 4226
rect 321 3706 648 3780
rect 2724 3768 3535 3918
rect 6455 3864 7266 4014
rect 9342 4002 9669 4076
rect 321 3556 1132 3706
rect 3208 3694 3535 3768
rect 5377 3747 5704 3821
rect 7780 3809 8591 3959
rect 1259 3462 1586 3536
rect 3804 3486 4615 3636
rect 5377 3597 6188 3747
rect 8264 3735 8591 3809
rect 1259 3312 2070 3462
rect 4288 3412 4615 3486
rect 6315 3503 6642 3577
rect 8860 3527 9671 3677
rect 6315 3353 7126 3503
rect 9344 3453 9671 3527
rect 320 3152 647 3226
rect 2865 3176 3676 3326
rect 320 3002 1131 3152
rect 3349 3102 3676 3176
rect 5376 3193 5703 3267
rect 7921 3217 8732 3367
rect 1369 2883 1696 2957
rect 3803 2932 4614 3082
rect 5376 3043 6187 3193
rect 8405 3143 8732 3217
rect 1369 2733 2180 2883
rect 4287 2858 4614 2932
rect 6425 2924 6752 2998
rect 8859 2973 9670 3123
rect 321 2603 648 2677
rect 2755 2652 3566 2802
rect 6425 2774 7236 2924
rect 9343 2899 9670 2973
rect 321 2453 1132 2603
rect 3239 2578 3566 2652
rect 5377 2644 5704 2718
rect 7811 2693 8622 2843
rect 1259 2359 1586 2433
rect 3804 2383 4615 2533
rect 5377 2494 6188 2644
rect 8295 2619 8622 2693
rect 1259 2209 2070 2359
rect 4288 2309 4615 2383
rect 6315 2400 6642 2474
rect 8860 2424 9671 2574
rect 6315 2250 7126 2400
rect 9344 2350 9671 2424
rect 320 2049 647 2123
rect 2865 2073 3676 2223
rect 320 1899 1131 2049
rect 3349 1999 3676 2073
rect 5376 2090 5703 2164
rect 7921 2114 8732 2264
rect 1400 1767 1727 1841
rect 3803 1829 4614 1979
rect 5376 1940 6187 2090
rect 8405 2040 8732 2114
rect 1400 1617 2211 1767
rect 4287 1755 4614 1829
rect 6456 1808 6783 1882
rect 8859 1870 9670 2020
rect 322 1500 649 1574
rect 2725 1562 3536 1712
rect 6456 1658 7267 1808
rect 9343 1796 9670 1870
rect 322 1350 1133 1500
rect 3209 1488 3536 1562
rect 5378 1541 5705 1615
rect 7781 1603 8592 1753
rect 1260 1256 1587 1330
rect 3805 1280 4616 1430
rect 5378 1391 6189 1541
rect 8265 1529 8592 1603
rect 1260 1106 2071 1256
rect 4289 1206 4616 1280
rect 6316 1297 6643 1371
rect 8861 1321 9672 1471
rect 6316 1147 7127 1297
rect 9345 1247 9672 1321
rect 321 946 648 1020
rect 2866 970 3677 1120
rect 321 796 1132 946
rect 3350 896 3677 970
rect 5377 987 5704 1061
rect 7922 1011 8733 1161
rect 3804 726 4615 876
rect 5377 837 6188 987
rect 8406 937 8733 1011
rect 8860 767 9671 917
rect 4288 652 4615 726
rect 9344 693 9671 767
rect 1568 387 1895 461
rect 1568 237 2379 387
rect 4518 367 4845 441
rect 6624 428 6951 502
rect 4518 217 5329 367
rect 6624 278 7435 428
<< nmos >>
rect 3869 9210 3919 9252
rect 4077 9210 4127 9252
rect 4285 9210 4335 9252
rect 4498 9210 4548 9252
rect 8925 9251 8975 9293
rect 9133 9251 9183 9293
rect 9341 9251 9391 9293
rect 9554 9251 9604 9293
rect 382 8970 432 9012
rect 595 8970 645 9012
rect 803 8970 853 9012
rect 1011 8970 1061 9012
rect 5438 9011 5488 9053
rect 5651 9011 5701 9053
rect 5859 9011 5909 9053
rect 6067 9011 6117 9053
rect 2930 8900 2980 8942
rect 3138 8900 3188 8942
rect 3346 8900 3396 8942
rect 3559 8900 3609 8942
rect 1320 8726 1370 8768
rect 1533 8726 1583 8768
rect 1741 8726 1791 8768
rect 1949 8726 1999 8768
rect 7986 8941 8036 8983
rect 8194 8941 8244 8983
rect 8402 8941 8452 8983
rect 8615 8941 8665 8983
rect 6376 8767 6426 8809
rect 6589 8767 6639 8809
rect 6797 8767 6847 8809
rect 7005 8767 7055 8809
rect 3868 8656 3918 8698
rect 4076 8656 4126 8698
rect 4284 8656 4334 8698
rect 4497 8656 4547 8698
rect 8924 8697 8974 8739
rect 9132 8697 9182 8739
rect 9340 8697 9390 8739
rect 9553 8697 9603 8739
rect 381 8416 431 8458
rect 594 8416 644 8458
rect 802 8416 852 8458
rect 1010 8416 1060 8458
rect 2790 8389 2840 8431
rect 2998 8389 3048 8431
rect 3206 8389 3256 8431
rect 3419 8389 3469 8431
rect 5437 8457 5487 8499
rect 5650 8457 5700 8499
rect 5858 8457 5908 8499
rect 6066 8457 6116 8499
rect 7846 8430 7896 8472
rect 8054 8430 8104 8472
rect 8262 8430 8312 8472
rect 8475 8430 8525 8472
rect 1461 8134 1511 8176
rect 1674 8134 1724 8176
rect 1882 8134 1932 8176
rect 2090 8134 2140 8176
rect 3870 8107 3920 8149
rect 4078 8107 4128 8149
rect 4286 8107 4336 8149
rect 4499 8107 4549 8149
rect 6517 8175 6567 8217
rect 6730 8175 6780 8217
rect 6938 8175 6988 8217
rect 7146 8175 7196 8217
rect 8926 8148 8976 8190
rect 9134 8148 9184 8190
rect 9342 8148 9392 8190
rect 9555 8148 9605 8190
rect 383 7867 433 7909
rect 596 7867 646 7909
rect 804 7867 854 7909
rect 1012 7867 1062 7909
rect 5439 7908 5489 7950
rect 5652 7908 5702 7950
rect 5860 7908 5910 7950
rect 6068 7908 6118 7950
rect 2931 7797 2981 7839
rect 3139 7797 3189 7839
rect 3347 7797 3397 7839
rect 3560 7797 3610 7839
rect 1321 7623 1371 7665
rect 1534 7623 1584 7665
rect 1742 7623 1792 7665
rect 1950 7623 2000 7665
rect 7987 7838 8037 7880
rect 8195 7838 8245 7880
rect 8403 7838 8453 7880
rect 8616 7838 8666 7880
rect 6377 7664 6427 7706
rect 6590 7664 6640 7706
rect 6798 7664 6848 7706
rect 7006 7664 7056 7706
rect 3869 7553 3919 7595
rect 4077 7553 4127 7595
rect 4285 7553 4335 7595
rect 4498 7553 4548 7595
rect 8925 7594 8975 7636
rect 9133 7594 9183 7636
rect 9341 7594 9391 7636
rect 9554 7594 9604 7636
rect 382 7313 432 7355
rect 595 7313 645 7355
rect 803 7313 853 7355
rect 1011 7313 1061 7355
rect 2821 7273 2871 7315
rect 3029 7273 3079 7315
rect 3237 7273 3287 7315
rect 3450 7273 3500 7315
rect 5438 7354 5488 7396
rect 5651 7354 5701 7396
rect 5859 7354 5909 7396
rect 6067 7354 6117 7396
rect 7877 7314 7927 7356
rect 8085 7314 8135 7356
rect 8293 7314 8343 7356
rect 8506 7314 8556 7356
rect 1431 7044 1481 7086
rect 1644 7044 1694 7086
rect 1852 7044 1902 7086
rect 2060 7044 2110 7086
rect 3870 7004 3920 7046
rect 4078 7004 4128 7046
rect 4286 7004 4336 7046
rect 4499 7004 4549 7046
rect 6487 7085 6537 7127
rect 6700 7085 6750 7127
rect 6908 7085 6958 7127
rect 7116 7085 7166 7127
rect 8926 7045 8976 7087
rect 9134 7045 9184 7087
rect 9342 7045 9392 7087
rect 9555 7045 9605 7087
rect 383 6764 433 6806
rect 596 6764 646 6806
rect 804 6764 854 6806
rect 1012 6764 1062 6806
rect 5439 6805 5489 6847
rect 5652 6805 5702 6847
rect 5860 6805 5910 6847
rect 6068 6805 6118 6847
rect 2931 6694 2981 6736
rect 3139 6694 3189 6736
rect 3347 6694 3397 6736
rect 3560 6694 3610 6736
rect 1321 6520 1371 6562
rect 1534 6520 1584 6562
rect 1742 6520 1792 6562
rect 1950 6520 2000 6562
rect 7987 6735 8037 6777
rect 8195 6735 8245 6777
rect 8403 6735 8453 6777
rect 8616 6735 8666 6777
rect 6377 6561 6427 6603
rect 6590 6561 6640 6603
rect 6798 6561 6848 6603
rect 7006 6561 7056 6603
rect 3869 6450 3919 6492
rect 4077 6450 4127 6492
rect 4285 6450 4335 6492
rect 4498 6450 4548 6492
rect 8925 6491 8975 6533
rect 9133 6491 9183 6533
rect 9341 6491 9391 6533
rect 9554 6491 9604 6533
rect 382 6210 432 6252
rect 595 6210 645 6252
rect 803 6210 853 6252
rect 1011 6210 1061 6252
rect 2791 6183 2841 6225
rect 2999 6183 3049 6225
rect 3207 6183 3257 6225
rect 3420 6183 3470 6225
rect 5438 6251 5488 6293
rect 5651 6251 5701 6293
rect 5859 6251 5909 6293
rect 6067 6251 6117 6293
rect 7847 6224 7897 6266
rect 8055 6224 8105 6266
rect 8263 6224 8313 6266
rect 8476 6224 8526 6266
rect 1462 5928 1512 5970
rect 1675 5928 1725 5970
rect 1883 5928 1933 5970
rect 2091 5928 2141 5970
rect 3871 5901 3921 5943
rect 4079 5901 4129 5943
rect 4287 5901 4337 5943
rect 4500 5901 4550 5943
rect 6518 5969 6568 6011
rect 6731 5969 6781 6011
rect 6939 5969 6989 6011
rect 7147 5969 7197 6011
rect 8927 5942 8977 5984
rect 9135 5942 9185 5984
rect 9343 5942 9393 5984
rect 9556 5942 9606 5984
rect 384 5661 434 5703
rect 597 5661 647 5703
rect 805 5661 855 5703
rect 1013 5661 1063 5703
rect 5440 5702 5490 5744
rect 5653 5702 5703 5744
rect 5861 5702 5911 5744
rect 6069 5702 6119 5744
rect 2932 5591 2982 5633
rect 3140 5591 3190 5633
rect 3348 5591 3398 5633
rect 3561 5591 3611 5633
rect 1322 5417 1372 5459
rect 1535 5417 1585 5459
rect 1743 5417 1793 5459
rect 1951 5417 2001 5459
rect 7988 5632 8038 5674
rect 8196 5632 8246 5674
rect 8404 5632 8454 5674
rect 8617 5632 8667 5674
rect 6378 5458 6428 5500
rect 6591 5458 6641 5500
rect 6799 5458 6849 5500
rect 7007 5458 7057 5500
rect 3870 5347 3920 5389
rect 4078 5347 4128 5389
rect 4286 5347 4336 5389
rect 4499 5347 4549 5389
rect 8926 5388 8976 5430
rect 9134 5388 9184 5430
rect 9342 5388 9392 5430
rect 9555 5388 9605 5430
rect 383 5107 433 5149
rect 596 5107 646 5149
rect 804 5107 854 5149
rect 1012 5107 1062 5149
rect 2823 5061 2873 5103
rect 3031 5061 3081 5103
rect 3239 5061 3289 5103
rect 3452 5061 3502 5103
rect 5439 5148 5489 5190
rect 5652 5148 5702 5190
rect 5860 5148 5910 5190
rect 6068 5148 6118 5190
rect 7879 5102 7929 5144
rect 8087 5102 8137 5144
rect 8295 5102 8345 5144
rect 8508 5102 8558 5144
rect 1431 4844 1481 4886
rect 1644 4844 1694 4886
rect 1852 4844 1902 4886
rect 2060 4844 2110 4886
rect 3871 4798 3921 4840
rect 4079 4798 4129 4840
rect 4287 4798 4337 4840
rect 4500 4798 4550 4840
rect 6487 4885 6537 4927
rect 6700 4885 6750 4927
rect 6908 4885 6958 4927
rect 7116 4885 7166 4927
rect 8927 4839 8977 4881
rect 9135 4839 9185 4881
rect 9343 4839 9393 4881
rect 9556 4839 9606 4881
rect 384 4558 434 4600
rect 597 4558 647 4600
rect 805 4558 855 4600
rect 1013 4558 1063 4600
rect 5440 4599 5490 4641
rect 5653 4599 5703 4641
rect 5861 4599 5911 4641
rect 6069 4599 6119 4641
rect 2932 4488 2982 4530
rect 3140 4488 3190 4530
rect 3348 4488 3398 4530
rect 3561 4488 3611 4530
rect 1322 4314 1372 4356
rect 1535 4314 1585 4356
rect 1743 4314 1793 4356
rect 1951 4314 2001 4356
rect 7988 4529 8038 4571
rect 8196 4529 8246 4571
rect 8404 4529 8454 4571
rect 8617 4529 8667 4571
rect 6378 4355 6428 4397
rect 6591 4355 6641 4397
rect 6799 4355 6849 4397
rect 7007 4355 7057 4397
rect 3870 4244 3920 4286
rect 4078 4244 4128 4286
rect 4286 4244 4336 4286
rect 4499 4244 4549 4286
rect 8926 4285 8976 4327
rect 9134 4285 9184 4327
rect 9342 4285 9392 4327
rect 9555 4285 9605 4327
rect 383 4004 433 4046
rect 596 4004 646 4046
rect 804 4004 854 4046
rect 1012 4004 1062 4046
rect 2792 3977 2842 4019
rect 3000 3977 3050 4019
rect 3208 3977 3258 4019
rect 3421 3977 3471 4019
rect 5439 4045 5489 4087
rect 5652 4045 5702 4087
rect 5860 4045 5910 4087
rect 6068 4045 6118 4087
rect 7848 4018 7898 4060
rect 8056 4018 8106 4060
rect 8264 4018 8314 4060
rect 8477 4018 8527 4060
rect 1463 3722 1513 3764
rect 1676 3722 1726 3764
rect 1884 3722 1934 3764
rect 2092 3722 2142 3764
rect 3872 3695 3922 3737
rect 4080 3695 4130 3737
rect 4288 3695 4338 3737
rect 4501 3695 4551 3737
rect 6519 3763 6569 3805
rect 6732 3763 6782 3805
rect 6940 3763 6990 3805
rect 7148 3763 7198 3805
rect 8928 3736 8978 3778
rect 9136 3736 9186 3778
rect 9344 3736 9394 3778
rect 9557 3736 9607 3778
rect 385 3455 435 3497
rect 598 3455 648 3497
rect 806 3455 856 3497
rect 1014 3455 1064 3497
rect 5441 3496 5491 3538
rect 5654 3496 5704 3538
rect 5862 3496 5912 3538
rect 6070 3496 6120 3538
rect 2933 3385 2983 3427
rect 3141 3385 3191 3427
rect 3349 3385 3399 3427
rect 3562 3385 3612 3427
rect 1323 3211 1373 3253
rect 1536 3211 1586 3253
rect 1744 3211 1794 3253
rect 1952 3211 2002 3253
rect 7989 3426 8039 3468
rect 8197 3426 8247 3468
rect 8405 3426 8455 3468
rect 8618 3426 8668 3468
rect 6379 3252 6429 3294
rect 6592 3252 6642 3294
rect 6800 3252 6850 3294
rect 7008 3252 7058 3294
rect 3871 3141 3921 3183
rect 4079 3141 4129 3183
rect 4287 3141 4337 3183
rect 4500 3141 4550 3183
rect 8927 3182 8977 3224
rect 9135 3182 9185 3224
rect 9343 3182 9393 3224
rect 9556 3182 9606 3224
rect 384 2901 434 2943
rect 597 2901 647 2943
rect 805 2901 855 2943
rect 1013 2901 1063 2943
rect 2823 2861 2873 2903
rect 3031 2861 3081 2903
rect 3239 2861 3289 2903
rect 3452 2861 3502 2903
rect 5440 2942 5490 2984
rect 5653 2942 5703 2984
rect 5861 2942 5911 2984
rect 6069 2942 6119 2984
rect 7879 2902 7929 2944
rect 8087 2902 8137 2944
rect 8295 2902 8345 2944
rect 8508 2902 8558 2944
rect 1433 2632 1483 2674
rect 1646 2632 1696 2674
rect 1854 2632 1904 2674
rect 2062 2632 2112 2674
rect 3872 2592 3922 2634
rect 4080 2592 4130 2634
rect 4288 2592 4338 2634
rect 4501 2592 4551 2634
rect 6489 2673 6539 2715
rect 6702 2673 6752 2715
rect 6910 2673 6960 2715
rect 7118 2673 7168 2715
rect 8928 2633 8978 2675
rect 9136 2633 9186 2675
rect 9344 2633 9394 2675
rect 9557 2633 9607 2675
rect 385 2352 435 2394
rect 598 2352 648 2394
rect 806 2352 856 2394
rect 1014 2352 1064 2394
rect 5441 2393 5491 2435
rect 5654 2393 5704 2435
rect 5862 2393 5912 2435
rect 6070 2393 6120 2435
rect 2933 2282 2983 2324
rect 3141 2282 3191 2324
rect 3349 2282 3399 2324
rect 3562 2282 3612 2324
rect 1323 2108 1373 2150
rect 1536 2108 1586 2150
rect 1744 2108 1794 2150
rect 1952 2108 2002 2150
rect 7989 2323 8039 2365
rect 8197 2323 8247 2365
rect 8405 2323 8455 2365
rect 8618 2323 8668 2365
rect 6379 2149 6429 2191
rect 6592 2149 6642 2191
rect 6800 2149 6850 2191
rect 7008 2149 7058 2191
rect 3871 2038 3921 2080
rect 4079 2038 4129 2080
rect 4287 2038 4337 2080
rect 4500 2038 4550 2080
rect 8927 2079 8977 2121
rect 9135 2079 9185 2121
rect 9343 2079 9393 2121
rect 9556 2079 9606 2121
rect 384 1798 434 1840
rect 597 1798 647 1840
rect 805 1798 855 1840
rect 1013 1798 1063 1840
rect 2793 1771 2843 1813
rect 3001 1771 3051 1813
rect 3209 1771 3259 1813
rect 3422 1771 3472 1813
rect 5440 1839 5490 1881
rect 5653 1839 5703 1881
rect 5861 1839 5911 1881
rect 6069 1839 6119 1881
rect 7849 1812 7899 1854
rect 8057 1812 8107 1854
rect 8265 1812 8315 1854
rect 8478 1812 8528 1854
rect 1464 1516 1514 1558
rect 1677 1516 1727 1558
rect 1885 1516 1935 1558
rect 2093 1516 2143 1558
rect 3873 1489 3923 1531
rect 4081 1489 4131 1531
rect 4289 1489 4339 1531
rect 4502 1489 4552 1531
rect 6520 1557 6570 1599
rect 6733 1557 6783 1599
rect 6941 1557 6991 1599
rect 7149 1557 7199 1599
rect 8929 1530 8979 1572
rect 9137 1530 9187 1572
rect 9345 1530 9395 1572
rect 9558 1530 9608 1572
rect 386 1249 436 1291
rect 599 1249 649 1291
rect 807 1249 857 1291
rect 1015 1249 1065 1291
rect 5442 1290 5492 1332
rect 5655 1290 5705 1332
rect 5863 1290 5913 1332
rect 6071 1290 6121 1332
rect 2934 1179 2984 1221
rect 3142 1179 3192 1221
rect 3350 1179 3400 1221
rect 3563 1179 3613 1221
rect 1324 1005 1374 1047
rect 1537 1005 1587 1047
rect 1745 1005 1795 1047
rect 1953 1005 2003 1047
rect 7990 1220 8040 1262
rect 8198 1220 8248 1262
rect 8406 1220 8456 1262
rect 8619 1220 8669 1262
rect 6380 1046 6430 1088
rect 6593 1046 6643 1088
rect 6801 1046 6851 1088
rect 7009 1046 7059 1088
rect 3872 935 3922 977
rect 4080 935 4130 977
rect 4288 935 4338 977
rect 4501 935 4551 977
rect 8928 976 8978 1018
rect 9136 976 9186 1018
rect 9344 976 9394 1018
rect 9557 976 9607 1018
rect 385 695 435 737
rect 598 695 648 737
rect 806 695 856 737
rect 1014 695 1064 737
rect 5441 736 5491 778
rect 5654 736 5704 778
rect 5862 736 5912 778
rect 6070 736 6120 778
rect 1632 136 1682 178
rect 1845 136 1895 178
rect 2053 136 2103 178
rect 2261 136 2311 178
rect 6688 177 6738 219
rect 6901 177 6951 219
rect 7109 177 7159 219
rect 7317 177 7367 219
rect 4582 116 4632 158
rect 4795 116 4845 158
rect 5003 116 5053 158
rect 5211 116 5261 158
<< pmos >>
rect 382 9089 432 9189
rect 595 9089 645 9189
rect 803 9089 853 9189
rect 1011 9089 1061 9189
rect 3869 9033 3919 9133
rect 4077 9033 4127 9133
rect 4285 9033 4335 9133
rect 4498 9033 4548 9133
rect 5438 9130 5488 9230
rect 5651 9130 5701 9230
rect 5859 9130 5909 9230
rect 6067 9130 6117 9230
rect 8925 9074 8975 9174
rect 9133 9074 9183 9174
rect 9341 9074 9391 9174
rect 9554 9074 9604 9174
rect 1320 8845 1370 8945
rect 1533 8845 1583 8945
rect 1741 8845 1791 8945
rect 1949 8845 1999 8945
rect 2930 8723 2980 8823
rect 3138 8723 3188 8823
rect 3346 8723 3396 8823
rect 3559 8723 3609 8823
rect 6376 8886 6426 8986
rect 6589 8886 6639 8986
rect 6797 8886 6847 8986
rect 7005 8886 7055 8986
rect 7986 8764 8036 8864
rect 8194 8764 8244 8864
rect 8402 8764 8452 8864
rect 8615 8764 8665 8864
rect 381 8535 431 8635
rect 594 8535 644 8635
rect 802 8535 852 8635
rect 1010 8535 1060 8635
rect 3868 8479 3918 8579
rect 4076 8479 4126 8579
rect 4284 8479 4334 8579
rect 4497 8479 4547 8579
rect 5437 8576 5487 8676
rect 5650 8576 5700 8676
rect 5858 8576 5908 8676
rect 6066 8576 6116 8676
rect 8924 8520 8974 8620
rect 9132 8520 9182 8620
rect 9340 8520 9390 8620
rect 9553 8520 9603 8620
rect 1461 8253 1511 8353
rect 1674 8253 1724 8353
rect 1882 8253 1932 8353
rect 2090 8253 2140 8353
rect 2790 8212 2840 8312
rect 2998 8212 3048 8312
rect 3206 8212 3256 8312
rect 3419 8212 3469 8312
rect 6517 8294 6567 8394
rect 6730 8294 6780 8394
rect 6938 8294 6988 8394
rect 7146 8294 7196 8394
rect 7846 8253 7896 8353
rect 8054 8253 8104 8353
rect 8262 8253 8312 8353
rect 8475 8253 8525 8353
rect 383 7986 433 8086
rect 596 7986 646 8086
rect 804 7986 854 8086
rect 1012 7986 1062 8086
rect 3870 7930 3920 8030
rect 4078 7930 4128 8030
rect 4286 7930 4336 8030
rect 4499 7930 4549 8030
rect 5439 8027 5489 8127
rect 5652 8027 5702 8127
rect 5860 8027 5910 8127
rect 6068 8027 6118 8127
rect 8926 7971 8976 8071
rect 9134 7971 9184 8071
rect 9342 7971 9392 8071
rect 9555 7971 9605 8071
rect 1321 7742 1371 7842
rect 1534 7742 1584 7842
rect 1742 7742 1792 7842
rect 1950 7742 2000 7842
rect 2931 7620 2981 7720
rect 3139 7620 3189 7720
rect 3347 7620 3397 7720
rect 3560 7620 3610 7720
rect 6377 7783 6427 7883
rect 6590 7783 6640 7883
rect 6798 7783 6848 7883
rect 7006 7783 7056 7883
rect 7987 7661 8037 7761
rect 8195 7661 8245 7761
rect 8403 7661 8453 7761
rect 8616 7661 8666 7761
rect 382 7432 432 7532
rect 595 7432 645 7532
rect 803 7432 853 7532
rect 1011 7432 1061 7532
rect 3869 7376 3919 7476
rect 4077 7376 4127 7476
rect 4285 7376 4335 7476
rect 4498 7376 4548 7476
rect 5438 7473 5488 7573
rect 5651 7473 5701 7573
rect 5859 7473 5909 7573
rect 6067 7473 6117 7573
rect 8925 7417 8975 7517
rect 9133 7417 9183 7517
rect 9341 7417 9391 7517
rect 9554 7417 9604 7517
rect 1431 7163 1481 7263
rect 1644 7163 1694 7263
rect 1852 7163 1902 7263
rect 2060 7163 2110 7263
rect 6487 7204 6537 7304
rect 6700 7204 6750 7304
rect 6908 7204 6958 7304
rect 7116 7204 7166 7304
rect 2821 7096 2871 7196
rect 3029 7096 3079 7196
rect 3237 7096 3287 7196
rect 3450 7096 3500 7196
rect 7877 7137 7927 7237
rect 8085 7137 8135 7237
rect 8293 7137 8343 7237
rect 8506 7137 8556 7237
rect 383 6883 433 6983
rect 596 6883 646 6983
rect 804 6883 854 6983
rect 1012 6883 1062 6983
rect 3870 6827 3920 6927
rect 4078 6827 4128 6927
rect 4286 6827 4336 6927
rect 4499 6827 4549 6927
rect 5439 6924 5489 7024
rect 5652 6924 5702 7024
rect 5860 6924 5910 7024
rect 6068 6924 6118 7024
rect 8926 6868 8976 6968
rect 9134 6868 9184 6968
rect 9342 6868 9392 6968
rect 9555 6868 9605 6968
rect 1321 6639 1371 6739
rect 1534 6639 1584 6739
rect 1742 6639 1792 6739
rect 1950 6639 2000 6739
rect 2931 6517 2981 6617
rect 3139 6517 3189 6617
rect 3347 6517 3397 6617
rect 3560 6517 3610 6617
rect 6377 6680 6427 6780
rect 6590 6680 6640 6780
rect 6798 6680 6848 6780
rect 7006 6680 7056 6780
rect 7987 6558 8037 6658
rect 8195 6558 8245 6658
rect 8403 6558 8453 6658
rect 8616 6558 8666 6658
rect 382 6329 432 6429
rect 595 6329 645 6429
rect 803 6329 853 6429
rect 1011 6329 1061 6429
rect 3869 6273 3919 6373
rect 4077 6273 4127 6373
rect 4285 6273 4335 6373
rect 4498 6273 4548 6373
rect 5438 6370 5488 6470
rect 5651 6370 5701 6470
rect 5859 6370 5909 6470
rect 6067 6370 6117 6470
rect 8925 6314 8975 6414
rect 9133 6314 9183 6414
rect 9341 6314 9391 6414
rect 9554 6314 9604 6414
rect 1462 6047 1512 6147
rect 1675 6047 1725 6147
rect 1883 6047 1933 6147
rect 2091 6047 2141 6147
rect 2791 6006 2841 6106
rect 2999 6006 3049 6106
rect 3207 6006 3257 6106
rect 3420 6006 3470 6106
rect 6518 6088 6568 6188
rect 6731 6088 6781 6188
rect 6939 6088 6989 6188
rect 7147 6088 7197 6188
rect 7847 6047 7897 6147
rect 8055 6047 8105 6147
rect 8263 6047 8313 6147
rect 8476 6047 8526 6147
rect 384 5780 434 5880
rect 597 5780 647 5880
rect 805 5780 855 5880
rect 1013 5780 1063 5880
rect 3871 5724 3921 5824
rect 4079 5724 4129 5824
rect 4287 5724 4337 5824
rect 4500 5724 4550 5824
rect 5440 5821 5490 5921
rect 5653 5821 5703 5921
rect 5861 5821 5911 5921
rect 6069 5821 6119 5921
rect 8927 5765 8977 5865
rect 9135 5765 9185 5865
rect 9343 5765 9393 5865
rect 9556 5765 9606 5865
rect 1322 5536 1372 5636
rect 1535 5536 1585 5636
rect 1743 5536 1793 5636
rect 1951 5536 2001 5636
rect 2932 5414 2982 5514
rect 3140 5414 3190 5514
rect 3348 5414 3398 5514
rect 3561 5414 3611 5514
rect 6378 5577 6428 5677
rect 6591 5577 6641 5677
rect 6799 5577 6849 5677
rect 7007 5577 7057 5677
rect 7988 5455 8038 5555
rect 8196 5455 8246 5555
rect 8404 5455 8454 5555
rect 8617 5455 8667 5555
rect 383 5226 433 5326
rect 596 5226 646 5326
rect 804 5226 854 5326
rect 1012 5226 1062 5326
rect 3870 5170 3920 5270
rect 4078 5170 4128 5270
rect 4286 5170 4336 5270
rect 4499 5170 4549 5270
rect 5439 5267 5489 5367
rect 5652 5267 5702 5367
rect 5860 5267 5910 5367
rect 6068 5267 6118 5367
rect 8926 5211 8976 5311
rect 9134 5211 9184 5311
rect 9342 5211 9392 5311
rect 9555 5211 9605 5311
rect 1431 4963 1481 5063
rect 1644 4963 1694 5063
rect 1852 4963 1902 5063
rect 2060 4963 2110 5063
rect 6487 5004 6537 5104
rect 6700 5004 6750 5104
rect 6908 5004 6958 5104
rect 7116 5004 7166 5104
rect 2823 4884 2873 4984
rect 3031 4884 3081 4984
rect 3239 4884 3289 4984
rect 3452 4884 3502 4984
rect 7879 4925 7929 5025
rect 8087 4925 8137 5025
rect 8295 4925 8345 5025
rect 8508 4925 8558 5025
rect 384 4677 434 4777
rect 597 4677 647 4777
rect 805 4677 855 4777
rect 1013 4677 1063 4777
rect 3871 4621 3921 4721
rect 4079 4621 4129 4721
rect 4287 4621 4337 4721
rect 4500 4621 4550 4721
rect 5440 4718 5490 4818
rect 5653 4718 5703 4818
rect 5861 4718 5911 4818
rect 6069 4718 6119 4818
rect 8927 4662 8977 4762
rect 9135 4662 9185 4762
rect 9343 4662 9393 4762
rect 9556 4662 9606 4762
rect 1322 4433 1372 4533
rect 1535 4433 1585 4533
rect 1743 4433 1793 4533
rect 1951 4433 2001 4533
rect 2932 4311 2982 4411
rect 3140 4311 3190 4411
rect 3348 4311 3398 4411
rect 3561 4311 3611 4411
rect 6378 4474 6428 4574
rect 6591 4474 6641 4574
rect 6799 4474 6849 4574
rect 7007 4474 7057 4574
rect 7988 4352 8038 4452
rect 8196 4352 8246 4452
rect 8404 4352 8454 4452
rect 8617 4352 8667 4452
rect 383 4123 433 4223
rect 596 4123 646 4223
rect 804 4123 854 4223
rect 1012 4123 1062 4223
rect 3870 4067 3920 4167
rect 4078 4067 4128 4167
rect 4286 4067 4336 4167
rect 4499 4067 4549 4167
rect 5439 4164 5489 4264
rect 5652 4164 5702 4264
rect 5860 4164 5910 4264
rect 6068 4164 6118 4264
rect 8926 4108 8976 4208
rect 9134 4108 9184 4208
rect 9342 4108 9392 4208
rect 9555 4108 9605 4208
rect 1463 3841 1513 3941
rect 1676 3841 1726 3941
rect 1884 3841 1934 3941
rect 2092 3841 2142 3941
rect 2792 3800 2842 3900
rect 3000 3800 3050 3900
rect 3208 3800 3258 3900
rect 3421 3800 3471 3900
rect 6519 3882 6569 3982
rect 6732 3882 6782 3982
rect 6940 3882 6990 3982
rect 7148 3882 7198 3982
rect 7848 3841 7898 3941
rect 8056 3841 8106 3941
rect 8264 3841 8314 3941
rect 8477 3841 8527 3941
rect 385 3574 435 3674
rect 598 3574 648 3674
rect 806 3574 856 3674
rect 1014 3574 1064 3674
rect 3872 3518 3922 3618
rect 4080 3518 4130 3618
rect 4288 3518 4338 3618
rect 4501 3518 4551 3618
rect 5441 3615 5491 3715
rect 5654 3615 5704 3715
rect 5862 3615 5912 3715
rect 6070 3615 6120 3715
rect 8928 3559 8978 3659
rect 9136 3559 9186 3659
rect 9344 3559 9394 3659
rect 9557 3559 9607 3659
rect 1323 3330 1373 3430
rect 1536 3330 1586 3430
rect 1744 3330 1794 3430
rect 1952 3330 2002 3430
rect 2933 3208 2983 3308
rect 3141 3208 3191 3308
rect 3349 3208 3399 3308
rect 3562 3208 3612 3308
rect 6379 3371 6429 3471
rect 6592 3371 6642 3471
rect 6800 3371 6850 3471
rect 7008 3371 7058 3471
rect 7989 3249 8039 3349
rect 8197 3249 8247 3349
rect 8405 3249 8455 3349
rect 8618 3249 8668 3349
rect 384 3020 434 3120
rect 597 3020 647 3120
rect 805 3020 855 3120
rect 1013 3020 1063 3120
rect 3871 2964 3921 3064
rect 4079 2964 4129 3064
rect 4287 2964 4337 3064
rect 4500 2964 4550 3064
rect 5440 3061 5490 3161
rect 5653 3061 5703 3161
rect 5861 3061 5911 3161
rect 6069 3061 6119 3161
rect 8927 3005 8977 3105
rect 9135 3005 9185 3105
rect 9343 3005 9393 3105
rect 9556 3005 9606 3105
rect 1433 2751 1483 2851
rect 1646 2751 1696 2851
rect 1854 2751 1904 2851
rect 2062 2751 2112 2851
rect 6489 2792 6539 2892
rect 6702 2792 6752 2892
rect 6910 2792 6960 2892
rect 7118 2792 7168 2892
rect 2823 2684 2873 2784
rect 3031 2684 3081 2784
rect 3239 2684 3289 2784
rect 3452 2684 3502 2784
rect 7879 2725 7929 2825
rect 8087 2725 8137 2825
rect 8295 2725 8345 2825
rect 8508 2725 8558 2825
rect 385 2471 435 2571
rect 598 2471 648 2571
rect 806 2471 856 2571
rect 1014 2471 1064 2571
rect 3872 2415 3922 2515
rect 4080 2415 4130 2515
rect 4288 2415 4338 2515
rect 4501 2415 4551 2515
rect 5441 2512 5491 2612
rect 5654 2512 5704 2612
rect 5862 2512 5912 2612
rect 6070 2512 6120 2612
rect 8928 2456 8978 2556
rect 9136 2456 9186 2556
rect 9344 2456 9394 2556
rect 9557 2456 9607 2556
rect 1323 2227 1373 2327
rect 1536 2227 1586 2327
rect 1744 2227 1794 2327
rect 1952 2227 2002 2327
rect 2933 2105 2983 2205
rect 3141 2105 3191 2205
rect 3349 2105 3399 2205
rect 3562 2105 3612 2205
rect 6379 2268 6429 2368
rect 6592 2268 6642 2368
rect 6800 2268 6850 2368
rect 7008 2268 7058 2368
rect 7989 2146 8039 2246
rect 8197 2146 8247 2246
rect 8405 2146 8455 2246
rect 8618 2146 8668 2246
rect 384 1917 434 2017
rect 597 1917 647 2017
rect 805 1917 855 2017
rect 1013 1917 1063 2017
rect 3871 1861 3921 1961
rect 4079 1861 4129 1961
rect 4287 1861 4337 1961
rect 4500 1861 4550 1961
rect 5440 1958 5490 2058
rect 5653 1958 5703 2058
rect 5861 1958 5911 2058
rect 6069 1958 6119 2058
rect 8927 1902 8977 2002
rect 9135 1902 9185 2002
rect 9343 1902 9393 2002
rect 9556 1902 9606 2002
rect 1464 1635 1514 1735
rect 1677 1635 1727 1735
rect 1885 1635 1935 1735
rect 2093 1635 2143 1735
rect 2793 1594 2843 1694
rect 3001 1594 3051 1694
rect 3209 1594 3259 1694
rect 3422 1594 3472 1694
rect 6520 1676 6570 1776
rect 6733 1676 6783 1776
rect 6941 1676 6991 1776
rect 7149 1676 7199 1776
rect 7849 1635 7899 1735
rect 8057 1635 8107 1735
rect 8265 1635 8315 1735
rect 8478 1635 8528 1735
rect 386 1368 436 1468
rect 599 1368 649 1468
rect 807 1368 857 1468
rect 1015 1368 1065 1468
rect 3873 1312 3923 1412
rect 4081 1312 4131 1412
rect 4289 1312 4339 1412
rect 4502 1312 4552 1412
rect 5442 1409 5492 1509
rect 5655 1409 5705 1509
rect 5863 1409 5913 1509
rect 6071 1409 6121 1509
rect 8929 1353 8979 1453
rect 9137 1353 9187 1453
rect 9345 1353 9395 1453
rect 9558 1353 9608 1453
rect 1324 1124 1374 1224
rect 1537 1124 1587 1224
rect 1745 1124 1795 1224
rect 1953 1124 2003 1224
rect 2934 1002 2984 1102
rect 3142 1002 3192 1102
rect 3350 1002 3400 1102
rect 3563 1002 3613 1102
rect 6380 1165 6430 1265
rect 6593 1165 6643 1265
rect 6801 1165 6851 1265
rect 7009 1165 7059 1265
rect 7990 1043 8040 1143
rect 8198 1043 8248 1143
rect 8406 1043 8456 1143
rect 8619 1043 8669 1143
rect 385 814 435 914
rect 598 814 648 914
rect 806 814 856 914
rect 1014 814 1064 914
rect 3872 758 3922 858
rect 4080 758 4130 858
rect 4288 758 4338 858
rect 4501 758 4551 858
rect 5441 855 5491 955
rect 5654 855 5704 955
rect 5862 855 5912 955
rect 6070 855 6120 955
rect 8928 799 8978 899
rect 9136 799 9186 899
rect 9344 799 9394 899
rect 9557 799 9607 899
rect 1632 255 1682 355
rect 1845 255 1895 355
rect 2053 255 2103 355
rect 2261 255 2311 355
rect 4582 235 4632 335
rect 4795 235 4845 335
rect 5003 235 5053 335
rect 5211 235 5261 335
rect 6688 296 6738 396
rect 6901 296 6951 396
rect 7109 296 7159 396
rect 7317 296 7367 396
<< ndiff >>
rect 3820 9240 3869 9252
rect 3820 9220 3831 9240
rect 3851 9220 3869 9240
rect 3820 9210 3869 9220
rect 3919 9236 3963 9252
rect 3919 9216 3934 9236
rect 3954 9216 3963 9236
rect 3919 9210 3963 9216
rect 4033 9236 4077 9252
rect 4033 9216 4042 9236
rect 4062 9216 4077 9236
rect 4033 9210 4077 9216
rect 4127 9240 4176 9252
rect 4127 9220 4145 9240
rect 4165 9220 4176 9240
rect 4127 9210 4176 9220
rect 4241 9236 4285 9252
rect 4241 9216 4250 9236
rect 4270 9216 4285 9236
rect 4241 9210 4285 9216
rect 4335 9240 4384 9252
rect 4335 9220 4353 9240
rect 4373 9220 4384 9240
rect 4335 9210 4384 9220
rect 4454 9236 4498 9252
rect 4454 9216 4463 9236
rect 4483 9216 4498 9236
rect 4454 9210 4498 9216
rect 4548 9240 4597 9252
rect 8876 9281 8925 9293
rect 8876 9261 8887 9281
rect 8907 9261 8925 9281
rect 8876 9251 8925 9261
rect 8975 9277 9019 9293
rect 8975 9257 8990 9277
rect 9010 9257 9019 9277
rect 8975 9251 9019 9257
rect 9089 9277 9133 9293
rect 9089 9257 9098 9277
rect 9118 9257 9133 9277
rect 9089 9251 9133 9257
rect 9183 9281 9232 9293
rect 9183 9261 9201 9281
rect 9221 9261 9232 9281
rect 9183 9251 9232 9261
rect 9297 9277 9341 9293
rect 9297 9257 9306 9277
rect 9326 9257 9341 9277
rect 9297 9251 9341 9257
rect 9391 9281 9440 9293
rect 9391 9261 9409 9281
rect 9429 9261 9440 9281
rect 9391 9251 9440 9261
rect 9510 9277 9554 9293
rect 9510 9257 9519 9277
rect 9539 9257 9554 9277
rect 9510 9251 9554 9257
rect 9604 9281 9653 9293
rect 9604 9261 9622 9281
rect 9642 9261 9653 9281
rect 9604 9251 9653 9261
rect 4548 9220 4566 9240
rect 4586 9220 4597 9240
rect 4548 9210 4597 9220
rect 333 9002 382 9012
rect 333 8982 344 9002
rect 364 8982 382 9002
rect 333 8970 382 8982
rect 432 9006 476 9012
rect 432 8986 447 9006
rect 467 8986 476 9006
rect 432 8970 476 8986
rect 546 9002 595 9012
rect 546 8982 557 9002
rect 577 8982 595 9002
rect 546 8970 595 8982
rect 645 9006 689 9012
rect 645 8986 660 9006
rect 680 8986 689 9006
rect 645 8970 689 8986
rect 754 9002 803 9012
rect 754 8982 765 9002
rect 785 8982 803 9002
rect 754 8970 803 8982
rect 853 9006 897 9012
rect 853 8986 868 9006
rect 888 8986 897 9006
rect 853 8970 897 8986
rect 967 9006 1011 9012
rect 967 8986 976 9006
rect 996 8986 1011 9006
rect 967 8970 1011 8986
rect 1061 9002 1110 9012
rect 1061 8982 1079 9002
rect 1099 8982 1110 9002
rect 1061 8970 1110 8982
rect 5389 9043 5438 9053
rect 5389 9023 5400 9043
rect 5420 9023 5438 9043
rect 5389 9011 5438 9023
rect 5488 9047 5532 9053
rect 5488 9027 5503 9047
rect 5523 9027 5532 9047
rect 5488 9011 5532 9027
rect 5602 9043 5651 9053
rect 5602 9023 5613 9043
rect 5633 9023 5651 9043
rect 5602 9011 5651 9023
rect 5701 9047 5745 9053
rect 5701 9027 5716 9047
rect 5736 9027 5745 9047
rect 5701 9011 5745 9027
rect 5810 9043 5859 9053
rect 5810 9023 5821 9043
rect 5841 9023 5859 9043
rect 5810 9011 5859 9023
rect 5909 9047 5953 9053
rect 5909 9027 5924 9047
rect 5944 9027 5953 9047
rect 5909 9011 5953 9027
rect 6023 9047 6067 9053
rect 6023 9027 6032 9047
rect 6052 9027 6067 9047
rect 6023 9011 6067 9027
rect 6117 9043 6166 9053
rect 6117 9023 6135 9043
rect 6155 9023 6166 9043
rect 6117 9011 6166 9023
rect 2881 8930 2930 8942
rect 2881 8910 2892 8930
rect 2912 8910 2930 8930
rect 2881 8900 2930 8910
rect 2980 8926 3024 8942
rect 2980 8906 2995 8926
rect 3015 8906 3024 8926
rect 2980 8900 3024 8906
rect 3094 8926 3138 8942
rect 3094 8906 3103 8926
rect 3123 8906 3138 8926
rect 3094 8900 3138 8906
rect 3188 8930 3237 8942
rect 3188 8910 3206 8930
rect 3226 8910 3237 8930
rect 3188 8900 3237 8910
rect 3302 8926 3346 8942
rect 3302 8906 3311 8926
rect 3331 8906 3346 8926
rect 3302 8900 3346 8906
rect 3396 8930 3445 8942
rect 3396 8910 3414 8930
rect 3434 8910 3445 8930
rect 3396 8900 3445 8910
rect 3515 8926 3559 8942
rect 3515 8906 3524 8926
rect 3544 8906 3559 8926
rect 3515 8900 3559 8906
rect 3609 8930 3658 8942
rect 3609 8910 3627 8930
rect 3647 8910 3658 8930
rect 3609 8900 3658 8910
rect 1271 8758 1320 8768
rect 1271 8738 1282 8758
rect 1302 8738 1320 8758
rect 1271 8726 1320 8738
rect 1370 8762 1414 8768
rect 1370 8742 1385 8762
rect 1405 8742 1414 8762
rect 1370 8726 1414 8742
rect 1484 8758 1533 8768
rect 1484 8738 1495 8758
rect 1515 8738 1533 8758
rect 1484 8726 1533 8738
rect 1583 8762 1627 8768
rect 1583 8742 1598 8762
rect 1618 8742 1627 8762
rect 1583 8726 1627 8742
rect 1692 8758 1741 8768
rect 1692 8738 1703 8758
rect 1723 8738 1741 8758
rect 1692 8726 1741 8738
rect 1791 8762 1835 8768
rect 1791 8742 1806 8762
rect 1826 8742 1835 8762
rect 1791 8726 1835 8742
rect 1905 8762 1949 8768
rect 1905 8742 1914 8762
rect 1934 8742 1949 8762
rect 1905 8726 1949 8742
rect 1999 8758 2048 8768
rect 1999 8738 2017 8758
rect 2037 8738 2048 8758
rect 1999 8726 2048 8738
rect 7937 8971 7986 8983
rect 7937 8951 7948 8971
rect 7968 8951 7986 8971
rect 7937 8941 7986 8951
rect 8036 8967 8080 8983
rect 8036 8947 8051 8967
rect 8071 8947 8080 8967
rect 8036 8941 8080 8947
rect 8150 8967 8194 8983
rect 8150 8947 8159 8967
rect 8179 8947 8194 8967
rect 8150 8941 8194 8947
rect 8244 8971 8293 8983
rect 8244 8951 8262 8971
rect 8282 8951 8293 8971
rect 8244 8941 8293 8951
rect 8358 8967 8402 8983
rect 8358 8947 8367 8967
rect 8387 8947 8402 8967
rect 8358 8941 8402 8947
rect 8452 8971 8501 8983
rect 8452 8951 8470 8971
rect 8490 8951 8501 8971
rect 8452 8941 8501 8951
rect 8571 8967 8615 8983
rect 8571 8947 8580 8967
rect 8600 8947 8615 8967
rect 8571 8941 8615 8947
rect 8665 8971 8714 8983
rect 8665 8951 8683 8971
rect 8703 8951 8714 8971
rect 8665 8941 8714 8951
rect 6327 8799 6376 8809
rect 6327 8779 6338 8799
rect 6358 8779 6376 8799
rect 6327 8767 6376 8779
rect 6426 8803 6470 8809
rect 6426 8783 6441 8803
rect 6461 8783 6470 8803
rect 6426 8767 6470 8783
rect 6540 8799 6589 8809
rect 6540 8779 6551 8799
rect 6571 8779 6589 8799
rect 6540 8767 6589 8779
rect 6639 8803 6683 8809
rect 6639 8783 6654 8803
rect 6674 8783 6683 8803
rect 6639 8767 6683 8783
rect 6748 8799 6797 8809
rect 6748 8779 6759 8799
rect 6779 8779 6797 8799
rect 6748 8767 6797 8779
rect 6847 8803 6891 8809
rect 6847 8783 6862 8803
rect 6882 8783 6891 8803
rect 6847 8767 6891 8783
rect 6961 8803 7005 8809
rect 6961 8783 6970 8803
rect 6990 8783 7005 8803
rect 6961 8767 7005 8783
rect 7055 8799 7104 8809
rect 7055 8779 7073 8799
rect 7093 8779 7104 8799
rect 7055 8767 7104 8779
rect 3819 8686 3868 8698
rect 3819 8666 3830 8686
rect 3850 8666 3868 8686
rect 3819 8656 3868 8666
rect 3918 8682 3962 8698
rect 3918 8662 3933 8682
rect 3953 8662 3962 8682
rect 3918 8656 3962 8662
rect 4032 8682 4076 8698
rect 4032 8662 4041 8682
rect 4061 8662 4076 8682
rect 4032 8656 4076 8662
rect 4126 8686 4175 8698
rect 4126 8666 4144 8686
rect 4164 8666 4175 8686
rect 4126 8656 4175 8666
rect 4240 8682 4284 8698
rect 4240 8662 4249 8682
rect 4269 8662 4284 8682
rect 4240 8656 4284 8662
rect 4334 8686 4383 8698
rect 4334 8666 4352 8686
rect 4372 8666 4383 8686
rect 4334 8656 4383 8666
rect 4453 8682 4497 8698
rect 4453 8662 4462 8682
rect 4482 8662 4497 8682
rect 4453 8656 4497 8662
rect 4547 8686 4596 8698
rect 4547 8666 4565 8686
rect 4585 8666 4596 8686
rect 4547 8656 4596 8666
rect 8875 8727 8924 8739
rect 8875 8707 8886 8727
rect 8906 8707 8924 8727
rect 8875 8697 8924 8707
rect 8974 8723 9018 8739
rect 8974 8703 8989 8723
rect 9009 8703 9018 8723
rect 8974 8697 9018 8703
rect 9088 8723 9132 8739
rect 9088 8703 9097 8723
rect 9117 8703 9132 8723
rect 9088 8697 9132 8703
rect 9182 8727 9231 8739
rect 9182 8707 9200 8727
rect 9220 8707 9231 8727
rect 9182 8697 9231 8707
rect 9296 8723 9340 8739
rect 9296 8703 9305 8723
rect 9325 8703 9340 8723
rect 9296 8697 9340 8703
rect 9390 8727 9439 8739
rect 9390 8707 9408 8727
rect 9428 8707 9439 8727
rect 9390 8697 9439 8707
rect 9509 8723 9553 8739
rect 9509 8703 9518 8723
rect 9538 8703 9553 8723
rect 9509 8697 9553 8703
rect 9603 8727 9652 8739
rect 9603 8707 9621 8727
rect 9641 8707 9652 8727
rect 9603 8697 9652 8707
rect 5388 8489 5437 8499
rect 5388 8469 5399 8489
rect 5419 8469 5437 8489
rect 332 8448 381 8458
rect 332 8428 343 8448
rect 363 8428 381 8448
rect 332 8416 381 8428
rect 431 8452 475 8458
rect 431 8432 446 8452
rect 466 8432 475 8452
rect 431 8416 475 8432
rect 545 8448 594 8458
rect 545 8428 556 8448
rect 576 8428 594 8448
rect 545 8416 594 8428
rect 644 8452 688 8458
rect 644 8432 659 8452
rect 679 8432 688 8452
rect 644 8416 688 8432
rect 753 8448 802 8458
rect 753 8428 764 8448
rect 784 8428 802 8448
rect 753 8416 802 8428
rect 852 8452 896 8458
rect 852 8432 867 8452
rect 887 8432 896 8452
rect 852 8416 896 8432
rect 966 8452 1010 8458
rect 966 8432 975 8452
rect 995 8432 1010 8452
rect 966 8416 1010 8432
rect 1060 8448 1109 8458
rect 1060 8428 1078 8448
rect 1098 8428 1109 8448
rect 1060 8416 1109 8428
rect 2741 8419 2790 8431
rect 2741 8399 2752 8419
rect 2772 8399 2790 8419
rect 2741 8389 2790 8399
rect 2840 8415 2884 8431
rect 2840 8395 2855 8415
rect 2875 8395 2884 8415
rect 2840 8389 2884 8395
rect 2954 8415 2998 8431
rect 2954 8395 2963 8415
rect 2983 8395 2998 8415
rect 2954 8389 2998 8395
rect 3048 8419 3097 8431
rect 3048 8399 3066 8419
rect 3086 8399 3097 8419
rect 3048 8389 3097 8399
rect 3162 8415 3206 8431
rect 3162 8395 3171 8415
rect 3191 8395 3206 8415
rect 3162 8389 3206 8395
rect 3256 8419 3305 8431
rect 3256 8399 3274 8419
rect 3294 8399 3305 8419
rect 3256 8389 3305 8399
rect 3375 8415 3419 8431
rect 3375 8395 3384 8415
rect 3404 8395 3419 8415
rect 3375 8389 3419 8395
rect 3469 8419 3518 8431
rect 3469 8399 3487 8419
rect 3507 8399 3518 8419
rect 3469 8389 3518 8399
rect 5388 8457 5437 8469
rect 5487 8493 5531 8499
rect 5487 8473 5502 8493
rect 5522 8473 5531 8493
rect 5487 8457 5531 8473
rect 5601 8489 5650 8499
rect 5601 8469 5612 8489
rect 5632 8469 5650 8489
rect 5601 8457 5650 8469
rect 5700 8493 5744 8499
rect 5700 8473 5715 8493
rect 5735 8473 5744 8493
rect 5700 8457 5744 8473
rect 5809 8489 5858 8499
rect 5809 8469 5820 8489
rect 5840 8469 5858 8489
rect 5809 8457 5858 8469
rect 5908 8493 5952 8499
rect 5908 8473 5923 8493
rect 5943 8473 5952 8493
rect 5908 8457 5952 8473
rect 6022 8493 6066 8499
rect 6022 8473 6031 8493
rect 6051 8473 6066 8493
rect 6022 8457 6066 8473
rect 6116 8489 6165 8499
rect 6116 8469 6134 8489
rect 6154 8469 6165 8489
rect 6116 8457 6165 8469
rect 7797 8460 7846 8472
rect 7797 8440 7808 8460
rect 7828 8440 7846 8460
rect 7797 8430 7846 8440
rect 7896 8456 7940 8472
rect 7896 8436 7911 8456
rect 7931 8436 7940 8456
rect 7896 8430 7940 8436
rect 8010 8456 8054 8472
rect 8010 8436 8019 8456
rect 8039 8436 8054 8456
rect 8010 8430 8054 8436
rect 8104 8460 8153 8472
rect 8104 8440 8122 8460
rect 8142 8440 8153 8460
rect 8104 8430 8153 8440
rect 8218 8456 8262 8472
rect 8218 8436 8227 8456
rect 8247 8436 8262 8456
rect 8218 8430 8262 8436
rect 8312 8460 8361 8472
rect 8312 8440 8330 8460
rect 8350 8440 8361 8460
rect 8312 8430 8361 8440
rect 8431 8456 8475 8472
rect 8431 8436 8440 8456
rect 8460 8436 8475 8456
rect 8431 8430 8475 8436
rect 8525 8460 8574 8472
rect 8525 8440 8543 8460
rect 8563 8440 8574 8460
rect 8525 8430 8574 8440
rect 1412 8166 1461 8176
rect 1412 8146 1423 8166
rect 1443 8146 1461 8166
rect 1412 8134 1461 8146
rect 1511 8170 1555 8176
rect 1511 8150 1526 8170
rect 1546 8150 1555 8170
rect 1511 8134 1555 8150
rect 1625 8166 1674 8176
rect 1625 8146 1636 8166
rect 1656 8146 1674 8166
rect 1625 8134 1674 8146
rect 1724 8170 1768 8176
rect 1724 8150 1739 8170
rect 1759 8150 1768 8170
rect 1724 8134 1768 8150
rect 1833 8166 1882 8176
rect 1833 8146 1844 8166
rect 1864 8146 1882 8166
rect 1833 8134 1882 8146
rect 1932 8170 1976 8176
rect 1932 8150 1947 8170
rect 1967 8150 1976 8170
rect 1932 8134 1976 8150
rect 2046 8170 2090 8176
rect 2046 8150 2055 8170
rect 2075 8150 2090 8170
rect 2046 8134 2090 8150
rect 2140 8166 2189 8176
rect 2140 8146 2158 8166
rect 2178 8146 2189 8166
rect 2140 8134 2189 8146
rect 3821 8137 3870 8149
rect 3821 8117 3832 8137
rect 3852 8117 3870 8137
rect 3821 8107 3870 8117
rect 3920 8133 3964 8149
rect 3920 8113 3935 8133
rect 3955 8113 3964 8133
rect 3920 8107 3964 8113
rect 4034 8133 4078 8149
rect 4034 8113 4043 8133
rect 4063 8113 4078 8133
rect 4034 8107 4078 8113
rect 4128 8137 4177 8149
rect 4128 8117 4146 8137
rect 4166 8117 4177 8137
rect 4128 8107 4177 8117
rect 4242 8133 4286 8149
rect 4242 8113 4251 8133
rect 4271 8113 4286 8133
rect 4242 8107 4286 8113
rect 4336 8137 4385 8149
rect 4336 8117 4354 8137
rect 4374 8117 4385 8137
rect 4336 8107 4385 8117
rect 4455 8133 4499 8149
rect 4455 8113 4464 8133
rect 4484 8113 4499 8133
rect 4455 8107 4499 8113
rect 4549 8137 4598 8149
rect 6468 8207 6517 8217
rect 6468 8187 6479 8207
rect 6499 8187 6517 8207
rect 6468 8175 6517 8187
rect 6567 8211 6611 8217
rect 6567 8191 6582 8211
rect 6602 8191 6611 8211
rect 6567 8175 6611 8191
rect 6681 8207 6730 8217
rect 6681 8187 6692 8207
rect 6712 8187 6730 8207
rect 6681 8175 6730 8187
rect 6780 8211 6824 8217
rect 6780 8191 6795 8211
rect 6815 8191 6824 8211
rect 6780 8175 6824 8191
rect 6889 8207 6938 8217
rect 6889 8187 6900 8207
rect 6920 8187 6938 8207
rect 6889 8175 6938 8187
rect 6988 8211 7032 8217
rect 6988 8191 7003 8211
rect 7023 8191 7032 8211
rect 6988 8175 7032 8191
rect 7102 8211 7146 8217
rect 7102 8191 7111 8211
rect 7131 8191 7146 8211
rect 7102 8175 7146 8191
rect 7196 8207 7245 8217
rect 7196 8187 7214 8207
rect 7234 8187 7245 8207
rect 7196 8175 7245 8187
rect 8877 8178 8926 8190
rect 8877 8158 8888 8178
rect 8908 8158 8926 8178
rect 8877 8148 8926 8158
rect 8976 8174 9020 8190
rect 8976 8154 8991 8174
rect 9011 8154 9020 8174
rect 8976 8148 9020 8154
rect 9090 8174 9134 8190
rect 9090 8154 9099 8174
rect 9119 8154 9134 8174
rect 9090 8148 9134 8154
rect 9184 8178 9233 8190
rect 9184 8158 9202 8178
rect 9222 8158 9233 8178
rect 9184 8148 9233 8158
rect 9298 8174 9342 8190
rect 9298 8154 9307 8174
rect 9327 8154 9342 8174
rect 9298 8148 9342 8154
rect 9392 8178 9441 8190
rect 9392 8158 9410 8178
rect 9430 8158 9441 8178
rect 9392 8148 9441 8158
rect 9511 8174 9555 8190
rect 9511 8154 9520 8174
rect 9540 8154 9555 8174
rect 9511 8148 9555 8154
rect 9605 8178 9654 8190
rect 9605 8158 9623 8178
rect 9643 8158 9654 8178
rect 9605 8148 9654 8158
rect 4549 8117 4567 8137
rect 4587 8117 4598 8137
rect 4549 8107 4598 8117
rect 334 7899 383 7909
rect 334 7879 345 7899
rect 365 7879 383 7899
rect 334 7867 383 7879
rect 433 7903 477 7909
rect 433 7883 448 7903
rect 468 7883 477 7903
rect 433 7867 477 7883
rect 547 7899 596 7909
rect 547 7879 558 7899
rect 578 7879 596 7899
rect 547 7867 596 7879
rect 646 7903 690 7909
rect 646 7883 661 7903
rect 681 7883 690 7903
rect 646 7867 690 7883
rect 755 7899 804 7909
rect 755 7879 766 7899
rect 786 7879 804 7899
rect 755 7867 804 7879
rect 854 7903 898 7909
rect 854 7883 869 7903
rect 889 7883 898 7903
rect 854 7867 898 7883
rect 968 7903 1012 7909
rect 968 7883 977 7903
rect 997 7883 1012 7903
rect 968 7867 1012 7883
rect 1062 7899 1111 7909
rect 1062 7879 1080 7899
rect 1100 7879 1111 7899
rect 1062 7867 1111 7879
rect 5390 7940 5439 7950
rect 5390 7920 5401 7940
rect 5421 7920 5439 7940
rect 5390 7908 5439 7920
rect 5489 7944 5533 7950
rect 5489 7924 5504 7944
rect 5524 7924 5533 7944
rect 5489 7908 5533 7924
rect 5603 7940 5652 7950
rect 5603 7920 5614 7940
rect 5634 7920 5652 7940
rect 5603 7908 5652 7920
rect 5702 7944 5746 7950
rect 5702 7924 5717 7944
rect 5737 7924 5746 7944
rect 5702 7908 5746 7924
rect 5811 7940 5860 7950
rect 5811 7920 5822 7940
rect 5842 7920 5860 7940
rect 5811 7908 5860 7920
rect 5910 7944 5954 7950
rect 5910 7924 5925 7944
rect 5945 7924 5954 7944
rect 5910 7908 5954 7924
rect 6024 7944 6068 7950
rect 6024 7924 6033 7944
rect 6053 7924 6068 7944
rect 6024 7908 6068 7924
rect 6118 7940 6167 7950
rect 6118 7920 6136 7940
rect 6156 7920 6167 7940
rect 6118 7908 6167 7920
rect 2882 7827 2931 7839
rect 2882 7807 2893 7827
rect 2913 7807 2931 7827
rect 2882 7797 2931 7807
rect 2981 7823 3025 7839
rect 2981 7803 2996 7823
rect 3016 7803 3025 7823
rect 2981 7797 3025 7803
rect 3095 7823 3139 7839
rect 3095 7803 3104 7823
rect 3124 7803 3139 7823
rect 3095 7797 3139 7803
rect 3189 7827 3238 7839
rect 3189 7807 3207 7827
rect 3227 7807 3238 7827
rect 3189 7797 3238 7807
rect 3303 7823 3347 7839
rect 3303 7803 3312 7823
rect 3332 7803 3347 7823
rect 3303 7797 3347 7803
rect 3397 7827 3446 7839
rect 3397 7807 3415 7827
rect 3435 7807 3446 7827
rect 3397 7797 3446 7807
rect 3516 7823 3560 7839
rect 3516 7803 3525 7823
rect 3545 7803 3560 7823
rect 3516 7797 3560 7803
rect 3610 7827 3659 7839
rect 3610 7807 3628 7827
rect 3648 7807 3659 7827
rect 3610 7797 3659 7807
rect 1272 7655 1321 7665
rect 1272 7635 1283 7655
rect 1303 7635 1321 7655
rect 1272 7623 1321 7635
rect 1371 7659 1415 7665
rect 1371 7639 1386 7659
rect 1406 7639 1415 7659
rect 1371 7623 1415 7639
rect 1485 7655 1534 7665
rect 1485 7635 1496 7655
rect 1516 7635 1534 7655
rect 1485 7623 1534 7635
rect 1584 7659 1628 7665
rect 1584 7639 1599 7659
rect 1619 7639 1628 7659
rect 1584 7623 1628 7639
rect 1693 7655 1742 7665
rect 1693 7635 1704 7655
rect 1724 7635 1742 7655
rect 1693 7623 1742 7635
rect 1792 7659 1836 7665
rect 1792 7639 1807 7659
rect 1827 7639 1836 7659
rect 1792 7623 1836 7639
rect 1906 7659 1950 7665
rect 1906 7639 1915 7659
rect 1935 7639 1950 7659
rect 1906 7623 1950 7639
rect 2000 7655 2049 7665
rect 2000 7635 2018 7655
rect 2038 7635 2049 7655
rect 2000 7623 2049 7635
rect 7938 7868 7987 7880
rect 7938 7848 7949 7868
rect 7969 7848 7987 7868
rect 7938 7838 7987 7848
rect 8037 7864 8081 7880
rect 8037 7844 8052 7864
rect 8072 7844 8081 7864
rect 8037 7838 8081 7844
rect 8151 7864 8195 7880
rect 8151 7844 8160 7864
rect 8180 7844 8195 7864
rect 8151 7838 8195 7844
rect 8245 7868 8294 7880
rect 8245 7848 8263 7868
rect 8283 7848 8294 7868
rect 8245 7838 8294 7848
rect 8359 7864 8403 7880
rect 8359 7844 8368 7864
rect 8388 7844 8403 7864
rect 8359 7838 8403 7844
rect 8453 7868 8502 7880
rect 8453 7848 8471 7868
rect 8491 7848 8502 7868
rect 8453 7838 8502 7848
rect 8572 7864 8616 7880
rect 8572 7844 8581 7864
rect 8601 7844 8616 7864
rect 8572 7838 8616 7844
rect 8666 7868 8715 7880
rect 8666 7848 8684 7868
rect 8704 7848 8715 7868
rect 8666 7838 8715 7848
rect 6328 7696 6377 7706
rect 6328 7676 6339 7696
rect 6359 7676 6377 7696
rect 6328 7664 6377 7676
rect 6427 7700 6471 7706
rect 6427 7680 6442 7700
rect 6462 7680 6471 7700
rect 6427 7664 6471 7680
rect 6541 7696 6590 7706
rect 6541 7676 6552 7696
rect 6572 7676 6590 7696
rect 6541 7664 6590 7676
rect 6640 7700 6684 7706
rect 6640 7680 6655 7700
rect 6675 7680 6684 7700
rect 6640 7664 6684 7680
rect 6749 7696 6798 7706
rect 6749 7676 6760 7696
rect 6780 7676 6798 7696
rect 6749 7664 6798 7676
rect 6848 7700 6892 7706
rect 6848 7680 6863 7700
rect 6883 7680 6892 7700
rect 6848 7664 6892 7680
rect 6962 7700 7006 7706
rect 6962 7680 6971 7700
rect 6991 7680 7006 7700
rect 6962 7664 7006 7680
rect 7056 7696 7105 7706
rect 7056 7676 7074 7696
rect 7094 7676 7105 7696
rect 7056 7664 7105 7676
rect 3820 7583 3869 7595
rect 3820 7563 3831 7583
rect 3851 7563 3869 7583
rect 3820 7553 3869 7563
rect 3919 7579 3963 7595
rect 3919 7559 3934 7579
rect 3954 7559 3963 7579
rect 3919 7553 3963 7559
rect 4033 7579 4077 7595
rect 4033 7559 4042 7579
rect 4062 7559 4077 7579
rect 4033 7553 4077 7559
rect 4127 7583 4176 7595
rect 4127 7563 4145 7583
rect 4165 7563 4176 7583
rect 4127 7553 4176 7563
rect 4241 7579 4285 7595
rect 4241 7559 4250 7579
rect 4270 7559 4285 7579
rect 4241 7553 4285 7559
rect 4335 7583 4384 7595
rect 4335 7563 4353 7583
rect 4373 7563 4384 7583
rect 4335 7553 4384 7563
rect 4454 7579 4498 7595
rect 4454 7559 4463 7579
rect 4483 7559 4498 7579
rect 4454 7553 4498 7559
rect 4548 7583 4597 7595
rect 4548 7563 4566 7583
rect 4586 7563 4597 7583
rect 4548 7553 4597 7563
rect 8876 7624 8925 7636
rect 8876 7604 8887 7624
rect 8907 7604 8925 7624
rect 8876 7594 8925 7604
rect 8975 7620 9019 7636
rect 8975 7600 8990 7620
rect 9010 7600 9019 7620
rect 8975 7594 9019 7600
rect 9089 7620 9133 7636
rect 9089 7600 9098 7620
rect 9118 7600 9133 7620
rect 9089 7594 9133 7600
rect 9183 7624 9232 7636
rect 9183 7604 9201 7624
rect 9221 7604 9232 7624
rect 9183 7594 9232 7604
rect 9297 7620 9341 7636
rect 9297 7600 9306 7620
rect 9326 7600 9341 7620
rect 9297 7594 9341 7600
rect 9391 7624 9440 7636
rect 9391 7604 9409 7624
rect 9429 7604 9440 7624
rect 9391 7594 9440 7604
rect 9510 7620 9554 7636
rect 9510 7600 9519 7620
rect 9539 7600 9554 7620
rect 9510 7594 9554 7600
rect 9604 7624 9653 7636
rect 9604 7604 9622 7624
rect 9642 7604 9653 7624
rect 9604 7594 9653 7604
rect 5389 7386 5438 7396
rect 5389 7366 5400 7386
rect 5420 7366 5438 7386
rect 333 7345 382 7355
rect 333 7325 344 7345
rect 364 7325 382 7345
rect 333 7313 382 7325
rect 432 7349 476 7355
rect 432 7329 447 7349
rect 467 7329 476 7349
rect 432 7313 476 7329
rect 546 7345 595 7355
rect 546 7325 557 7345
rect 577 7325 595 7345
rect 546 7313 595 7325
rect 645 7349 689 7355
rect 645 7329 660 7349
rect 680 7329 689 7349
rect 645 7313 689 7329
rect 754 7345 803 7355
rect 754 7325 765 7345
rect 785 7325 803 7345
rect 754 7313 803 7325
rect 853 7349 897 7355
rect 853 7329 868 7349
rect 888 7329 897 7349
rect 853 7313 897 7329
rect 967 7349 1011 7355
rect 967 7329 976 7349
rect 996 7329 1011 7349
rect 967 7313 1011 7329
rect 1061 7345 1110 7355
rect 1061 7325 1079 7345
rect 1099 7325 1110 7345
rect 1061 7313 1110 7325
rect 2772 7303 2821 7315
rect 2772 7283 2783 7303
rect 2803 7283 2821 7303
rect 2772 7273 2821 7283
rect 2871 7299 2915 7315
rect 2871 7279 2886 7299
rect 2906 7279 2915 7299
rect 2871 7273 2915 7279
rect 2985 7299 3029 7315
rect 2985 7279 2994 7299
rect 3014 7279 3029 7299
rect 2985 7273 3029 7279
rect 3079 7303 3128 7315
rect 3079 7283 3097 7303
rect 3117 7283 3128 7303
rect 3079 7273 3128 7283
rect 3193 7299 3237 7315
rect 3193 7279 3202 7299
rect 3222 7279 3237 7299
rect 3193 7273 3237 7279
rect 3287 7303 3336 7315
rect 3287 7283 3305 7303
rect 3325 7283 3336 7303
rect 3287 7273 3336 7283
rect 3406 7299 3450 7315
rect 3406 7279 3415 7299
rect 3435 7279 3450 7299
rect 3406 7273 3450 7279
rect 3500 7303 3549 7315
rect 3500 7283 3518 7303
rect 3538 7283 3549 7303
rect 5389 7354 5438 7366
rect 5488 7390 5532 7396
rect 5488 7370 5503 7390
rect 5523 7370 5532 7390
rect 5488 7354 5532 7370
rect 5602 7386 5651 7396
rect 5602 7366 5613 7386
rect 5633 7366 5651 7386
rect 5602 7354 5651 7366
rect 5701 7390 5745 7396
rect 5701 7370 5716 7390
rect 5736 7370 5745 7390
rect 5701 7354 5745 7370
rect 5810 7386 5859 7396
rect 5810 7366 5821 7386
rect 5841 7366 5859 7386
rect 5810 7354 5859 7366
rect 5909 7390 5953 7396
rect 5909 7370 5924 7390
rect 5944 7370 5953 7390
rect 5909 7354 5953 7370
rect 6023 7390 6067 7396
rect 6023 7370 6032 7390
rect 6052 7370 6067 7390
rect 6023 7354 6067 7370
rect 6117 7386 6166 7396
rect 6117 7366 6135 7386
rect 6155 7366 6166 7386
rect 6117 7354 6166 7366
rect 7828 7344 7877 7356
rect 7828 7324 7839 7344
rect 7859 7324 7877 7344
rect 3500 7273 3549 7283
rect 7828 7314 7877 7324
rect 7927 7340 7971 7356
rect 7927 7320 7942 7340
rect 7962 7320 7971 7340
rect 7927 7314 7971 7320
rect 8041 7340 8085 7356
rect 8041 7320 8050 7340
rect 8070 7320 8085 7340
rect 8041 7314 8085 7320
rect 8135 7344 8184 7356
rect 8135 7324 8153 7344
rect 8173 7324 8184 7344
rect 8135 7314 8184 7324
rect 8249 7340 8293 7356
rect 8249 7320 8258 7340
rect 8278 7320 8293 7340
rect 8249 7314 8293 7320
rect 8343 7344 8392 7356
rect 8343 7324 8361 7344
rect 8381 7324 8392 7344
rect 8343 7314 8392 7324
rect 8462 7340 8506 7356
rect 8462 7320 8471 7340
rect 8491 7320 8506 7340
rect 8462 7314 8506 7320
rect 8556 7344 8605 7356
rect 8556 7324 8574 7344
rect 8594 7324 8605 7344
rect 8556 7314 8605 7324
rect 1382 7076 1431 7086
rect 1382 7056 1393 7076
rect 1413 7056 1431 7076
rect 1382 7044 1431 7056
rect 1481 7080 1525 7086
rect 1481 7060 1496 7080
rect 1516 7060 1525 7080
rect 1481 7044 1525 7060
rect 1595 7076 1644 7086
rect 1595 7056 1606 7076
rect 1626 7056 1644 7076
rect 1595 7044 1644 7056
rect 1694 7080 1738 7086
rect 1694 7060 1709 7080
rect 1729 7060 1738 7080
rect 1694 7044 1738 7060
rect 1803 7076 1852 7086
rect 1803 7056 1814 7076
rect 1834 7056 1852 7076
rect 1803 7044 1852 7056
rect 1902 7080 1946 7086
rect 1902 7060 1917 7080
rect 1937 7060 1946 7080
rect 1902 7044 1946 7060
rect 2016 7080 2060 7086
rect 2016 7060 2025 7080
rect 2045 7060 2060 7080
rect 2016 7044 2060 7060
rect 2110 7076 2159 7086
rect 6438 7117 6487 7127
rect 2110 7056 2128 7076
rect 2148 7056 2159 7076
rect 2110 7044 2159 7056
rect 3821 7034 3870 7046
rect 3821 7014 3832 7034
rect 3852 7014 3870 7034
rect 3821 7004 3870 7014
rect 3920 7030 3964 7046
rect 3920 7010 3935 7030
rect 3955 7010 3964 7030
rect 3920 7004 3964 7010
rect 4034 7030 4078 7046
rect 4034 7010 4043 7030
rect 4063 7010 4078 7030
rect 4034 7004 4078 7010
rect 4128 7034 4177 7046
rect 4128 7014 4146 7034
rect 4166 7014 4177 7034
rect 4128 7004 4177 7014
rect 4242 7030 4286 7046
rect 4242 7010 4251 7030
rect 4271 7010 4286 7030
rect 4242 7004 4286 7010
rect 4336 7034 4385 7046
rect 4336 7014 4354 7034
rect 4374 7014 4385 7034
rect 4336 7004 4385 7014
rect 4455 7030 4499 7046
rect 4455 7010 4464 7030
rect 4484 7010 4499 7030
rect 4455 7004 4499 7010
rect 4549 7034 4598 7046
rect 6438 7097 6449 7117
rect 6469 7097 6487 7117
rect 6438 7085 6487 7097
rect 6537 7121 6581 7127
rect 6537 7101 6552 7121
rect 6572 7101 6581 7121
rect 6537 7085 6581 7101
rect 6651 7117 6700 7127
rect 6651 7097 6662 7117
rect 6682 7097 6700 7117
rect 6651 7085 6700 7097
rect 6750 7121 6794 7127
rect 6750 7101 6765 7121
rect 6785 7101 6794 7121
rect 6750 7085 6794 7101
rect 6859 7117 6908 7127
rect 6859 7097 6870 7117
rect 6890 7097 6908 7117
rect 6859 7085 6908 7097
rect 6958 7121 7002 7127
rect 6958 7101 6973 7121
rect 6993 7101 7002 7121
rect 6958 7085 7002 7101
rect 7072 7121 7116 7127
rect 7072 7101 7081 7121
rect 7101 7101 7116 7121
rect 7072 7085 7116 7101
rect 7166 7117 7215 7127
rect 7166 7097 7184 7117
rect 7204 7097 7215 7117
rect 7166 7085 7215 7097
rect 8877 7075 8926 7087
rect 8877 7055 8888 7075
rect 8908 7055 8926 7075
rect 8877 7045 8926 7055
rect 8976 7071 9020 7087
rect 8976 7051 8991 7071
rect 9011 7051 9020 7071
rect 8976 7045 9020 7051
rect 9090 7071 9134 7087
rect 9090 7051 9099 7071
rect 9119 7051 9134 7071
rect 9090 7045 9134 7051
rect 9184 7075 9233 7087
rect 9184 7055 9202 7075
rect 9222 7055 9233 7075
rect 9184 7045 9233 7055
rect 9298 7071 9342 7087
rect 9298 7051 9307 7071
rect 9327 7051 9342 7071
rect 9298 7045 9342 7051
rect 9392 7075 9441 7087
rect 9392 7055 9410 7075
rect 9430 7055 9441 7075
rect 9392 7045 9441 7055
rect 9511 7071 9555 7087
rect 9511 7051 9520 7071
rect 9540 7051 9555 7071
rect 9511 7045 9555 7051
rect 9605 7075 9654 7087
rect 9605 7055 9623 7075
rect 9643 7055 9654 7075
rect 9605 7045 9654 7055
rect 4549 7014 4567 7034
rect 4587 7014 4598 7034
rect 4549 7004 4598 7014
rect 334 6796 383 6806
rect 334 6776 345 6796
rect 365 6776 383 6796
rect 334 6764 383 6776
rect 433 6800 477 6806
rect 433 6780 448 6800
rect 468 6780 477 6800
rect 433 6764 477 6780
rect 547 6796 596 6806
rect 547 6776 558 6796
rect 578 6776 596 6796
rect 547 6764 596 6776
rect 646 6800 690 6806
rect 646 6780 661 6800
rect 681 6780 690 6800
rect 646 6764 690 6780
rect 755 6796 804 6806
rect 755 6776 766 6796
rect 786 6776 804 6796
rect 755 6764 804 6776
rect 854 6800 898 6806
rect 854 6780 869 6800
rect 889 6780 898 6800
rect 854 6764 898 6780
rect 968 6800 1012 6806
rect 968 6780 977 6800
rect 997 6780 1012 6800
rect 968 6764 1012 6780
rect 1062 6796 1111 6806
rect 1062 6776 1080 6796
rect 1100 6776 1111 6796
rect 1062 6764 1111 6776
rect 5390 6837 5439 6847
rect 5390 6817 5401 6837
rect 5421 6817 5439 6837
rect 5390 6805 5439 6817
rect 5489 6841 5533 6847
rect 5489 6821 5504 6841
rect 5524 6821 5533 6841
rect 5489 6805 5533 6821
rect 5603 6837 5652 6847
rect 5603 6817 5614 6837
rect 5634 6817 5652 6837
rect 5603 6805 5652 6817
rect 5702 6841 5746 6847
rect 5702 6821 5717 6841
rect 5737 6821 5746 6841
rect 5702 6805 5746 6821
rect 5811 6837 5860 6847
rect 5811 6817 5822 6837
rect 5842 6817 5860 6837
rect 5811 6805 5860 6817
rect 5910 6841 5954 6847
rect 5910 6821 5925 6841
rect 5945 6821 5954 6841
rect 5910 6805 5954 6821
rect 6024 6841 6068 6847
rect 6024 6821 6033 6841
rect 6053 6821 6068 6841
rect 6024 6805 6068 6821
rect 6118 6837 6167 6847
rect 6118 6817 6136 6837
rect 6156 6817 6167 6837
rect 6118 6805 6167 6817
rect 2882 6724 2931 6736
rect 2882 6704 2893 6724
rect 2913 6704 2931 6724
rect 2882 6694 2931 6704
rect 2981 6720 3025 6736
rect 2981 6700 2996 6720
rect 3016 6700 3025 6720
rect 2981 6694 3025 6700
rect 3095 6720 3139 6736
rect 3095 6700 3104 6720
rect 3124 6700 3139 6720
rect 3095 6694 3139 6700
rect 3189 6724 3238 6736
rect 3189 6704 3207 6724
rect 3227 6704 3238 6724
rect 3189 6694 3238 6704
rect 3303 6720 3347 6736
rect 3303 6700 3312 6720
rect 3332 6700 3347 6720
rect 3303 6694 3347 6700
rect 3397 6724 3446 6736
rect 3397 6704 3415 6724
rect 3435 6704 3446 6724
rect 3397 6694 3446 6704
rect 3516 6720 3560 6736
rect 3516 6700 3525 6720
rect 3545 6700 3560 6720
rect 3516 6694 3560 6700
rect 3610 6724 3659 6736
rect 3610 6704 3628 6724
rect 3648 6704 3659 6724
rect 3610 6694 3659 6704
rect 1272 6552 1321 6562
rect 1272 6532 1283 6552
rect 1303 6532 1321 6552
rect 1272 6520 1321 6532
rect 1371 6556 1415 6562
rect 1371 6536 1386 6556
rect 1406 6536 1415 6556
rect 1371 6520 1415 6536
rect 1485 6552 1534 6562
rect 1485 6532 1496 6552
rect 1516 6532 1534 6552
rect 1485 6520 1534 6532
rect 1584 6556 1628 6562
rect 1584 6536 1599 6556
rect 1619 6536 1628 6556
rect 1584 6520 1628 6536
rect 1693 6552 1742 6562
rect 1693 6532 1704 6552
rect 1724 6532 1742 6552
rect 1693 6520 1742 6532
rect 1792 6556 1836 6562
rect 1792 6536 1807 6556
rect 1827 6536 1836 6556
rect 1792 6520 1836 6536
rect 1906 6556 1950 6562
rect 1906 6536 1915 6556
rect 1935 6536 1950 6556
rect 1906 6520 1950 6536
rect 2000 6552 2049 6562
rect 2000 6532 2018 6552
rect 2038 6532 2049 6552
rect 2000 6520 2049 6532
rect 7938 6765 7987 6777
rect 7938 6745 7949 6765
rect 7969 6745 7987 6765
rect 7938 6735 7987 6745
rect 8037 6761 8081 6777
rect 8037 6741 8052 6761
rect 8072 6741 8081 6761
rect 8037 6735 8081 6741
rect 8151 6761 8195 6777
rect 8151 6741 8160 6761
rect 8180 6741 8195 6761
rect 8151 6735 8195 6741
rect 8245 6765 8294 6777
rect 8245 6745 8263 6765
rect 8283 6745 8294 6765
rect 8245 6735 8294 6745
rect 8359 6761 8403 6777
rect 8359 6741 8368 6761
rect 8388 6741 8403 6761
rect 8359 6735 8403 6741
rect 8453 6765 8502 6777
rect 8453 6745 8471 6765
rect 8491 6745 8502 6765
rect 8453 6735 8502 6745
rect 8572 6761 8616 6777
rect 8572 6741 8581 6761
rect 8601 6741 8616 6761
rect 8572 6735 8616 6741
rect 8666 6765 8715 6777
rect 8666 6745 8684 6765
rect 8704 6745 8715 6765
rect 8666 6735 8715 6745
rect 6328 6593 6377 6603
rect 6328 6573 6339 6593
rect 6359 6573 6377 6593
rect 6328 6561 6377 6573
rect 6427 6597 6471 6603
rect 6427 6577 6442 6597
rect 6462 6577 6471 6597
rect 6427 6561 6471 6577
rect 6541 6593 6590 6603
rect 6541 6573 6552 6593
rect 6572 6573 6590 6593
rect 6541 6561 6590 6573
rect 6640 6597 6684 6603
rect 6640 6577 6655 6597
rect 6675 6577 6684 6597
rect 6640 6561 6684 6577
rect 6749 6593 6798 6603
rect 6749 6573 6760 6593
rect 6780 6573 6798 6593
rect 6749 6561 6798 6573
rect 6848 6597 6892 6603
rect 6848 6577 6863 6597
rect 6883 6577 6892 6597
rect 6848 6561 6892 6577
rect 6962 6597 7006 6603
rect 6962 6577 6971 6597
rect 6991 6577 7006 6597
rect 6962 6561 7006 6577
rect 7056 6593 7105 6603
rect 7056 6573 7074 6593
rect 7094 6573 7105 6593
rect 7056 6561 7105 6573
rect 3820 6480 3869 6492
rect 3820 6460 3831 6480
rect 3851 6460 3869 6480
rect 3820 6450 3869 6460
rect 3919 6476 3963 6492
rect 3919 6456 3934 6476
rect 3954 6456 3963 6476
rect 3919 6450 3963 6456
rect 4033 6476 4077 6492
rect 4033 6456 4042 6476
rect 4062 6456 4077 6476
rect 4033 6450 4077 6456
rect 4127 6480 4176 6492
rect 4127 6460 4145 6480
rect 4165 6460 4176 6480
rect 4127 6450 4176 6460
rect 4241 6476 4285 6492
rect 4241 6456 4250 6476
rect 4270 6456 4285 6476
rect 4241 6450 4285 6456
rect 4335 6480 4384 6492
rect 4335 6460 4353 6480
rect 4373 6460 4384 6480
rect 4335 6450 4384 6460
rect 4454 6476 4498 6492
rect 4454 6456 4463 6476
rect 4483 6456 4498 6476
rect 4454 6450 4498 6456
rect 4548 6480 4597 6492
rect 4548 6460 4566 6480
rect 4586 6460 4597 6480
rect 4548 6450 4597 6460
rect 8876 6521 8925 6533
rect 8876 6501 8887 6521
rect 8907 6501 8925 6521
rect 8876 6491 8925 6501
rect 8975 6517 9019 6533
rect 8975 6497 8990 6517
rect 9010 6497 9019 6517
rect 8975 6491 9019 6497
rect 9089 6517 9133 6533
rect 9089 6497 9098 6517
rect 9118 6497 9133 6517
rect 9089 6491 9133 6497
rect 9183 6521 9232 6533
rect 9183 6501 9201 6521
rect 9221 6501 9232 6521
rect 9183 6491 9232 6501
rect 9297 6517 9341 6533
rect 9297 6497 9306 6517
rect 9326 6497 9341 6517
rect 9297 6491 9341 6497
rect 9391 6521 9440 6533
rect 9391 6501 9409 6521
rect 9429 6501 9440 6521
rect 9391 6491 9440 6501
rect 9510 6517 9554 6533
rect 9510 6497 9519 6517
rect 9539 6497 9554 6517
rect 9510 6491 9554 6497
rect 9604 6521 9653 6533
rect 9604 6501 9622 6521
rect 9642 6501 9653 6521
rect 9604 6491 9653 6501
rect 5389 6283 5438 6293
rect 5389 6263 5400 6283
rect 5420 6263 5438 6283
rect 333 6242 382 6252
rect 333 6222 344 6242
rect 364 6222 382 6242
rect 333 6210 382 6222
rect 432 6246 476 6252
rect 432 6226 447 6246
rect 467 6226 476 6246
rect 432 6210 476 6226
rect 546 6242 595 6252
rect 546 6222 557 6242
rect 577 6222 595 6242
rect 546 6210 595 6222
rect 645 6246 689 6252
rect 645 6226 660 6246
rect 680 6226 689 6246
rect 645 6210 689 6226
rect 754 6242 803 6252
rect 754 6222 765 6242
rect 785 6222 803 6242
rect 754 6210 803 6222
rect 853 6246 897 6252
rect 853 6226 868 6246
rect 888 6226 897 6246
rect 853 6210 897 6226
rect 967 6246 1011 6252
rect 967 6226 976 6246
rect 996 6226 1011 6246
rect 967 6210 1011 6226
rect 1061 6242 1110 6252
rect 1061 6222 1079 6242
rect 1099 6222 1110 6242
rect 1061 6210 1110 6222
rect 2742 6213 2791 6225
rect 2742 6193 2753 6213
rect 2773 6193 2791 6213
rect 2742 6183 2791 6193
rect 2841 6209 2885 6225
rect 2841 6189 2856 6209
rect 2876 6189 2885 6209
rect 2841 6183 2885 6189
rect 2955 6209 2999 6225
rect 2955 6189 2964 6209
rect 2984 6189 2999 6209
rect 2955 6183 2999 6189
rect 3049 6213 3098 6225
rect 3049 6193 3067 6213
rect 3087 6193 3098 6213
rect 3049 6183 3098 6193
rect 3163 6209 3207 6225
rect 3163 6189 3172 6209
rect 3192 6189 3207 6209
rect 3163 6183 3207 6189
rect 3257 6213 3306 6225
rect 3257 6193 3275 6213
rect 3295 6193 3306 6213
rect 3257 6183 3306 6193
rect 3376 6209 3420 6225
rect 3376 6189 3385 6209
rect 3405 6189 3420 6209
rect 3376 6183 3420 6189
rect 3470 6213 3519 6225
rect 3470 6193 3488 6213
rect 3508 6193 3519 6213
rect 3470 6183 3519 6193
rect 5389 6251 5438 6263
rect 5488 6287 5532 6293
rect 5488 6267 5503 6287
rect 5523 6267 5532 6287
rect 5488 6251 5532 6267
rect 5602 6283 5651 6293
rect 5602 6263 5613 6283
rect 5633 6263 5651 6283
rect 5602 6251 5651 6263
rect 5701 6287 5745 6293
rect 5701 6267 5716 6287
rect 5736 6267 5745 6287
rect 5701 6251 5745 6267
rect 5810 6283 5859 6293
rect 5810 6263 5821 6283
rect 5841 6263 5859 6283
rect 5810 6251 5859 6263
rect 5909 6287 5953 6293
rect 5909 6267 5924 6287
rect 5944 6267 5953 6287
rect 5909 6251 5953 6267
rect 6023 6287 6067 6293
rect 6023 6267 6032 6287
rect 6052 6267 6067 6287
rect 6023 6251 6067 6267
rect 6117 6283 6166 6293
rect 6117 6263 6135 6283
rect 6155 6263 6166 6283
rect 6117 6251 6166 6263
rect 7798 6254 7847 6266
rect 7798 6234 7809 6254
rect 7829 6234 7847 6254
rect 7798 6224 7847 6234
rect 7897 6250 7941 6266
rect 7897 6230 7912 6250
rect 7932 6230 7941 6250
rect 7897 6224 7941 6230
rect 8011 6250 8055 6266
rect 8011 6230 8020 6250
rect 8040 6230 8055 6250
rect 8011 6224 8055 6230
rect 8105 6254 8154 6266
rect 8105 6234 8123 6254
rect 8143 6234 8154 6254
rect 8105 6224 8154 6234
rect 8219 6250 8263 6266
rect 8219 6230 8228 6250
rect 8248 6230 8263 6250
rect 8219 6224 8263 6230
rect 8313 6254 8362 6266
rect 8313 6234 8331 6254
rect 8351 6234 8362 6254
rect 8313 6224 8362 6234
rect 8432 6250 8476 6266
rect 8432 6230 8441 6250
rect 8461 6230 8476 6250
rect 8432 6224 8476 6230
rect 8526 6254 8575 6266
rect 8526 6234 8544 6254
rect 8564 6234 8575 6254
rect 8526 6224 8575 6234
rect 1413 5960 1462 5970
rect 1413 5940 1424 5960
rect 1444 5940 1462 5960
rect 1413 5928 1462 5940
rect 1512 5964 1556 5970
rect 1512 5944 1527 5964
rect 1547 5944 1556 5964
rect 1512 5928 1556 5944
rect 1626 5960 1675 5970
rect 1626 5940 1637 5960
rect 1657 5940 1675 5960
rect 1626 5928 1675 5940
rect 1725 5964 1769 5970
rect 1725 5944 1740 5964
rect 1760 5944 1769 5964
rect 1725 5928 1769 5944
rect 1834 5960 1883 5970
rect 1834 5940 1845 5960
rect 1865 5940 1883 5960
rect 1834 5928 1883 5940
rect 1933 5964 1977 5970
rect 1933 5944 1948 5964
rect 1968 5944 1977 5964
rect 1933 5928 1977 5944
rect 2047 5964 2091 5970
rect 2047 5944 2056 5964
rect 2076 5944 2091 5964
rect 2047 5928 2091 5944
rect 2141 5960 2190 5970
rect 2141 5940 2159 5960
rect 2179 5940 2190 5960
rect 2141 5928 2190 5940
rect 3822 5931 3871 5943
rect 3822 5911 3833 5931
rect 3853 5911 3871 5931
rect 3822 5901 3871 5911
rect 3921 5927 3965 5943
rect 3921 5907 3936 5927
rect 3956 5907 3965 5927
rect 3921 5901 3965 5907
rect 4035 5927 4079 5943
rect 4035 5907 4044 5927
rect 4064 5907 4079 5927
rect 4035 5901 4079 5907
rect 4129 5931 4178 5943
rect 4129 5911 4147 5931
rect 4167 5911 4178 5931
rect 4129 5901 4178 5911
rect 4243 5927 4287 5943
rect 4243 5907 4252 5927
rect 4272 5907 4287 5927
rect 4243 5901 4287 5907
rect 4337 5931 4386 5943
rect 4337 5911 4355 5931
rect 4375 5911 4386 5931
rect 4337 5901 4386 5911
rect 4456 5927 4500 5943
rect 4456 5907 4465 5927
rect 4485 5907 4500 5927
rect 4456 5901 4500 5907
rect 4550 5931 4599 5943
rect 6469 6001 6518 6011
rect 6469 5981 6480 6001
rect 6500 5981 6518 6001
rect 6469 5969 6518 5981
rect 6568 6005 6612 6011
rect 6568 5985 6583 6005
rect 6603 5985 6612 6005
rect 6568 5969 6612 5985
rect 6682 6001 6731 6011
rect 6682 5981 6693 6001
rect 6713 5981 6731 6001
rect 6682 5969 6731 5981
rect 6781 6005 6825 6011
rect 6781 5985 6796 6005
rect 6816 5985 6825 6005
rect 6781 5969 6825 5985
rect 6890 6001 6939 6011
rect 6890 5981 6901 6001
rect 6921 5981 6939 6001
rect 6890 5969 6939 5981
rect 6989 6005 7033 6011
rect 6989 5985 7004 6005
rect 7024 5985 7033 6005
rect 6989 5969 7033 5985
rect 7103 6005 7147 6011
rect 7103 5985 7112 6005
rect 7132 5985 7147 6005
rect 7103 5969 7147 5985
rect 7197 6001 7246 6011
rect 7197 5981 7215 6001
rect 7235 5981 7246 6001
rect 7197 5969 7246 5981
rect 8878 5972 8927 5984
rect 8878 5952 8889 5972
rect 8909 5952 8927 5972
rect 8878 5942 8927 5952
rect 8977 5968 9021 5984
rect 8977 5948 8992 5968
rect 9012 5948 9021 5968
rect 8977 5942 9021 5948
rect 9091 5968 9135 5984
rect 9091 5948 9100 5968
rect 9120 5948 9135 5968
rect 9091 5942 9135 5948
rect 9185 5972 9234 5984
rect 9185 5952 9203 5972
rect 9223 5952 9234 5972
rect 9185 5942 9234 5952
rect 9299 5968 9343 5984
rect 9299 5948 9308 5968
rect 9328 5948 9343 5968
rect 9299 5942 9343 5948
rect 9393 5972 9442 5984
rect 9393 5952 9411 5972
rect 9431 5952 9442 5972
rect 9393 5942 9442 5952
rect 9512 5968 9556 5984
rect 9512 5948 9521 5968
rect 9541 5948 9556 5968
rect 9512 5942 9556 5948
rect 9606 5972 9655 5984
rect 9606 5952 9624 5972
rect 9644 5952 9655 5972
rect 9606 5942 9655 5952
rect 4550 5911 4568 5931
rect 4588 5911 4599 5931
rect 4550 5901 4599 5911
rect 335 5693 384 5703
rect 335 5673 346 5693
rect 366 5673 384 5693
rect 335 5661 384 5673
rect 434 5697 478 5703
rect 434 5677 449 5697
rect 469 5677 478 5697
rect 434 5661 478 5677
rect 548 5693 597 5703
rect 548 5673 559 5693
rect 579 5673 597 5693
rect 548 5661 597 5673
rect 647 5697 691 5703
rect 647 5677 662 5697
rect 682 5677 691 5697
rect 647 5661 691 5677
rect 756 5693 805 5703
rect 756 5673 767 5693
rect 787 5673 805 5693
rect 756 5661 805 5673
rect 855 5697 899 5703
rect 855 5677 870 5697
rect 890 5677 899 5697
rect 855 5661 899 5677
rect 969 5697 1013 5703
rect 969 5677 978 5697
rect 998 5677 1013 5697
rect 969 5661 1013 5677
rect 1063 5693 1112 5703
rect 1063 5673 1081 5693
rect 1101 5673 1112 5693
rect 1063 5661 1112 5673
rect 5391 5734 5440 5744
rect 5391 5714 5402 5734
rect 5422 5714 5440 5734
rect 5391 5702 5440 5714
rect 5490 5738 5534 5744
rect 5490 5718 5505 5738
rect 5525 5718 5534 5738
rect 5490 5702 5534 5718
rect 5604 5734 5653 5744
rect 5604 5714 5615 5734
rect 5635 5714 5653 5734
rect 5604 5702 5653 5714
rect 5703 5738 5747 5744
rect 5703 5718 5718 5738
rect 5738 5718 5747 5738
rect 5703 5702 5747 5718
rect 5812 5734 5861 5744
rect 5812 5714 5823 5734
rect 5843 5714 5861 5734
rect 5812 5702 5861 5714
rect 5911 5738 5955 5744
rect 5911 5718 5926 5738
rect 5946 5718 5955 5738
rect 5911 5702 5955 5718
rect 6025 5738 6069 5744
rect 6025 5718 6034 5738
rect 6054 5718 6069 5738
rect 6025 5702 6069 5718
rect 6119 5734 6168 5744
rect 6119 5714 6137 5734
rect 6157 5714 6168 5734
rect 6119 5702 6168 5714
rect 2883 5621 2932 5633
rect 2883 5601 2894 5621
rect 2914 5601 2932 5621
rect 2883 5591 2932 5601
rect 2982 5617 3026 5633
rect 2982 5597 2997 5617
rect 3017 5597 3026 5617
rect 2982 5591 3026 5597
rect 3096 5617 3140 5633
rect 3096 5597 3105 5617
rect 3125 5597 3140 5617
rect 3096 5591 3140 5597
rect 3190 5621 3239 5633
rect 3190 5601 3208 5621
rect 3228 5601 3239 5621
rect 3190 5591 3239 5601
rect 3304 5617 3348 5633
rect 3304 5597 3313 5617
rect 3333 5597 3348 5617
rect 3304 5591 3348 5597
rect 3398 5621 3447 5633
rect 3398 5601 3416 5621
rect 3436 5601 3447 5621
rect 3398 5591 3447 5601
rect 3517 5617 3561 5633
rect 3517 5597 3526 5617
rect 3546 5597 3561 5617
rect 3517 5591 3561 5597
rect 3611 5621 3660 5633
rect 3611 5601 3629 5621
rect 3649 5601 3660 5621
rect 3611 5591 3660 5601
rect 1273 5449 1322 5459
rect 1273 5429 1284 5449
rect 1304 5429 1322 5449
rect 1273 5417 1322 5429
rect 1372 5453 1416 5459
rect 1372 5433 1387 5453
rect 1407 5433 1416 5453
rect 1372 5417 1416 5433
rect 1486 5449 1535 5459
rect 1486 5429 1497 5449
rect 1517 5429 1535 5449
rect 1486 5417 1535 5429
rect 1585 5453 1629 5459
rect 1585 5433 1600 5453
rect 1620 5433 1629 5453
rect 1585 5417 1629 5433
rect 1694 5449 1743 5459
rect 1694 5429 1705 5449
rect 1725 5429 1743 5449
rect 1694 5417 1743 5429
rect 1793 5453 1837 5459
rect 1793 5433 1808 5453
rect 1828 5433 1837 5453
rect 1793 5417 1837 5433
rect 1907 5453 1951 5459
rect 1907 5433 1916 5453
rect 1936 5433 1951 5453
rect 1907 5417 1951 5433
rect 2001 5449 2050 5459
rect 2001 5429 2019 5449
rect 2039 5429 2050 5449
rect 2001 5417 2050 5429
rect 7939 5662 7988 5674
rect 7939 5642 7950 5662
rect 7970 5642 7988 5662
rect 7939 5632 7988 5642
rect 8038 5658 8082 5674
rect 8038 5638 8053 5658
rect 8073 5638 8082 5658
rect 8038 5632 8082 5638
rect 8152 5658 8196 5674
rect 8152 5638 8161 5658
rect 8181 5638 8196 5658
rect 8152 5632 8196 5638
rect 8246 5662 8295 5674
rect 8246 5642 8264 5662
rect 8284 5642 8295 5662
rect 8246 5632 8295 5642
rect 8360 5658 8404 5674
rect 8360 5638 8369 5658
rect 8389 5638 8404 5658
rect 8360 5632 8404 5638
rect 8454 5662 8503 5674
rect 8454 5642 8472 5662
rect 8492 5642 8503 5662
rect 8454 5632 8503 5642
rect 8573 5658 8617 5674
rect 8573 5638 8582 5658
rect 8602 5638 8617 5658
rect 8573 5632 8617 5638
rect 8667 5662 8716 5674
rect 8667 5642 8685 5662
rect 8705 5642 8716 5662
rect 8667 5632 8716 5642
rect 6329 5490 6378 5500
rect 6329 5470 6340 5490
rect 6360 5470 6378 5490
rect 6329 5458 6378 5470
rect 6428 5494 6472 5500
rect 6428 5474 6443 5494
rect 6463 5474 6472 5494
rect 6428 5458 6472 5474
rect 6542 5490 6591 5500
rect 6542 5470 6553 5490
rect 6573 5470 6591 5490
rect 6542 5458 6591 5470
rect 6641 5494 6685 5500
rect 6641 5474 6656 5494
rect 6676 5474 6685 5494
rect 6641 5458 6685 5474
rect 6750 5490 6799 5500
rect 6750 5470 6761 5490
rect 6781 5470 6799 5490
rect 6750 5458 6799 5470
rect 6849 5494 6893 5500
rect 6849 5474 6864 5494
rect 6884 5474 6893 5494
rect 6849 5458 6893 5474
rect 6963 5494 7007 5500
rect 6963 5474 6972 5494
rect 6992 5474 7007 5494
rect 6963 5458 7007 5474
rect 7057 5490 7106 5500
rect 7057 5470 7075 5490
rect 7095 5470 7106 5490
rect 7057 5458 7106 5470
rect 3821 5377 3870 5389
rect 3821 5357 3832 5377
rect 3852 5357 3870 5377
rect 3821 5347 3870 5357
rect 3920 5373 3964 5389
rect 3920 5353 3935 5373
rect 3955 5353 3964 5373
rect 3920 5347 3964 5353
rect 4034 5373 4078 5389
rect 4034 5353 4043 5373
rect 4063 5353 4078 5373
rect 4034 5347 4078 5353
rect 4128 5377 4177 5389
rect 4128 5357 4146 5377
rect 4166 5357 4177 5377
rect 4128 5347 4177 5357
rect 4242 5373 4286 5389
rect 4242 5353 4251 5373
rect 4271 5353 4286 5373
rect 4242 5347 4286 5353
rect 4336 5377 4385 5389
rect 4336 5357 4354 5377
rect 4374 5357 4385 5377
rect 4336 5347 4385 5357
rect 4455 5373 4499 5389
rect 4455 5353 4464 5373
rect 4484 5353 4499 5373
rect 4455 5347 4499 5353
rect 4549 5377 4598 5389
rect 4549 5357 4567 5377
rect 4587 5357 4598 5377
rect 4549 5347 4598 5357
rect 8877 5418 8926 5430
rect 8877 5398 8888 5418
rect 8908 5398 8926 5418
rect 8877 5388 8926 5398
rect 8976 5414 9020 5430
rect 8976 5394 8991 5414
rect 9011 5394 9020 5414
rect 8976 5388 9020 5394
rect 9090 5414 9134 5430
rect 9090 5394 9099 5414
rect 9119 5394 9134 5414
rect 9090 5388 9134 5394
rect 9184 5418 9233 5430
rect 9184 5398 9202 5418
rect 9222 5398 9233 5418
rect 9184 5388 9233 5398
rect 9298 5414 9342 5430
rect 9298 5394 9307 5414
rect 9327 5394 9342 5414
rect 9298 5388 9342 5394
rect 9392 5418 9441 5430
rect 9392 5398 9410 5418
rect 9430 5398 9441 5418
rect 9392 5388 9441 5398
rect 9511 5414 9555 5430
rect 9511 5394 9520 5414
rect 9540 5394 9555 5414
rect 9511 5388 9555 5394
rect 9605 5418 9654 5430
rect 9605 5398 9623 5418
rect 9643 5398 9654 5418
rect 9605 5388 9654 5398
rect 334 5139 383 5149
rect 334 5119 345 5139
rect 365 5119 383 5139
rect 334 5107 383 5119
rect 433 5143 477 5149
rect 433 5123 448 5143
rect 468 5123 477 5143
rect 433 5107 477 5123
rect 547 5139 596 5149
rect 547 5119 558 5139
rect 578 5119 596 5139
rect 547 5107 596 5119
rect 646 5143 690 5149
rect 646 5123 661 5143
rect 681 5123 690 5143
rect 646 5107 690 5123
rect 755 5139 804 5149
rect 755 5119 766 5139
rect 786 5119 804 5139
rect 755 5107 804 5119
rect 854 5143 898 5149
rect 854 5123 869 5143
rect 889 5123 898 5143
rect 854 5107 898 5123
rect 968 5143 1012 5149
rect 968 5123 977 5143
rect 997 5123 1012 5143
rect 968 5107 1012 5123
rect 1062 5139 1111 5149
rect 1062 5119 1080 5139
rect 1100 5119 1111 5139
rect 1062 5107 1111 5119
rect 5390 5180 5439 5190
rect 5390 5160 5401 5180
rect 5421 5160 5439 5180
rect 2774 5091 2823 5103
rect 2774 5071 2785 5091
rect 2805 5071 2823 5091
rect 2774 5061 2823 5071
rect 2873 5087 2917 5103
rect 2873 5067 2888 5087
rect 2908 5067 2917 5087
rect 2873 5061 2917 5067
rect 2987 5087 3031 5103
rect 2987 5067 2996 5087
rect 3016 5067 3031 5087
rect 2987 5061 3031 5067
rect 3081 5091 3130 5103
rect 3081 5071 3099 5091
rect 3119 5071 3130 5091
rect 3081 5061 3130 5071
rect 3195 5087 3239 5103
rect 3195 5067 3204 5087
rect 3224 5067 3239 5087
rect 3195 5061 3239 5067
rect 3289 5091 3338 5103
rect 3289 5071 3307 5091
rect 3327 5071 3338 5091
rect 3289 5061 3338 5071
rect 3408 5087 3452 5103
rect 3408 5067 3417 5087
rect 3437 5067 3452 5087
rect 3408 5061 3452 5067
rect 3502 5091 3551 5103
rect 3502 5071 3520 5091
rect 3540 5071 3551 5091
rect 5390 5148 5439 5160
rect 5489 5184 5533 5190
rect 5489 5164 5504 5184
rect 5524 5164 5533 5184
rect 5489 5148 5533 5164
rect 5603 5180 5652 5190
rect 5603 5160 5614 5180
rect 5634 5160 5652 5180
rect 5603 5148 5652 5160
rect 5702 5184 5746 5190
rect 5702 5164 5717 5184
rect 5737 5164 5746 5184
rect 5702 5148 5746 5164
rect 5811 5180 5860 5190
rect 5811 5160 5822 5180
rect 5842 5160 5860 5180
rect 5811 5148 5860 5160
rect 5910 5184 5954 5190
rect 5910 5164 5925 5184
rect 5945 5164 5954 5184
rect 5910 5148 5954 5164
rect 6024 5184 6068 5190
rect 6024 5164 6033 5184
rect 6053 5164 6068 5184
rect 6024 5148 6068 5164
rect 6118 5180 6167 5190
rect 6118 5160 6136 5180
rect 6156 5160 6167 5180
rect 6118 5148 6167 5160
rect 7830 5132 7879 5144
rect 3502 5061 3551 5071
rect 7830 5112 7841 5132
rect 7861 5112 7879 5132
rect 7830 5102 7879 5112
rect 7929 5128 7973 5144
rect 7929 5108 7944 5128
rect 7964 5108 7973 5128
rect 7929 5102 7973 5108
rect 8043 5128 8087 5144
rect 8043 5108 8052 5128
rect 8072 5108 8087 5128
rect 8043 5102 8087 5108
rect 8137 5132 8186 5144
rect 8137 5112 8155 5132
rect 8175 5112 8186 5132
rect 8137 5102 8186 5112
rect 8251 5128 8295 5144
rect 8251 5108 8260 5128
rect 8280 5108 8295 5128
rect 8251 5102 8295 5108
rect 8345 5132 8394 5144
rect 8345 5112 8363 5132
rect 8383 5112 8394 5132
rect 8345 5102 8394 5112
rect 8464 5128 8508 5144
rect 8464 5108 8473 5128
rect 8493 5108 8508 5128
rect 8464 5102 8508 5108
rect 8558 5132 8607 5144
rect 8558 5112 8576 5132
rect 8596 5112 8607 5132
rect 8558 5102 8607 5112
rect 1382 4876 1431 4886
rect 1382 4856 1393 4876
rect 1413 4856 1431 4876
rect 1382 4844 1431 4856
rect 1481 4880 1525 4886
rect 1481 4860 1496 4880
rect 1516 4860 1525 4880
rect 1481 4844 1525 4860
rect 1595 4876 1644 4886
rect 1595 4856 1606 4876
rect 1626 4856 1644 4876
rect 1595 4844 1644 4856
rect 1694 4880 1738 4886
rect 1694 4860 1709 4880
rect 1729 4860 1738 4880
rect 1694 4844 1738 4860
rect 1803 4876 1852 4886
rect 1803 4856 1814 4876
rect 1834 4856 1852 4876
rect 1803 4844 1852 4856
rect 1902 4880 1946 4886
rect 1902 4860 1917 4880
rect 1937 4860 1946 4880
rect 1902 4844 1946 4860
rect 2016 4880 2060 4886
rect 2016 4860 2025 4880
rect 2045 4860 2060 4880
rect 2016 4844 2060 4860
rect 2110 4876 2159 4886
rect 2110 4856 2128 4876
rect 2148 4856 2159 4876
rect 6438 4917 6487 4927
rect 2110 4844 2159 4856
rect 3822 4828 3871 4840
rect 3822 4808 3833 4828
rect 3853 4808 3871 4828
rect 3822 4798 3871 4808
rect 3921 4824 3965 4840
rect 3921 4804 3936 4824
rect 3956 4804 3965 4824
rect 3921 4798 3965 4804
rect 4035 4824 4079 4840
rect 4035 4804 4044 4824
rect 4064 4804 4079 4824
rect 4035 4798 4079 4804
rect 4129 4828 4178 4840
rect 4129 4808 4147 4828
rect 4167 4808 4178 4828
rect 4129 4798 4178 4808
rect 4243 4824 4287 4840
rect 4243 4804 4252 4824
rect 4272 4804 4287 4824
rect 4243 4798 4287 4804
rect 4337 4828 4386 4840
rect 4337 4808 4355 4828
rect 4375 4808 4386 4828
rect 4337 4798 4386 4808
rect 4456 4824 4500 4840
rect 4456 4804 4465 4824
rect 4485 4804 4500 4824
rect 4456 4798 4500 4804
rect 4550 4828 4599 4840
rect 6438 4897 6449 4917
rect 6469 4897 6487 4917
rect 6438 4885 6487 4897
rect 6537 4921 6581 4927
rect 6537 4901 6552 4921
rect 6572 4901 6581 4921
rect 6537 4885 6581 4901
rect 6651 4917 6700 4927
rect 6651 4897 6662 4917
rect 6682 4897 6700 4917
rect 6651 4885 6700 4897
rect 6750 4921 6794 4927
rect 6750 4901 6765 4921
rect 6785 4901 6794 4921
rect 6750 4885 6794 4901
rect 6859 4917 6908 4927
rect 6859 4897 6870 4917
rect 6890 4897 6908 4917
rect 6859 4885 6908 4897
rect 6958 4921 7002 4927
rect 6958 4901 6973 4921
rect 6993 4901 7002 4921
rect 6958 4885 7002 4901
rect 7072 4921 7116 4927
rect 7072 4901 7081 4921
rect 7101 4901 7116 4921
rect 7072 4885 7116 4901
rect 7166 4917 7215 4927
rect 7166 4897 7184 4917
rect 7204 4897 7215 4917
rect 7166 4885 7215 4897
rect 4550 4808 4568 4828
rect 4588 4808 4599 4828
rect 4550 4798 4599 4808
rect 8878 4869 8927 4881
rect 8878 4849 8889 4869
rect 8909 4849 8927 4869
rect 8878 4839 8927 4849
rect 8977 4865 9021 4881
rect 8977 4845 8992 4865
rect 9012 4845 9021 4865
rect 8977 4839 9021 4845
rect 9091 4865 9135 4881
rect 9091 4845 9100 4865
rect 9120 4845 9135 4865
rect 9091 4839 9135 4845
rect 9185 4869 9234 4881
rect 9185 4849 9203 4869
rect 9223 4849 9234 4869
rect 9185 4839 9234 4849
rect 9299 4865 9343 4881
rect 9299 4845 9308 4865
rect 9328 4845 9343 4865
rect 9299 4839 9343 4845
rect 9393 4869 9442 4881
rect 9393 4849 9411 4869
rect 9431 4849 9442 4869
rect 9393 4839 9442 4849
rect 9512 4865 9556 4881
rect 9512 4845 9521 4865
rect 9541 4845 9556 4865
rect 9512 4839 9556 4845
rect 9606 4869 9655 4881
rect 9606 4849 9624 4869
rect 9644 4849 9655 4869
rect 9606 4839 9655 4849
rect 335 4590 384 4600
rect 335 4570 346 4590
rect 366 4570 384 4590
rect 335 4558 384 4570
rect 434 4594 478 4600
rect 434 4574 449 4594
rect 469 4574 478 4594
rect 434 4558 478 4574
rect 548 4590 597 4600
rect 548 4570 559 4590
rect 579 4570 597 4590
rect 548 4558 597 4570
rect 647 4594 691 4600
rect 647 4574 662 4594
rect 682 4574 691 4594
rect 647 4558 691 4574
rect 756 4590 805 4600
rect 756 4570 767 4590
rect 787 4570 805 4590
rect 756 4558 805 4570
rect 855 4594 899 4600
rect 855 4574 870 4594
rect 890 4574 899 4594
rect 855 4558 899 4574
rect 969 4594 1013 4600
rect 969 4574 978 4594
rect 998 4574 1013 4594
rect 969 4558 1013 4574
rect 1063 4590 1112 4600
rect 1063 4570 1081 4590
rect 1101 4570 1112 4590
rect 1063 4558 1112 4570
rect 5391 4631 5440 4641
rect 5391 4611 5402 4631
rect 5422 4611 5440 4631
rect 5391 4599 5440 4611
rect 5490 4635 5534 4641
rect 5490 4615 5505 4635
rect 5525 4615 5534 4635
rect 5490 4599 5534 4615
rect 5604 4631 5653 4641
rect 5604 4611 5615 4631
rect 5635 4611 5653 4631
rect 5604 4599 5653 4611
rect 5703 4635 5747 4641
rect 5703 4615 5718 4635
rect 5738 4615 5747 4635
rect 5703 4599 5747 4615
rect 5812 4631 5861 4641
rect 5812 4611 5823 4631
rect 5843 4611 5861 4631
rect 5812 4599 5861 4611
rect 5911 4635 5955 4641
rect 5911 4615 5926 4635
rect 5946 4615 5955 4635
rect 5911 4599 5955 4615
rect 6025 4635 6069 4641
rect 6025 4615 6034 4635
rect 6054 4615 6069 4635
rect 6025 4599 6069 4615
rect 6119 4631 6168 4641
rect 6119 4611 6137 4631
rect 6157 4611 6168 4631
rect 6119 4599 6168 4611
rect 2883 4518 2932 4530
rect 2883 4498 2894 4518
rect 2914 4498 2932 4518
rect 2883 4488 2932 4498
rect 2982 4514 3026 4530
rect 2982 4494 2997 4514
rect 3017 4494 3026 4514
rect 2982 4488 3026 4494
rect 3096 4514 3140 4530
rect 3096 4494 3105 4514
rect 3125 4494 3140 4514
rect 3096 4488 3140 4494
rect 3190 4518 3239 4530
rect 3190 4498 3208 4518
rect 3228 4498 3239 4518
rect 3190 4488 3239 4498
rect 3304 4514 3348 4530
rect 3304 4494 3313 4514
rect 3333 4494 3348 4514
rect 3304 4488 3348 4494
rect 3398 4518 3447 4530
rect 3398 4498 3416 4518
rect 3436 4498 3447 4518
rect 3398 4488 3447 4498
rect 3517 4514 3561 4530
rect 3517 4494 3526 4514
rect 3546 4494 3561 4514
rect 3517 4488 3561 4494
rect 3611 4518 3660 4530
rect 3611 4498 3629 4518
rect 3649 4498 3660 4518
rect 3611 4488 3660 4498
rect 1273 4346 1322 4356
rect 1273 4326 1284 4346
rect 1304 4326 1322 4346
rect 1273 4314 1322 4326
rect 1372 4350 1416 4356
rect 1372 4330 1387 4350
rect 1407 4330 1416 4350
rect 1372 4314 1416 4330
rect 1486 4346 1535 4356
rect 1486 4326 1497 4346
rect 1517 4326 1535 4346
rect 1486 4314 1535 4326
rect 1585 4350 1629 4356
rect 1585 4330 1600 4350
rect 1620 4330 1629 4350
rect 1585 4314 1629 4330
rect 1694 4346 1743 4356
rect 1694 4326 1705 4346
rect 1725 4326 1743 4346
rect 1694 4314 1743 4326
rect 1793 4350 1837 4356
rect 1793 4330 1808 4350
rect 1828 4330 1837 4350
rect 1793 4314 1837 4330
rect 1907 4350 1951 4356
rect 1907 4330 1916 4350
rect 1936 4330 1951 4350
rect 1907 4314 1951 4330
rect 2001 4346 2050 4356
rect 2001 4326 2019 4346
rect 2039 4326 2050 4346
rect 2001 4314 2050 4326
rect 7939 4559 7988 4571
rect 7939 4539 7950 4559
rect 7970 4539 7988 4559
rect 7939 4529 7988 4539
rect 8038 4555 8082 4571
rect 8038 4535 8053 4555
rect 8073 4535 8082 4555
rect 8038 4529 8082 4535
rect 8152 4555 8196 4571
rect 8152 4535 8161 4555
rect 8181 4535 8196 4555
rect 8152 4529 8196 4535
rect 8246 4559 8295 4571
rect 8246 4539 8264 4559
rect 8284 4539 8295 4559
rect 8246 4529 8295 4539
rect 8360 4555 8404 4571
rect 8360 4535 8369 4555
rect 8389 4535 8404 4555
rect 8360 4529 8404 4535
rect 8454 4559 8503 4571
rect 8454 4539 8472 4559
rect 8492 4539 8503 4559
rect 8454 4529 8503 4539
rect 8573 4555 8617 4571
rect 8573 4535 8582 4555
rect 8602 4535 8617 4555
rect 8573 4529 8617 4535
rect 8667 4559 8716 4571
rect 8667 4539 8685 4559
rect 8705 4539 8716 4559
rect 8667 4529 8716 4539
rect 6329 4387 6378 4397
rect 6329 4367 6340 4387
rect 6360 4367 6378 4387
rect 6329 4355 6378 4367
rect 6428 4391 6472 4397
rect 6428 4371 6443 4391
rect 6463 4371 6472 4391
rect 6428 4355 6472 4371
rect 6542 4387 6591 4397
rect 6542 4367 6553 4387
rect 6573 4367 6591 4387
rect 6542 4355 6591 4367
rect 6641 4391 6685 4397
rect 6641 4371 6656 4391
rect 6676 4371 6685 4391
rect 6641 4355 6685 4371
rect 6750 4387 6799 4397
rect 6750 4367 6761 4387
rect 6781 4367 6799 4387
rect 6750 4355 6799 4367
rect 6849 4391 6893 4397
rect 6849 4371 6864 4391
rect 6884 4371 6893 4391
rect 6849 4355 6893 4371
rect 6963 4391 7007 4397
rect 6963 4371 6972 4391
rect 6992 4371 7007 4391
rect 6963 4355 7007 4371
rect 7057 4387 7106 4397
rect 7057 4367 7075 4387
rect 7095 4367 7106 4387
rect 7057 4355 7106 4367
rect 3821 4274 3870 4286
rect 3821 4254 3832 4274
rect 3852 4254 3870 4274
rect 3821 4244 3870 4254
rect 3920 4270 3964 4286
rect 3920 4250 3935 4270
rect 3955 4250 3964 4270
rect 3920 4244 3964 4250
rect 4034 4270 4078 4286
rect 4034 4250 4043 4270
rect 4063 4250 4078 4270
rect 4034 4244 4078 4250
rect 4128 4274 4177 4286
rect 4128 4254 4146 4274
rect 4166 4254 4177 4274
rect 4128 4244 4177 4254
rect 4242 4270 4286 4286
rect 4242 4250 4251 4270
rect 4271 4250 4286 4270
rect 4242 4244 4286 4250
rect 4336 4274 4385 4286
rect 4336 4254 4354 4274
rect 4374 4254 4385 4274
rect 4336 4244 4385 4254
rect 4455 4270 4499 4286
rect 4455 4250 4464 4270
rect 4484 4250 4499 4270
rect 4455 4244 4499 4250
rect 4549 4274 4598 4286
rect 4549 4254 4567 4274
rect 4587 4254 4598 4274
rect 4549 4244 4598 4254
rect 8877 4315 8926 4327
rect 8877 4295 8888 4315
rect 8908 4295 8926 4315
rect 8877 4285 8926 4295
rect 8976 4311 9020 4327
rect 8976 4291 8991 4311
rect 9011 4291 9020 4311
rect 8976 4285 9020 4291
rect 9090 4311 9134 4327
rect 9090 4291 9099 4311
rect 9119 4291 9134 4311
rect 9090 4285 9134 4291
rect 9184 4315 9233 4327
rect 9184 4295 9202 4315
rect 9222 4295 9233 4315
rect 9184 4285 9233 4295
rect 9298 4311 9342 4327
rect 9298 4291 9307 4311
rect 9327 4291 9342 4311
rect 9298 4285 9342 4291
rect 9392 4315 9441 4327
rect 9392 4295 9410 4315
rect 9430 4295 9441 4315
rect 9392 4285 9441 4295
rect 9511 4311 9555 4327
rect 9511 4291 9520 4311
rect 9540 4291 9555 4311
rect 9511 4285 9555 4291
rect 9605 4315 9654 4327
rect 9605 4295 9623 4315
rect 9643 4295 9654 4315
rect 9605 4285 9654 4295
rect 5390 4077 5439 4087
rect 5390 4057 5401 4077
rect 5421 4057 5439 4077
rect 334 4036 383 4046
rect 334 4016 345 4036
rect 365 4016 383 4036
rect 334 4004 383 4016
rect 433 4040 477 4046
rect 433 4020 448 4040
rect 468 4020 477 4040
rect 433 4004 477 4020
rect 547 4036 596 4046
rect 547 4016 558 4036
rect 578 4016 596 4036
rect 547 4004 596 4016
rect 646 4040 690 4046
rect 646 4020 661 4040
rect 681 4020 690 4040
rect 646 4004 690 4020
rect 755 4036 804 4046
rect 755 4016 766 4036
rect 786 4016 804 4036
rect 755 4004 804 4016
rect 854 4040 898 4046
rect 854 4020 869 4040
rect 889 4020 898 4040
rect 854 4004 898 4020
rect 968 4040 1012 4046
rect 968 4020 977 4040
rect 997 4020 1012 4040
rect 968 4004 1012 4020
rect 1062 4036 1111 4046
rect 1062 4016 1080 4036
rect 1100 4016 1111 4036
rect 1062 4004 1111 4016
rect 2743 4007 2792 4019
rect 2743 3987 2754 4007
rect 2774 3987 2792 4007
rect 2743 3977 2792 3987
rect 2842 4003 2886 4019
rect 2842 3983 2857 4003
rect 2877 3983 2886 4003
rect 2842 3977 2886 3983
rect 2956 4003 3000 4019
rect 2956 3983 2965 4003
rect 2985 3983 3000 4003
rect 2956 3977 3000 3983
rect 3050 4007 3099 4019
rect 3050 3987 3068 4007
rect 3088 3987 3099 4007
rect 3050 3977 3099 3987
rect 3164 4003 3208 4019
rect 3164 3983 3173 4003
rect 3193 3983 3208 4003
rect 3164 3977 3208 3983
rect 3258 4007 3307 4019
rect 3258 3987 3276 4007
rect 3296 3987 3307 4007
rect 3258 3977 3307 3987
rect 3377 4003 3421 4019
rect 3377 3983 3386 4003
rect 3406 3983 3421 4003
rect 3377 3977 3421 3983
rect 3471 4007 3520 4019
rect 3471 3987 3489 4007
rect 3509 3987 3520 4007
rect 3471 3977 3520 3987
rect 5390 4045 5439 4057
rect 5489 4081 5533 4087
rect 5489 4061 5504 4081
rect 5524 4061 5533 4081
rect 5489 4045 5533 4061
rect 5603 4077 5652 4087
rect 5603 4057 5614 4077
rect 5634 4057 5652 4077
rect 5603 4045 5652 4057
rect 5702 4081 5746 4087
rect 5702 4061 5717 4081
rect 5737 4061 5746 4081
rect 5702 4045 5746 4061
rect 5811 4077 5860 4087
rect 5811 4057 5822 4077
rect 5842 4057 5860 4077
rect 5811 4045 5860 4057
rect 5910 4081 5954 4087
rect 5910 4061 5925 4081
rect 5945 4061 5954 4081
rect 5910 4045 5954 4061
rect 6024 4081 6068 4087
rect 6024 4061 6033 4081
rect 6053 4061 6068 4081
rect 6024 4045 6068 4061
rect 6118 4077 6167 4087
rect 6118 4057 6136 4077
rect 6156 4057 6167 4077
rect 6118 4045 6167 4057
rect 7799 4048 7848 4060
rect 7799 4028 7810 4048
rect 7830 4028 7848 4048
rect 7799 4018 7848 4028
rect 7898 4044 7942 4060
rect 7898 4024 7913 4044
rect 7933 4024 7942 4044
rect 7898 4018 7942 4024
rect 8012 4044 8056 4060
rect 8012 4024 8021 4044
rect 8041 4024 8056 4044
rect 8012 4018 8056 4024
rect 8106 4048 8155 4060
rect 8106 4028 8124 4048
rect 8144 4028 8155 4048
rect 8106 4018 8155 4028
rect 8220 4044 8264 4060
rect 8220 4024 8229 4044
rect 8249 4024 8264 4044
rect 8220 4018 8264 4024
rect 8314 4048 8363 4060
rect 8314 4028 8332 4048
rect 8352 4028 8363 4048
rect 8314 4018 8363 4028
rect 8433 4044 8477 4060
rect 8433 4024 8442 4044
rect 8462 4024 8477 4044
rect 8433 4018 8477 4024
rect 8527 4048 8576 4060
rect 8527 4028 8545 4048
rect 8565 4028 8576 4048
rect 8527 4018 8576 4028
rect 1414 3754 1463 3764
rect 1414 3734 1425 3754
rect 1445 3734 1463 3754
rect 1414 3722 1463 3734
rect 1513 3758 1557 3764
rect 1513 3738 1528 3758
rect 1548 3738 1557 3758
rect 1513 3722 1557 3738
rect 1627 3754 1676 3764
rect 1627 3734 1638 3754
rect 1658 3734 1676 3754
rect 1627 3722 1676 3734
rect 1726 3758 1770 3764
rect 1726 3738 1741 3758
rect 1761 3738 1770 3758
rect 1726 3722 1770 3738
rect 1835 3754 1884 3764
rect 1835 3734 1846 3754
rect 1866 3734 1884 3754
rect 1835 3722 1884 3734
rect 1934 3758 1978 3764
rect 1934 3738 1949 3758
rect 1969 3738 1978 3758
rect 1934 3722 1978 3738
rect 2048 3758 2092 3764
rect 2048 3738 2057 3758
rect 2077 3738 2092 3758
rect 2048 3722 2092 3738
rect 2142 3754 2191 3764
rect 2142 3734 2160 3754
rect 2180 3734 2191 3754
rect 2142 3722 2191 3734
rect 3823 3725 3872 3737
rect 3823 3705 3834 3725
rect 3854 3705 3872 3725
rect 3823 3695 3872 3705
rect 3922 3721 3966 3737
rect 3922 3701 3937 3721
rect 3957 3701 3966 3721
rect 3922 3695 3966 3701
rect 4036 3721 4080 3737
rect 4036 3701 4045 3721
rect 4065 3701 4080 3721
rect 4036 3695 4080 3701
rect 4130 3725 4179 3737
rect 4130 3705 4148 3725
rect 4168 3705 4179 3725
rect 4130 3695 4179 3705
rect 4244 3721 4288 3737
rect 4244 3701 4253 3721
rect 4273 3701 4288 3721
rect 4244 3695 4288 3701
rect 4338 3725 4387 3737
rect 4338 3705 4356 3725
rect 4376 3705 4387 3725
rect 4338 3695 4387 3705
rect 4457 3721 4501 3737
rect 4457 3701 4466 3721
rect 4486 3701 4501 3721
rect 4457 3695 4501 3701
rect 4551 3725 4600 3737
rect 6470 3795 6519 3805
rect 6470 3775 6481 3795
rect 6501 3775 6519 3795
rect 6470 3763 6519 3775
rect 6569 3799 6613 3805
rect 6569 3779 6584 3799
rect 6604 3779 6613 3799
rect 6569 3763 6613 3779
rect 6683 3795 6732 3805
rect 6683 3775 6694 3795
rect 6714 3775 6732 3795
rect 6683 3763 6732 3775
rect 6782 3799 6826 3805
rect 6782 3779 6797 3799
rect 6817 3779 6826 3799
rect 6782 3763 6826 3779
rect 6891 3795 6940 3805
rect 6891 3775 6902 3795
rect 6922 3775 6940 3795
rect 6891 3763 6940 3775
rect 6990 3799 7034 3805
rect 6990 3779 7005 3799
rect 7025 3779 7034 3799
rect 6990 3763 7034 3779
rect 7104 3799 7148 3805
rect 7104 3779 7113 3799
rect 7133 3779 7148 3799
rect 7104 3763 7148 3779
rect 7198 3795 7247 3805
rect 7198 3775 7216 3795
rect 7236 3775 7247 3795
rect 7198 3763 7247 3775
rect 8879 3766 8928 3778
rect 8879 3746 8890 3766
rect 8910 3746 8928 3766
rect 8879 3736 8928 3746
rect 8978 3762 9022 3778
rect 8978 3742 8993 3762
rect 9013 3742 9022 3762
rect 8978 3736 9022 3742
rect 9092 3762 9136 3778
rect 9092 3742 9101 3762
rect 9121 3742 9136 3762
rect 9092 3736 9136 3742
rect 9186 3766 9235 3778
rect 9186 3746 9204 3766
rect 9224 3746 9235 3766
rect 9186 3736 9235 3746
rect 9300 3762 9344 3778
rect 9300 3742 9309 3762
rect 9329 3742 9344 3762
rect 9300 3736 9344 3742
rect 9394 3766 9443 3778
rect 9394 3746 9412 3766
rect 9432 3746 9443 3766
rect 9394 3736 9443 3746
rect 9513 3762 9557 3778
rect 9513 3742 9522 3762
rect 9542 3742 9557 3762
rect 9513 3736 9557 3742
rect 9607 3766 9656 3778
rect 9607 3746 9625 3766
rect 9645 3746 9656 3766
rect 9607 3736 9656 3746
rect 4551 3705 4569 3725
rect 4589 3705 4600 3725
rect 4551 3695 4600 3705
rect 336 3487 385 3497
rect 336 3467 347 3487
rect 367 3467 385 3487
rect 336 3455 385 3467
rect 435 3491 479 3497
rect 435 3471 450 3491
rect 470 3471 479 3491
rect 435 3455 479 3471
rect 549 3487 598 3497
rect 549 3467 560 3487
rect 580 3467 598 3487
rect 549 3455 598 3467
rect 648 3491 692 3497
rect 648 3471 663 3491
rect 683 3471 692 3491
rect 648 3455 692 3471
rect 757 3487 806 3497
rect 757 3467 768 3487
rect 788 3467 806 3487
rect 757 3455 806 3467
rect 856 3491 900 3497
rect 856 3471 871 3491
rect 891 3471 900 3491
rect 856 3455 900 3471
rect 970 3491 1014 3497
rect 970 3471 979 3491
rect 999 3471 1014 3491
rect 970 3455 1014 3471
rect 1064 3487 1113 3497
rect 1064 3467 1082 3487
rect 1102 3467 1113 3487
rect 1064 3455 1113 3467
rect 5392 3528 5441 3538
rect 5392 3508 5403 3528
rect 5423 3508 5441 3528
rect 5392 3496 5441 3508
rect 5491 3532 5535 3538
rect 5491 3512 5506 3532
rect 5526 3512 5535 3532
rect 5491 3496 5535 3512
rect 5605 3528 5654 3538
rect 5605 3508 5616 3528
rect 5636 3508 5654 3528
rect 5605 3496 5654 3508
rect 5704 3532 5748 3538
rect 5704 3512 5719 3532
rect 5739 3512 5748 3532
rect 5704 3496 5748 3512
rect 5813 3528 5862 3538
rect 5813 3508 5824 3528
rect 5844 3508 5862 3528
rect 5813 3496 5862 3508
rect 5912 3532 5956 3538
rect 5912 3512 5927 3532
rect 5947 3512 5956 3532
rect 5912 3496 5956 3512
rect 6026 3532 6070 3538
rect 6026 3512 6035 3532
rect 6055 3512 6070 3532
rect 6026 3496 6070 3512
rect 6120 3528 6169 3538
rect 6120 3508 6138 3528
rect 6158 3508 6169 3528
rect 6120 3496 6169 3508
rect 2884 3415 2933 3427
rect 2884 3395 2895 3415
rect 2915 3395 2933 3415
rect 2884 3385 2933 3395
rect 2983 3411 3027 3427
rect 2983 3391 2998 3411
rect 3018 3391 3027 3411
rect 2983 3385 3027 3391
rect 3097 3411 3141 3427
rect 3097 3391 3106 3411
rect 3126 3391 3141 3411
rect 3097 3385 3141 3391
rect 3191 3415 3240 3427
rect 3191 3395 3209 3415
rect 3229 3395 3240 3415
rect 3191 3385 3240 3395
rect 3305 3411 3349 3427
rect 3305 3391 3314 3411
rect 3334 3391 3349 3411
rect 3305 3385 3349 3391
rect 3399 3415 3448 3427
rect 3399 3395 3417 3415
rect 3437 3395 3448 3415
rect 3399 3385 3448 3395
rect 3518 3411 3562 3427
rect 3518 3391 3527 3411
rect 3547 3391 3562 3411
rect 3518 3385 3562 3391
rect 3612 3415 3661 3427
rect 3612 3395 3630 3415
rect 3650 3395 3661 3415
rect 3612 3385 3661 3395
rect 1274 3243 1323 3253
rect 1274 3223 1285 3243
rect 1305 3223 1323 3243
rect 1274 3211 1323 3223
rect 1373 3247 1417 3253
rect 1373 3227 1388 3247
rect 1408 3227 1417 3247
rect 1373 3211 1417 3227
rect 1487 3243 1536 3253
rect 1487 3223 1498 3243
rect 1518 3223 1536 3243
rect 1487 3211 1536 3223
rect 1586 3247 1630 3253
rect 1586 3227 1601 3247
rect 1621 3227 1630 3247
rect 1586 3211 1630 3227
rect 1695 3243 1744 3253
rect 1695 3223 1706 3243
rect 1726 3223 1744 3243
rect 1695 3211 1744 3223
rect 1794 3247 1838 3253
rect 1794 3227 1809 3247
rect 1829 3227 1838 3247
rect 1794 3211 1838 3227
rect 1908 3247 1952 3253
rect 1908 3227 1917 3247
rect 1937 3227 1952 3247
rect 1908 3211 1952 3227
rect 2002 3243 2051 3253
rect 2002 3223 2020 3243
rect 2040 3223 2051 3243
rect 2002 3211 2051 3223
rect 7940 3456 7989 3468
rect 7940 3436 7951 3456
rect 7971 3436 7989 3456
rect 7940 3426 7989 3436
rect 8039 3452 8083 3468
rect 8039 3432 8054 3452
rect 8074 3432 8083 3452
rect 8039 3426 8083 3432
rect 8153 3452 8197 3468
rect 8153 3432 8162 3452
rect 8182 3432 8197 3452
rect 8153 3426 8197 3432
rect 8247 3456 8296 3468
rect 8247 3436 8265 3456
rect 8285 3436 8296 3456
rect 8247 3426 8296 3436
rect 8361 3452 8405 3468
rect 8361 3432 8370 3452
rect 8390 3432 8405 3452
rect 8361 3426 8405 3432
rect 8455 3456 8504 3468
rect 8455 3436 8473 3456
rect 8493 3436 8504 3456
rect 8455 3426 8504 3436
rect 8574 3452 8618 3468
rect 8574 3432 8583 3452
rect 8603 3432 8618 3452
rect 8574 3426 8618 3432
rect 8668 3456 8717 3468
rect 8668 3436 8686 3456
rect 8706 3436 8717 3456
rect 8668 3426 8717 3436
rect 6330 3284 6379 3294
rect 6330 3264 6341 3284
rect 6361 3264 6379 3284
rect 6330 3252 6379 3264
rect 6429 3288 6473 3294
rect 6429 3268 6444 3288
rect 6464 3268 6473 3288
rect 6429 3252 6473 3268
rect 6543 3284 6592 3294
rect 6543 3264 6554 3284
rect 6574 3264 6592 3284
rect 6543 3252 6592 3264
rect 6642 3288 6686 3294
rect 6642 3268 6657 3288
rect 6677 3268 6686 3288
rect 6642 3252 6686 3268
rect 6751 3284 6800 3294
rect 6751 3264 6762 3284
rect 6782 3264 6800 3284
rect 6751 3252 6800 3264
rect 6850 3288 6894 3294
rect 6850 3268 6865 3288
rect 6885 3268 6894 3288
rect 6850 3252 6894 3268
rect 6964 3288 7008 3294
rect 6964 3268 6973 3288
rect 6993 3268 7008 3288
rect 6964 3252 7008 3268
rect 7058 3284 7107 3294
rect 7058 3264 7076 3284
rect 7096 3264 7107 3284
rect 7058 3252 7107 3264
rect 3822 3171 3871 3183
rect 3822 3151 3833 3171
rect 3853 3151 3871 3171
rect 3822 3141 3871 3151
rect 3921 3167 3965 3183
rect 3921 3147 3936 3167
rect 3956 3147 3965 3167
rect 3921 3141 3965 3147
rect 4035 3167 4079 3183
rect 4035 3147 4044 3167
rect 4064 3147 4079 3167
rect 4035 3141 4079 3147
rect 4129 3171 4178 3183
rect 4129 3151 4147 3171
rect 4167 3151 4178 3171
rect 4129 3141 4178 3151
rect 4243 3167 4287 3183
rect 4243 3147 4252 3167
rect 4272 3147 4287 3167
rect 4243 3141 4287 3147
rect 4337 3171 4386 3183
rect 4337 3151 4355 3171
rect 4375 3151 4386 3171
rect 4337 3141 4386 3151
rect 4456 3167 4500 3183
rect 4456 3147 4465 3167
rect 4485 3147 4500 3167
rect 4456 3141 4500 3147
rect 4550 3171 4599 3183
rect 4550 3151 4568 3171
rect 4588 3151 4599 3171
rect 4550 3141 4599 3151
rect 8878 3212 8927 3224
rect 8878 3192 8889 3212
rect 8909 3192 8927 3212
rect 8878 3182 8927 3192
rect 8977 3208 9021 3224
rect 8977 3188 8992 3208
rect 9012 3188 9021 3208
rect 8977 3182 9021 3188
rect 9091 3208 9135 3224
rect 9091 3188 9100 3208
rect 9120 3188 9135 3208
rect 9091 3182 9135 3188
rect 9185 3212 9234 3224
rect 9185 3192 9203 3212
rect 9223 3192 9234 3212
rect 9185 3182 9234 3192
rect 9299 3208 9343 3224
rect 9299 3188 9308 3208
rect 9328 3188 9343 3208
rect 9299 3182 9343 3188
rect 9393 3212 9442 3224
rect 9393 3192 9411 3212
rect 9431 3192 9442 3212
rect 9393 3182 9442 3192
rect 9512 3208 9556 3224
rect 9512 3188 9521 3208
rect 9541 3188 9556 3208
rect 9512 3182 9556 3188
rect 9606 3212 9655 3224
rect 9606 3192 9624 3212
rect 9644 3192 9655 3212
rect 9606 3182 9655 3192
rect 5391 2974 5440 2984
rect 5391 2954 5402 2974
rect 5422 2954 5440 2974
rect 335 2933 384 2943
rect 335 2913 346 2933
rect 366 2913 384 2933
rect 335 2901 384 2913
rect 434 2937 478 2943
rect 434 2917 449 2937
rect 469 2917 478 2937
rect 434 2901 478 2917
rect 548 2933 597 2943
rect 548 2913 559 2933
rect 579 2913 597 2933
rect 548 2901 597 2913
rect 647 2937 691 2943
rect 647 2917 662 2937
rect 682 2917 691 2937
rect 647 2901 691 2917
rect 756 2933 805 2943
rect 756 2913 767 2933
rect 787 2913 805 2933
rect 756 2901 805 2913
rect 855 2937 899 2943
rect 855 2917 870 2937
rect 890 2917 899 2937
rect 855 2901 899 2917
rect 969 2937 1013 2943
rect 969 2917 978 2937
rect 998 2917 1013 2937
rect 969 2901 1013 2917
rect 1063 2933 1112 2943
rect 1063 2913 1081 2933
rect 1101 2913 1112 2933
rect 1063 2901 1112 2913
rect 2774 2891 2823 2903
rect 2774 2871 2785 2891
rect 2805 2871 2823 2891
rect 2774 2861 2823 2871
rect 2873 2887 2917 2903
rect 2873 2867 2888 2887
rect 2908 2867 2917 2887
rect 2873 2861 2917 2867
rect 2987 2887 3031 2903
rect 2987 2867 2996 2887
rect 3016 2867 3031 2887
rect 2987 2861 3031 2867
rect 3081 2891 3130 2903
rect 3081 2871 3099 2891
rect 3119 2871 3130 2891
rect 3081 2861 3130 2871
rect 3195 2887 3239 2903
rect 3195 2867 3204 2887
rect 3224 2867 3239 2887
rect 3195 2861 3239 2867
rect 3289 2891 3338 2903
rect 3289 2871 3307 2891
rect 3327 2871 3338 2891
rect 3289 2861 3338 2871
rect 3408 2887 3452 2903
rect 3408 2867 3417 2887
rect 3437 2867 3452 2887
rect 3408 2861 3452 2867
rect 3502 2891 3551 2903
rect 3502 2871 3520 2891
rect 3540 2871 3551 2891
rect 5391 2942 5440 2954
rect 5490 2978 5534 2984
rect 5490 2958 5505 2978
rect 5525 2958 5534 2978
rect 5490 2942 5534 2958
rect 5604 2974 5653 2984
rect 5604 2954 5615 2974
rect 5635 2954 5653 2974
rect 5604 2942 5653 2954
rect 5703 2978 5747 2984
rect 5703 2958 5718 2978
rect 5738 2958 5747 2978
rect 5703 2942 5747 2958
rect 5812 2974 5861 2984
rect 5812 2954 5823 2974
rect 5843 2954 5861 2974
rect 5812 2942 5861 2954
rect 5911 2978 5955 2984
rect 5911 2958 5926 2978
rect 5946 2958 5955 2978
rect 5911 2942 5955 2958
rect 6025 2978 6069 2984
rect 6025 2958 6034 2978
rect 6054 2958 6069 2978
rect 6025 2942 6069 2958
rect 6119 2974 6168 2984
rect 6119 2954 6137 2974
rect 6157 2954 6168 2974
rect 6119 2942 6168 2954
rect 7830 2932 7879 2944
rect 7830 2912 7841 2932
rect 7861 2912 7879 2932
rect 3502 2861 3551 2871
rect 7830 2902 7879 2912
rect 7929 2928 7973 2944
rect 7929 2908 7944 2928
rect 7964 2908 7973 2928
rect 7929 2902 7973 2908
rect 8043 2928 8087 2944
rect 8043 2908 8052 2928
rect 8072 2908 8087 2928
rect 8043 2902 8087 2908
rect 8137 2932 8186 2944
rect 8137 2912 8155 2932
rect 8175 2912 8186 2932
rect 8137 2902 8186 2912
rect 8251 2928 8295 2944
rect 8251 2908 8260 2928
rect 8280 2908 8295 2928
rect 8251 2902 8295 2908
rect 8345 2932 8394 2944
rect 8345 2912 8363 2932
rect 8383 2912 8394 2932
rect 8345 2902 8394 2912
rect 8464 2928 8508 2944
rect 8464 2908 8473 2928
rect 8493 2908 8508 2928
rect 8464 2902 8508 2908
rect 8558 2932 8607 2944
rect 8558 2912 8576 2932
rect 8596 2912 8607 2932
rect 8558 2902 8607 2912
rect 1384 2664 1433 2674
rect 1384 2644 1395 2664
rect 1415 2644 1433 2664
rect 1384 2632 1433 2644
rect 1483 2668 1527 2674
rect 1483 2648 1498 2668
rect 1518 2648 1527 2668
rect 1483 2632 1527 2648
rect 1597 2664 1646 2674
rect 1597 2644 1608 2664
rect 1628 2644 1646 2664
rect 1597 2632 1646 2644
rect 1696 2668 1740 2674
rect 1696 2648 1711 2668
rect 1731 2648 1740 2668
rect 1696 2632 1740 2648
rect 1805 2664 1854 2674
rect 1805 2644 1816 2664
rect 1836 2644 1854 2664
rect 1805 2632 1854 2644
rect 1904 2668 1948 2674
rect 1904 2648 1919 2668
rect 1939 2648 1948 2668
rect 1904 2632 1948 2648
rect 2018 2668 2062 2674
rect 2018 2648 2027 2668
rect 2047 2648 2062 2668
rect 2018 2632 2062 2648
rect 2112 2664 2161 2674
rect 6440 2705 6489 2715
rect 2112 2644 2130 2664
rect 2150 2644 2161 2664
rect 2112 2632 2161 2644
rect 3823 2622 3872 2634
rect 3823 2602 3834 2622
rect 3854 2602 3872 2622
rect 3823 2592 3872 2602
rect 3922 2618 3966 2634
rect 3922 2598 3937 2618
rect 3957 2598 3966 2618
rect 3922 2592 3966 2598
rect 4036 2618 4080 2634
rect 4036 2598 4045 2618
rect 4065 2598 4080 2618
rect 4036 2592 4080 2598
rect 4130 2622 4179 2634
rect 4130 2602 4148 2622
rect 4168 2602 4179 2622
rect 4130 2592 4179 2602
rect 4244 2618 4288 2634
rect 4244 2598 4253 2618
rect 4273 2598 4288 2618
rect 4244 2592 4288 2598
rect 4338 2622 4387 2634
rect 4338 2602 4356 2622
rect 4376 2602 4387 2622
rect 4338 2592 4387 2602
rect 4457 2618 4501 2634
rect 4457 2598 4466 2618
rect 4486 2598 4501 2618
rect 4457 2592 4501 2598
rect 4551 2622 4600 2634
rect 6440 2685 6451 2705
rect 6471 2685 6489 2705
rect 6440 2673 6489 2685
rect 6539 2709 6583 2715
rect 6539 2689 6554 2709
rect 6574 2689 6583 2709
rect 6539 2673 6583 2689
rect 6653 2705 6702 2715
rect 6653 2685 6664 2705
rect 6684 2685 6702 2705
rect 6653 2673 6702 2685
rect 6752 2709 6796 2715
rect 6752 2689 6767 2709
rect 6787 2689 6796 2709
rect 6752 2673 6796 2689
rect 6861 2705 6910 2715
rect 6861 2685 6872 2705
rect 6892 2685 6910 2705
rect 6861 2673 6910 2685
rect 6960 2709 7004 2715
rect 6960 2689 6975 2709
rect 6995 2689 7004 2709
rect 6960 2673 7004 2689
rect 7074 2709 7118 2715
rect 7074 2689 7083 2709
rect 7103 2689 7118 2709
rect 7074 2673 7118 2689
rect 7168 2705 7217 2715
rect 7168 2685 7186 2705
rect 7206 2685 7217 2705
rect 7168 2673 7217 2685
rect 8879 2663 8928 2675
rect 8879 2643 8890 2663
rect 8910 2643 8928 2663
rect 8879 2633 8928 2643
rect 8978 2659 9022 2675
rect 8978 2639 8993 2659
rect 9013 2639 9022 2659
rect 8978 2633 9022 2639
rect 9092 2659 9136 2675
rect 9092 2639 9101 2659
rect 9121 2639 9136 2659
rect 9092 2633 9136 2639
rect 9186 2663 9235 2675
rect 9186 2643 9204 2663
rect 9224 2643 9235 2663
rect 9186 2633 9235 2643
rect 9300 2659 9344 2675
rect 9300 2639 9309 2659
rect 9329 2639 9344 2659
rect 9300 2633 9344 2639
rect 9394 2663 9443 2675
rect 9394 2643 9412 2663
rect 9432 2643 9443 2663
rect 9394 2633 9443 2643
rect 9513 2659 9557 2675
rect 9513 2639 9522 2659
rect 9542 2639 9557 2659
rect 9513 2633 9557 2639
rect 9607 2663 9656 2675
rect 9607 2643 9625 2663
rect 9645 2643 9656 2663
rect 9607 2633 9656 2643
rect 4551 2602 4569 2622
rect 4589 2602 4600 2622
rect 4551 2592 4600 2602
rect 336 2384 385 2394
rect 336 2364 347 2384
rect 367 2364 385 2384
rect 336 2352 385 2364
rect 435 2388 479 2394
rect 435 2368 450 2388
rect 470 2368 479 2388
rect 435 2352 479 2368
rect 549 2384 598 2394
rect 549 2364 560 2384
rect 580 2364 598 2384
rect 549 2352 598 2364
rect 648 2388 692 2394
rect 648 2368 663 2388
rect 683 2368 692 2388
rect 648 2352 692 2368
rect 757 2384 806 2394
rect 757 2364 768 2384
rect 788 2364 806 2384
rect 757 2352 806 2364
rect 856 2388 900 2394
rect 856 2368 871 2388
rect 891 2368 900 2388
rect 856 2352 900 2368
rect 970 2388 1014 2394
rect 970 2368 979 2388
rect 999 2368 1014 2388
rect 970 2352 1014 2368
rect 1064 2384 1113 2394
rect 1064 2364 1082 2384
rect 1102 2364 1113 2384
rect 1064 2352 1113 2364
rect 5392 2425 5441 2435
rect 5392 2405 5403 2425
rect 5423 2405 5441 2425
rect 5392 2393 5441 2405
rect 5491 2429 5535 2435
rect 5491 2409 5506 2429
rect 5526 2409 5535 2429
rect 5491 2393 5535 2409
rect 5605 2425 5654 2435
rect 5605 2405 5616 2425
rect 5636 2405 5654 2425
rect 5605 2393 5654 2405
rect 5704 2429 5748 2435
rect 5704 2409 5719 2429
rect 5739 2409 5748 2429
rect 5704 2393 5748 2409
rect 5813 2425 5862 2435
rect 5813 2405 5824 2425
rect 5844 2405 5862 2425
rect 5813 2393 5862 2405
rect 5912 2429 5956 2435
rect 5912 2409 5927 2429
rect 5947 2409 5956 2429
rect 5912 2393 5956 2409
rect 6026 2429 6070 2435
rect 6026 2409 6035 2429
rect 6055 2409 6070 2429
rect 6026 2393 6070 2409
rect 6120 2425 6169 2435
rect 6120 2405 6138 2425
rect 6158 2405 6169 2425
rect 6120 2393 6169 2405
rect 2884 2312 2933 2324
rect 2884 2292 2895 2312
rect 2915 2292 2933 2312
rect 2884 2282 2933 2292
rect 2983 2308 3027 2324
rect 2983 2288 2998 2308
rect 3018 2288 3027 2308
rect 2983 2282 3027 2288
rect 3097 2308 3141 2324
rect 3097 2288 3106 2308
rect 3126 2288 3141 2308
rect 3097 2282 3141 2288
rect 3191 2312 3240 2324
rect 3191 2292 3209 2312
rect 3229 2292 3240 2312
rect 3191 2282 3240 2292
rect 3305 2308 3349 2324
rect 3305 2288 3314 2308
rect 3334 2288 3349 2308
rect 3305 2282 3349 2288
rect 3399 2312 3448 2324
rect 3399 2292 3417 2312
rect 3437 2292 3448 2312
rect 3399 2282 3448 2292
rect 3518 2308 3562 2324
rect 3518 2288 3527 2308
rect 3547 2288 3562 2308
rect 3518 2282 3562 2288
rect 3612 2312 3661 2324
rect 3612 2292 3630 2312
rect 3650 2292 3661 2312
rect 3612 2282 3661 2292
rect 1274 2140 1323 2150
rect 1274 2120 1285 2140
rect 1305 2120 1323 2140
rect 1274 2108 1323 2120
rect 1373 2144 1417 2150
rect 1373 2124 1388 2144
rect 1408 2124 1417 2144
rect 1373 2108 1417 2124
rect 1487 2140 1536 2150
rect 1487 2120 1498 2140
rect 1518 2120 1536 2140
rect 1487 2108 1536 2120
rect 1586 2144 1630 2150
rect 1586 2124 1601 2144
rect 1621 2124 1630 2144
rect 1586 2108 1630 2124
rect 1695 2140 1744 2150
rect 1695 2120 1706 2140
rect 1726 2120 1744 2140
rect 1695 2108 1744 2120
rect 1794 2144 1838 2150
rect 1794 2124 1809 2144
rect 1829 2124 1838 2144
rect 1794 2108 1838 2124
rect 1908 2144 1952 2150
rect 1908 2124 1917 2144
rect 1937 2124 1952 2144
rect 1908 2108 1952 2124
rect 2002 2140 2051 2150
rect 2002 2120 2020 2140
rect 2040 2120 2051 2140
rect 2002 2108 2051 2120
rect 7940 2353 7989 2365
rect 7940 2333 7951 2353
rect 7971 2333 7989 2353
rect 7940 2323 7989 2333
rect 8039 2349 8083 2365
rect 8039 2329 8054 2349
rect 8074 2329 8083 2349
rect 8039 2323 8083 2329
rect 8153 2349 8197 2365
rect 8153 2329 8162 2349
rect 8182 2329 8197 2349
rect 8153 2323 8197 2329
rect 8247 2353 8296 2365
rect 8247 2333 8265 2353
rect 8285 2333 8296 2353
rect 8247 2323 8296 2333
rect 8361 2349 8405 2365
rect 8361 2329 8370 2349
rect 8390 2329 8405 2349
rect 8361 2323 8405 2329
rect 8455 2353 8504 2365
rect 8455 2333 8473 2353
rect 8493 2333 8504 2353
rect 8455 2323 8504 2333
rect 8574 2349 8618 2365
rect 8574 2329 8583 2349
rect 8603 2329 8618 2349
rect 8574 2323 8618 2329
rect 8668 2353 8717 2365
rect 8668 2333 8686 2353
rect 8706 2333 8717 2353
rect 8668 2323 8717 2333
rect 6330 2181 6379 2191
rect 6330 2161 6341 2181
rect 6361 2161 6379 2181
rect 6330 2149 6379 2161
rect 6429 2185 6473 2191
rect 6429 2165 6444 2185
rect 6464 2165 6473 2185
rect 6429 2149 6473 2165
rect 6543 2181 6592 2191
rect 6543 2161 6554 2181
rect 6574 2161 6592 2181
rect 6543 2149 6592 2161
rect 6642 2185 6686 2191
rect 6642 2165 6657 2185
rect 6677 2165 6686 2185
rect 6642 2149 6686 2165
rect 6751 2181 6800 2191
rect 6751 2161 6762 2181
rect 6782 2161 6800 2181
rect 6751 2149 6800 2161
rect 6850 2185 6894 2191
rect 6850 2165 6865 2185
rect 6885 2165 6894 2185
rect 6850 2149 6894 2165
rect 6964 2185 7008 2191
rect 6964 2165 6973 2185
rect 6993 2165 7008 2185
rect 6964 2149 7008 2165
rect 7058 2181 7107 2191
rect 7058 2161 7076 2181
rect 7096 2161 7107 2181
rect 7058 2149 7107 2161
rect 3822 2068 3871 2080
rect 3822 2048 3833 2068
rect 3853 2048 3871 2068
rect 3822 2038 3871 2048
rect 3921 2064 3965 2080
rect 3921 2044 3936 2064
rect 3956 2044 3965 2064
rect 3921 2038 3965 2044
rect 4035 2064 4079 2080
rect 4035 2044 4044 2064
rect 4064 2044 4079 2064
rect 4035 2038 4079 2044
rect 4129 2068 4178 2080
rect 4129 2048 4147 2068
rect 4167 2048 4178 2068
rect 4129 2038 4178 2048
rect 4243 2064 4287 2080
rect 4243 2044 4252 2064
rect 4272 2044 4287 2064
rect 4243 2038 4287 2044
rect 4337 2068 4386 2080
rect 4337 2048 4355 2068
rect 4375 2048 4386 2068
rect 4337 2038 4386 2048
rect 4456 2064 4500 2080
rect 4456 2044 4465 2064
rect 4485 2044 4500 2064
rect 4456 2038 4500 2044
rect 4550 2068 4599 2080
rect 4550 2048 4568 2068
rect 4588 2048 4599 2068
rect 4550 2038 4599 2048
rect 8878 2109 8927 2121
rect 8878 2089 8889 2109
rect 8909 2089 8927 2109
rect 8878 2079 8927 2089
rect 8977 2105 9021 2121
rect 8977 2085 8992 2105
rect 9012 2085 9021 2105
rect 8977 2079 9021 2085
rect 9091 2105 9135 2121
rect 9091 2085 9100 2105
rect 9120 2085 9135 2105
rect 9091 2079 9135 2085
rect 9185 2109 9234 2121
rect 9185 2089 9203 2109
rect 9223 2089 9234 2109
rect 9185 2079 9234 2089
rect 9299 2105 9343 2121
rect 9299 2085 9308 2105
rect 9328 2085 9343 2105
rect 9299 2079 9343 2085
rect 9393 2109 9442 2121
rect 9393 2089 9411 2109
rect 9431 2089 9442 2109
rect 9393 2079 9442 2089
rect 9512 2105 9556 2121
rect 9512 2085 9521 2105
rect 9541 2085 9556 2105
rect 9512 2079 9556 2085
rect 9606 2109 9655 2121
rect 9606 2089 9624 2109
rect 9644 2089 9655 2109
rect 9606 2079 9655 2089
rect 5391 1871 5440 1881
rect 5391 1851 5402 1871
rect 5422 1851 5440 1871
rect 335 1830 384 1840
rect 335 1810 346 1830
rect 366 1810 384 1830
rect 335 1798 384 1810
rect 434 1834 478 1840
rect 434 1814 449 1834
rect 469 1814 478 1834
rect 434 1798 478 1814
rect 548 1830 597 1840
rect 548 1810 559 1830
rect 579 1810 597 1830
rect 548 1798 597 1810
rect 647 1834 691 1840
rect 647 1814 662 1834
rect 682 1814 691 1834
rect 647 1798 691 1814
rect 756 1830 805 1840
rect 756 1810 767 1830
rect 787 1810 805 1830
rect 756 1798 805 1810
rect 855 1834 899 1840
rect 855 1814 870 1834
rect 890 1814 899 1834
rect 855 1798 899 1814
rect 969 1834 1013 1840
rect 969 1814 978 1834
rect 998 1814 1013 1834
rect 969 1798 1013 1814
rect 1063 1830 1112 1840
rect 1063 1810 1081 1830
rect 1101 1810 1112 1830
rect 1063 1798 1112 1810
rect 2744 1801 2793 1813
rect 2744 1781 2755 1801
rect 2775 1781 2793 1801
rect 2744 1771 2793 1781
rect 2843 1797 2887 1813
rect 2843 1777 2858 1797
rect 2878 1777 2887 1797
rect 2843 1771 2887 1777
rect 2957 1797 3001 1813
rect 2957 1777 2966 1797
rect 2986 1777 3001 1797
rect 2957 1771 3001 1777
rect 3051 1801 3100 1813
rect 3051 1781 3069 1801
rect 3089 1781 3100 1801
rect 3051 1771 3100 1781
rect 3165 1797 3209 1813
rect 3165 1777 3174 1797
rect 3194 1777 3209 1797
rect 3165 1771 3209 1777
rect 3259 1801 3308 1813
rect 3259 1781 3277 1801
rect 3297 1781 3308 1801
rect 3259 1771 3308 1781
rect 3378 1797 3422 1813
rect 3378 1777 3387 1797
rect 3407 1777 3422 1797
rect 3378 1771 3422 1777
rect 3472 1801 3521 1813
rect 3472 1781 3490 1801
rect 3510 1781 3521 1801
rect 3472 1771 3521 1781
rect 5391 1839 5440 1851
rect 5490 1875 5534 1881
rect 5490 1855 5505 1875
rect 5525 1855 5534 1875
rect 5490 1839 5534 1855
rect 5604 1871 5653 1881
rect 5604 1851 5615 1871
rect 5635 1851 5653 1871
rect 5604 1839 5653 1851
rect 5703 1875 5747 1881
rect 5703 1855 5718 1875
rect 5738 1855 5747 1875
rect 5703 1839 5747 1855
rect 5812 1871 5861 1881
rect 5812 1851 5823 1871
rect 5843 1851 5861 1871
rect 5812 1839 5861 1851
rect 5911 1875 5955 1881
rect 5911 1855 5926 1875
rect 5946 1855 5955 1875
rect 5911 1839 5955 1855
rect 6025 1875 6069 1881
rect 6025 1855 6034 1875
rect 6054 1855 6069 1875
rect 6025 1839 6069 1855
rect 6119 1871 6168 1881
rect 6119 1851 6137 1871
rect 6157 1851 6168 1871
rect 6119 1839 6168 1851
rect 7800 1842 7849 1854
rect 7800 1822 7811 1842
rect 7831 1822 7849 1842
rect 7800 1812 7849 1822
rect 7899 1838 7943 1854
rect 7899 1818 7914 1838
rect 7934 1818 7943 1838
rect 7899 1812 7943 1818
rect 8013 1838 8057 1854
rect 8013 1818 8022 1838
rect 8042 1818 8057 1838
rect 8013 1812 8057 1818
rect 8107 1842 8156 1854
rect 8107 1822 8125 1842
rect 8145 1822 8156 1842
rect 8107 1812 8156 1822
rect 8221 1838 8265 1854
rect 8221 1818 8230 1838
rect 8250 1818 8265 1838
rect 8221 1812 8265 1818
rect 8315 1842 8364 1854
rect 8315 1822 8333 1842
rect 8353 1822 8364 1842
rect 8315 1812 8364 1822
rect 8434 1838 8478 1854
rect 8434 1818 8443 1838
rect 8463 1818 8478 1838
rect 8434 1812 8478 1818
rect 8528 1842 8577 1854
rect 8528 1822 8546 1842
rect 8566 1822 8577 1842
rect 8528 1812 8577 1822
rect 1415 1548 1464 1558
rect 1415 1528 1426 1548
rect 1446 1528 1464 1548
rect 1415 1516 1464 1528
rect 1514 1552 1558 1558
rect 1514 1532 1529 1552
rect 1549 1532 1558 1552
rect 1514 1516 1558 1532
rect 1628 1548 1677 1558
rect 1628 1528 1639 1548
rect 1659 1528 1677 1548
rect 1628 1516 1677 1528
rect 1727 1552 1771 1558
rect 1727 1532 1742 1552
rect 1762 1532 1771 1552
rect 1727 1516 1771 1532
rect 1836 1548 1885 1558
rect 1836 1528 1847 1548
rect 1867 1528 1885 1548
rect 1836 1516 1885 1528
rect 1935 1552 1979 1558
rect 1935 1532 1950 1552
rect 1970 1532 1979 1552
rect 1935 1516 1979 1532
rect 2049 1552 2093 1558
rect 2049 1532 2058 1552
rect 2078 1532 2093 1552
rect 2049 1516 2093 1532
rect 2143 1548 2192 1558
rect 2143 1528 2161 1548
rect 2181 1528 2192 1548
rect 2143 1516 2192 1528
rect 3824 1519 3873 1531
rect 3824 1499 3835 1519
rect 3855 1499 3873 1519
rect 3824 1489 3873 1499
rect 3923 1515 3967 1531
rect 3923 1495 3938 1515
rect 3958 1495 3967 1515
rect 3923 1489 3967 1495
rect 4037 1515 4081 1531
rect 4037 1495 4046 1515
rect 4066 1495 4081 1515
rect 4037 1489 4081 1495
rect 4131 1519 4180 1531
rect 4131 1499 4149 1519
rect 4169 1499 4180 1519
rect 4131 1489 4180 1499
rect 4245 1515 4289 1531
rect 4245 1495 4254 1515
rect 4274 1495 4289 1515
rect 4245 1489 4289 1495
rect 4339 1519 4388 1531
rect 4339 1499 4357 1519
rect 4377 1499 4388 1519
rect 4339 1489 4388 1499
rect 4458 1515 4502 1531
rect 4458 1495 4467 1515
rect 4487 1495 4502 1515
rect 4458 1489 4502 1495
rect 4552 1519 4601 1531
rect 6471 1589 6520 1599
rect 6471 1569 6482 1589
rect 6502 1569 6520 1589
rect 6471 1557 6520 1569
rect 6570 1593 6614 1599
rect 6570 1573 6585 1593
rect 6605 1573 6614 1593
rect 6570 1557 6614 1573
rect 6684 1589 6733 1599
rect 6684 1569 6695 1589
rect 6715 1569 6733 1589
rect 6684 1557 6733 1569
rect 6783 1593 6827 1599
rect 6783 1573 6798 1593
rect 6818 1573 6827 1593
rect 6783 1557 6827 1573
rect 6892 1589 6941 1599
rect 6892 1569 6903 1589
rect 6923 1569 6941 1589
rect 6892 1557 6941 1569
rect 6991 1593 7035 1599
rect 6991 1573 7006 1593
rect 7026 1573 7035 1593
rect 6991 1557 7035 1573
rect 7105 1593 7149 1599
rect 7105 1573 7114 1593
rect 7134 1573 7149 1593
rect 7105 1557 7149 1573
rect 7199 1589 7248 1599
rect 7199 1569 7217 1589
rect 7237 1569 7248 1589
rect 7199 1557 7248 1569
rect 8880 1560 8929 1572
rect 8880 1540 8891 1560
rect 8911 1540 8929 1560
rect 8880 1530 8929 1540
rect 8979 1556 9023 1572
rect 8979 1536 8994 1556
rect 9014 1536 9023 1556
rect 8979 1530 9023 1536
rect 9093 1556 9137 1572
rect 9093 1536 9102 1556
rect 9122 1536 9137 1556
rect 9093 1530 9137 1536
rect 9187 1560 9236 1572
rect 9187 1540 9205 1560
rect 9225 1540 9236 1560
rect 9187 1530 9236 1540
rect 9301 1556 9345 1572
rect 9301 1536 9310 1556
rect 9330 1536 9345 1556
rect 9301 1530 9345 1536
rect 9395 1560 9444 1572
rect 9395 1540 9413 1560
rect 9433 1540 9444 1560
rect 9395 1530 9444 1540
rect 9514 1556 9558 1572
rect 9514 1536 9523 1556
rect 9543 1536 9558 1556
rect 9514 1530 9558 1536
rect 9608 1560 9657 1572
rect 9608 1540 9626 1560
rect 9646 1540 9657 1560
rect 9608 1530 9657 1540
rect 4552 1499 4570 1519
rect 4590 1499 4601 1519
rect 4552 1489 4601 1499
rect 337 1281 386 1291
rect 337 1261 348 1281
rect 368 1261 386 1281
rect 337 1249 386 1261
rect 436 1285 480 1291
rect 436 1265 451 1285
rect 471 1265 480 1285
rect 436 1249 480 1265
rect 550 1281 599 1291
rect 550 1261 561 1281
rect 581 1261 599 1281
rect 550 1249 599 1261
rect 649 1285 693 1291
rect 649 1265 664 1285
rect 684 1265 693 1285
rect 649 1249 693 1265
rect 758 1281 807 1291
rect 758 1261 769 1281
rect 789 1261 807 1281
rect 758 1249 807 1261
rect 857 1285 901 1291
rect 857 1265 872 1285
rect 892 1265 901 1285
rect 857 1249 901 1265
rect 971 1285 1015 1291
rect 971 1265 980 1285
rect 1000 1265 1015 1285
rect 971 1249 1015 1265
rect 1065 1281 1114 1291
rect 1065 1261 1083 1281
rect 1103 1261 1114 1281
rect 1065 1249 1114 1261
rect 5393 1322 5442 1332
rect 5393 1302 5404 1322
rect 5424 1302 5442 1322
rect 5393 1290 5442 1302
rect 5492 1326 5536 1332
rect 5492 1306 5507 1326
rect 5527 1306 5536 1326
rect 5492 1290 5536 1306
rect 5606 1322 5655 1332
rect 5606 1302 5617 1322
rect 5637 1302 5655 1322
rect 5606 1290 5655 1302
rect 5705 1326 5749 1332
rect 5705 1306 5720 1326
rect 5740 1306 5749 1326
rect 5705 1290 5749 1306
rect 5814 1322 5863 1332
rect 5814 1302 5825 1322
rect 5845 1302 5863 1322
rect 5814 1290 5863 1302
rect 5913 1326 5957 1332
rect 5913 1306 5928 1326
rect 5948 1306 5957 1326
rect 5913 1290 5957 1306
rect 6027 1326 6071 1332
rect 6027 1306 6036 1326
rect 6056 1306 6071 1326
rect 6027 1290 6071 1306
rect 6121 1322 6170 1332
rect 6121 1302 6139 1322
rect 6159 1302 6170 1322
rect 6121 1290 6170 1302
rect 2885 1209 2934 1221
rect 2885 1189 2896 1209
rect 2916 1189 2934 1209
rect 2885 1179 2934 1189
rect 2984 1205 3028 1221
rect 2984 1185 2999 1205
rect 3019 1185 3028 1205
rect 2984 1179 3028 1185
rect 3098 1205 3142 1221
rect 3098 1185 3107 1205
rect 3127 1185 3142 1205
rect 3098 1179 3142 1185
rect 3192 1209 3241 1221
rect 3192 1189 3210 1209
rect 3230 1189 3241 1209
rect 3192 1179 3241 1189
rect 3306 1205 3350 1221
rect 3306 1185 3315 1205
rect 3335 1185 3350 1205
rect 3306 1179 3350 1185
rect 3400 1209 3449 1221
rect 3400 1189 3418 1209
rect 3438 1189 3449 1209
rect 3400 1179 3449 1189
rect 3519 1205 3563 1221
rect 3519 1185 3528 1205
rect 3548 1185 3563 1205
rect 3519 1179 3563 1185
rect 3613 1209 3662 1221
rect 3613 1189 3631 1209
rect 3651 1189 3662 1209
rect 3613 1179 3662 1189
rect 1275 1037 1324 1047
rect 1275 1017 1286 1037
rect 1306 1017 1324 1037
rect 1275 1005 1324 1017
rect 1374 1041 1418 1047
rect 1374 1021 1389 1041
rect 1409 1021 1418 1041
rect 1374 1005 1418 1021
rect 1488 1037 1537 1047
rect 1488 1017 1499 1037
rect 1519 1017 1537 1037
rect 1488 1005 1537 1017
rect 1587 1041 1631 1047
rect 1587 1021 1602 1041
rect 1622 1021 1631 1041
rect 1587 1005 1631 1021
rect 1696 1037 1745 1047
rect 1696 1017 1707 1037
rect 1727 1017 1745 1037
rect 1696 1005 1745 1017
rect 1795 1041 1839 1047
rect 1795 1021 1810 1041
rect 1830 1021 1839 1041
rect 1795 1005 1839 1021
rect 1909 1041 1953 1047
rect 1909 1021 1918 1041
rect 1938 1021 1953 1041
rect 1909 1005 1953 1021
rect 2003 1037 2052 1047
rect 2003 1017 2021 1037
rect 2041 1017 2052 1037
rect 2003 1005 2052 1017
rect 7941 1250 7990 1262
rect 7941 1230 7952 1250
rect 7972 1230 7990 1250
rect 7941 1220 7990 1230
rect 8040 1246 8084 1262
rect 8040 1226 8055 1246
rect 8075 1226 8084 1246
rect 8040 1220 8084 1226
rect 8154 1246 8198 1262
rect 8154 1226 8163 1246
rect 8183 1226 8198 1246
rect 8154 1220 8198 1226
rect 8248 1250 8297 1262
rect 8248 1230 8266 1250
rect 8286 1230 8297 1250
rect 8248 1220 8297 1230
rect 8362 1246 8406 1262
rect 8362 1226 8371 1246
rect 8391 1226 8406 1246
rect 8362 1220 8406 1226
rect 8456 1250 8505 1262
rect 8456 1230 8474 1250
rect 8494 1230 8505 1250
rect 8456 1220 8505 1230
rect 8575 1246 8619 1262
rect 8575 1226 8584 1246
rect 8604 1226 8619 1246
rect 8575 1220 8619 1226
rect 8669 1250 8718 1262
rect 8669 1230 8687 1250
rect 8707 1230 8718 1250
rect 8669 1220 8718 1230
rect 6331 1078 6380 1088
rect 6331 1058 6342 1078
rect 6362 1058 6380 1078
rect 6331 1046 6380 1058
rect 6430 1082 6474 1088
rect 6430 1062 6445 1082
rect 6465 1062 6474 1082
rect 6430 1046 6474 1062
rect 6544 1078 6593 1088
rect 6544 1058 6555 1078
rect 6575 1058 6593 1078
rect 6544 1046 6593 1058
rect 6643 1082 6687 1088
rect 6643 1062 6658 1082
rect 6678 1062 6687 1082
rect 6643 1046 6687 1062
rect 6752 1078 6801 1088
rect 6752 1058 6763 1078
rect 6783 1058 6801 1078
rect 6752 1046 6801 1058
rect 6851 1082 6895 1088
rect 6851 1062 6866 1082
rect 6886 1062 6895 1082
rect 6851 1046 6895 1062
rect 6965 1082 7009 1088
rect 6965 1062 6974 1082
rect 6994 1062 7009 1082
rect 6965 1046 7009 1062
rect 7059 1078 7108 1088
rect 7059 1058 7077 1078
rect 7097 1058 7108 1078
rect 7059 1046 7108 1058
rect 3823 965 3872 977
rect 3823 945 3834 965
rect 3854 945 3872 965
rect 3823 935 3872 945
rect 3922 961 3966 977
rect 3922 941 3937 961
rect 3957 941 3966 961
rect 3922 935 3966 941
rect 4036 961 4080 977
rect 4036 941 4045 961
rect 4065 941 4080 961
rect 4036 935 4080 941
rect 4130 965 4179 977
rect 4130 945 4148 965
rect 4168 945 4179 965
rect 4130 935 4179 945
rect 4244 961 4288 977
rect 4244 941 4253 961
rect 4273 941 4288 961
rect 4244 935 4288 941
rect 4338 965 4387 977
rect 4338 945 4356 965
rect 4376 945 4387 965
rect 4338 935 4387 945
rect 4457 961 4501 977
rect 4457 941 4466 961
rect 4486 941 4501 961
rect 4457 935 4501 941
rect 4551 965 4600 977
rect 4551 945 4569 965
rect 4589 945 4600 965
rect 4551 935 4600 945
rect 8879 1006 8928 1018
rect 8879 986 8890 1006
rect 8910 986 8928 1006
rect 8879 976 8928 986
rect 8978 1002 9022 1018
rect 8978 982 8993 1002
rect 9013 982 9022 1002
rect 8978 976 9022 982
rect 9092 1002 9136 1018
rect 9092 982 9101 1002
rect 9121 982 9136 1002
rect 9092 976 9136 982
rect 9186 1006 9235 1018
rect 9186 986 9204 1006
rect 9224 986 9235 1006
rect 9186 976 9235 986
rect 9300 1002 9344 1018
rect 9300 982 9309 1002
rect 9329 982 9344 1002
rect 9300 976 9344 982
rect 9394 1006 9443 1018
rect 9394 986 9412 1006
rect 9432 986 9443 1006
rect 9394 976 9443 986
rect 9513 1002 9557 1018
rect 9513 982 9522 1002
rect 9542 982 9557 1002
rect 9513 976 9557 982
rect 9607 1006 9656 1018
rect 9607 986 9625 1006
rect 9645 986 9656 1006
rect 9607 976 9656 986
rect 5392 768 5441 778
rect 5392 748 5403 768
rect 5423 748 5441 768
rect 336 727 385 737
rect 336 707 347 727
rect 367 707 385 727
rect 336 695 385 707
rect 435 731 479 737
rect 435 711 450 731
rect 470 711 479 731
rect 435 695 479 711
rect 549 727 598 737
rect 549 707 560 727
rect 580 707 598 727
rect 549 695 598 707
rect 648 731 692 737
rect 648 711 663 731
rect 683 711 692 731
rect 648 695 692 711
rect 757 727 806 737
rect 757 707 768 727
rect 788 707 806 727
rect 757 695 806 707
rect 856 731 900 737
rect 856 711 871 731
rect 891 711 900 731
rect 856 695 900 711
rect 970 731 1014 737
rect 970 711 979 731
rect 999 711 1014 731
rect 970 695 1014 711
rect 1064 727 1113 737
rect 1064 707 1082 727
rect 1102 707 1113 727
rect 1064 695 1113 707
rect 5392 736 5441 748
rect 5491 772 5535 778
rect 5491 752 5506 772
rect 5526 752 5535 772
rect 5491 736 5535 752
rect 5605 768 5654 778
rect 5605 748 5616 768
rect 5636 748 5654 768
rect 5605 736 5654 748
rect 5704 772 5748 778
rect 5704 752 5719 772
rect 5739 752 5748 772
rect 5704 736 5748 752
rect 5813 768 5862 778
rect 5813 748 5824 768
rect 5844 748 5862 768
rect 5813 736 5862 748
rect 5912 772 5956 778
rect 5912 752 5927 772
rect 5947 752 5956 772
rect 5912 736 5956 752
rect 6026 772 6070 778
rect 6026 752 6035 772
rect 6055 752 6070 772
rect 6026 736 6070 752
rect 6120 768 6169 778
rect 6120 748 6138 768
rect 6158 748 6169 768
rect 6120 736 6169 748
rect 1583 168 1632 178
rect 1583 148 1594 168
rect 1614 148 1632 168
rect 1583 136 1632 148
rect 1682 172 1726 178
rect 1682 152 1697 172
rect 1717 152 1726 172
rect 1682 136 1726 152
rect 1796 168 1845 178
rect 1796 148 1807 168
rect 1827 148 1845 168
rect 1796 136 1845 148
rect 1895 172 1939 178
rect 1895 152 1910 172
rect 1930 152 1939 172
rect 1895 136 1939 152
rect 2004 168 2053 178
rect 2004 148 2015 168
rect 2035 148 2053 168
rect 2004 136 2053 148
rect 2103 172 2147 178
rect 2103 152 2118 172
rect 2138 152 2147 172
rect 2103 136 2147 152
rect 2217 172 2261 178
rect 2217 152 2226 172
rect 2246 152 2261 172
rect 2217 136 2261 152
rect 2311 168 2360 178
rect 2311 148 2329 168
rect 2349 148 2360 168
rect 6639 209 6688 219
rect 6639 189 6650 209
rect 6670 189 6688 209
rect 6639 177 6688 189
rect 6738 213 6782 219
rect 6738 193 6753 213
rect 6773 193 6782 213
rect 6738 177 6782 193
rect 6852 209 6901 219
rect 6852 189 6863 209
rect 6883 189 6901 209
rect 6852 177 6901 189
rect 6951 213 6995 219
rect 6951 193 6966 213
rect 6986 193 6995 213
rect 6951 177 6995 193
rect 7060 209 7109 219
rect 7060 189 7071 209
rect 7091 189 7109 209
rect 7060 177 7109 189
rect 7159 213 7203 219
rect 7159 193 7174 213
rect 7194 193 7203 213
rect 7159 177 7203 193
rect 7273 213 7317 219
rect 7273 193 7282 213
rect 7302 193 7317 213
rect 7273 177 7317 193
rect 7367 209 7416 219
rect 7367 189 7385 209
rect 7405 189 7416 209
rect 7367 177 7416 189
rect 2311 136 2360 148
rect 4533 148 4582 158
rect 4533 128 4544 148
rect 4564 128 4582 148
rect 4533 116 4582 128
rect 4632 152 4676 158
rect 4632 132 4647 152
rect 4667 132 4676 152
rect 4632 116 4676 132
rect 4746 148 4795 158
rect 4746 128 4757 148
rect 4777 128 4795 148
rect 4746 116 4795 128
rect 4845 152 4889 158
rect 4845 132 4860 152
rect 4880 132 4889 152
rect 4845 116 4889 132
rect 4954 148 5003 158
rect 4954 128 4965 148
rect 4985 128 5003 148
rect 4954 116 5003 128
rect 5053 152 5097 158
rect 5053 132 5068 152
rect 5088 132 5097 152
rect 5053 116 5097 132
rect 5167 152 5211 158
rect 5167 132 5176 152
rect 5196 132 5211 152
rect 5167 116 5211 132
rect 5261 148 5310 158
rect 5261 128 5279 148
rect 5299 128 5310 148
rect 5261 116 5310 128
<< pdiff >>
rect 338 9151 382 9189
rect 338 9131 350 9151
rect 370 9131 382 9151
rect 338 9089 382 9131
rect 432 9151 474 9189
rect 432 9131 446 9151
rect 466 9131 474 9151
rect 432 9089 474 9131
rect 551 9151 595 9189
rect 551 9131 563 9151
rect 583 9131 595 9151
rect 551 9089 595 9131
rect 645 9151 687 9189
rect 645 9131 659 9151
rect 679 9131 687 9151
rect 645 9089 687 9131
rect 759 9151 803 9189
rect 759 9131 771 9151
rect 791 9131 803 9151
rect 759 9089 803 9131
rect 853 9151 895 9189
rect 853 9131 867 9151
rect 887 9131 895 9151
rect 853 9089 895 9131
rect 969 9151 1011 9189
rect 969 9131 977 9151
rect 997 9131 1011 9151
rect 969 9089 1011 9131
rect 1061 9158 1106 9189
rect 1061 9151 1105 9158
rect 1061 9131 1073 9151
rect 1093 9131 1105 9151
rect 5394 9192 5438 9230
rect 5394 9172 5406 9192
rect 5426 9172 5438 9192
rect 1061 9089 1105 9131
rect 3825 9091 3869 9133
rect 3825 9071 3837 9091
rect 3857 9071 3869 9091
rect 3825 9064 3869 9071
rect 3824 9033 3869 9064
rect 3919 9091 3961 9133
rect 3919 9071 3933 9091
rect 3953 9071 3961 9091
rect 3919 9033 3961 9071
rect 4035 9091 4077 9133
rect 4035 9071 4043 9091
rect 4063 9071 4077 9091
rect 4035 9033 4077 9071
rect 4127 9091 4171 9133
rect 4127 9071 4139 9091
rect 4159 9071 4171 9091
rect 4127 9033 4171 9071
rect 4243 9091 4285 9133
rect 4243 9071 4251 9091
rect 4271 9071 4285 9091
rect 4243 9033 4285 9071
rect 4335 9091 4379 9133
rect 4335 9071 4347 9091
rect 4367 9071 4379 9091
rect 4335 9033 4379 9071
rect 4456 9091 4498 9133
rect 4456 9071 4464 9091
rect 4484 9071 4498 9091
rect 4456 9033 4498 9071
rect 4548 9091 4592 9133
rect 5394 9130 5438 9172
rect 5488 9192 5530 9230
rect 5488 9172 5502 9192
rect 5522 9172 5530 9192
rect 5488 9130 5530 9172
rect 5607 9192 5651 9230
rect 5607 9172 5619 9192
rect 5639 9172 5651 9192
rect 5607 9130 5651 9172
rect 5701 9192 5743 9230
rect 5701 9172 5715 9192
rect 5735 9172 5743 9192
rect 5701 9130 5743 9172
rect 5815 9192 5859 9230
rect 5815 9172 5827 9192
rect 5847 9172 5859 9192
rect 5815 9130 5859 9172
rect 5909 9192 5951 9230
rect 5909 9172 5923 9192
rect 5943 9172 5951 9192
rect 5909 9130 5951 9172
rect 6025 9192 6067 9230
rect 6025 9172 6033 9192
rect 6053 9172 6067 9192
rect 6025 9130 6067 9172
rect 6117 9199 6162 9230
rect 6117 9192 6161 9199
rect 6117 9172 6129 9192
rect 6149 9172 6161 9192
rect 6117 9130 6161 9172
rect 8881 9132 8925 9174
rect 4548 9071 4560 9091
rect 4580 9071 4592 9091
rect 4548 9033 4592 9071
rect 8881 9112 8893 9132
rect 8913 9112 8925 9132
rect 8881 9105 8925 9112
rect 8880 9074 8925 9105
rect 8975 9132 9017 9174
rect 8975 9112 8989 9132
rect 9009 9112 9017 9132
rect 8975 9074 9017 9112
rect 9091 9132 9133 9174
rect 9091 9112 9099 9132
rect 9119 9112 9133 9132
rect 9091 9074 9133 9112
rect 9183 9132 9227 9174
rect 9183 9112 9195 9132
rect 9215 9112 9227 9132
rect 9183 9074 9227 9112
rect 9299 9132 9341 9174
rect 9299 9112 9307 9132
rect 9327 9112 9341 9132
rect 9299 9074 9341 9112
rect 9391 9132 9435 9174
rect 9391 9112 9403 9132
rect 9423 9112 9435 9132
rect 9391 9074 9435 9112
rect 9512 9132 9554 9174
rect 9512 9112 9520 9132
rect 9540 9112 9554 9132
rect 9512 9074 9554 9112
rect 9604 9132 9648 9174
rect 9604 9112 9616 9132
rect 9636 9112 9648 9132
rect 9604 9074 9648 9112
rect 1276 8907 1320 8945
rect 1276 8887 1288 8907
rect 1308 8887 1320 8907
rect 1276 8845 1320 8887
rect 1370 8907 1412 8945
rect 1370 8887 1384 8907
rect 1404 8887 1412 8907
rect 1370 8845 1412 8887
rect 1489 8907 1533 8945
rect 1489 8887 1501 8907
rect 1521 8887 1533 8907
rect 1489 8845 1533 8887
rect 1583 8907 1625 8945
rect 1583 8887 1597 8907
rect 1617 8887 1625 8907
rect 1583 8845 1625 8887
rect 1697 8907 1741 8945
rect 1697 8887 1709 8907
rect 1729 8887 1741 8907
rect 1697 8845 1741 8887
rect 1791 8907 1833 8945
rect 1791 8887 1805 8907
rect 1825 8887 1833 8907
rect 1791 8845 1833 8887
rect 1907 8907 1949 8945
rect 1907 8887 1915 8907
rect 1935 8887 1949 8907
rect 1907 8845 1949 8887
rect 1999 8914 2044 8945
rect 1999 8907 2043 8914
rect 1999 8887 2011 8907
rect 2031 8887 2043 8907
rect 1999 8845 2043 8887
rect 6332 8948 6376 8986
rect 6332 8928 6344 8948
rect 6364 8928 6376 8948
rect 2886 8781 2930 8823
rect 2886 8761 2898 8781
rect 2918 8761 2930 8781
rect 2886 8754 2930 8761
rect 2885 8723 2930 8754
rect 2980 8781 3022 8823
rect 2980 8761 2994 8781
rect 3014 8761 3022 8781
rect 2980 8723 3022 8761
rect 3096 8781 3138 8823
rect 3096 8761 3104 8781
rect 3124 8761 3138 8781
rect 3096 8723 3138 8761
rect 3188 8781 3232 8823
rect 3188 8761 3200 8781
rect 3220 8761 3232 8781
rect 3188 8723 3232 8761
rect 3304 8781 3346 8823
rect 3304 8761 3312 8781
rect 3332 8761 3346 8781
rect 3304 8723 3346 8761
rect 3396 8781 3440 8823
rect 3396 8761 3408 8781
rect 3428 8761 3440 8781
rect 3396 8723 3440 8761
rect 3517 8781 3559 8823
rect 3517 8761 3525 8781
rect 3545 8761 3559 8781
rect 3517 8723 3559 8761
rect 3609 8781 3653 8823
rect 6332 8886 6376 8928
rect 6426 8948 6468 8986
rect 6426 8928 6440 8948
rect 6460 8928 6468 8948
rect 6426 8886 6468 8928
rect 6545 8948 6589 8986
rect 6545 8928 6557 8948
rect 6577 8928 6589 8948
rect 6545 8886 6589 8928
rect 6639 8948 6681 8986
rect 6639 8928 6653 8948
rect 6673 8928 6681 8948
rect 6639 8886 6681 8928
rect 6753 8948 6797 8986
rect 6753 8928 6765 8948
rect 6785 8928 6797 8948
rect 6753 8886 6797 8928
rect 6847 8948 6889 8986
rect 6847 8928 6861 8948
rect 6881 8928 6889 8948
rect 6847 8886 6889 8928
rect 6963 8948 7005 8986
rect 6963 8928 6971 8948
rect 6991 8928 7005 8948
rect 6963 8886 7005 8928
rect 7055 8955 7100 8986
rect 7055 8948 7099 8955
rect 7055 8928 7067 8948
rect 7087 8928 7099 8948
rect 7055 8886 7099 8928
rect 3609 8761 3621 8781
rect 3641 8761 3653 8781
rect 3609 8723 3653 8761
rect 7942 8822 7986 8864
rect 7942 8802 7954 8822
rect 7974 8802 7986 8822
rect 7942 8795 7986 8802
rect 7941 8764 7986 8795
rect 8036 8822 8078 8864
rect 8036 8802 8050 8822
rect 8070 8802 8078 8822
rect 8036 8764 8078 8802
rect 8152 8822 8194 8864
rect 8152 8802 8160 8822
rect 8180 8802 8194 8822
rect 8152 8764 8194 8802
rect 8244 8822 8288 8864
rect 8244 8802 8256 8822
rect 8276 8802 8288 8822
rect 8244 8764 8288 8802
rect 8360 8822 8402 8864
rect 8360 8802 8368 8822
rect 8388 8802 8402 8822
rect 8360 8764 8402 8802
rect 8452 8822 8496 8864
rect 8452 8802 8464 8822
rect 8484 8802 8496 8822
rect 8452 8764 8496 8802
rect 8573 8822 8615 8864
rect 8573 8802 8581 8822
rect 8601 8802 8615 8822
rect 8573 8764 8615 8802
rect 8665 8822 8709 8864
rect 8665 8802 8677 8822
rect 8697 8802 8709 8822
rect 8665 8764 8709 8802
rect 337 8597 381 8635
rect 337 8577 349 8597
rect 369 8577 381 8597
rect 337 8535 381 8577
rect 431 8597 473 8635
rect 431 8577 445 8597
rect 465 8577 473 8597
rect 431 8535 473 8577
rect 550 8597 594 8635
rect 550 8577 562 8597
rect 582 8577 594 8597
rect 550 8535 594 8577
rect 644 8597 686 8635
rect 644 8577 658 8597
rect 678 8577 686 8597
rect 644 8535 686 8577
rect 758 8597 802 8635
rect 758 8577 770 8597
rect 790 8577 802 8597
rect 758 8535 802 8577
rect 852 8597 894 8635
rect 852 8577 866 8597
rect 886 8577 894 8597
rect 852 8535 894 8577
rect 968 8597 1010 8635
rect 968 8577 976 8597
rect 996 8577 1010 8597
rect 968 8535 1010 8577
rect 1060 8604 1105 8635
rect 1060 8597 1104 8604
rect 1060 8577 1072 8597
rect 1092 8577 1104 8597
rect 5393 8638 5437 8676
rect 5393 8618 5405 8638
rect 5425 8618 5437 8638
rect 1060 8535 1104 8577
rect 3824 8537 3868 8579
rect 3824 8517 3836 8537
rect 3856 8517 3868 8537
rect 3824 8510 3868 8517
rect 3823 8479 3868 8510
rect 3918 8537 3960 8579
rect 3918 8517 3932 8537
rect 3952 8517 3960 8537
rect 3918 8479 3960 8517
rect 4034 8537 4076 8579
rect 4034 8517 4042 8537
rect 4062 8517 4076 8537
rect 4034 8479 4076 8517
rect 4126 8537 4170 8579
rect 4126 8517 4138 8537
rect 4158 8517 4170 8537
rect 4126 8479 4170 8517
rect 4242 8537 4284 8579
rect 4242 8517 4250 8537
rect 4270 8517 4284 8537
rect 4242 8479 4284 8517
rect 4334 8537 4378 8579
rect 4334 8517 4346 8537
rect 4366 8517 4378 8537
rect 4334 8479 4378 8517
rect 4455 8537 4497 8579
rect 4455 8517 4463 8537
rect 4483 8517 4497 8537
rect 4455 8479 4497 8517
rect 4547 8537 4591 8579
rect 5393 8576 5437 8618
rect 5487 8638 5529 8676
rect 5487 8618 5501 8638
rect 5521 8618 5529 8638
rect 5487 8576 5529 8618
rect 5606 8638 5650 8676
rect 5606 8618 5618 8638
rect 5638 8618 5650 8638
rect 5606 8576 5650 8618
rect 5700 8638 5742 8676
rect 5700 8618 5714 8638
rect 5734 8618 5742 8638
rect 5700 8576 5742 8618
rect 5814 8638 5858 8676
rect 5814 8618 5826 8638
rect 5846 8618 5858 8638
rect 5814 8576 5858 8618
rect 5908 8638 5950 8676
rect 5908 8618 5922 8638
rect 5942 8618 5950 8638
rect 5908 8576 5950 8618
rect 6024 8638 6066 8676
rect 6024 8618 6032 8638
rect 6052 8618 6066 8638
rect 6024 8576 6066 8618
rect 6116 8645 6161 8676
rect 6116 8638 6160 8645
rect 6116 8618 6128 8638
rect 6148 8618 6160 8638
rect 6116 8576 6160 8618
rect 8880 8578 8924 8620
rect 4547 8517 4559 8537
rect 4579 8517 4591 8537
rect 4547 8479 4591 8517
rect 8880 8558 8892 8578
rect 8912 8558 8924 8578
rect 8880 8551 8924 8558
rect 8879 8520 8924 8551
rect 8974 8578 9016 8620
rect 8974 8558 8988 8578
rect 9008 8558 9016 8578
rect 8974 8520 9016 8558
rect 9090 8578 9132 8620
rect 9090 8558 9098 8578
rect 9118 8558 9132 8578
rect 9090 8520 9132 8558
rect 9182 8578 9226 8620
rect 9182 8558 9194 8578
rect 9214 8558 9226 8578
rect 9182 8520 9226 8558
rect 9298 8578 9340 8620
rect 9298 8558 9306 8578
rect 9326 8558 9340 8578
rect 9298 8520 9340 8558
rect 9390 8578 9434 8620
rect 9390 8558 9402 8578
rect 9422 8558 9434 8578
rect 9390 8520 9434 8558
rect 9511 8578 9553 8620
rect 9511 8558 9519 8578
rect 9539 8558 9553 8578
rect 9511 8520 9553 8558
rect 9603 8578 9647 8620
rect 9603 8558 9615 8578
rect 9635 8558 9647 8578
rect 9603 8520 9647 8558
rect 1417 8315 1461 8353
rect 1417 8295 1429 8315
rect 1449 8295 1461 8315
rect 1417 8253 1461 8295
rect 1511 8315 1553 8353
rect 1511 8295 1525 8315
rect 1545 8295 1553 8315
rect 1511 8253 1553 8295
rect 1630 8315 1674 8353
rect 1630 8295 1642 8315
rect 1662 8295 1674 8315
rect 1630 8253 1674 8295
rect 1724 8315 1766 8353
rect 1724 8295 1738 8315
rect 1758 8295 1766 8315
rect 1724 8253 1766 8295
rect 1838 8315 1882 8353
rect 1838 8295 1850 8315
rect 1870 8295 1882 8315
rect 1838 8253 1882 8295
rect 1932 8315 1974 8353
rect 1932 8295 1946 8315
rect 1966 8295 1974 8315
rect 1932 8253 1974 8295
rect 2048 8315 2090 8353
rect 2048 8295 2056 8315
rect 2076 8295 2090 8315
rect 2048 8253 2090 8295
rect 2140 8322 2185 8353
rect 2140 8315 2184 8322
rect 2140 8295 2152 8315
rect 2172 8295 2184 8315
rect 6473 8356 6517 8394
rect 6473 8336 6485 8356
rect 6505 8336 6517 8356
rect 2140 8253 2184 8295
rect 2746 8270 2790 8312
rect 2746 8250 2758 8270
rect 2778 8250 2790 8270
rect 2746 8243 2790 8250
rect 2745 8212 2790 8243
rect 2840 8270 2882 8312
rect 2840 8250 2854 8270
rect 2874 8250 2882 8270
rect 2840 8212 2882 8250
rect 2956 8270 2998 8312
rect 2956 8250 2964 8270
rect 2984 8250 2998 8270
rect 2956 8212 2998 8250
rect 3048 8270 3092 8312
rect 3048 8250 3060 8270
rect 3080 8250 3092 8270
rect 3048 8212 3092 8250
rect 3164 8270 3206 8312
rect 3164 8250 3172 8270
rect 3192 8250 3206 8270
rect 3164 8212 3206 8250
rect 3256 8270 3300 8312
rect 3256 8250 3268 8270
rect 3288 8250 3300 8270
rect 3256 8212 3300 8250
rect 3377 8270 3419 8312
rect 3377 8250 3385 8270
rect 3405 8250 3419 8270
rect 3377 8212 3419 8250
rect 3469 8270 3513 8312
rect 6473 8294 6517 8336
rect 6567 8356 6609 8394
rect 6567 8336 6581 8356
rect 6601 8336 6609 8356
rect 6567 8294 6609 8336
rect 6686 8356 6730 8394
rect 6686 8336 6698 8356
rect 6718 8336 6730 8356
rect 6686 8294 6730 8336
rect 6780 8356 6822 8394
rect 6780 8336 6794 8356
rect 6814 8336 6822 8356
rect 6780 8294 6822 8336
rect 6894 8356 6938 8394
rect 6894 8336 6906 8356
rect 6926 8336 6938 8356
rect 6894 8294 6938 8336
rect 6988 8356 7030 8394
rect 6988 8336 7002 8356
rect 7022 8336 7030 8356
rect 6988 8294 7030 8336
rect 7104 8356 7146 8394
rect 7104 8336 7112 8356
rect 7132 8336 7146 8356
rect 7104 8294 7146 8336
rect 7196 8363 7241 8394
rect 7196 8356 7240 8363
rect 7196 8336 7208 8356
rect 7228 8336 7240 8356
rect 7196 8294 7240 8336
rect 7802 8311 7846 8353
rect 3469 8250 3481 8270
rect 3501 8250 3513 8270
rect 3469 8212 3513 8250
rect 7802 8291 7814 8311
rect 7834 8291 7846 8311
rect 7802 8284 7846 8291
rect 7801 8253 7846 8284
rect 7896 8311 7938 8353
rect 7896 8291 7910 8311
rect 7930 8291 7938 8311
rect 7896 8253 7938 8291
rect 8012 8311 8054 8353
rect 8012 8291 8020 8311
rect 8040 8291 8054 8311
rect 8012 8253 8054 8291
rect 8104 8311 8148 8353
rect 8104 8291 8116 8311
rect 8136 8291 8148 8311
rect 8104 8253 8148 8291
rect 8220 8311 8262 8353
rect 8220 8291 8228 8311
rect 8248 8291 8262 8311
rect 8220 8253 8262 8291
rect 8312 8311 8356 8353
rect 8312 8291 8324 8311
rect 8344 8291 8356 8311
rect 8312 8253 8356 8291
rect 8433 8311 8475 8353
rect 8433 8291 8441 8311
rect 8461 8291 8475 8311
rect 8433 8253 8475 8291
rect 8525 8311 8569 8353
rect 8525 8291 8537 8311
rect 8557 8291 8569 8311
rect 8525 8253 8569 8291
rect 339 8048 383 8086
rect 339 8028 351 8048
rect 371 8028 383 8048
rect 339 7986 383 8028
rect 433 8048 475 8086
rect 433 8028 447 8048
rect 467 8028 475 8048
rect 433 7986 475 8028
rect 552 8048 596 8086
rect 552 8028 564 8048
rect 584 8028 596 8048
rect 552 7986 596 8028
rect 646 8048 688 8086
rect 646 8028 660 8048
rect 680 8028 688 8048
rect 646 7986 688 8028
rect 760 8048 804 8086
rect 760 8028 772 8048
rect 792 8028 804 8048
rect 760 7986 804 8028
rect 854 8048 896 8086
rect 854 8028 868 8048
rect 888 8028 896 8048
rect 854 7986 896 8028
rect 970 8048 1012 8086
rect 970 8028 978 8048
rect 998 8028 1012 8048
rect 970 7986 1012 8028
rect 1062 8055 1107 8086
rect 1062 8048 1106 8055
rect 1062 8028 1074 8048
rect 1094 8028 1106 8048
rect 5395 8089 5439 8127
rect 5395 8069 5407 8089
rect 5427 8069 5439 8089
rect 1062 7986 1106 8028
rect 3826 7988 3870 8030
rect 3826 7968 3838 7988
rect 3858 7968 3870 7988
rect 3826 7961 3870 7968
rect 3825 7930 3870 7961
rect 3920 7988 3962 8030
rect 3920 7968 3934 7988
rect 3954 7968 3962 7988
rect 3920 7930 3962 7968
rect 4036 7988 4078 8030
rect 4036 7968 4044 7988
rect 4064 7968 4078 7988
rect 4036 7930 4078 7968
rect 4128 7988 4172 8030
rect 4128 7968 4140 7988
rect 4160 7968 4172 7988
rect 4128 7930 4172 7968
rect 4244 7988 4286 8030
rect 4244 7968 4252 7988
rect 4272 7968 4286 7988
rect 4244 7930 4286 7968
rect 4336 7988 4380 8030
rect 4336 7968 4348 7988
rect 4368 7968 4380 7988
rect 4336 7930 4380 7968
rect 4457 7988 4499 8030
rect 4457 7968 4465 7988
rect 4485 7968 4499 7988
rect 4457 7930 4499 7968
rect 4549 7988 4593 8030
rect 5395 8027 5439 8069
rect 5489 8089 5531 8127
rect 5489 8069 5503 8089
rect 5523 8069 5531 8089
rect 5489 8027 5531 8069
rect 5608 8089 5652 8127
rect 5608 8069 5620 8089
rect 5640 8069 5652 8089
rect 5608 8027 5652 8069
rect 5702 8089 5744 8127
rect 5702 8069 5716 8089
rect 5736 8069 5744 8089
rect 5702 8027 5744 8069
rect 5816 8089 5860 8127
rect 5816 8069 5828 8089
rect 5848 8069 5860 8089
rect 5816 8027 5860 8069
rect 5910 8089 5952 8127
rect 5910 8069 5924 8089
rect 5944 8069 5952 8089
rect 5910 8027 5952 8069
rect 6026 8089 6068 8127
rect 6026 8069 6034 8089
rect 6054 8069 6068 8089
rect 6026 8027 6068 8069
rect 6118 8096 6163 8127
rect 6118 8089 6162 8096
rect 6118 8069 6130 8089
rect 6150 8069 6162 8089
rect 6118 8027 6162 8069
rect 8882 8029 8926 8071
rect 4549 7968 4561 7988
rect 4581 7968 4593 7988
rect 4549 7930 4593 7968
rect 8882 8009 8894 8029
rect 8914 8009 8926 8029
rect 8882 8002 8926 8009
rect 8881 7971 8926 8002
rect 8976 8029 9018 8071
rect 8976 8009 8990 8029
rect 9010 8009 9018 8029
rect 8976 7971 9018 8009
rect 9092 8029 9134 8071
rect 9092 8009 9100 8029
rect 9120 8009 9134 8029
rect 9092 7971 9134 8009
rect 9184 8029 9228 8071
rect 9184 8009 9196 8029
rect 9216 8009 9228 8029
rect 9184 7971 9228 8009
rect 9300 8029 9342 8071
rect 9300 8009 9308 8029
rect 9328 8009 9342 8029
rect 9300 7971 9342 8009
rect 9392 8029 9436 8071
rect 9392 8009 9404 8029
rect 9424 8009 9436 8029
rect 9392 7971 9436 8009
rect 9513 8029 9555 8071
rect 9513 8009 9521 8029
rect 9541 8009 9555 8029
rect 9513 7971 9555 8009
rect 9605 8029 9649 8071
rect 9605 8009 9617 8029
rect 9637 8009 9649 8029
rect 9605 7971 9649 8009
rect 1277 7804 1321 7842
rect 1277 7784 1289 7804
rect 1309 7784 1321 7804
rect 1277 7742 1321 7784
rect 1371 7804 1413 7842
rect 1371 7784 1385 7804
rect 1405 7784 1413 7804
rect 1371 7742 1413 7784
rect 1490 7804 1534 7842
rect 1490 7784 1502 7804
rect 1522 7784 1534 7804
rect 1490 7742 1534 7784
rect 1584 7804 1626 7842
rect 1584 7784 1598 7804
rect 1618 7784 1626 7804
rect 1584 7742 1626 7784
rect 1698 7804 1742 7842
rect 1698 7784 1710 7804
rect 1730 7784 1742 7804
rect 1698 7742 1742 7784
rect 1792 7804 1834 7842
rect 1792 7784 1806 7804
rect 1826 7784 1834 7804
rect 1792 7742 1834 7784
rect 1908 7804 1950 7842
rect 1908 7784 1916 7804
rect 1936 7784 1950 7804
rect 1908 7742 1950 7784
rect 2000 7811 2045 7842
rect 2000 7804 2044 7811
rect 2000 7784 2012 7804
rect 2032 7784 2044 7804
rect 2000 7742 2044 7784
rect 6333 7845 6377 7883
rect 6333 7825 6345 7845
rect 6365 7825 6377 7845
rect 2887 7678 2931 7720
rect 2887 7658 2899 7678
rect 2919 7658 2931 7678
rect 2887 7651 2931 7658
rect 2886 7620 2931 7651
rect 2981 7678 3023 7720
rect 2981 7658 2995 7678
rect 3015 7658 3023 7678
rect 2981 7620 3023 7658
rect 3097 7678 3139 7720
rect 3097 7658 3105 7678
rect 3125 7658 3139 7678
rect 3097 7620 3139 7658
rect 3189 7678 3233 7720
rect 3189 7658 3201 7678
rect 3221 7658 3233 7678
rect 3189 7620 3233 7658
rect 3305 7678 3347 7720
rect 3305 7658 3313 7678
rect 3333 7658 3347 7678
rect 3305 7620 3347 7658
rect 3397 7678 3441 7720
rect 3397 7658 3409 7678
rect 3429 7658 3441 7678
rect 3397 7620 3441 7658
rect 3518 7678 3560 7720
rect 3518 7658 3526 7678
rect 3546 7658 3560 7678
rect 3518 7620 3560 7658
rect 3610 7678 3654 7720
rect 6333 7783 6377 7825
rect 6427 7845 6469 7883
rect 6427 7825 6441 7845
rect 6461 7825 6469 7845
rect 6427 7783 6469 7825
rect 6546 7845 6590 7883
rect 6546 7825 6558 7845
rect 6578 7825 6590 7845
rect 6546 7783 6590 7825
rect 6640 7845 6682 7883
rect 6640 7825 6654 7845
rect 6674 7825 6682 7845
rect 6640 7783 6682 7825
rect 6754 7845 6798 7883
rect 6754 7825 6766 7845
rect 6786 7825 6798 7845
rect 6754 7783 6798 7825
rect 6848 7845 6890 7883
rect 6848 7825 6862 7845
rect 6882 7825 6890 7845
rect 6848 7783 6890 7825
rect 6964 7845 7006 7883
rect 6964 7825 6972 7845
rect 6992 7825 7006 7845
rect 6964 7783 7006 7825
rect 7056 7852 7101 7883
rect 7056 7845 7100 7852
rect 7056 7825 7068 7845
rect 7088 7825 7100 7845
rect 7056 7783 7100 7825
rect 3610 7658 3622 7678
rect 3642 7658 3654 7678
rect 3610 7620 3654 7658
rect 7943 7719 7987 7761
rect 7943 7699 7955 7719
rect 7975 7699 7987 7719
rect 7943 7692 7987 7699
rect 7942 7661 7987 7692
rect 8037 7719 8079 7761
rect 8037 7699 8051 7719
rect 8071 7699 8079 7719
rect 8037 7661 8079 7699
rect 8153 7719 8195 7761
rect 8153 7699 8161 7719
rect 8181 7699 8195 7719
rect 8153 7661 8195 7699
rect 8245 7719 8289 7761
rect 8245 7699 8257 7719
rect 8277 7699 8289 7719
rect 8245 7661 8289 7699
rect 8361 7719 8403 7761
rect 8361 7699 8369 7719
rect 8389 7699 8403 7719
rect 8361 7661 8403 7699
rect 8453 7719 8497 7761
rect 8453 7699 8465 7719
rect 8485 7699 8497 7719
rect 8453 7661 8497 7699
rect 8574 7719 8616 7761
rect 8574 7699 8582 7719
rect 8602 7699 8616 7719
rect 8574 7661 8616 7699
rect 8666 7719 8710 7761
rect 8666 7699 8678 7719
rect 8698 7699 8710 7719
rect 8666 7661 8710 7699
rect 338 7494 382 7532
rect 338 7474 350 7494
rect 370 7474 382 7494
rect 338 7432 382 7474
rect 432 7494 474 7532
rect 432 7474 446 7494
rect 466 7474 474 7494
rect 432 7432 474 7474
rect 551 7494 595 7532
rect 551 7474 563 7494
rect 583 7474 595 7494
rect 551 7432 595 7474
rect 645 7494 687 7532
rect 645 7474 659 7494
rect 679 7474 687 7494
rect 645 7432 687 7474
rect 759 7494 803 7532
rect 759 7474 771 7494
rect 791 7474 803 7494
rect 759 7432 803 7474
rect 853 7494 895 7532
rect 853 7474 867 7494
rect 887 7474 895 7494
rect 853 7432 895 7474
rect 969 7494 1011 7532
rect 969 7474 977 7494
rect 997 7474 1011 7494
rect 969 7432 1011 7474
rect 1061 7501 1106 7532
rect 1061 7494 1105 7501
rect 1061 7474 1073 7494
rect 1093 7474 1105 7494
rect 5394 7535 5438 7573
rect 5394 7515 5406 7535
rect 5426 7515 5438 7535
rect 1061 7432 1105 7474
rect 3825 7434 3869 7476
rect 3825 7414 3837 7434
rect 3857 7414 3869 7434
rect 3825 7407 3869 7414
rect 3824 7376 3869 7407
rect 3919 7434 3961 7476
rect 3919 7414 3933 7434
rect 3953 7414 3961 7434
rect 3919 7376 3961 7414
rect 4035 7434 4077 7476
rect 4035 7414 4043 7434
rect 4063 7414 4077 7434
rect 4035 7376 4077 7414
rect 4127 7434 4171 7476
rect 4127 7414 4139 7434
rect 4159 7414 4171 7434
rect 4127 7376 4171 7414
rect 4243 7434 4285 7476
rect 4243 7414 4251 7434
rect 4271 7414 4285 7434
rect 4243 7376 4285 7414
rect 4335 7434 4379 7476
rect 4335 7414 4347 7434
rect 4367 7414 4379 7434
rect 4335 7376 4379 7414
rect 4456 7434 4498 7476
rect 4456 7414 4464 7434
rect 4484 7414 4498 7434
rect 4456 7376 4498 7414
rect 4548 7434 4592 7476
rect 5394 7473 5438 7515
rect 5488 7535 5530 7573
rect 5488 7515 5502 7535
rect 5522 7515 5530 7535
rect 5488 7473 5530 7515
rect 5607 7535 5651 7573
rect 5607 7515 5619 7535
rect 5639 7515 5651 7535
rect 5607 7473 5651 7515
rect 5701 7535 5743 7573
rect 5701 7515 5715 7535
rect 5735 7515 5743 7535
rect 5701 7473 5743 7515
rect 5815 7535 5859 7573
rect 5815 7515 5827 7535
rect 5847 7515 5859 7535
rect 5815 7473 5859 7515
rect 5909 7535 5951 7573
rect 5909 7515 5923 7535
rect 5943 7515 5951 7535
rect 5909 7473 5951 7515
rect 6025 7535 6067 7573
rect 6025 7515 6033 7535
rect 6053 7515 6067 7535
rect 6025 7473 6067 7515
rect 6117 7542 6162 7573
rect 6117 7535 6161 7542
rect 6117 7515 6129 7535
rect 6149 7515 6161 7535
rect 6117 7473 6161 7515
rect 8881 7475 8925 7517
rect 4548 7414 4560 7434
rect 4580 7414 4592 7434
rect 4548 7376 4592 7414
rect 8881 7455 8893 7475
rect 8913 7455 8925 7475
rect 8881 7448 8925 7455
rect 8880 7417 8925 7448
rect 8975 7475 9017 7517
rect 8975 7455 8989 7475
rect 9009 7455 9017 7475
rect 8975 7417 9017 7455
rect 9091 7475 9133 7517
rect 9091 7455 9099 7475
rect 9119 7455 9133 7475
rect 9091 7417 9133 7455
rect 9183 7475 9227 7517
rect 9183 7455 9195 7475
rect 9215 7455 9227 7475
rect 9183 7417 9227 7455
rect 9299 7475 9341 7517
rect 9299 7455 9307 7475
rect 9327 7455 9341 7475
rect 9299 7417 9341 7455
rect 9391 7475 9435 7517
rect 9391 7455 9403 7475
rect 9423 7455 9435 7475
rect 9391 7417 9435 7455
rect 9512 7475 9554 7517
rect 9512 7455 9520 7475
rect 9540 7455 9554 7475
rect 9512 7417 9554 7455
rect 9604 7475 9648 7517
rect 9604 7455 9616 7475
rect 9636 7455 9648 7475
rect 9604 7417 9648 7455
rect 1387 7225 1431 7263
rect 1387 7205 1399 7225
rect 1419 7205 1431 7225
rect 1387 7163 1431 7205
rect 1481 7225 1523 7263
rect 1481 7205 1495 7225
rect 1515 7205 1523 7225
rect 1481 7163 1523 7205
rect 1600 7225 1644 7263
rect 1600 7205 1612 7225
rect 1632 7205 1644 7225
rect 1600 7163 1644 7205
rect 1694 7225 1736 7263
rect 1694 7205 1708 7225
rect 1728 7205 1736 7225
rect 1694 7163 1736 7205
rect 1808 7225 1852 7263
rect 1808 7205 1820 7225
rect 1840 7205 1852 7225
rect 1808 7163 1852 7205
rect 1902 7225 1944 7263
rect 1902 7205 1916 7225
rect 1936 7205 1944 7225
rect 1902 7163 1944 7205
rect 2018 7225 2060 7263
rect 2018 7205 2026 7225
rect 2046 7205 2060 7225
rect 2018 7163 2060 7205
rect 2110 7232 2155 7263
rect 2110 7225 2154 7232
rect 2110 7205 2122 7225
rect 2142 7205 2154 7225
rect 2110 7163 2154 7205
rect 6443 7266 6487 7304
rect 6443 7246 6455 7266
rect 6475 7246 6487 7266
rect 6443 7204 6487 7246
rect 6537 7266 6579 7304
rect 6537 7246 6551 7266
rect 6571 7246 6579 7266
rect 6537 7204 6579 7246
rect 6656 7266 6700 7304
rect 6656 7246 6668 7266
rect 6688 7246 6700 7266
rect 6656 7204 6700 7246
rect 6750 7266 6792 7304
rect 6750 7246 6764 7266
rect 6784 7246 6792 7266
rect 6750 7204 6792 7246
rect 6864 7266 6908 7304
rect 6864 7246 6876 7266
rect 6896 7246 6908 7266
rect 6864 7204 6908 7246
rect 6958 7266 7000 7304
rect 6958 7246 6972 7266
rect 6992 7246 7000 7266
rect 6958 7204 7000 7246
rect 7074 7266 7116 7304
rect 7074 7246 7082 7266
rect 7102 7246 7116 7266
rect 7074 7204 7116 7246
rect 7166 7273 7211 7304
rect 7166 7266 7210 7273
rect 7166 7246 7178 7266
rect 7198 7246 7210 7266
rect 7166 7204 7210 7246
rect 2777 7154 2821 7196
rect 2777 7134 2789 7154
rect 2809 7134 2821 7154
rect 2777 7127 2821 7134
rect 2776 7096 2821 7127
rect 2871 7154 2913 7196
rect 2871 7134 2885 7154
rect 2905 7134 2913 7154
rect 2871 7096 2913 7134
rect 2987 7154 3029 7196
rect 2987 7134 2995 7154
rect 3015 7134 3029 7154
rect 2987 7096 3029 7134
rect 3079 7154 3123 7196
rect 3079 7134 3091 7154
rect 3111 7134 3123 7154
rect 3079 7096 3123 7134
rect 3195 7154 3237 7196
rect 3195 7134 3203 7154
rect 3223 7134 3237 7154
rect 3195 7096 3237 7134
rect 3287 7154 3331 7196
rect 3287 7134 3299 7154
rect 3319 7134 3331 7154
rect 3287 7096 3331 7134
rect 3408 7154 3450 7196
rect 3408 7134 3416 7154
rect 3436 7134 3450 7154
rect 3408 7096 3450 7134
rect 3500 7154 3544 7196
rect 3500 7134 3512 7154
rect 3532 7134 3544 7154
rect 3500 7096 3544 7134
rect 7833 7195 7877 7237
rect 7833 7175 7845 7195
rect 7865 7175 7877 7195
rect 7833 7168 7877 7175
rect 7832 7137 7877 7168
rect 7927 7195 7969 7237
rect 7927 7175 7941 7195
rect 7961 7175 7969 7195
rect 7927 7137 7969 7175
rect 8043 7195 8085 7237
rect 8043 7175 8051 7195
rect 8071 7175 8085 7195
rect 8043 7137 8085 7175
rect 8135 7195 8179 7237
rect 8135 7175 8147 7195
rect 8167 7175 8179 7195
rect 8135 7137 8179 7175
rect 8251 7195 8293 7237
rect 8251 7175 8259 7195
rect 8279 7175 8293 7195
rect 8251 7137 8293 7175
rect 8343 7195 8387 7237
rect 8343 7175 8355 7195
rect 8375 7175 8387 7195
rect 8343 7137 8387 7175
rect 8464 7195 8506 7237
rect 8464 7175 8472 7195
rect 8492 7175 8506 7195
rect 8464 7137 8506 7175
rect 8556 7195 8600 7237
rect 8556 7175 8568 7195
rect 8588 7175 8600 7195
rect 8556 7137 8600 7175
rect 339 6945 383 6983
rect 339 6925 351 6945
rect 371 6925 383 6945
rect 339 6883 383 6925
rect 433 6945 475 6983
rect 433 6925 447 6945
rect 467 6925 475 6945
rect 433 6883 475 6925
rect 552 6945 596 6983
rect 552 6925 564 6945
rect 584 6925 596 6945
rect 552 6883 596 6925
rect 646 6945 688 6983
rect 646 6925 660 6945
rect 680 6925 688 6945
rect 646 6883 688 6925
rect 760 6945 804 6983
rect 760 6925 772 6945
rect 792 6925 804 6945
rect 760 6883 804 6925
rect 854 6945 896 6983
rect 854 6925 868 6945
rect 888 6925 896 6945
rect 854 6883 896 6925
rect 970 6945 1012 6983
rect 970 6925 978 6945
rect 998 6925 1012 6945
rect 970 6883 1012 6925
rect 1062 6952 1107 6983
rect 1062 6945 1106 6952
rect 1062 6925 1074 6945
rect 1094 6925 1106 6945
rect 5395 6986 5439 7024
rect 5395 6966 5407 6986
rect 5427 6966 5439 6986
rect 1062 6883 1106 6925
rect 3826 6885 3870 6927
rect 3826 6865 3838 6885
rect 3858 6865 3870 6885
rect 3826 6858 3870 6865
rect 3825 6827 3870 6858
rect 3920 6885 3962 6927
rect 3920 6865 3934 6885
rect 3954 6865 3962 6885
rect 3920 6827 3962 6865
rect 4036 6885 4078 6927
rect 4036 6865 4044 6885
rect 4064 6865 4078 6885
rect 4036 6827 4078 6865
rect 4128 6885 4172 6927
rect 4128 6865 4140 6885
rect 4160 6865 4172 6885
rect 4128 6827 4172 6865
rect 4244 6885 4286 6927
rect 4244 6865 4252 6885
rect 4272 6865 4286 6885
rect 4244 6827 4286 6865
rect 4336 6885 4380 6927
rect 4336 6865 4348 6885
rect 4368 6865 4380 6885
rect 4336 6827 4380 6865
rect 4457 6885 4499 6927
rect 4457 6865 4465 6885
rect 4485 6865 4499 6885
rect 4457 6827 4499 6865
rect 4549 6885 4593 6927
rect 5395 6924 5439 6966
rect 5489 6986 5531 7024
rect 5489 6966 5503 6986
rect 5523 6966 5531 6986
rect 5489 6924 5531 6966
rect 5608 6986 5652 7024
rect 5608 6966 5620 6986
rect 5640 6966 5652 6986
rect 5608 6924 5652 6966
rect 5702 6986 5744 7024
rect 5702 6966 5716 6986
rect 5736 6966 5744 6986
rect 5702 6924 5744 6966
rect 5816 6986 5860 7024
rect 5816 6966 5828 6986
rect 5848 6966 5860 6986
rect 5816 6924 5860 6966
rect 5910 6986 5952 7024
rect 5910 6966 5924 6986
rect 5944 6966 5952 6986
rect 5910 6924 5952 6966
rect 6026 6986 6068 7024
rect 6026 6966 6034 6986
rect 6054 6966 6068 6986
rect 6026 6924 6068 6966
rect 6118 6993 6163 7024
rect 6118 6986 6162 6993
rect 6118 6966 6130 6986
rect 6150 6966 6162 6986
rect 6118 6924 6162 6966
rect 8882 6926 8926 6968
rect 4549 6865 4561 6885
rect 4581 6865 4593 6885
rect 4549 6827 4593 6865
rect 8882 6906 8894 6926
rect 8914 6906 8926 6926
rect 8882 6899 8926 6906
rect 8881 6868 8926 6899
rect 8976 6926 9018 6968
rect 8976 6906 8990 6926
rect 9010 6906 9018 6926
rect 8976 6868 9018 6906
rect 9092 6926 9134 6968
rect 9092 6906 9100 6926
rect 9120 6906 9134 6926
rect 9092 6868 9134 6906
rect 9184 6926 9228 6968
rect 9184 6906 9196 6926
rect 9216 6906 9228 6926
rect 9184 6868 9228 6906
rect 9300 6926 9342 6968
rect 9300 6906 9308 6926
rect 9328 6906 9342 6926
rect 9300 6868 9342 6906
rect 9392 6926 9436 6968
rect 9392 6906 9404 6926
rect 9424 6906 9436 6926
rect 9392 6868 9436 6906
rect 9513 6926 9555 6968
rect 9513 6906 9521 6926
rect 9541 6906 9555 6926
rect 9513 6868 9555 6906
rect 9605 6926 9649 6968
rect 9605 6906 9617 6926
rect 9637 6906 9649 6926
rect 9605 6868 9649 6906
rect 1277 6701 1321 6739
rect 1277 6681 1289 6701
rect 1309 6681 1321 6701
rect 1277 6639 1321 6681
rect 1371 6701 1413 6739
rect 1371 6681 1385 6701
rect 1405 6681 1413 6701
rect 1371 6639 1413 6681
rect 1490 6701 1534 6739
rect 1490 6681 1502 6701
rect 1522 6681 1534 6701
rect 1490 6639 1534 6681
rect 1584 6701 1626 6739
rect 1584 6681 1598 6701
rect 1618 6681 1626 6701
rect 1584 6639 1626 6681
rect 1698 6701 1742 6739
rect 1698 6681 1710 6701
rect 1730 6681 1742 6701
rect 1698 6639 1742 6681
rect 1792 6701 1834 6739
rect 1792 6681 1806 6701
rect 1826 6681 1834 6701
rect 1792 6639 1834 6681
rect 1908 6701 1950 6739
rect 1908 6681 1916 6701
rect 1936 6681 1950 6701
rect 1908 6639 1950 6681
rect 2000 6708 2045 6739
rect 2000 6701 2044 6708
rect 2000 6681 2012 6701
rect 2032 6681 2044 6701
rect 2000 6639 2044 6681
rect 6333 6742 6377 6780
rect 6333 6722 6345 6742
rect 6365 6722 6377 6742
rect 2887 6575 2931 6617
rect 2887 6555 2899 6575
rect 2919 6555 2931 6575
rect 2887 6548 2931 6555
rect 2886 6517 2931 6548
rect 2981 6575 3023 6617
rect 2981 6555 2995 6575
rect 3015 6555 3023 6575
rect 2981 6517 3023 6555
rect 3097 6575 3139 6617
rect 3097 6555 3105 6575
rect 3125 6555 3139 6575
rect 3097 6517 3139 6555
rect 3189 6575 3233 6617
rect 3189 6555 3201 6575
rect 3221 6555 3233 6575
rect 3189 6517 3233 6555
rect 3305 6575 3347 6617
rect 3305 6555 3313 6575
rect 3333 6555 3347 6575
rect 3305 6517 3347 6555
rect 3397 6575 3441 6617
rect 3397 6555 3409 6575
rect 3429 6555 3441 6575
rect 3397 6517 3441 6555
rect 3518 6575 3560 6617
rect 3518 6555 3526 6575
rect 3546 6555 3560 6575
rect 3518 6517 3560 6555
rect 3610 6575 3654 6617
rect 6333 6680 6377 6722
rect 6427 6742 6469 6780
rect 6427 6722 6441 6742
rect 6461 6722 6469 6742
rect 6427 6680 6469 6722
rect 6546 6742 6590 6780
rect 6546 6722 6558 6742
rect 6578 6722 6590 6742
rect 6546 6680 6590 6722
rect 6640 6742 6682 6780
rect 6640 6722 6654 6742
rect 6674 6722 6682 6742
rect 6640 6680 6682 6722
rect 6754 6742 6798 6780
rect 6754 6722 6766 6742
rect 6786 6722 6798 6742
rect 6754 6680 6798 6722
rect 6848 6742 6890 6780
rect 6848 6722 6862 6742
rect 6882 6722 6890 6742
rect 6848 6680 6890 6722
rect 6964 6742 7006 6780
rect 6964 6722 6972 6742
rect 6992 6722 7006 6742
rect 6964 6680 7006 6722
rect 7056 6749 7101 6780
rect 7056 6742 7100 6749
rect 7056 6722 7068 6742
rect 7088 6722 7100 6742
rect 7056 6680 7100 6722
rect 3610 6555 3622 6575
rect 3642 6555 3654 6575
rect 3610 6517 3654 6555
rect 7943 6616 7987 6658
rect 7943 6596 7955 6616
rect 7975 6596 7987 6616
rect 7943 6589 7987 6596
rect 7942 6558 7987 6589
rect 8037 6616 8079 6658
rect 8037 6596 8051 6616
rect 8071 6596 8079 6616
rect 8037 6558 8079 6596
rect 8153 6616 8195 6658
rect 8153 6596 8161 6616
rect 8181 6596 8195 6616
rect 8153 6558 8195 6596
rect 8245 6616 8289 6658
rect 8245 6596 8257 6616
rect 8277 6596 8289 6616
rect 8245 6558 8289 6596
rect 8361 6616 8403 6658
rect 8361 6596 8369 6616
rect 8389 6596 8403 6616
rect 8361 6558 8403 6596
rect 8453 6616 8497 6658
rect 8453 6596 8465 6616
rect 8485 6596 8497 6616
rect 8453 6558 8497 6596
rect 8574 6616 8616 6658
rect 8574 6596 8582 6616
rect 8602 6596 8616 6616
rect 8574 6558 8616 6596
rect 8666 6616 8710 6658
rect 8666 6596 8678 6616
rect 8698 6596 8710 6616
rect 8666 6558 8710 6596
rect 338 6391 382 6429
rect 338 6371 350 6391
rect 370 6371 382 6391
rect 338 6329 382 6371
rect 432 6391 474 6429
rect 432 6371 446 6391
rect 466 6371 474 6391
rect 432 6329 474 6371
rect 551 6391 595 6429
rect 551 6371 563 6391
rect 583 6371 595 6391
rect 551 6329 595 6371
rect 645 6391 687 6429
rect 645 6371 659 6391
rect 679 6371 687 6391
rect 645 6329 687 6371
rect 759 6391 803 6429
rect 759 6371 771 6391
rect 791 6371 803 6391
rect 759 6329 803 6371
rect 853 6391 895 6429
rect 853 6371 867 6391
rect 887 6371 895 6391
rect 853 6329 895 6371
rect 969 6391 1011 6429
rect 969 6371 977 6391
rect 997 6371 1011 6391
rect 969 6329 1011 6371
rect 1061 6398 1106 6429
rect 1061 6391 1105 6398
rect 1061 6371 1073 6391
rect 1093 6371 1105 6391
rect 5394 6432 5438 6470
rect 5394 6412 5406 6432
rect 5426 6412 5438 6432
rect 1061 6329 1105 6371
rect 3825 6331 3869 6373
rect 3825 6311 3837 6331
rect 3857 6311 3869 6331
rect 3825 6304 3869 6311
rect 3824 6273 3869 6304
rect 3919 6331 3961 6373
rect 3919 6311 3933 6331
rect 3953 6311 3961 6331
rect 3919 6273 3961 6311
rect 4035 6331 4077 6373
rect 4035 6311 4043 6331
rect 4063 6311 4077 6331
rect 4035 6273 4077 6311
rect 4127 6331 4171 6373
rect 4127 6311 4139 6331
rect 4159 6311 4171 6331
rect 4127 6273 4171 6311
rect 4243 6331 4285 6373
rect 4243 6311 4251 6331
rect 4271 6311 4285 6331
rect 4243 6273 4285 6311
rect 4335 6331 4379 6373
rect 4335 6311 4347 6331
rect 4367 6311 4379 6331
rect 4335 6273 4379 6311
rect 4456 6331 4498 6373
rect 4456 6311 4464 6331
rect 4484 6311 4498 6331
rect 4456 6273 4498 6311
rect 4548 6331 4592 6373
rect 5394 6370 5438 6412
rect 5488 6432 5530 6470
rect 5488 6412 5502 6432
rect 5522 6412 5530 6432
rect 5488 6370 5530 6412
rect 5607 6432 5651 6470
rect 5607 6412 5619 6432
rect 5639 6412 5651 6432
rect 5607 6370 5651 6412
rect 5701 6432 5743 6470
rect 5701 6412 5715 6432
rect 5735 6412 5743 6432
rect 5701 6370 5743 6412
rect 5815 6432 5859 6470
rect 5815 6412 5827 6432
rect 5847 6412 5859 6432
rect 5815 6370 5859 6412
rect 5909 6432 5951 6470
rect 5909 6412 5923 6432
rect 5943 6412 5951 6432
rect 5909 6370 5951 6412
rect 6025 6432 6067 6470
rect 6025 6412 6033 6432
rect 6053 6412 6067 6432
rect 6025 6370 6067 6412
rect 6117 6439 6162 6470
rect 6117 6432 6161 6439
rect 6117 6412 6129 6432
rect 6149 6412 6161 6432
rect 6117 6370 6161 6412
rect 8881 6372 8925 6414
rect 4548 6311 4560 6331
rect 4580 6311 4592 6331
rect 4548 6273 4592 6311
rect 8881 6352 8893 6372
rect 8913 6352 8925 6372
rect 8881 6345 8925 6352
rect 8880 6314 8925 6345
rect 8975 6372 9017 6414
rect 8975 6352 8989 6372
rect 9009 6352 9017 6372
rect 8975 6314 9017 6352
rect 9091 6372 9133 6414
rect 9091 6352 9099 6372
rect 9119 6352 9133 6372
rect 9091 6314 9133 6352
rect 9183 6372 9227 6414
rect 9183 6352 9195 6372
rect 9215 6352 9227 6372
rect 9183 6314 9227 6352
rect 9299 6372 9341 6414
rect 9299 6352 9307 6372
rect 9327 6352 9341 6372
rect 9299 6314 9341 6352
rect 9391 6372 9435 6414
rect 9391 6352 9403 6372
rect 9423 6352 9435 6372
rect 9391 6314 9435 6352
rect 9512 6372 9554 6414
rect 9512 6352 9520 6372
rect 9540 6352 9554 6372
rect 9512 6314 9554 6352
rect 9604 6372 9648 6414
rect 9604 6352 9616 6372
rect 9636 6352 9648 6372
rect 9604 6314 9648 6352
rect 1418 6109 1462 6147
rect 1418 6089 1430 6109
rect 1450 6089 1462 6109
rect 1418 6047 1462 6089
rect 1512 6109 1554 6147
rect 1512 6089 1526 6109
rect 1546 6089 1554 6109
rect 1512 6047 1554 6089
rect 1631 6109 1675 6147
rect 1631 6089 1643 6109
rect 1663 6089 1675 6109
rect 1631 6047 1675 6089
rect 1725 6109 1767 6147
rect 1725 6089 1739 6109
rect 1759 6089 1767 6109
rect 1725 6047 1767 6089
rect 1839 6109 1883 6147
rect 1839 6089 1851 6109
rect 1871 6089 1883 6109
rect 1839 6047 1883 6089
rect 1933 6109 1975 6147
rect 1933 6089 1947 6109
rect 1967 6089 1975 6109
rect 1933 6047 1975 6089
rect 2049 6109 2091 6147
rect 2049 6089 2057 6109
rect 2077 6089 2091 6109
rect 2049 6047 2091 6089
rect 2141 6116 2186 6147
rect 2141 6109 2185 6116
rect 2141 6089 2153 6109
rect 2173 6089 2185 6109
rect 6474 6150 6518 6188
rect 6474 6130 6486 6150
rect 6506 6130 6518 6150
rect 2141 6047 2185 6089
rect 2747 6064 2791 6106
rect 2747 6044 2759 6064
rect 2779 6044 2791 6064
rect 2747 6037 2791 6044
rect 2746 6006 2791 6037
rect 2841 6064 2883 6106
rect 2841 6044 2855 6064
rect 2875 6044 2883 6064
rect 2841 6006 2883 6044
rect 2957 6064 2999 6106
rect 2957 6044 2965 6064
rect 2985 6044 2999 6064
rect 2957 6006 2999 6044
rect 3049 6064 3093 6106
rect 3049 6044 3061 6064
rect 3081 6044 3093 6064
rect 3049 6006 3093 6044
rect 3165 6064 3207 6106
rect 3165 6044 3173 6064
rect 3193 6044 3207 6064
rect 3165 6006 3207 6044
rect 3257 6064 3301 6106
rect 3257 6044 3269 6064
rect 3289 6044 3301 6064
rect 3257 6006 3301 6044
rect 3378 6064 3420 6106
rect 3378 6044 3386 6064
rect 3406 6044 3420 6064
rect 3378 6006 3420 6044
rect 3470 6064 3514 6106
rect 6474 6088 6518 6130
rect 6568 6150 6610 6188
rect 6568 6130 6582 6150
rect 6602 6130 6610 6150
rect 6568 6088 6610 6130
rect 6687 6150 6731 6188
rect 6687 6130 6699 6150
rect 6719 6130 6731 6150
rect 6687 6088 6731 6130
rect 6781 6150 6823 6188
rect 6781 6130 6795 6150
rect 6815 6130 6823 6150
rect 6781 6088 6823 6130
rect 6895 6150 6939 6188
rect 6895 6130 6907 6150
rect 6927 6130 6939 6150
rect 6895 6088 6939 6130
rect 6989 6150 7031 6188
rect 6989 6130 7003 6150
rect 7023 6130 7031 6150
rect 6989 6088 7031 6130
rect 7105 6150 7147 6188
rect 7105 6130 7113 6150
rect 7133 6130 7147 6150
rect 7105 6088 7147 6130
rect 7197 6157 7242 6188
rect 7197 6150 7241 6157
rect 7197 6130 7209 6150
rect 7229 6130 7241 6150
rect 7197 6088 7241 6130
rect 7803 6105 7847 6147
rect 3470 6044 3482 6064
rect 3502 6044 3514 6064
rect 3470 6006 3514 6044
rect 7803 6085 7815 6105
rect 7835 6085 7847 6105
rect 7803 6078 7847 6085
rect 7802 6047 7847 6078
rect 7897 6105 7939 6147
rect 7897 6085 7911 6105
rect 7931 6085 7939 6105
rect 7897 6047 7939 6085
rect 8013 6105 8055 6147
rect 8013 6085 8021 6105
rect 8041 6085 8055 6105
rect 8013 6047 8055 6085
rect 8105 6105 8149 6147
rect 8105 6085 8117 6105
rect 8137 6085 8149 6105
rect 8105 6047 8149 6085
rect 8221 6105 8263 6147
rect 8221 6085 8229 6105
rect 8249 6085 8263 6105
rect 8221 6047 8263 6085
rect 8313 6105 8357 6147
rect 8313 6085 8325 6105
rect 8345 6085 8357 6105
rect 8313 6047 8357 6085
rect 8434 6105 8476 6147
rect 8434 6085 8442 6105
rect 8462 6085 8476 6105
rect 8434 6047 8476 6085
rect 8526 6105 8570 6147
rect 8526 6085 8538 6105
rect 8558 6085 8570 6105
rect 8526 6047 8570 6085
rect 340 5842 384 5880
rect 340 5822 352 5842
rect 372 5822 384 5842
rect 340 5780 384 5822
rect 434 5842 476 5880
rect 434 5822 448 5842
rect 468 5822 476 5842
rect 434 5780 476 5822
rect 553 5842 597 5880
rect 553 5822 565 5842
rect 585 5822 597 5842
rect 553 5780 597 5822
rect 647 5842 689 5880
rect 647 5822 661 5842
rect 681 5822 689 5842
rect 647 5780 689 5822
rect 761 5842 805 5880
rect 761 5822 773 5842
rect 793 5822 805 5842
rect 761 5780 805 5822
rect 855 5842 897 5880
rect 855 5822 869 5842
rect 889 5822 897 5842
rect 855 5780 897 5822
rect 971 5842 1013 5880
rect 971 5822 979 5842
rect 999 5822 1013 5842
rect 971 5780 1013 5822
rect 1063 5849 1108 5880
rect 1063 5842 1107 5849
rect 1063 5822 1075 5842
rect 1095 5822 1107 5842
rect 5396 5883 5440 5921
rect 5396 5863 5408 5883
rect 5428 5863 5440 5883
rect 1063 5780 1107 5822
rect 3827 5782 3871 5824
rect 3827 5762 3839 5782
rect 3859 5762 3871 5782
rect 3827 5755 3871 5762
rect 3826 5724 3871 5755
rect 3921 5782 3963 5824
rect 3921 5762 3935 5782
rect 3955 5762 3963 5782
rect 3921 5724 3963 5762
rect 4037 5782 4079 5824
rect 4037 5762 4045 5782
rect 4065 5762 4079 5782
rect 4037 5724 4079 5762
rect 4129 5782 4173 5824
rect 4129 5762 4141 5782
rect 4161 5762 4173 5782
rect 4129 5724 4173 5762
rect 4245 5782 4287 5824
rect 4245 5762 4253 5782
rect 4273 5762 4287 5782
rect 4245 5724 4287 5762
rect 4337 5782 4381 5824
rect 4337 5762 4349 5782
rect 4369 5762 4381 5782
rect 4337 5724 4381 5762
rect 4458 5782 4500 5824
rect 4458 5762 4466 5782
rect 4486 5762 4500 5782
rect 4458 5724 4500 5762
rect 4550 5782 4594 5824
rect 5396 5821 5440 5863
rect 5490 5883 5532 5921
rect 5490 5863 5504 5883
rect 5524 5863 5532 5883
rect 5490 5821 5532 5863
rect 5609 5883 5653 5921
rect 5609 5863 5621 5883
rect 5641 5863 5653 5883
rect 5609 5821 5653 5863
rect 5703 5883 5745 5921
rect 5703 5863 5717 5883
rect 5737 5863 5745 5883
rect 5703 5821 5745 5863
rect 5817 5883 5861 5921
rect 5817 5863 5829 5883
rect 5849 5863 5861 5883
rect 5817 5821 5861 5863
rect 5911 5883 5953 5921
rect 5911 5863 5925 5883
rect 5945 5863 5953 5883
rect 5911 5821 5953 5863
rect 6027 5883 6069 5921
rect 6027 5863 6035 5883
rect 6055 5863 6069 5883
rect 6027 5821 6069 5863
rect 6119 5890 6164 5921
rect 6119 5883 6163 5890
rect 6119 5863 6131 5883
rect 6151 5863 6163 5883
rect 6119 5821 6163 5863
rect 8883 5823 8927 5865
rect 4550 5762 4562 5782
rect 4582 5762 4594 5782
rect 4550 5724 4594 5762
rect 8883 5803 8895 5823
rect 8915 5803 8927 5823
rect 8883 5796 8927 5803
rect 8882 5765 8927 5796
rect 8977 5823 9019 5865
rect 8977 5803 8991 5823
rect 9011 5803 9019 5823
rect 8977 5765 9019 5803
rect 9093 5823 9135 5865
rect 9093 5803 9101 5823
rect 9121 5803 9135 5823
rect 9093 5765 9135 5803
rect 9185 5823 9229 5865
rect 9185 5803 9197 5823
rect 9217 5803 9229 5823
rect 9185 5765 9229 5803
rect 9301 5823 9343 5865
rect 9301 5803 9309 5823
rect 9329 5803 9343 5823
rect 9301 5765 9343 5803
rect 9393 5823 9437 5865
rect 9393 5803 9405 5823
rect 9425 5803 9437 5823
rect 9393 5765 9437 5803
rect 9514 5823 9556 5865
rect 9514 5803 9522 5823
rect 9542 5803 9556 5823
rect 9514 5765 9556 5803
rect 9606 5823 9650 5865
rect 9606 5803 9618 5823
rect 9638 5803 9650 5823
rect 9606 5765 9650 5803
rect 1278 5598 1322 5636
rect 1278 5578 1290 5598
rect 1310 5578 1322 5598
rect 1278 5536 1322 5578
rect 1372 5598 1414 5636
rect 1372 5578 1386 5598
rect 1406 5578 1414 5598
rect 1372 5536 1414 5578
rect 1491 5598 1535 5636
rect 1491 5578 1503 5598
rect 1523 5578 1535 5598
rect 1491 5536 1535 5578
rect 1585 5598 1627 5636
rect 1585 5578 1599 5598
rect 1619 5578 1627 5598
rect 1585 5536 1627 5578
rect 1699 5598 1743 5636
rect 1699 5578 1711 5598
rect 1731 5578 1743 5598
rect 1699 5536 1743 5578
rect 1793 5598 1835 5636
rect 1793 5578 1807 5598
rect 1827 5578 1835 5598
rect 1793 5536 1835 5578
rect 1909 5598 1951 5636
rect 1909 5578 1917 5598
rect 1937 5578 1951 5598
rect 1909 5536 1951 5578
rect 2001 5605 2046 5636
rect 2001 5598 2045 5605
rect 2001 5578 2013 5598
rect 2033 5578 2045 5598
rect 2001 5536 2045 5578
rect 6334 5639 6378 5677
rect 6334 5619 6346 5639
rect 6366 5619 6378 5639
rect 2888 5472 2932 5514
rect 2888 5452 2900 5472
rect 2920 5452 2932 5472
rect 2888 5445 2932 5452
rect 2887 5414 2932 5445
rect 2982 5472 3024 5514
rect 2982 5452 2996 5472
rect 3016 5452 3024 5472
rect 2982 5414 3024 5452
rect 3098 5472 3140 5514
rect 3098 5452 3106 5472
rect 3126 5452 3140 5472
rect 3098 5414 3140 5452
rect 3190 5472 3234 5514
rect 3190 5452 3202 5472
rect 3222 5452 3234 5472
rect 3190 5414 3234 5452
rect 3306 5472 3348 5514
rect 3306 5452 3314 5472
rect 3334 5452 3348 5472
rect 3306 5414 3348 5452
rect 3398 5472 3442 5514
rect 3398 5452 3410 5472
rect 3430 5452 3442 5472
rect 3398 5414 3442 5452
rect 3519 5472 3561 5514
rect 3519 5452 3527 5472
rect 3547 5452 3561 5472
rect 3519 5414 3561 5452
rect 3611 5472 3655 5514
rect 6334 5577 6378 5619
rect 6428 5639 6470 5677
rect 6428 5619 6442 5639
rect 6462 5619 6470 5639
rect 6428 5577 6470 5619
rect 6547 5639 6591 5677
rect 6547 5619 6559 5639
rect 6579 5619 6591 5639
rect 6547 5577 6591 5619
rect 6641 5639 6683 5677
rect 6641 5619 6655 5639
rect 6675 5619 6683 5639
rect 6641 5577 6683 5619
rect 6755 5639 6799 5677
rect 6755 5619 6767 5639
rect 6787 5619 6799 5639
rect 6755 5577 6799 5619
rect 6849 5639 6891 5677
rect 6849 5619 6863 5639
rect 6883 5619 6891 5639
rect 6849 5577 6891 5619
rect 6965 5639 7007 5677
rect 6965 5619 6973 5639
rect 6993 5619 7007 5639
rect 6965 5577 7007 5619
rect 7057 5646 7102 5677
rect 7057 5639 7101 5646
rect 7057 5619 7069 5639
rect 7089 5619 7101 5639
rect 7057 5577 7101 5619
rect 3611 5452 3623 5472
rect 3643 5452 3655 5472
rect 3611 5414 3655 5452
rect 7944 5513 7988 5555
rect 7944 5493 7956 5513
rect 7976 5493 7988 5513
rect 7944 5486 7988 5493
rect 7943 5455 7988 5486
rect 8038 5513 8080 5555
rect 8038 5493 8052 5513
rect 8072 5493 8080 5513
rect 8038 5455 8080 5493
rect 8154 5513 8196 5555
rect 8154 5493 8162 5513
rect 8182 5493 8196 5513
rect 8154 5455 8196 5493
rect 8246 5513 8290 5555
rect 8246 5493 8258 5513
rect 8278 5493 8290 5513
rect 8246 5455 8290 5493
rect 8362 5513 8404 5555
rect 8362 5493 8370 5513
rect 8390 5493 8404 5513
rect 8362 5455 8404 5493
rect 8454 5513 8498 5555
rect 8454 5493 8466 5513
rect 8486 5493 8498 5513
rect 8454 5455 8498 5493
rect 8575 5513 8617 5555
rect 8575 5493 8583 5513
rect 8603 5493 8617 5513
rect 8575 5455 8617 5493
rect 8667 5513 8711 5555
rect 8667 5493 8679 5513
rect 8699 5493 8711 5513
rect 8667 5455 8711 5493
rect 339 5288 383 5326
rect 339 5268 351 5288
rect 371 5268 383 5288
rect 339 5226 383 5268
rect 433 5288 475 5326
rect 433 5268 447 5288
rect 467 5268 475 5288
rect 433 5226 475 5268
rect 552 5288 596 5326
rect 552 5268 564 5288
rect 584 5268 596 5288
rect 552 5226 596 5268
rect 646 5288 688 5326
rect 646 5268 660 5288
rect 680 5268 688 5288
rect 646 5226 688 5268
rect 760 5288 804 5326
rect 760 5268 772 5288
rect 792 5268 804 5288
rect 760 5226 804 5268
rect 854 5288 896 5326
rect 854 5268 868 5288
rect 888 5268 896 5288
rect 854 5226 896 5268
rect 970 5288 1012 5326
rect 970 5268 978 5288
rect 998 5268 1012 5288
rect 970 5226 1012 5268
rect 1062 5295 1107 5326
rect 1062 5288 1106 5295
rect 1062 5268 1074 5288
rect 1094 5268 1106 5288
rect 5395 5329 5439 5367
rect 5395 5309 5407 5329
rect 5427 5309 5439 5329
rect 1062 5226 1106 5268
rect 3826 5228 3870 5270
rect 3826 5208 3838 5228
rect 3858 5208 3870 5228
rect 3826 5201 3870 5208
rect 3825 5170 3870 5201
rect 3920 5228 3962 5270
rect 3920 5208 3934 5228
rect 3954 5208 3962 5228
rect 3920 5170 3962 5208
rect 4036 5228 4078 5270
rect 4036 5208 4044 5228
rect 4064 5208 4078 5228
rect 4036 5170 4078 5208
rect 4128 5228 4172 5270
rect 4128 5208 4140 5228
rect 4160 5208 4172 5228
rect 4128 5170 4172 5208
rect 4244 5228 4286 5270
rect 4244 5208 4252 5228
rect 4272 5208 4286 5228
rect 4244 5170 4286 5208
rect 4336 5228 4380 5270
rect 4336 5208 4348 5228
rect 4368 5208 4380 5228
rect 4336 5170 4380 5208
rect 4457 5228 4499 5270
rect 4457 5208 4465 5228
rect 4485 5208 4499 5228
rect 4457 5170 4499 5208
rect 4549 5228 4593 5270
rect 5395 5267 5439 5309
rect 5489 5329 5531 5367
rect 5489 5309 5503 5329
rect 5523 5309 5531 5329
rect 5489 5267 5531 5309
rect 5608 5329 5652 5367
rect 5608 5309 5620 5329
rect 5640 5309 5652 5329
rect 5608 5267 5652 5309
rect 5702 5329 5744 5367
rect 5702 5309 5716 5329
rect 5736 5309 5744 5329
rect 5702 5267 5744 5309
rect 5816 5329 5860 5367
rect 5816 5309 5828 5329
rect 5848 5309 5860 5329
rect 5816 5267 5860 5309
rect 5910 5329 5952 5367
rect 5910 5309 5924 5329
rect 5944 5309 5952 5329
rect 5910 5267 5952 5309
rect 6026 5329 6068 5367
rect 6026 5309 6034 5329
rect 6054 5309 6068 5329
rect 6026 5267 6068 5309
rect 6118 5336 6163 5367
rect 6118 5329 6162 5336
rect 6118 5309 6130 5329
rect 6150 5309 6162 5329
rect 6118 5267 6162 5309
rect 8882 5269 8926 5311
rect 4549 5208 4561 5228
rect 4581 5208 4593 5228
rect 4549 5170 4593 5208
rect 8882 5249 8894 5269
rect 8914 5249 8926 5269
rect 8882 5242 8926 5249
rect 8881 5211 8926 5242
rect 8976 5269 9018 5311
rect 8976 5249 8990 5269
rect 9010 5249 9018 5269
rect 8976 5211 9018 5249
rect 9092 5269 9134 5311
rect 9092 5249 9100 5269
rect 9120 5249 9134 5269
rect 9092 5211 9134 5249
rect 9184 5269 9228 5311
rect 9184 5249 9196 5269
rect 9216 5249 9228 5269
rect 9184 5211 9228 5249
rect 9300 5269 9342 5311
rect 9300 5249 9308 5269
rect 9328 5249 9342 5269
rect 9300 5211 9342 5249
rect 9392 5269 9436 5311
rect 9392 5249 9404 5269
rect 9424 5249 9436 5269
rect 9392 5211 9436 5249
rect 9513 5269 9555 5311
rect 9513 5249 9521 5269
rect 9541 5249 9555 5269
rect 9513 5211 9555 5249
rect 9605 5269 9649 5311
rect 9605 5249 9617 5269
rect 9637 5249 9649 5269
rect 9605 5211 9649 5249
rect 1387 5025 1431 5063
rect 1387 5005 1399 5025
rect 1419 5005 1431 5025
rect 1387 4963 1431 5005
rect 1481 5025 1523 5063
rect 1481 5005 1495 5025
rect 1515 5005 1523 5025
rect 1481 4963 1523 5005
rect 1600 5025 1644 5063
rect 1600 5005 1612 5025
rect 1632 5005 1644 5025
rect 1600 4963 1644 5005
rect 1694 5025 1736 5063
rect 1694 5005 1708 5025
rect 1728 5005 1736 5025
rect 1694 4963 1736 5005
rect 1808 5025 1852 5063
rect 1808 5005 1820 5025
rect 1840 5005 1852 5025
rect 1808 4963 1852 5005
rect 1902 5025 1944 5063
rect 1902 5005 1916 5025
rect 1936 5005 1944 5025
rect 1902 4963 1944 5005
rect 2018 5025 2060 5063
rect 2018 5005 2026 5025
rect 2046 5005 2060 5025
rect 2018 4963 2060 5005
rect 2110 5032 2155 5063
rect 2110 5025 2154 5032
rect 2110 5005 2122 5025
rect 2142 5005 2154 5025
rect 2110 4963 2154 5005
rect 6443 5066 6487 5104
rect 6443 5046 6455 5066
rect 6475 5046 6487 5066
rect 6443 5004 6487 5046
rect 6537 5066 6579 5104
rect 6537 5046 6551 5066
rect 6571 5046 6579 5066
rect 6537 5004 6579 5046
rect 6656 5066 6700 5104
rect 6656 5046 6668 5066
rect 6688 5046 6700 5066
rect 6656 5004 6700 5046
rect 6750 5066 6792 5104
rect 6750 5046 6764 5066
rect 6784 5046 6792 5066
rect 6750 5004 6792 5046
rect 6864 5066 6908 5104
rect 6864 5046 6876 5066
rect 6896 5046 6908 5066
rect 6864 5004 6908 5046
rect 6958 5066 7000 5104
rect 6958 5046 6972 5066
rect 6992 5046 7000 5066
rect 6958 5004 7000 5046
rect 7074 5066 7116 5104
rect 7074 5046 7082 5066
rect 7102 5046 7116 5066
rect 7074 5004 7116 5046
rect 7166 5073 7211 5104
rect 7166 5066 7210 5073
rect 7166 5046 7178 5066
rect 7198 5046 7210 5066
rect 7166 5004 7210 5046
rect 2779 4942 2823 4984
rect 2779 4922 2791 4942
rect 2811 4922 2823 4942
rect 2779 4915 2823 4922
rect 2778 4884 2823 4915
rect 2873 4942 2915 4984
rect 2873 4922 2887 4942
rect 2907 4922 2915 4942
rect 2873 4884 2915 4922
rect 2989 4942 3031 4984
rect 2989 4922 2997 4942
rect 3017 4922 3031 4942
rect 2989 4884 3031 4922
rect 3081 4942 3125 4984
rect 3081 4922 3093 4942
rect 3113 4922 3125 4942
rect 3081 4884 3125 4922
rect 3197 4942 3239 4984
rect 3197 4922 3205 4942
rect 3225 4922 3239 4942
rect 3197 4884 3239 4922
rect 3289 4942 3333 4984
rect 3289 4922 3301 4942
rect 3321 4922 3333 4942
rect 3289 4884 3333 4922
rect 3410 4942 3452 4984
rect 3410 4922 3418 4942
rect 3438 4922 3452 4942
rect 3410 4884 3452 4922
rect 3502 4942 3546 4984
rect 3502 4922 3514 4942
rect 3534 4922 3546 4942
rect 3502 4884 3546 4922
rect 7835 4983 7879 5025
rect 7835 4963 7847 4983
rect 7867 4963 7879 4983
rect 7835 4956 7879 4963
rect 7834 4925 7879 4956
rect 7929 4983 7971 5025
rect 7929 4963 7943 4983
rect 7963 4963 7971 4983
rect 7929 4925 7971 4963
rect 8045 4983 8087 5025
rect 8045 4963 8053 4983
rect 8073 4963 8087 4983
rect 8045 4925 8087 4963
rect 8137 4983 8181 5025
rect 8137 4963 8149 4983
rect 8169 4963 8181 4983
rect 8137 4925 8181 4963
rect 8253 4983 8295 5025
rect 8253 4963 8261 4983
rect 8281 4963 8295 4983
rect 8253 4925 8295 4963
rect 8345 4983 8389 5025
rect 8345 4963 8357 4983
rect 8377 4963 8389 4983
rect 8345 4925 8389 4963
rect 8466 4983 8508 5025
rect 8466 4963 8474 4983
rect 8494 4963 8508 4983
rect 8466 4925 8508 4963
rect 8558 4983 8602 5025
rect 8558 4963 8570 4983
rect 8590 4963 8602 4983
rect 8558 4925 8602 4963
rect 340 4739 384 4777
rect 340 4719 352 4739
rect 372 4719 384 4739
rect 340 4677 384 4719
rect 434 4739 476 4777
rect 434 4719 448 4739
rect 468 4719 476 4739
rect 434 4677 476 4719
rect 553 4739 597 4777
rect 553 4719 565 4739
rect 585 4719 597 4739
rect 553 4677 597 4719
rect 647 4739 689 4777
rect 647 4719 661 4739
rect 681 4719 689 4739
rect 647 4677 689 4719
rect 761 4739 805 4777
rect 761 4719 773 4739
rect 793 4719 805 4739
rect 761 4677 805 4719
rect 855 4739 897 4777
rect 855 4719 869 4739
rect 889 4719 897 4739
rect 855 4677 897 4719
rect 971 4739 1013 4777
rect 971 4719 979 4739
rect 999 4719 1013 4739
rect 971 4677 1013 4719
rect 1063 4746 1108 4777
rect 1063 4739 1107 4746
rect 1063 4719 1075 4739
rect 1095 4719 1107 4739
rect 5396 4780 5440 4818
rect 5396 4760 5408 4780
rect 5428 4760 5440 4780
rect 1063 4677 1107 4719
rect 3827 4679 3871 4721
rect 3827 4659 3839 4679
rect 3859 4659 3871 4679
rect 3827 4652 3871 4659
rect 3826 4621 3871 4652
rect 3921 4679 3963 4721
rect 3921 4659 3935 4679
rect 3955 4659 3963 4679
rect 3921 4621 3963 4659
rect 4037 4679 4079 4721
rect 4037 4659 4045 4679
rect 4065 4659 4079 4679
rect 4037 4621 4079 4659
rect 4129 4679 4173 4721
rect 4129 4659 4141 4679
rect 4161 4659 4173 4679
rect 4129 4621 4173 4659
rect 4245 4679 4287 4721
rect 4245 4659 4253 4679
rect 4273 4659 4287 4679
rect 4245 4621 4287 4659
rect 4337 4679 4381 4721
rect 4337 4659 4349 4679
rect 4369 4659 4381 4679
rect 4337 4621 4381 4659
rect 4458 4679 4500 4721
rect 4458 4659 4466 4679
rect 4486 4659 4500 4679
rect 4458 4621 4500 4659
rect 4550 4679 4594 4721
rect 5396 4718 5440 4760
rect 5490 4780 5532 4818
rect 5490 4760 5504 4780
rect 5524 4760 5532 4780
rect 5490 4718 5532 4760
rect 5609 4780 5653 4818
rect 5609 4760 5621 4780
rect 5641 4760 5653 4780
rect 5609 4718 5653 4760
rect 5703 4780 5745 4818
rect 5703 4760 5717 4780
rect 5737 4760 5745 4780
rect 5703 4718 5745 4760
rect 5817 4780 5861 4818
rect 5817 4760 5829 4780
rect 5849 4760 5861 4780
rect 5817 4718 5861 4760
rect 5911 4780 5953 4818
rect 5911 4760 5925 4780
rect 5945 4760 5953 4780
rect 5911 4718 5953 4760
rect 6027 4780 6069 4818
rect 6027 4760 6035 4780
rect 6055 4760 6069 4780
rect 6027 4718 6069 4760
rect 6119 4787 6164 4818
rect 6119 4780 6163 4787
rect 6119 4760 6131 4780
rect 6151 4760 6163 4780
rect 6119 4718 6163 4760
rect 8883 4720 8927 4762
rect 4550 4659 4562 4679
rect 4582 4659 4594 4679
rect 4550 4621 4594 4659
rect 8883 4700 8895 4720
rect 8915 4700 8927 4720
rect 8883 4693 8927 4700
rect 8882 4662 8927 4693
rect 8977 4720 9019 4762
rect 8977 4700 8991 4720
rect 9011 4700 9019 4720
rect 8977 4662 9019 4700
rect 9093 4720 9135 4762
rect 9093 4700 9101 4720
rect 9121 4700 9135 4720
rect 9093 4662 9135 4700
rect 9185 4720 9229 4762
rect 9185 4700 9197 4720
rect 9217 4700 9229 4720
rect 9185 4662 9229 4700
rect 9301 4720 9343 4762
rect 9301 4700 9309 4720
rect 9329 4700 9343 4720
rect 9301 4662 9343 4700
rect 9393 4720 9437 4762
rect 9393 4700 9405 4720
rect 9425 4700 9437 4720
rect 9393 4662 9437 4700
rect 9514 4720 9556 4762
rect 9514 4700 9522 4720
rect 9542 4700 9556 4720
rect 9514 4662 9556 4700
rect 9606 4720 9650 4762
rect 9606 4700 9618 4720
rect 9638 4700 9650 4720
rect 9606 4662 9650 4700
rect 1278 4495 1322 4533
rect 1278 4475 1290 4495
rect 1310 4475 1322 4495
rect 1278 4433 1322 4475
rect 1372 4495 1414 4533
rect 1372 4475 1386 4495
rect 1406 4475 1414 4495
rect 1372 4433 1414 4475
rect 1491 4495 1535 4533
rect 1491 4475 1503 4495
rect 1523 4475 1535 4495
rect 1491 4433 1535 4475
rect 1585 4495 1627 4533
rect 1585 4475 1599 4495
rect 1619 4475 1627 4495
rect 1585 4433 1627 4475
rect 1699 4495 1743 4533
rect 1699 4475 1711 4495
rect 1731 4475 1743 4495
rect 1699 4433 1743 4475
rect 1793 4495 1835 4533
rect 1793 4475 1807 4495
rect 1827 4475 1835 4495
rect 1793 4433 1835 4475
rect 1909 4495 1951 4533
rect 1909 4475 1917 4495
rect 1937 4475 1951 4495
rect 1909 4433 1951 4475
rect 2001 4502 2046 4533
rect 2001 4495 2045 4502
rect 2001 4475 2013 4495
rect 2033 4475 2045 4495
rect 2001 4433 2045 4475
rect 6334 4536 6378 4574
rect 6334 4516 6346 4536
rect 6366 4516 6378 4536
rect 2888 4369 2932 4411
rect 2888 4349 2900 4369
rect 2920 4349 2932 4369
rect 2888 4342 2932 4349
rect 2887 4311 2932 4342
rect 2982 4369 3024 4411
rect 2982 4349 2996 4369
rect 3016 4349 3024 4369
rect 2982 4311 3024 4349
rect 3098 4369 3140 4411
rect 3098 4349 3106 4369
rect 3126 4349 3140 4369
rect 3098 4311 3140 4349
rect 3190 4369 3234 4411
rect 3190 4349 3202 4369
rect 3222 4349 3234 4369
rect 3190 4311 3234 4349
rect 3306 4369 3348 4411
rect 3306 4349 3314 4369
rect 3334 4349 3348 4369
rect 3306 4311 3348 4349
rect 3398 4369 3442 4411
rect 3398 4349 3410 4369
rect 3430 4349 3442 4369
rect 3398 4311 3442 4349
rect 3519 4369 3561 4411
rect 3519 4349 3527 4369
rect 3547 4349 3561 4369
rect 3519 4311 3561 4349
rect 3611 4369 3655 4411
rect 6334 4474 6378 4516
rect 6428 4536 6470 4574
rect 6428 4516 6442 4536
rect 6462 4516 6470 4536
rect 6428 4474 6470 4516
rect 6547 4536 6591 4574
rect 6547 4516 6559 4536
rect 6579 4516 6591 4536
rect 6547 4474 6591 4516
rect 6641 4536 6683 4574
rect 6641 4516 6655 4536
rect 6675 4516 6683 4536
rect 6641 4474 6683 4516
rect 6755 4536 6799 4574
rect 6755 4516 6767 4536
rect 6787 4516 6799 4536
rect 6755 4474 6799 4516
rect 6849 4536 6891 4574
rect 6849 4516 6863 4536
rect 6883 4516 6891 4536
rect 6849 4474 6891 4516
rect 6965 4536 7007 4574
rect 6965 4516 6973 4536
rect 6993 4516 7007 4536
rect 6965 4474 7007 4516
rect 7057 4543 7102 4574
rect 7057 4536 7101 4543
rect 7057 4516 7069 4536
rect 7089 4516 7101 4536
rect 7057 4474 7101 4516
rect 3611 4349 3623 4369
rect 3643 4349 3655 4369
rect 3611 4311 3655 4349
rect 7944 4410 7988 4452
rect 7944 4390 7956 4410
rect 7976 4390 7988 4410
rect 7944 4383 7988 4390
rect 7943 4352 7988 4383
rect 8038 4410 8080 4452
rect 8038 4390 8052 4410
rect 8072 4390 8080 4410
rect 8038 4352 8080 4390
rect 8154 4410 8196 4452
rect 8154 4390 8162 4410
rect 8182 4390 8196 4410
rect 8154 4352 8196 4390
rect 8246 4410 8290 4452
rect 8246 4390 8258 4410
rect 8278 4390 8290 4410
rect 8246 4352 8290 4390
rect 8362 4410 8404 4452
rect 8362 4390 8370 4410
rect 8390 4390 8404 4410
rect 8362 4352 8404 4390
rect 8454 4410 8498 4452
rect 8454 4390 8466 4410
rect 8486 4390 8498 4410
rect 8454 4352 8498 4390
rect 8575 4410 8617 4452
rect 8575 4390 8583 4410
rect 8603 4390 8617 4410
rect 8575 4352 8617 4390
rect 8667 4410 8711 4452
rect 8667 4390 8679 4410
rect 8699 4390 8711 4410
rect 8667 4352 8711 4390
rect 339 4185 383 4223
rect 339 4165 351 4185
rect 371 4165 383 4185
rect 339 4123 383 4165
rect 433 4185 475 4223
rect 433 4165 447 4185
rect 467 4165 475 4185
rect 433 4123 475 4165
rect 552 4185 596 4223
rect 552 4165 564 4185
rect 584 4165 596 4185
rect 552 4123 596 4165
rect 646 4185 688 4223
rect 646 4165 660 4185
rect 680 4165 688 4185
rect 646 4123 688 4165
rect 760 4185 804 4223
rect 760 4165 772 4185
rect 792 4165 804 4185
rect 760 4123 804 4165
rect 854 4185 896 4223
rect 854 4165 868 4185
rect 888 4165 896 4185
rect 854 4123 896 4165
rect 970 4185 1012 4223
rect 970 4165 978 4185
rect 998 4165 1012 4185
rect 970 4123 1012 4165
rect 1062 4192 1107 4223
rect 1062 4185 1106 4192
rect 1062 4165 1074 4185
rect 1094 4165 1106 4185
rect 5395 4226 5439 4264
rect 5395 4206 5407 4226
rect 5427 4206 5439 4226
rect 1062 4123 1106 4165
rect 3826 4125 3870 4167
rect 3826 4105 3838 4125
rect 3858 4105 3870 4125
rect 3826 4098 3870 4105
rect 3825 4067 3870 4098
rect 3920 4125 3962 4167
rect 3920 4105 3934 4125
rect 3954 4105 3962 4125
rect 3920 4067 3962 4105
rect 4036 4125 4078 4167
rect 4036 4105 4044 4125
rect 4064 4105 4078 4125
rect 4036 4067 4078 4105
rect 4128 4125 4172 4167
rect 4128 4105 4140 4125
rect 4160 4105 4172 4125
rect 4128 4067 4172 4105
rect 4244 4125 4286 4167
rect 4244 4105 4252 4125
rect 4272 4105 4286 4125
rect 4244 4067 4286 4105
rect 4336 4125 4380 4167
rect 4336 4105 4348 4125
rect 4368 4105 4380 4125
rect 4336 4067 4380 4105
rect 4457 4125 4499 4167
rect 4457 4105 4465 4125
rect 4485 4105 4499 4125
rect 4457 4067 4499 4105
rect 4549 4125 4593 4167
rect 5395 4164 5439 4206
rect 5489 4226 5531 4264
rect 5489 4206 5503 4226
rect 5523 4206 5531 4226
rect 5489 4164 5531 4206
rect 5608 4226 5652 4264
rect 5608 4206 5620 4226
rect 5640 4206 5652 4226
rect 5608 4164 5652 4206
rect 5702 4226 5744 4264
rect 5702 4206 5716 4226
rect 5736 4206 5744 4226
rect 5702 4164 5744 4206
rect 5816 4226 5860 4264
rect 5816 4206 5828 4226
rect 5848 4206 5860 4226
rect 5816 4164 5860 4206
rect 5910 4226 5952 4264
rect 5910 4206 5924 4226
rect 5944 4206 5952 4226
rect 5910 4164 5952 4206
rect 6026 4226 6068 4264
rect 6026 4206 6034 4226
rect 6054 4206 6068 4226
rect 6026 4164 6068 4206
rect 6118 4233 6163 4264
rect 6118 4226 6162 4233
rect 6118 4206 6130 4226
rect 6150 4206 6162 4226
rect 6118 4164 6162 4206
rect 8882 4166 8926 4208
rect 4549 4105 4561 4125
rect 4581 4105 4593 4125
rect 4549 4067 4593 4105
rect 8882 4146 8894 4166
rect 8914 4146 8926 4166
rect 8882 4139 8926 4146
rect 8881 4108 8926 4139
rect 8976 4166 9018 4208
rect 8976 4146 8990 4166
rect 9010 4146 9018 4166
rect 8976 4108 9018 4146
rect 9092 4166 9134 4208
rect 9092 4146 9100 4166
rect 9120 4146 9134 4166
rect 9092 4108 9134 4146
rect 9184 4166 9228 4208
rect 9184 4146 9196 4166
rect 9216 4146 9228 4166
rect 9184 4108 9228 4146
rect 9300 4166 9342 4208
rect 9300 4146 9308 4166
rect 9328 4146 9342 4166
rect 9300 4108 9342 4146
rect 9392 4166 9436 4208
rect 9392 4146 9404 4166
rect 9424 4146 9436 4166
rect 9392 4108 9436 4146
rect 9513 4166 9555 4208
rect 9513 4146 9521 4166
rect 9541 4146 9555 4166
rect 9513 4108 9555 4146
rect 9605 4166 9649 4208
rect 9605 4146 9617 4166
rect 9637 4146 9649 4166
rect 9605 4108 9649 4146
rect 1419 3903 1463 3941
rect 1419 3883 1431 3903
rect 1451 3883 1463 3903
rect 1419 3841 1463 3883
rect 1513 3903 1555 3941
rect 1513 3883 1527 3903
rect 1547 3883 1555 3903
rect 1513 3841 1555 3883
rect 1632 3903 1676 3941
rect 1632 3883 1644 3903
rect 1664 3883 1676 3903
rect 1632 3841 1676 3883
rect 1726 3903 1768 3941
rect 1726 3883 1740 3903
rect 1760 3883 1768 3903
rect 1726 3841 1768 3883
rect 1840 3903 1884 3941
rect 1840 3883 1852 3903
rect 1872 3883 1884 3903
rect 1840 3841 1884 3883
rect 1934 3903 1976 3941
rect 1934 3883 1948 3903
rect 1968 3883 1976 3903
rect 1934 3841 1976 3883
rect 2050 3903 2092 3941
rect 2050 3883 2058 3903
rect 2078 3883 2092 3903
rect 2050 3841 2092 3883
rect 2142 3910 2187 3941
rect 2142 3903 2186 3910
rect 2142 3883 2154 3903
rect 2174 3883 2186 3903
rect 6475 3944 6519 3982
rect 6475 3924 6487 3944
rect 6507 3924 6519 3944
rect 2142 3841 2186 3883
rect 2748 3858 2792 3900
rect 2748 3838 2760 3858
rect 2780 3838 2792 3858
rect 2748 3831 2792 3838
rect 2747 3800 2792 3831
rect 2842 3858 2884 3900
rect 2842 3838 2856 3858
rect 2876 3838 2884 3858
rect 2842 3800 2884 3838
rect 2958 3858 3000 3900
rect 2958 3838 2966 3858
rect 2986 3838 3000 3858
rect 2958 3800 3000 3838
rect 3050 3858 3094 3900
rect 3050 3838 3062 3858
rect 3082 3838 3094 3858
rect 3050 3800 3094 3838
rect 3166 3858 3208 3900
rect 3166 3838 3174 3858
rect 3194 3838 3208 3858
rect 3166 3800 3208 3838
rect 3258 3858 3302 3900
rect 3258 3838 3270 3858
rect 3290 3838 3302 3858
rect 3258 3800 3302 3838
rect 3379 3858 3421 3900
rect 3379 3838 3387 3858
rect 3407 3838 3421 3858
rect 3379 3800 3421 3838
rect 3471 3858 3515 3900
rect 6475 3882 6519 3924
rect 6569 3944 6611 3982
rect 6569 3924 6583 3944
rect 6603 3924 6611 3944
rect 6569 3882 6611 3924
rect 6688 3944 6732 3982
rect 6688 3924 6700 3944
rect 6720 3924 6732 3944
rect 6688 3882 6732 3924
rect 6782 3944 6824 3982
rect 6782 3924 6796 3944
rect 6816 3924 6824 3944
rect 6782 3882 6824 3924
rect 6896 3944 6940 3982
rect 6896 3924 6908 3944
rect 6928 3924 6940 3944
rect 6896 3882 6940 3924
rect 6990 3944 7032 3982
rect 6990 3924 7004 3944
rect 7024 3924 7032 3944
rect 6990 3882 7032 3924
rect 7106 3944 7148 3982
rect 7106 3924 7114 3944
rect 7134 3924 7148 3944
rect 7106 3882 7148 3924
rect 7198 3951 7243 3982
rect 7198 3944 7242 3951
rect 7198 3924 7210 3944
rect 7230 3924 7242 3944
rect 7198 3882 7242 3924
rect 7804 3899 7848 3941
rect 3471 3838 3483 3858
rect 3503 3838 3515 3858
rect 3471 3800 3515 3838
rect 7804 3879 7816 3899
rect 7836 3879 7848 3899
rect 7804 3872 7848 3879
rect 7803 3841 7848 3872
rect 7898 3899 7940 3941
rect 7898 3879 7912 3899
rect 7932 3879 7940 3899
rect 7898 3841 7940 3879
rect 8014 3899 8056 3941
rect 8014 3879 8022 3899
rect 8042 3879 8056 3899
rect 8014 3841 8056 3879
rect 8106 3899 8150 3941
rect 8106 3879 8118 3899
rect 8138 3879 8150 3899
rect 8106 3841 8150 3879
rect 8222 3899 8264 3941
rect 8222 3879 8230 3899
rect 8250 3879 8264 3899
rect 8222 3841 8264 3879
rect 8314 3899 8358 3941
rect 8314 3879 8326 3899
rect 8346 3879 8358 3899
rect 8314 3841 8358 3879
rect 8435 3899 8477 3941
rect 8435 3879 8443 3899
rect 8463 3879 8477 3899
rect 8435 3841 8477 3879
rect 8527 3899 8571 3941
rect 8527 3879 8539 3899
rect 8559 3879 8571 3899
rect 8527 3841 8571 3879
rect 341 3636 385 3674
rect 341 3616 353 3636
rect 373 3616 385 3636
rect 341 3574 385 3616
rect 435 3636 477 3674
rect 435 3616 449 3636
rect 469 3616 477 3636
rect 435 3574 477 3616
rect 554 3636 598 3674
rect 554 3616 566 3636
rect 586 3616 598 3636
rect 554 3574 598 3616
rect 648 3636 690 3674
rect 648 3616 662 3636
rect 682 3616 690 3636
rect 648 3574 690 3616
rect 762 3636 806 3674
rect 762 3616 774 3636
rect 794 3616 806 3636
rect 762 3574 806 3616
rect 856 3636 898 3674
rect 856 3616 870 3636
rect 890 3616 898 3636
rect 856 3574 898 3616
rect 972 3636 1014 3674
rect 972 3616 980 3636
rect 1000 3616 1014 3636
rect 972 3574 1014 3616
rect 1064 3643 1109 3674
rect 1064 3636 1108 3643
rect 1064 3616 1076 3636
rect 1096 3616 1108 3636
rect 5397 3677 5441 3715
rect 5397 3657 5409 3677
rect 5429 3657 5441 3677
rect 1064 3574 1108 3616
rect 3828 3576 3872 3618
rect 3828 3556 3840 3576
rect 3860 3556 3872 3576
rect 3828 3549 3872 3556
rect 3827 3518 3872 3549
rect 3922 3576 3964 3618
rect 3922 3556 3936 3576
rect 3956 3556 3964 3576
rect 3922 3518 3964 3556
rect 4038 3576 4080 3618
rect 4038 3556 4046 3576
rect 4066 3556 4080 3576
rect 4038 3518 4080 3556
rect 4130 3576 4174 3618
rect 4130 3556 4142 3576
rect 4162 3556 4174 3576
rect 4130 3518 4174 3556
rect 4246 3576 4288 3618
rect 4246 3556 4254 3576
rect 4274 3556 4288 3576
rect 4246 3518 4288 3556
rect 4338 3576 4382 3618
rect 4338 3556 4350 3576
rect 4370 3556 4382 3576
rect 4338 3518 4382 3556
rect 4459 3576 4501 3618
rect 4459 3556 4467 3576
rect 4487 3556 4501 3576
rect 4459 3518 4501 3556
rect 4551 3576 4595 3618
rect 5397 3615 5441 3657
rect 5491 3677 5533 3715
rect 5491 3657 5505 3677
rect 5525 3657 5533 3677
rect 5491 3615 5533 3657
rect 5610 3677 5654 3715
rect 5610 3657 5622 3677
rect 5642 3657 5654 3677
rect 5610 3615 5654 3657
rect 5704 3677 5746 3715
rect 5704 3657 5718 3677
rect 5738 3657 5746 3677
rect 5704 3615 5746 3657
rect 5818 3677 5862 3715
rect 5818 3657 5830 3677
rect 5850 3657 5862 3677
rect 5818 3615 5862 3657
rect 5912 3677 5954 3715
rect 5912 3657 5926 3677
rect 5946 3657 5954 3677
rect 5912 3615 5954 3657
rect 6028 3677 6070 3715
rect 6028 3657 6036 3677
rect 6056 3657 6070 3677
rect 6028 3615 6070 3657
rect 6120 3684 6165 3715
rect 6120 3677 6164 3684
rect 6120 3657 6132 3677
rect 6152 3657 6164 3677
rect 6120 3615 6164 3657
rect 8884 3617 8928 3659
rect 4551 3556 4563 3576
rect 4583 3556 4595 3576
rect 4551 3518 4595 3556
rect 8884 3597 8896 3617
rect 8916 3597 8928 3617
rect 8884 3590 8928 3597
rect 8883 3559 8928 3590
rect 8978 3617 9020 3659
rect 8978 3597 8992 3617
rect 9012 3597 9020 3617
rect 8978 3559 9020 3597
rect 9094 3617 9136 3659
rect 9094 3597 9102 3617
rect 9122 3597 9136 3617
rect 9094 3559 9136 3597
rect 9186 3617 9230 3659
rect 9186 3597 9198 3617
rect 9218 3597 9230 3617
rect 9186 3559 9230 3597
rect 9302 3617 9344 3659
rect 9302 3597 9310 3617
rect 9330 3597 9344 3617
rect 9302 3559 9344 3597
rect 9394 3617 9438 3659
rect 9394 3597 9406 3617
rect 9426 3597 9438 3617
rect 9394 3559 9438 3597
rect 9515 3617 9557 3659
rect 9515 3597 9523 3617
rect 9543 3597 9557 3617
rect 9515 3559 9557 3597
rect 9607 3617 9651 3659
rect 9607 3597 9619 3617
rect 9639 3597 9651 3617
rect 9607 3559 9651 3597
rect 1279 3392 1323 3430
rect 1279 3372 1291 3392
rect 1311 3372 1323 3392
rect 1279 3330 1323 3372
rect 1373 3392 1415 3430
rect 1373 3372 1387 3392
rect 1407 3372 1415 3392
rect 1373 3330 1415 3372
rect 1492 3392 1536 3430
rect 1492 3372 1504 3392
rect 1524 3372 1536 3392
rect 1492 3330 1536 3372
rect 1586 3392 1628 3430
rect 1586 3372 1600 3392
rect 1620 3372 1628 3392
rect 1586 3330 1628 3372
rect 1700 3392 1744 3430
rect 1700 3372 1712 3392
rect 1732 3372 1744 3392
rect 1700 3330 1744 3372
rect 1794 3392 1836 3430
rect 1794 3372 1808 3392
rect 1828 3372 1836 3392
rect 1794 3330 1836 3372
rect 1910 3392 1952 3430
rect 1910 3372 1918 3392
rect 1938 3372 1952 3392
rect 1910 3330 1952 3372
rect 2002 3399 2047 3430
rect 2002 3392 2046 3399
rect 2002 3372 2014 3392
rect 2034 3372 2046 3392
rect 2002 3330 2046 3372
rect 6335 3433 6379 3471
rect 6335 3413 6347 3433
rect 6367 3413 6379 3433
rect 2889 3266 2933 3308
rect 2889 3246 2901 3266
rect 2921 3246 2933 3266
rect 2889 3239 2933 3246
rect 2888 3208 2933 3239
rect 2983 3266 3025 3308
rect 2983 3246 2997 3266
rect 3017 3246 3025 3266
rect 2983 3208 3025 3246
rect 3099 3266 3141 3308
rect 3099 3246 3107 3266
rect 3127 3246 3141 3266
rect 3099 3208 3141 3246
rect 3191 3266 3235 3308
rect 3191 3246 3203 3266
rect 3223 3246 3235 3266
rect 3191 3208 3235 3246
rect 3307 3266 3349 3308
rect 3307 3246 3315 3266
rect 3335 3246 3349 3266
rect 3307 3208 3349 3246
rect 3399 3266 3443 3308
rect 3399 3246 3411 3266
rect 3431 3246 3443 3266
rect 3399 3208 3443 3246
rect 3520 3266 3562 3308
rect 3520 3246 3528 3266
rect 3548 3246 3562 3266
rect 3520 3208 3562 3246
rect 3612 3266 3656 3308
rect 6335 3371 6379 3413
rect 6429 3433 6471 3471
rect 6429 3413 6443 3433
rect 6463 3413 6471 3433
rect 6429 3371 6471 3413
rect 6548 3433 6592 3471
rect 6548 3413 6560 3433
rect 6580 3413 6592 3433
rect 6548 3371 6592 3413
rect 6642 3433 6684 3471
rect 6642 3413 6656 3433
rect 6676 3413 6684 3433
rect 6642 3371 6684 3413
rect 6756 3433 6800 3471
rect 6756 3413 6768 3433
rect 6788 3413 6800 3433
rect 6756 3371 6800 3413
rect 6850 3433 6892 3471
rect 6850 3413 6864 3433
rect 6884 3413 6892 3433
rect 6850 3371 6892 3413
rect 6966 3433 7008 3471
rect 6966 3413 6974 3433
rect 6994 3413 7008 3433
rect 6966 3371 7008 3413
rect 7058 3440 7103 3471
rect 7058 3433 7102 3440
rect 7058 3413 7070 3433
rect 7090 3413 7102 3433
rect 7058 3371 7102 3413
rect 3612 3246 3624 3266
rect 3644 3246 3656 3266
rect 3612 3208 3656 3246
rect 7945 3307 7989 3349
rect 7945 3287 7957 3307
rect 7977 3287 7989 3307
rect 7945 3280 7989 3287
rect 7944 3249 7989 3280
rect 8039 3307 8081 3349
rect 8039 3287 8053 3307
rect 8073 3287 8081 3307
rect 8039 3249 8081 3287
rect 8155 3307 8197 3349
rect 8155 3287 8163 3307
rect 8183 3287 8197 3307
rect 8155 3249 8197 3287
rect 8247 3307 8291 3349
rect 8247 3287 8259 3307
rect 8279 3287 8291 3307
rect 8247 3249 8291 3287
rect 8363 3307 8405 3349
rect 8363 3287 8371 3307
rect 8391 3287 8405 3307
rect 8363 3249 8405 3287
rect 8455 3307 8499 3349
rect 8455 3287 8467 3307
rect 8487 3287 8499 3307
rect 8455 3249 8499 3287
rect 8576 3307 8618 3349
rect 8576 3287 8584 3307
rect 8604 3287 8618 3307
rect 8576 3249 8618 3287
rect 8668 3307 8712 3349
rect 8668 3287 8680 3307
rect 8700 3287 8712 3307
rect 8668 3249 8712 3287
rect 340 3082 384 3120
rect 340 3062 352 3082
rect 372 3062 384 3082
rect 340 3020 384 3062
rect 434 3082 476 3120
rect 434 3062 448 3082
rect 468 3062 476 3082
rect 434 3020 476 3062
rect 553 3082 597 3120
rect 553 3062 565 3082
rect 585 3062 597 3082
rect 553 3020 597 3062
rect 647 3082 689 3120
rect 647 3062 661 3082
rect 681 3062 689 3082
rect 647 3020 689 3062
rect 761 3082 805 3120
rect 761 3062 773 3082
rect 793 3062 805 3082
rect 761 3020 805 3062
rect 855 3082 897 3120
rect 855 3062 869 3082
rect 889 3062 897 3082
rect 855 3020 897 3062
rect 971 3082 1013 3120
rect 971 3062 979 3082
rect 999 3062 1013 3082
rect 971 3020 1013 3062
rect 1063 3089 1108 3120
rect 1063 3082 1107 3089
rect 1063 3062 1075 3082
rect 1095 3062 1107 3082
rect 5396 3123 5440 3161
rect 5396 3103 5408 3123
rect 5428 3103 5440 3123
rect 1063 3020 1107 3062
rect 3827 3022 3871 3064
rect 3827 3002 3839 3022
rect 3859 3002 3871 3022
rect 3827 2995 3871 3002
rect 3826 2964 3871 2995
rect 3921 3022 3963 3064
rect 3921 3002 3935 3022
rect 3955 3002 3963 3022
rect 3921 2964 3963 3002
rect 4037 3022 4079 3064
rect 4037 3002 4045 3022
rect 4065 3002 4079 3022
rect 4037 2964 4079 3002
rect 4129 3022 4173 3064
rect 4129 3002 4141 3022
rect 4161 3002 4173 3022
rect 4129 2964 4173 3002
rect 4245 3022 4287 3064
rect 4245 3002 4253 3022
rect 4273 3002 4287 3022
rect 4245 2964 4287 3002
rect 4337 3022 4381 3064
rect 4337 3002 4349 3022
rect 4369 3002 4381 3022
rect 4337 2964 4381 3002
rect 4458 3022 4500 3064
rect 4458 3002 4466 3022
rect 4486 3002 4500 3022
rect 4458 2964 4500 3002
rect 4550 3022 4594 3064
rect 5396 3061 5440 3103
rect 5490 3123 5532 3161
rect 5490 3103 5504 3123
rect 5524 3103 5532 3123
rect 5490 3061 5532 3103
rect 5609 3123 5653 3161
rect 5609 3103 5621 3123
rect 5641 3103 5653 3123
rect 5609 3061 5653 3103
rect 5703 3123 5745 3161
rect 5703 3103 5717 3123
rect 5737 3103 5745 3123
rect 5703 3061 5745 3103
rect 5817 3123 5861 3161
rect 5817 3103 5829 3123
rect 5849 3103 5861 3123
rect 5817 3061 5861 3103
rect 5911 3123 5953 3161
rect 5911 3103 5925 3123
rect 5945 3103 5953 3123
rect 5911 3061 5953 3103
rect 6027 3123 6069 3161
rect 6027 3103 6035 3123
rect 6055 3103 6069 3123
rect 6027 3061 6069 3103
rect 6119 3130 6164 3161
rect 6119 3123 6163 3130
rect 6119 3103 6131 3123
rect 6151 3103 6163 3123
rect 6119 3061 6163 3103
rect 8883 3063 8927 3105
rect 4550 3002 4562 3022
rect 4582 3002 4594 3022
rect 4550 2964 4594 3002
rect 8883 3043 8895 3063
rect 8915 3043 8927 3063
rect 8883 3036 8927 3043
rect 8882 3005 8927 3036
rect 8977 3063 9019 3105
rect 8977 3043 8991 3063
rect 9011 3043 9019 3063
rect 8977 3005 9019 3043
rect 9093 3063 9135 3105
rect 9093 3043 9101 3063
rect 9121 3043 9135 3063
rect 9093 3005 9135 3043
rect 9185 3063 9229 3105
rect 9185 3043 9197 3063
rect 9217 3043 9229 3063
rect 9185 3005 9229 3043
rect 9301 3063 9343 3105
rect 9301 3043 9309 3063
rect 9329 3043 9343 3063
rect 9301 3005 9343 3043
rect 9393 3063 9437 3105
rect 9393 3043 9405 3063
rect 9425 3043 9437 3063
rect 9393 3005 9437 3043
rect 9514 3063 9556 3105
rect 9514 3043 9522 3063
rect 9542 3043 9556 3063
rect 9514 3005 9556 3043
rect 9606 3063 9650 3105
rect 9606 3043 9618 3063
rect 9638 3043 9650 3063
rect 9606 3005 9650 3043
rect 1389 2813 1433 2851
rect 1389 2793 1401 2813
rect 1421 2793 1433 2813
rect 1389 2751 1433 2793
rect 1483 2813 1525 2851
rect 1483 2793 1497 2813
rect 1517 2793 1525 2813
rect 1483 2751 1525 2793
rect 1602 2813 1646 2851
rect 1602 2793 1614 2813
rect 1634 2793 1646 2813
rect 1602 2751 1646 2793
rect 1696 2813 1738 2851
rect 1696 2793 1710 2813
rect 1730 2793 1738 2813
rect 1696 2751 1738 2793
rect 1810 2813 1854 2851
rect 1810 2793 1822 2813
rect 1842 2793 1854 2813
rect 1810 2751 1854 2793
rect 1904 2813 1946 2851
rect 1904 2793 1918 2813
rect 1938 2793 1946 2813
rect 1904 2751 1946 2793
rect 2020 2813 2062 2851
rect 2020 2793 2028 2813
rect 2048 2793 2062 2813
rect 2020 2751 2062 2793
rect 2112 2820 2157 2851
rect 2112 2813 2156 2820
rect 2112 2793 2124 2813
rect 2144 2793 2156 2813
rect 2112 2751 2156 2793
rect 6445 2854 6489 2892
rect 6445 2834 6457 2854
rect 6477 2834 6489 2854
rect 6445 2792 6489 2834
rect 6539 2854 6581 2892
rect 6539 2834 6553 2854
rect 6573 2834 6581 2854
rect 6539 2792 6581 2834
rect 6658 2854 6702 2892
rect 6658 2834 6670 2854
rect 6690 2834 6702 2854
rect 6658 2792 6702 2834
rect 6752 2854 6794 2892
rect 6752 2834 6766 2854
rect 6786 2834 6794 2854
rect 6752 2792 6794 2834
rect 6866 2854 6910 2892
rect 6866 2834 6878 2854
rect 6898 2834 6910 2854
rect 6866 2792 6910 2834
rect 6960 2854 7002 2892
rect 6960 2834 6974 2854
rect 6994 2834 7002 2854
rect 6960 2792 7002 2834
rect 7076 2854 7118 2892
rect 7076 2834 7084 2854
rect 7104 2834 7118 2854
rect 7076 2792 7118 2834
rect 7168 2861 7213 2892
rect 7168 2854 7212 2861
rect 7168 2834 7180 2854
rect 7200 2834 7212 2854
rect 7168 2792 7212 2834
rect 2779 2742 2823 2784
rect 2779 2722 2791 2742
rect 2811 2722 2823 2742
rect 2779 2715 2823 2722
rect 2778 2684 2823 2715
rect 2873 2742 2915 2784
rect 2873 2722 2887 2742
rect 2907 2722 2915 2742
rect 2873 2684 2915 2722
rect 2989 2742 3031 2784
rect 2989 2722 2997 2742
rect 3017 2722 3031 2742
rect 2989 2684 3031 2722
rect 3081 2742 3125 2784
rect 3081 2722 3093 2742
rect 3113 2722 3125 2742
rect 3081 2684 3125 2722
rect 3197 2742 3239 2784
rect 3197 2722 3205 2742
rect 3225 2722 3239 2742
rect 3197 2684 3239 2722
rect 3289 2742 3333 2784
rect 3289 2722 3301 2742
rect 3321 2722 3333 2742
rect 3289 2684 3333 2722
rect 3410 2742 3452 2784
rect 3410 2722 3418 2742
rect 3438 2722 3452 2742
rect 3410 2684 3452 2722
rect 3502 2742 3546 2784
rect 3502 2722 3514 2742
rect 3534 2722 3546 2742
rect 3502 2684 3546 2722
rect 7835 2783 7879 2825
rect 7835 2763 7847 2783
rect 7867 2763 7879 2783
rect 7835 2756 7879 2763
rect 7834 2725 7879 2756
rect 7929 2783 7971 2825
rect 7929 2763 7943 2783
rect 7963 2763 7971 2783
rect 7929 2725 7971 2763
rect 8045 2783 8087 2825
rect 8045 2763 8053 2783
rect 8073 2763 8087 2783
rect 8045 2725 8087 2763
rect 8137 2783 8181 2825
rect 8137 2763 8149 2783
rect 8169 2763 8181 2783
rect 8137 2725 8181 2763
rect 8253 2783 8295 2825
rect 8253 2763 8261 2783
rect 8281 2763 8295 2783
rect 8253 2725 8295 2763
rect 8345 2783 8389 2825
rect 8345 2763 8357 2783
rect 8377 2763 8389 2783
rect 8345 2725 8389 2763
rect 8466 2783 8508 2825
rect 8466 2763 8474 2783
rect 8494 2763 8508 2783
rect 8466 2725 8508 2763
rect 8558 2783 8602 2825
rect 8558 2763 8570 2783
rect 8590 2763 8602 2783
rect 8558 2725 8602 2763
rect 341 2533 385 2571
rect 341 2513 353 2533
rect 373 2513 385 2533
rect 341 2471 385 2513
rect 435 2533 477 2571
rect 435 2513 449 2533
rect 469 2513 477 2533
rect 435 2471 477 2513
rect 554 2533 598 2571
rect 554 2513 566 2533
rect 586 2513 598 2533
rect 554 2471 598 2513
rect 648 2533 690 2571
rect 648 2513 662 2533
rect 682 2513 690 2533
rect 648 2471 690 2513
rect 762 2533 806 2571
rect 762 2513 774 2533
rect 794 2513 806 2533
rect 762 2471 806 2513
rect 856 2533 898 2571
rect 856 2513 870 2533
rect 890 2513 898 2533
rect 856 2471 898 2513
rect 972 2533 1014 2571
rect 972 2513 980 2533
rect 1000 2513 1014 2533
rect 972 2471 1014 2513
rect 1064 2540 1109 2571
rect 1064 2533 1108 2540
rect 1064 2513 1076 2533
rect 1096 2513 1108 2533
rect 5397 2574 5441 2612
rect 5397 2554 5409 2574
rect 5429 2554 5441 2574
rect 1064 2471 1108 2513
rect 3828 2473 3872 2515
rect 3828 2453 3840 2473
rect 3860 2453 3872 2473
rect 3828 2446 3872 2453
rect 3827 2415 3872 2446
rect 3922 2473 3964 2515
rect 3922 2453 3936 2473
rect 3956 2453 3964 2473
rect 3922 2415 3964 2453
rect 4038 2473 4080 2515
rect 4038 2453 4046 2473
rect 4066 2453 4080 2473
rect 4038 2415 4080 2453
rect 4130 2473 4174 2515
rect 4130 2453 4142 2473
rect 4162 2453 4174 2473
rect 4130 2415 4174 2453
rect 4246 2473 4288 2515
rect 4246 2453 4254 2473
rect 4274 2453 4288 2473
rect 4246 2415 4288 2453
rect 4338 2473 4382 2515
rect 4338 2453 4350 2473
rect 4370 2453 4382 2473
rect 4338 2415 4382 2453
rect 4459 2473 4501 2515
rect 4459 2453 4467 2473
rect 4487 2453 4501 2473
rect 4459 2415 4501 2453
rect 4551 2473 4595 2515
rect 5397 2512 5441 2554
rect 5491 2574 5533 2612
rect 5491 2554 5505 2574
rect 5525 2554 5533 2574
rect 5491 2512 5533 2554
rect 5610 2574 5654 2612
rect 5610 2554 5622 2574
rect 5642 2554 5654 2574
rect 5610 2512 5654 2554
rect 5704 2574 5746 2612
rect 5704 2554 5718 2574
rect 5738 2554 5746 2574
rect 5704 2512 5746 2554
rect 5818 2574 5862 2612
rect 5818 2554 5830 2574
rect 5850 2554 5862 2574
rect 5818 2512 5862 2554
rect 5912 2574 5954 2612
rect 5912 2554 5926 2574
rect 5946 2554 5954 2574
rect 5912 2512 5954 2554
rect 6028 2574 6070 2612
rect 6028 2554 6036 2574
rect 6056 2554 6070 2574
rect 6028 2512 6070 2554
rect 6120 2581 6165 2612
rect 6120 2574 6164 2581
rect 6120 2554 6132 2574
rect 6152 2554 6164 2574
rect 6120 2512 6164 2554
rect 8884 2514 8928 2556
rect 4551 2453 4563 2473
rect 4583 2453 4595 2473
rect 4551 2415 4595 2453
rect 8884 2494 8896 2514
rect 8916 2494 8928 2514
rect 8884 2487 8928 2494
rect 8883 2456 8928 2487
rect 8978 2514 9020 2556
rect 8978 2494 8992 2514
rect 9012 2494 9020 2514
rect 8978 2456 9020 2494
rect 9094 2514 9136 2556
rect 9094 2494 9102 2514
rect 9122 2494 9136 2514
rect 9094 2456 9136 2494
rect 9186 2514 9230 2556
rect 9186 2494 9198 2514
rect 9218 2494 9230 2514
rect 9186 2456 9230 2494
rect 9302 2514 9344 2556
rect 9302 2494 9310 2514
rect 9330 2494 9344 2514
rect 9302 2456 9344 2494
rect 9394 2514 9438 2556
rect 9394 2494 9406 2514
rect 9426 2494 9438 2514
rect 9394 2456 9438 2494
rect 9515 2514 9557 2556
rect 9515 2494 9523 2514
rect 9543 2494 9557 2514
rect 9515 2456 9557 2494
rect 9607 2514 9651 2556
rect 9607 2494 9619 2514
rect 9639 2494 9651 2514
rect 9607 2456 9651 2494
rect 1279 2289 1323 2327
rect 1279 2269 1291 2289
rect 1311 2269 1323 2289
rect 1279 2227 1323 2269
rect 1373 2289 1415 2327
rect 1373 2269 1387 2289
rect 1407 2269 1415 2289
rect 1373 2227 1415 2269
rect 1492 2289 1536 2327
rect 1492 2269 1504 2289
rect 1524 2269 1536 2289
rect 1492 2227 1536 2269
rect 1586 2289 1628 2327
rect 1586 2269 1600 2289
rect 1620 2269 1628 2289
rect 1586 2227 1628 2269
rect 1700 2289 1744 2327
rect 1700 2269 1712 2289
rect 1732 2269 1744 2289
rect 1700 2227 1744 2269
rect 1794 2289 1836 2327
rect 1794 2269 1808 2289
rect 1828 2269 1836 2289
rect 1794 2227 1836 2269
rect 1910 2289 1952 2327
rect 1910 2269 1918 2289
rect 1938 2269 1952 2289
rect 1910 2227 1952 2269
rect 2002 2296 2047 2327
rect 2002 2289 2046 2296
rect 2002 2269 2014 2289
rect 2034 2269 2046 2289
rect 2002 2227 2046 2269
rect 6335 2330 6379 2368
rect 6335 2310 6347 2330
rect 6367 2310 6379 2330
rect 2889 2163 2933 2205
rect 2889 2143 2901 2163
rect 2921 2143 2933 2163
rect 2889 2136 2933 2143
rect 2888 2105 2933 2136
rect 2983 2163 3025 2205
rect 2983 2143 2997 2163
rect 3017 2143 3025 2163
rect 2983 2105 3025 2143
rect 3099 2163 3141 2205
rect 3099 2143 3107 2163
rect 3127 2143 3141 2163
rect 3099 2105 3141 2143
rect 3191 2163 3235 2205
rect 3191 2143 3203 2163
rect 3223 2143 3235 2163
rect 3191 2105 3235 2143
rect 3307 2163 3349 2205
rect 3307 2143 3315 2163
rect 3335 2143 3349 2163
rect 3307 2105 3349 2143
rect 3399 2163 3443 2205
rect 3399 2143 3411 2163
rect 3431 2143 3443 2163
rect 3399 2105 3443 2143
rect 3520 2163 3562 2205
rect 3520 2143 3528 2163
rect 3548 2143 3562 2163
rect 3520 2105 3562 2143
rect 3612 2163 3656 2205
rect 6335 2268 6379 2310
rect 6429 2330 6471 2368
rect 6429 2310 6443 2330
rect 6463 2310 6471 2330
rect 6429 2268 6471 2310
rect 6548 2330 6592 2368
rect 6548 2310 6560 2330
rect 6580 2310 6592 2330
rect 6548 2268 6592 2310
rect 6642 2330 6684 2368
rect 6642 2310 6656 2330
rect 6676 2310 6684 2330
rect 6642 2268 6684 2310
rect 6756 2330 6800 2368
rect 6756 2310 6768 2330
rect 6788 2310 6800 2330
rect 6756 2268 6800 2310
rect 6850 2330 6892 2368
rect 6850 2310 6864 2330
rect 6884 2310 6892 2330
rect 6850 2268 6892 2310
rect 6966 2330 7008 2368
rect 6966 2310 6974 2330
rect 6994 2310 7008 2330
rect 6966 2268 7008 2310
rect 7058 2337 7103 2368
rect 7058 2330 7102 2337
rect 7058 2310 7070 2330
rect 7090 2310 7102 2330
rect 7058 2268 7102 2310
rect 3612 2143 3624 2163
rect 3644 2143 3656 2163
rect 3612 2105 3656 2143
rect 7945 2204 7989 2246
rect 7945 2184 7957 2204
rect 7977 2184 7989 2204
rect 7945 2177 7989 2184
rect 7944 2146 7989 2177
rect 8039 2204 8081 2246
rect 8039 2184 8053 2204
rect 8073 2184 8081 2204
rect 8039 2146 8081 2184
rect 8155 2204 8197 2246
rect 8155 2184 8163 2204
rect 8183 2184 8197 2204
rect 8155 2146 8197 2184
rect 8247 2204 8291 2246
rect 8247 2184 8259 2204
rect 8279 2184 8291 2204
rect 8247 2146 8291 2184
rect 8363 2204 8405 2246
rect 8363 2184 8371 2204
rect 8391 2184 8405 2204
rect 8363 2146 8405 2184
rect 8455 2204 8499 2246
rect 8455 2184 8467 2204
rect 8487 2184 8499 2204
rect 8455 2146 8499 2184
rect 8576 2204 8618 2246
rect 8576 2184 8584 2204
rect 8604 2184 8618 2204
rect 8576 2146 8618 2184
rect 8668 2204 8712 2246
rect 8668 2184 8680 2204
rect 8700 2184 8712 2204
rect 8668 2146 8712 2184
rect 340 1979 384 2017
rect 340 1959 352 1979
rect 372 1959 384 1979
rect 340 1917 384 1959
rect 434 1979 476 2017
rect 434 1959 448 1979
rect 468 1959 476 1979
rect 434 1917 476 1959
rect 553 1979 597 2017
rect 553 1959 565 1979
rect 585 1959 597 1979
rect 553 1917 597 1959
rect 647 1979 689 2017
rect 647 1959 661 1979
rect 681 1959 689 1979
rect 647 1917 689 1959
rect 761 1979 805 2017
rect 761 1959 773 1979
rect 793 1959 805 1979
rect 761 1917 805 1959
rect 855 1979 897 2017
rect 855 1959 869 1979
rect 889 1959 897 1979
rect 855 1917 897 1959
rect 971 1979 1013 2017
rect 971 1959 979 1979
rect 999 1959 1013 1979
rect 971 1917 1013 1959
rect 1063 1986 1108 2017
rect 1063 1979 1107 1986
rect 1063 1959 1075 1979
rect 1095 1959 1107 1979
rect 5396 2020 5440 2058
rect 5396 2000 5408 2020
rect 5428 2000 5440 2020
rect 1063 1917 1107 1959
rect 3827 1919 3871 1961
rect 3827 1899 3839 1919
rect 3859 1899 3871 1919
rect 3827 1892 3871 1899
rect 3826 1861 3871 1892
rect 3921 1919 3963 1961
rect 3921 1899 3935 1919
rect 3955 1899 3963 1919
rect 3921 1861 3963 1899
rect 4037 1919 4079 1961
rect 4037 1899 4045 1919
rect 4065 1899 4079 1919
rect 4037 1861 4079 1899
rect 4129 1919 4173 1961
rect 4129 1899 4141 1919
rect 4161 1899 4173 1919
rect 4129 1861 4173 1899
rect 4245 1919 4287 1961
rect 4245 1899 4253 1919
rect 4273 1899 4287 1919
rect 4245 1861 4287 1899
rect 4337 1919 4381 1961
rect 4337 1899 4349 1919
rect 4369 1899 4381 1919
rect 4337 1861 4381 1899
rect 4458 1919 4500 1961
rect 4458 1899 4466 1919
rect 4486 1899 4500 1919
rect 4458 1861 4500 1899
rect 4550 1919 4594 1961
rect 5396 1958 5440 2000
rect 5490 2020 5532 2058
rect 5490 2000 5504 2020
rect 5524 2000 5532 2020
rect 5490 1958 5532 2000
rect 5609 2020 5653 2058
rect 5609 2000 5621 2020
rect 5641 2000 5653 2020
rect 5609 1958 5653 2000
rect 5703 2020 5745 2058
rect 5703 2000 5717 2020
rect 5737 2000 5745 2020
rect 5703 1958 5745 2000
rect 5817 2020 5861 2058
rect 5817 2000 5829 2020
rect 5849 2000 5861 2020
rect 5817 1958 5861 2000
rect 5911 2020 5953 2058
rect 5911 2000 5925 2020
rect 5945 2000 5953 2020
rect 5911 1958 5953 2000
rect 6027 2020 6069 2058
rect 6027 2000 6035 2020
rect 6055 2000 6069 2020
rect 6027 1958 6069 2000
rect 6119 2027 6164 2058
rect 6119 2020 6163 2027
rect 6119 2000 6131 2020
rect 6151 2000 6163 2020
rect 6119 1958 6163 2000
rect 8883 1960 8927 2002
rect 4550 1899 4562 1919
rect 4582 1899 4594 1919
rect 4550 1861 4594 1899
rect 8883 1940 8895 1960
rect 8915 1940 8927 1960
rect 8883 1933 8927 1940
rect 8882 1902 8927 1933
rect 8977 1960 9019 2002
rect 8977 1940 8991 1960
rect 9011 1940 9019 1960
rect 8977 1902 9019 1940
rect 9093 1960 9135 2002
rect 9093 1940 9101 1960
rect 9121 1940 9135 1960
rect 9093 1902 9135 1940
rect 9185 1960 9229 2002
rect 9185 1940 9197 1960
rect 9217 1940 9229 1960
rect 9185 1902 9229 1940
rect 9301 1960 9343 2002
rect 9301 1940 9309 1960
rect 9329 1940 9343 1960
rect 9301 1902 9343 1940
rect 9393 1960 9437 2002
rect 9393 1940 9405 1960
rect 9425 1940 9437 1960
rect 9393 1902 9437 1940
rect 9514 1960 9556 2002
rect 9514 1940 9522 1960
rect 9542 1940 9556 1960
rect 9514 1902 9556 1940
rect 9606 1960 9650 2002
rect 9606 1940 9618 1960
rect 9638 1940 9650 1960
rect 9606 1902 9650 1940
rect 1420 1697 1464 1735
rect 1420 1677 1432 1697
rect 1452 1677 1464 1697
rect 1420 1635 1464 1677
rect 1514 1697 1556 1735
rect 1514 1677 1528 1697
rect 1548 1677 1556 1697
rect 1514 1635 1556 1677
rect 1633 1697 1677 1735
rect 1633 1677 1645 1697
rect 1665 1677 1677 1697
rect 1633 1635 1677 1677
rect 1727 1697 1769 1735
rect 1727 1677 1741 1697
rect 1761 1677 1769 1697
rect 1727 1635 1769 1677
rect 1841 1697 1885 1735
rect 1841 1677 1853 1697
rect 1873 1677 1885 1697
rect 1841 1635 1885 1677
rect 1935 1697 1977 1735
rect 1935 1677 1949 1697
rect 1969 1677 1977 1697
rect 1935 1635 1977 1677
rect 2051 1697 2093 1735
rect 2051 1677 2059 1697
rect 2079 1677 2093 1697
rect 2051 1635 2093 1677
rect 2143 1704 2188 1735
rect 2143 1697 2187 1704
rect 2143 1677 2155 1697
rect 2175 1677 2187 1697
rect 6476 1738 6520 1776
rect 6476 1718 6488 1738
rect 6508 1718 6520 1738
rect 2143 1635 2187 1677
rect 2749 1652 2793 1694
rect 2749 1632 2761 1652
rect 2781 1632 2793 1652
rect 2749 1625 2793 1632
rect 2748 1594 2793 1625
rect 2843 1652 2885 1694
rect 2843 1632 2857 1652
rect 2877 1632 2885 1652
rect 2843 1594 2885 1632
rect 2959 1652 3001 1694
rect 2959 1632 2967 1652
rect 2987 1632 3001 1652
rect 2959 1594 3001 1632
rect 3051 1652 3095 1694
rect 3051 1632 3063 1652
rect 3083 1632 3095 1652
rect 3051 1594 3095 1632
rect 3167 1652 3209 1694
rect 3167 1632 3175 1652
rect 3195 1632 3209 1652
rect 3167 1594 3209 1632
rect 3259 1652 3303 1694
rect 3259 1632 3271 1652
rect 3291 1632 3303 1652
rect 3259 1594 3303 1632
rect 3380 1652 3422 1694
rect 3380 1632 3388 1652
rect 3408 1632 3422 1652
rect 3380 1594 3422 1632
rect 3472 1652 3516 1694
rect 6476 1676 6520 1718
rect 6570 1738 6612 1776
rect 6570 1718 6584 1738
rect 6604 1718 6612 1738
rect 6570 1676 6612 1718
rect 6689 1738 6733 1776
rect 6689 1718 6701 1738
rect 6721 1718 6733 1738
rect 6689 1676 6733 1718
rect 6783 1738 6825 1776
rect 6783 1718 6797 1738
rect 6817 1718 6825 1738
rect 6783 1676 6825 1718
rect 6897 1738 6941 1776
rect 6897 1718 6909 1738
rect 6929 1718 6941 1738
rect 6897 1676 6941 1718
rect 6991 1738 7033 1776
rect 6991 1718 7005 1738
rect 7025 1718 7033 1738
rect 6991 1676 7033 1718
rect 7107 1738 7149 1776
rect 7107 1718 7115 1738
rect 7135 1718 7149 1738
rect 7107 1676 7149 1718
rect 7199 1745 7244 1776
rect 7199 1738 7243 1745
rect 7199 1718 7211 1738
rect 7231 1718 7243 1738
rect 7199 1676 7243 1718
rect 7805 1693 7849 1735
rect 3472 1632 3484 1652
rect 3504 1632 3516 1652
rect 3472 1594 3516 1632
rect 7805 1673 7817 1693
rect 7837 1673 7849 1693
rect 7805 1666 7849 1673
rect 7804 1635 7849 1666
rect 7899 1693 7941 1735
rect 7899 1673 7913 1693
rect 7933 1673 7941 1693
rect 7899 1635 7941 1673
rect 8015 1693 8057 1735
rect 8015 1673 8023 1693
rect 8043 1673 8057 1693
rect 8015 1635 8057 1673
rect 8107 1693 8151 1735
rect 8107 1673 8119 1693
rect 8139 1673 8151 1693
rect 8107 1635 8151 1673
rect 8223 1693 8265 1735
rect 8223 1673 8231 1693
rect 8251 1673 8265 1693
rect 8223 1635 8265 1673
rect 8315 1693 8359 1735
rect 8315 1673 8327 1693
rect 8347 1673 8359 1693
rect 8315 1635 8359 1673
rect 8436 1693 8478 1735
rect 8436 1673 8444 1693
rect 8464 1673 8478 1693
rect 8436 1635 8478 1673
rect 8528 1693 8572 1735
rect 8528 1673 8540 1693
rect 8560 1673 8572 1693
rect 8528 1635 8572 1673
rect 342 1430 386 1468
rect 342 1410 354 1430
rect 374 1410 386 1430
rect 342 1368 386 1410
rect 436 1430 478 1468
rect 436 1410 450 1430
rect 470 1410 478 1430
rect 436 1368 478 1410
rect 555 1430 599 1468
rect 555 1410 567 1430
rect 587 1410 599 1430
rect 555 1368 599 1410
rect 649 1430 691 1468
rect 649 1410 663 1430
rect 683 1410 691 1430
rect 649 1368 691 1410
rect 763 1430 807 1468
rect 763 1410 775 1430
rect 795 1410 807 1430
rect 763 1368 807 1410
rect 857 1430 899 1468
rect 857 1410 871 1430
rect 891 1410 899 1430
rect 857 1368 899 1410
rect 973 1430 1015 1468
rect 973 1410 981 1430
rect 1001 1410 1015 1430
rect 973 1368 1015 1410
rect 1065 1437 1110 1468
rect 1065 1430 1109 1437
rect 1065 1410 1077 1430
rect 1097 1410 1109 1430
rect 5398 1471 5442 1509
rect 5398 1451 5410 1471
rect 5430 1451 5442 1471
rect 1065 1368 1109 1410
rect 3829 1370 3873 1412
rect 3829 1350 3841 1370
rect 3861 1350 3873 1370
rect 3829 1343 3873 1350
rect 3828 1312 3873 1343
rect 3923 1370 3965 1412
rect 3923 1350 3937 1370
rect 3957 1350 3965 1370
rect 3923 1312 3965 1350
rect 4039 1370 4081 1412
rect 4039 1350 4047 1370
rect 4067 1350 4081 1370
rect 4039 1312 4081 1350
rect 4131 1370 4175 1412
rect 4131 1350 4143 1370
rect 4163 1350 4175 1370
rect 4131 1312 4175 1350
rect 4247 1370 4289 1412
rect 4247 1350 4255 1370
rect 4275 1350 4289 1370
rect 4247 1312 4289 1350
rect 4339 1370 4383 1412
rect 4339 1350 4351 1370
rect 4371 1350 4383 1370
rect 4339 1312 4383 1350
rect 4460 1370 4502 1412
rect 4460 1350 4468 1370
rect 4488 1350 4502 1370
rect 4460 1312 4502 1350
rect 4552 1370 4596 1412
rect 5398 1409 5442 1451
rect 5492 1471 5534 1509
rect 5492 1451 5506 1471
rect 5526 1451 5534 1471
rect 5492 1409 5534 1451
rect 5611 1471 5655 1509
rect 5611 1451 5623 1471
rect 5643 1451 5655 1471
rect 5611 1409 5655 1451
rect 5705 1471 5747 1509
rect 5705 1451 5719 1471
rect 5739 1451 5747 1471
rect 5705 1409 5747 1451
rect 5819 1471 5863 1509
rect 5819 1451 5831 1471
rect 5851 1451 5863 1471
rect 5819 1409 5863 1451
rect 5913 1471 5955 1509
rect 5913 1451 5927 1471
rect 5947 1451 5955 1471
rect 5913 1409 5955 1451
rect 6029 1471 6071 1509
rect 6029 1451 6037 1471
rect 6057 1451 6071 1471
rect 6029 1409 6071 1451
rect 6121 1478 6166 1509
rect 6121 1471 6165 1478
rect 6121 1451 6133 1471
rect 6153 1451 6165 1471
rect 6121 1409 6165 1451
rect 8885 1411 8929 1453
rect 4552 1350 4564 1370
rect 4584 1350 4596 1370
rect 4552 1312 4596 1350
rect 8885 1391 8897 1411
rect 8917 1391 8929 1411
rect 8885 1384 8929 1391
rect 8884 1353 8929 1384
rect 8979 1411 9021 1453
rect 8979 1391 8993 1411
rect 9013 1391 9021 1411
rect 8979 1353 9021 1391
rect 9095 1411 9137 1453
rect 9095 1391 9103 1411
rect 9123 1391 9137 1411
rect 9095 1353 9137 1391
rect 9187 1411 9231 1453
rect 9187 1391 9199 1411
rect 9219 1391 9231 1411
rect 9187 1353 9231 1391
rect 9303 1411 9345 1453
rect 9303 1391 9311 1411
rect 9331 1391 9345 1411
rect 9303 1353 9345 1391
rect 9395 1411 9439 1453
rect 9395 1391 9407 1411
rect 9427 1391 9439 1411
rect 9395 1353 9439 1391
rect 9516 1411 9558 1453
rect 9516 1391 9524 1411
rect 9544 1391 9558 1411
rect 9516 1353 9558 1391
rect 9608 1411 9652 1453
rect 9608 1391 9620 1411
rect 9640 1391 9652 1411
rect 9608 1353 9652 1391
rect 1280 1186 1324 1224
rect 1280 1166 1292 1186
rect 1312 1166 1324 1186
rect 1280 1124 1324 1166
rect 1374 1186 1416 1224
rect 1374 1166 1388 1186
rect 1408 1166 1416 1186
rect 1374 1124 1416 1166
rect 1493 1186 1537 1224
rect 1493 1166 1505 1186
rect 1525 1166 1537 1186
rect 1493 1124 1537 1166
rect 1587 1186 1629 1224
rect 1587 1166 1601 1186
rect 1621 1166 1629 1186
rect 1587 1124 1629 1166
rect 1701 1186 1745 1224
rect 1701 1166 1713 1186
rect 1733 1166 1745 1186
rect 1701 1124 1745 1166
rect 1795 1186 1837 1224
rect 1795 1166 1809 1186
rect 1829 1166 1837 1186
rect 1795 1124 1837 1166
rect 1911 1186 1953 1224
rect 1911 1166 1919 1186
rect 1939 1166 1953 1186
rect 1911 1124 1953 1166
rect 2003 1193 2048 1224
rect 2003 1186 2047 1193
rect 2003 1166 2015 1186
rect 2035 1166 2047 1186
rect 2003 1124 2047 1166
rect 6336 1227 6380 1265
rect 6336 1207 6348 1227
rect 6368 1207 6380 1227
rect 2890 1060 2934 1102
rect 2890 1040 2902 1060
rect 2922 1040 2934 1060
rect 2890 1033 2934 1040
rect 2889 1002 2934 1033
rect 2984 1060 3026 1102
rect 2984 1040 2998 1060
rect 3018 1040 3026 1060
rect 2984 1002 3026 1040
rect 3100 1060 3142 1102
rect 3100 1040 3108 1060
rect 3128 1040 3142 1060
rect 3100 1002 3142 1040
rect 3192 1060 3236 1102
rect 3192 1040 3204 1060
rect 3224 1040 3236 1060
rect 3192 1002 3236 1040
rect 3308 1060 3350 1102
rect 3308 1040 3316 1060
rect 3336 1040 3350 1060
rect 3308 1002 3350 1040
rect 3400 1060 3444 1102
rect 3400 1040 3412 1060
rect 3432 1040 3444 1060
rect 3400 1002 3444 1040
rect 3521 1060 3563 1102
rect 3521 1040 3529 1060
rect 3549 1040 3563 1060
rect 3521 1002 3563 1040
rect 3613 1060 3657 1102
rect 6336 1165 6380 1207
rect 6430 1227 6472 1265
rect 6430 1207 6444 1227
rect 6464 1207 6472 1227
rect 6430 1165 6472 1207
rect 6549 1227 6593 1265
rect 6549 1207 6561 1227
rect 6581 1207 6593 1227
rect 6549 1165 6593 1207
rect 6643 1227 6685 1265
rect 6643 1207 6657 1227
rect 6677 1207 6685 1227
rect 6643 1165 6685 1207
rect 6757 1227 6801 1265
rect 6757 1207 6769 1227
rect 6789 1207 6801 1227
rect 6757 1165 6801 1207
rect 6851 1227 6893 1265
rect 6851 1207 6865 1227
rect 6885 1207 6893 1227
rect 6851 1165 6893 1207
rect 6967 1227 7009 1265
rect 6967 1207 6975 1227
rect 6995 1207 7009 1227
rect 6967 1165 7009 1207
rect 7059 1234 7104 1265
rect 7059 1227 7103 1234
rect 7059 1207 7071 1227
rect 7091 1207 7103 1227
rect 7059 1165 7103 1207
rect 3613 1040 3625 1060
rect 3645 1040 3657 1060
rect 3613 1002 3657 1040
rect 7946 1101 7990 1143
rect 7946 1081 7958 1101
rect 7978 1081 7990 1101
rect 7946 1074 7990 1081
rect 7945 1043 7990 1074
rect 8040 1101 8082 1143
rect 8040 1081 8054 1101
rect 8074 1081 8082 1101
rect 8040 1043 8082 1081
rect 8156 1101 8198 1143
rect 8156 1081 8164 1101
rect 8184 1081 8198 1101
rect 8156 1043 8198 1081
rect 8248 1101 8292 1143
rect 8248 1081 8260 1101
rect 8280 1081 8292 1101
rect 8248 1043 8292 1081
rect 8364 1101 8406 1143
rect 8364 1081 8372 1101
rect 8392 1081 8406 1101
rect 8364 1043 8406 1081
rect 8456 1101 8500 1143
rect 8456 1081 8468 1101
rect 8488 1081 8500 1101
rect 8456 1043 8500 1081
rect 8577 1101 8619 1143
rect 8577 1081 8585 1101
rect 8605 1081 8619 1101
rect 8577 1043 8619 1081
rect 8669 1101 8713 1143
rect 8669 1081 8681 1101
rect 8701 1081 8713 1101
rect 8669 1043 8713 1081
rect 341 876 385 914
rect 341 856 353 876
rect 373 856 385 876
rect 341 814 385 856
rect 435 876 477 914
rect 435 856 449 876
rect 469 856 477 876
rect 435 814 477 856
rect 554 876 598 914
rect 554 856 566 876
rect 586 856 598 876
rect 554 814 598 856
rect 648 876 690 914
rect 648 856 662 876
rect 682 856 690 876
rect 648 814 690 856
rect 762 876 806 914
rect 762 856 774 876
rect 794 856 806 876
rect 762 814 806 856
rect 856 876 898 914
rect 856 856 870 876
rect 890 856 898 876
rect 856 814 898 856
rect 972 876 1014 914
rect 972 856 980 876
rect 1000 856 1014 876
rect 972 814 1014 856
rect 1064 883 1109 914
rect 1064 876 1108 883
rect 1064 856 1076 876
rect 1096 856 1108 876
rect 5397 917 5441 955
rect 5397 897 5409 917
rect 5429 897 5441 917
rect 1064 814 1108 856
rect 3828 816 3872 858
rect 3828 796 3840 816
rect 3860 796 3872 816
rect 3828 789 3872 796
rect 3827 758 3872 789
rect 3922 816 3964 858
rect 3922 796 3936 816
rect 3956 796 3964 816
rect 3922 758 3964 796
rect 4038 816 4080 858
rect 4038 796 4046 816
rect 4066 796 4080 816
rect 4038 758 4080 796
rect 4130 816 4174 858
rect 4130 796 4142 816
rect 4162 796 4174 816
rect 4130 758 4174 796
rect 4246 816 4288 858
rect 4246 796 4254 816
rect 4274 796 4288 816
rect 4246 758 4288 796
rect 4338 816 4382 858
rect 4338 796 4350 816
rect 4370 796 4382 816
rect 4338 758 4382 796
rect 4459 816 4501 858
rect 4459 796 4467 816
rect 4487 796 4501 816
rect 4459 758 4501 796
rect 4551 816 4595 858
rect 5397 855 5441 897
rect 5491 917 5533 955
rect 5491 897 5505 917
rect 5525 897 5533 917
rect 5491 855 5533 897
rect 5610 917 5654 955
rect 5610 897 5622 917
rect 5642 897 5654 917
rect 5610 855 5654 897
rect 5704 917 5746 955
rect 5704 897 5718 917
rect 5738 897 5746 917
rect 5704 855 5746 897
rect 5818 917 5862 955
rect 5818 897 5830 917
rect 5850 897 5862 917
rect 5818 855 5862 897
rect 5912 917 5954 955
rect 5912 897 5926 917
rect 5946 897 5954 917
rect 5912 855 5954 897
rect 6028 917 6070 955
rect 6028 897 6036 917
rect 6056 897 6070 917
rect 6028 855 6070 897
rect 6120 924 6165 955
rect 6120 917 6164 924
rect 6120 897 6132 917
rect 6152 897 6164 917
rect 6120 855 6164 897
rect 8884 857 8928 899
rect 4551 796 4563 816
rect 4583 796 4595 816
rect 4551 758 4595 796
rect 8884 837 8896 857
rect 8916 837 8928 857
rect 8884 830 8928 837
rect 8883 799 8928 830
rect 8978 857 9020 899
rect 8978 837 8992 857
rect 9012 837 9020 857
rect 8978 799 9020 837
rect 9094 857 9136 899
rect 9094 837 9102 857
rect 9122 837 9136 857
rect 9094 799 9136 837
rect 9186 857 9230 899
rect 9186 837 9198 857
rect 9218 837 9230 857
rect 9186 799 9230 837
rect 9302 857 9344 899
rect 9302 837 9310 857
rect 9330 837 9344 857
rect 9302 799 9344 837
rect 9394 857 9438 899
rect 9394 837 9406 857
rect 9426 837 9438 857
rect 9394 799 9438 837
rect 9515 857 9557 899
rect 9515 837 9523 857
rect 9543 837 9557 857
rect 9515 799 9557 837
rect 9607 857 9651 899
rect 9607 837 9619 857
rect 9639 837 9651 857
rect 9607 799 9651 837
rect 6644 358 6688 396
rect 1588 317 1632 355
rect 1588 297 1600 317
rect 1620 297 1632 317
rect 1588 255 1632 297
rect 1682 317 1724 355
rect 1682 297 1696 317
rect 1716 297 1724 317
rect 1682 255 1724 297
rect 1801 317 1845 355
rect 1801 297 1813 317
rect 1833 297 1845 317
rect 1801 255 1845 297
rect 1895 317 1937 355
rect 1895 297 1909 317
rect 1929 297 1937 317
rect 1895 255 1937 297
rect 2009 317 2053 355
rect 2009 297 2021 317
rect 2041 297 2053 317
rect 2009 255 2053 297
rect 2103 317 2145 355
rect 2103 297 2117 317
rect 2137 297 2145 317
rect 2103 255 2145 297
rect 2219 317 2261 355
rect 2219 297 2227 317
rect 2247 297 2261 317
rect 2219 255 2261 297
rect 2311 324 2356 355
rect 6644 338 6656 358
rect 6676 338 6688 358
rect 2311 317 2355 324
rect 2311 297 2323 317
rect 2343 297 2355 317
rect 2311 255 2355 297
rect 4538 297 4582 335
rect 4538 277 4550 297
rect 4570 277 4582 297
rect 4538 235 4582 277
rect 4632 297 4674 335
rect 4632 277 4646 297
rect 4666 277 4674 297
rect 4632 235 4674 277
rect 4751 297 4795 335
rect 4751 277 4763 297
rect 4783 277 4795 297
rect 4751 235 4795 277
rect 4845 297 4887 335
rect 4845 277 4859 297
rect 4879 277 4887 297
rect 4845 235 4887 277
rect 4959 297 5003 335
rect 4959 277 4971 297
rect 4991 277 5003 297
rect 4959 235 5003 277
rect 5053 297 5095 335
rect 5053 277 5067 297
rect 5087 277 5095 297
rect 5053 235 5095 277
rect 5169 297 5211 335
rect 5169 277 5177 297
rect 5197 277 5211 297
rect 5169 235 5211 277
rect 5261 304 5306 335
rect 5261 297 5305 304
rect 5261 277 5273 297
rect 5293 277 5305 297
rect 6644 296 6688 338
rect 6738 358 6780 396
rect 6738 338 6752 358
rect 6772 338 6780 358
rect 6738 296 6780 338
rect 6857 358 6901 396
rect 6857 338 6869 358
rect 6889 338 6901 358
rect 6857 296 6901 338
rect 6951 358 6993 396
rect 6951 338 6965 358
rect 6985 338 6993 358
rect 6951 296 6993 338
rect 7065 358 7109 396
rect 7065 338 7077 358
rect 7097 338 7109 358
rect 7065 296 7109 338
rect 7159 358 7201 396
rect 7159 338 7173 358
rect 7193 338 7201 358
rect 7159 296 7201 338
rect 7275 358 7317 396
rect 7275 338 7283 358
rect 7303 338 7317 358
rect 7275 296 7317 338
rect 7367 365 7412 396
rect 7367 358 7411 365
rect 7367 338 7379 358
rect 7399 338 7411 358
rect 7367 296 7411 338
rect 5261 235 5305 277
<< ndiffc >>
rect 5172 9308 5190 9326
rect 116 9267 134 9285
rect 3831 9220 3851 9240
rect 3934 9216 3954 9236
rect 4042 9216 4062 9236
rect 4145 9220 4165 9240
rect 4250 9216 4270 9236
rect 4353 9220 4373 9240
rect 4463 9216 4483 9236
rect 8887 9261 8907 9281
rect 8990 9257 9010 9277
rect 9098 9257 9118 9277
rect 9201 9261 9221 9281
rect 9306 9257 9326 9277
rect 9409 9261 9429 9281
rect 9519 9257 9539 9277
rect 9622 9261 9642 9281
rect 4566 9220 4586 9240
rect 118 9168 136 9186
rect 116 9080 134 9098
rect 5174 9209 5192 9227
rect 118 8981 136 8999
rect 344 8982 364 9002
rect 447 8986 467 9006
rect 557 8982 577 9002
rect 660 8986 680 9006
rect 765 8982 785 9002
rect 868 8986 888 9006
rect 976 8986 996 9006
rect 1079 8982 1099 9002
rect 4793 9128 4811 9146
rect 5172 9121 5190 9139
rect 4795 9029 4813 9047
rect 5174 9022 5192 9040
rect 5400 9023 5420 9043
rect 5503 9027 5523 9047
rect 5613 9023 5633 9043
rect 5716 9027 5736 9047
rect 5821 9023 5841 9043
rect 5924 9027 5944 9047
rect 6032 9027 6052 9047
rect 6135 9023 6155 9043
rect 9849 9169 9867 9187
rect 9851 9070 9869 9088
rect 116 8851 134 8869
rect 2892 8910 2912 8930
rect 2995 8906 3015 8926
rect 3103 8906 3123 8926
rect 3206 8910 3226 8930
rect 3311 8906 3331 8926
rect 3414 8910 3434 8930
rect 3524 8906 3544 8926
rect 3627 8910 3647 8930
rect 118 8752 136 8770
rect 4793 8898 4811 8916
rect 5172 8892 5190 8910
rect 1282 8738 1302 8758
rect 1385 8742 1405 8762
rect 1495 8738 1515 8758
rect 1598 8742 1618 8762
rect 1703 8738 1723 8758
rect 1806 8742 1826 8762
rect 1914 8742 1934 8762
rect 2017 8738 2037 8758
rect 7948 8951 7968 8971
rect 8051 8947 8071 8967
rect 8159 8947 8179 8967
rect 8262 8951 8282 8971
rect 8367 8947 8387 8967
rect 8470 8951 8490 8971
rect 8580 8947 8600 8967
rect 8683 8951 8703 8971
rect 4795 8799 4813 8817
rect 5174 8793 5192 8811
rect 9849 8939 9867 8957
rect 6338 8779 6358 8799
rect 6441 8783 6461 8803
rect 6551 8779 6571 8799
rect 6654 8783 6674 8803
rect 6759 8779 6779 8799
rect 6862 8783 6882 8803
rect 6970 8783 6990 8803
rect 7073 8779 7093 8799
rect 9851 8840 9869 8858
rect 116 8621 134 8639
rect 118 8522 136 8540
rect 3830 8666 3850 8686
rect 3933 8662 3953 8682
rect 4041 8662 4061 8682
rect 4144 8666 4164 8686
rect 4249 8662 4269 8682
rect 4352 8666 4372 8686
rect 4462 8662 4482 8682
rect 4565 8666 4585 8686
rect 4793 8669 4811 8687
rect 5172 8662 5190 8680
rect 4795 8570 4813 8588
rect 5174 8563 5192 8581
rect 8886 8707 8906 8727
rect 8989 8703 9009 8723
rect 9097 8703 9117 8723
rect 9200 8707 9220 8727
rect 9305 8703 9325 8723
rect 9408 8707 9428 8727
rect 9518 8703 9538 8723
rect 9621 8707 9641 8727
rect 9849 8710 9867 8728
rect 4793 8482 4811 8500
rect 9851 8611 9869 8629
rect 9849 8523 9867 8541
rect 5399 8469 5419 8489
rect 343 8428 363 8448
rect 446 8432 466 8452
rect 556 8428 576 8448
rect 659 8432 679 8452
rect 764 8428 784 8448
rect 867 8432 887 8452
rect 975 8432 995 8452
rect 1078 8428 1098 8448
rect 2752 8399 2772 8419
rect 2855 8395 2875 8415
rect 2963 8395 2983 8415
rect 3066 8399 3086 8419
rect 3171 8395 3191 8415
rect 3274 8399 3294 8419
rect 3384 8395 3404 8415
rect 3487 8399 3507 8419
rect 5502 8473 5522 8493
rect 5612 8469 5632 8489
rect 5715 8473 5735 8493
rect 5820 8469 5840 8489
rect 5923 8473 5943 8493
rect 6031 8473 6051 8493
rect 6134 8469 6154 8489
rect 7808 8440 7828 8460
rect 7911 8436 7931 8456
rect 8019 8436 8039 8456
rect 8122 8440 8142 8460
rect 8227 8436 8247 8456
rect 8330 8440 8350 8460
rect 8440 8436 8460 8456
rect 8543 8440 8563 8460
rect 4795 8383 4813 8401
rect 117 8164 135 8182
rect 9851 8424 9869 8442
rect 5173 8205 5191 8223
rect 1423 8146 1443 8166
rect 1526 8150 1546 8170
rect 1636 8146 1656 8166
rect 1739 8150 1759 8170
rect 1844 8146 1864 8166
rect 1947 8150 1967 8170
rect 2055 8150 2075 8170
rect 2158 8146 2178 8166
rect 3832 8117 3852 8137
rect 3935 8113 3955 8133
rect 4043 8113 4063 8133
rect 4146 8117 4166 8137
rect 4251 8113 4271 8133
rect 4354 8117 4374 8137
rect 4464 8113 4484 8133
rect 6479 8187 6499 8207
rect 6582 8191 6602 8211
rect 6692 8187 6712 8207
rect 6795 8191 6815 8211
rect 6900 8187 6920 8207
rect 7003 8191 7023 8211
rect 7111 8191 7131 8211
rect 7214 8187 7234 8207
rect 8888 8158 8908 8178
rect 8991 8154 9011 8174
rect 9099 8154 9119 8174
rect 9202 8158 9222 8178
rect 9307 8154 9327 8174
rect 9410 8158 9430 8178
rect 9520 8154 9540 8174
rect 9623 8158 9643 8178
rect 4567 8117 4587 8137
rect 119 8065 137 8083
rect 117 7977 135 7995
rect 5175 8106 5193 8124
rect 119 7878 137 7896
rect 345 7879 365 7899
rect 448 7883 468 7903
rect 558 7879 578 7899
rect 661 7883 681 7903
rect 766 7879 786 7899
rect 869 7883 889 7903
rect 977 7883 997 7903
rect 1080 7879 1100 7899
rect 4794 8025 4812 8043
rect 5173 8018 5191 8036
rect 4796 7926 4814 7944
rect 5175 7919 5193 7937
rect 5401 7920 5421 7940
rect 5504 7924 5524 7944
rect 5614 7920 5634 7940
rect 5717 7924 5737 7944
rect 5822 7920 5842 7940
rect 5925 7924 5945 7944
rect 6033 7924 6053 7944
rect 6136 7920 6156 7940
rect 9850 8066 9868 8084
rect 9852 7967 9870 7985
rect 117 7748 135 7766
rect 2893 7807 2913 7827
rect 2996 7803 3016 7823
rect 3104 7803 3124 7823
rect 3207 7807 3227 7827
rect 3312 7803 3332 7823
rect 3415 7807 3435 7827
rect 3525 7803 3545 7823
rect 3628 7807 3648 7827
rect 119 7649 137 7667
rect 4794 7795 4812 7813
rect 5173 7789 5191 7807
rect 1283 7635 1303 7655
rect 1386 7639 1406 7659
rect 1496 7635 1516 7655
rect 1599 7639 1619 7659
rect 1704 7635 1724 7655
rect 1807 7639 1827 7659
rect 1915 7639 1935 7659
rect 2018 7635 2038 7655
rect 7949 7848 7969 7868
rect 8052 7844 8072 7864
rect 8160 7844 8180 7864
rect 8263 7848 8283 7868
rect 8368 7844 8388 7864
rect 8471 7848 8491 7868
rect 8581 7844 8601 7864
rect 8684 7848 8704 7868
rect 4796 7696 4814 7714
rect 5175 7690 5193 7708
rect 9850 7836 9868 7854
rect 6339 7676 6359 7696
rect 6442 7680 6462 7700
rect 6552 7676 6572 7696
rect 6655 7680 6675 7700
rect 6760 7676 6780 7696
rect 6863 7680 6883 7700
rect 6971 7680 6991 7700
rect 7074 7676 7094 7696
rect 9852 7737 9870 7755
rect 117 7518 135 7536
rect 119 7419 137 7437
rect 3831 7563 3851 7583
rect 3934 7559 3954 7579
rect 4042 7559 4062 7579
rect 4145 7563 4165 7583
rect 4250 7559 4270 7579
rect 4353 7563 4373 7583
rect 4463 7559 4483 7579
rect 4566 7563 4586 7583
rect 4794 7566 4812 7584
rect 5173 7559 5191 7577
rect 4796 7467 4814 7485
rect 5175 7460 5193 7478
rect 8887 7604 8907 7624
rect 8990 7600 9010 7620
rect 9098 7600 9118 7620
rect 9201 7604 9221 7624
rect 9306 7600 9326 7620
rect 9409 7604 9429 7624
rect 9519 7600 9539 7620
rect 9622 7604 9642 7624
rect 9850 7607 9868 7625
rect 4794 7379 4812 7397
rect 9852 7508 9870 7526
rect 9850 7420 9868 7438
rect 5400 7366 5420 7386
rect 344 7325 364 7345
rect 447 7329 467 7349
rect 557 7325 577 7345
rect 660 7329 680 7349
rect 765 7325 785 7345
rect 868 7329 888 7349
rect 976 7329 996 7349
rect 1079 7325 1099 7345
rect 2783 7283 2803 7303
rect 2886 7279 2906 7299
rect 2994 7279 3014 7299
rect 3097 7283 3117 7303
rect 3202 7279 3222 7299
rect 3305 7283 3325 7303
rect 3415 7279 3435 7299
rect 3518 7283 3538 7303
rect 5503 7370 5523 7390
rect 5613 7366 5633 7386
rect 5716 7370 5736 7390
rect 5821 7366 5841 7386
rect 5924 7370 5944 7390
rect 6032 7370 6052 7390
rect 6135 7366 6155 7386
rect 7839 7324 7859 7344
rect 4796 7280 4814 7298
rect 7942 7320 7962 7340
rect 8050 7320 8070 7340
rect 8153 7324 8173 7344
rect 8258 7320 8278 7340
rect 8361 7324 8381 7344
rect 8471 7320 8491 7340
rect 8574 7324 8594 7344
rect 9852 7321 9870 7339
rect 117 7061 135 7079
rect 1393 7056 1413 7076
rect 1496 7060 1516 7080
rect 1606 7056 1626 7076
rect 1709 7060 1729 7080
rect 1814 7056 1834 7076
rect 1917 7060 1937 7080
rect 2025 7060 2045 7080
rect 5173 7102 5191 7120
rect 2128 7056 2148 7076
rect 3832 7014 3852 7034
rect 3935 7010 3955 7030
rect 4043 7010 4063 7030
rect 4146 7014 4166 7034
rect 4251 7010 4271 7030
rect 4354 7014 4374 7034
rect 4464 7010 4484 7030
rect 6449 7097 6469 7117
rect 6552 7101 6572 7121
rect 6662 7097 6682 7117
rect 6765 7101 6785 7121
rect 6870 7097 6890 7117
rect 6973 7101 6993 7121
rect 7081 7101 7101 7121
rect 7184 7097 7204 7117
rect 8888 7055 8908 7075
rect 8991 7051 9011 7071
rect 9099 7051 9119 7071
rect 9202 7055 9222 7075
rect 9307 7051 9327 7071
rect 9410 7055 9430 7075
rect 9520 7051 9540 7071
rect 9623 7055 9643 7075
rect 4567 7014 4587 7034
rect 119 6962 137 6980
rect 117 6874 135 6892
rect 5175 7003 5193 7021
rect 119 6775 137 6793
rect 345 6776 365 6796
rect 448 6780 468 6800
rect 558 6776 578 6796
rect 661 6780 681 6800
rect 766 6776 786 6796
rect 869 6780 889 6800
rect 977 6780 997 6800
rect 1080 6776 1100 6796
rect 4794 6922 4812 6940
rect 5173 6915 5191 6933
rect 4796 6823 4814 6841
rect 5175 6816 5193 6834
rect 5401 6817 5421 6837
rect 5504 6821 5524 6841
rect 5614 6817 5634 6837
rect 5717 6821 5737 6841
rect 5822 6817 5842 6837
rect 5925 6821 5945 6841
rect 6033 6821 6053 6841
rect 6136 6817 6156 6837
rect 9850 6963 9868 6981
rect 9852 6864 9870 6882
rect 117 6645 135 6663
rect 2893 6704 2913 6724
rect 2996 6700 3016 6720
rect 3104 6700 3124 6720
rect 3207 6704 3227 6724
rect 3312 6700 3332 6720
rect 3415 6704 3435 6724
rect 3525 6700 3545 6720
rect 3628 6704 3648 6724
rect 119 6546 137 6564
rect 4794 6692 4812 6710
rect 5173 6686 5191 6704
rect 1283 6532 1303 6552
rect 1386 6536 1406 6556
rect 1496 6532 1516 6552
rect 1599 6536 1619 6556
rect 1704 6532 1724 6552
rect 1807 6536 1827 6556
rect 1915 6536 1935 6556
rect 2018 6532 2038 6552
rect 7949 6745 7969 6765
rect 8052 6741 8072 6761
rect 8160 6741 8180 6761
rect 8263 6745 8283 6765
rect 8368 6741 8388 6761
rect 8471 6745 8491 6765
rect 8581 6741 8601 6761
rect 8684 6745 8704 6765
rect 4796 6593 4814 6611
rect 5175 6587 5193 6605
rect 9850 6733 9868 6751
rect 6339 6573 6359 6593
rect 6442 6577 6462 6597
rect 6552 6573 6572 6593
rect 6655 6577 6675 6597
rect 6760 6573 6780 6593
rect 6863 6577 6883 6597
rect 6971 6577 6991 6597
rect 7074 6573 7094 6593
rect 9852 6634 9870 6652
rect 117 6415 135 6433
rect 119 6316 137 6334
rect 3831 6460 3851 6480
rect 3934 6456 3954 6476
rect 4042 6456 4062 6476
rect 4145 6460 4165 6480
rect 4250 6456 4270 6476
rect 4353 6460 4373 6480
rect 4463 6456 4483 6476
rect 4566 6460 4586 6480
rect 4794 6463 4812 6481
rect 5173 6456 5191 6474
rect 4796 6364 4814 6382
rect 5175 6357 5193 6375
rect 8887 6501 8907 6521
rect 8990 6497 9010 6517
rect 9098 6497 9118 6517
rect 9201 6501 9221 6521
rect 9306 6497 9326 6517
rect 9409 6501 9429 6521
rect 9519 6497 9539 6517
rect 9622 6501 9642 6521
rect 9850 6504 9868 6522
rect 4794 6276 4812 6294
rect 9852 6405 9870 6423
rect 9850 6317 9868 6335
rect 5400 6263 5420 6283
rect 344 6222 364 6242
rect 447 6226 467 6246
rect 557 6222 577 6242
rect 660 6226 680 6246
rect 765 6222 785 6242
rect 868 6226 888 6246
rect 976 6226 996 6246
rect 1079 6222 1099 6242
rect 2753 6193 2773 6213
rect 2856 6189 2876 6209
rect 2964 6189 2984 6209
rect 3067 6193 3087 6213
rect 3172 6189 3192 6209
rect 3275 6193 3295 6213
rect 3385 6189 3405 6209
rect 3488 6193 3508 6213
rect 5503 6267 5523 6287
rect 5613 6263 5633 6283
rect 5716 6267 5736 6287
rect 5821 6263 5841 6283
rect 5924 6267 5944 6287
rect 6032 6267 6052 6287
rect 6135 6263 6155 6283
rect 7809 6234 7829 6254
rect 7912 6230 7932 6250
rect 8020 6230 8040 6250
rect 8123 6234 8143 6254
rect 8228 6230 8248 6250
rect 8331 6234 8351 6254
rect 8441 6230 8461 6250
rect 8544 6234 8564 6254
rect 4796 6177 4814 6195
rect 118 5958 136 5976
rect 9852 6218 9870 6236
rect 5174 5999 5192 6017
rect 1424 5940 1444 5960
rect 1527 5944 1547 5964
rect 1637 5940 1657 5960
rect 1740 5944 1760 5964
rect 1845 5940 1865 5960
rect 1948 5944 1968 5964
rect 2056 5944 2076 5964
rect 2159 5940 2179 5960
rect 3833 5911 3853 5931
rect 3936 5907 3956 5927
rect 4044 5907 4064 5927
rect 4147 5911 4167 5931
rect 4252 5907 4272 5927
rect 4355 5911 4375 5931
rect 4465 5907 4485 5927
rect 6480 5981 6500 6001
rect 6583 5985 6603 6005
rect 6693 5981 6713 6001
rect 6796 5985 6816 6005
rect 6901 5981 6921 6001
rect 7004 5985 7024 6005
rect 7112 5985 7132 6005
rect 7215 5981 7235 6001
rect 8889 5952 8909 5972
rect 8992 5948 9012 5968
rect 9100 5948 9120 5968
rect 9203 5952 9223 5972
rect 9308 5948 9328 5968
rect 9411 5952 9431 5972
rect 9521 5948 9541 5968
rect 9624 5952 9644 5972
rect 4568 5911 4588 5931
rect 120 5859 138 5877
rect 118 5771 136 5789
rect 5176 5900 5194 5918
rect 120 5672 138 5690
rect 346 5673 366 5693
rect 449 5677 469 5697
rect 559 5673 579 5693
rect 662 5677 682 5697
rect 767 5673 787 5693
rect 870 5677 890 5697
rect 978 5677 998 5697
rect 1081 5673 1101 5693
rect 4795 5819 4813 5837
rect 5174 5812 5192 5830
rect 4797 5720 4815 5738
rect 5176 5713 5194 5731
rect 5402 5714 5422 5734
rect 5505 5718 5525 5738
rect 5615 5714 5635 5734
rect 5718 5718 5738 5738
rect 5823 5714 5843 5734
rect 5926 5718 5946 5738
rect 6034 5718 6054 5738
rect 6137 5714 6157 5734
rect 9851 5860 9869 5878
rect 9853 5761 9871 5779
rect 118 5542 136 5560
rect 2894 5601 2914 5621
rect 2997 5597 3017 5617
rect 3105 5597 3125 5617
rect 3208 5601 3228 5621
rect 3313 5597 3333 5617
rect 3416 5601 3436 5621
rect 3526 5597 3546 5617
rect 3629 5601 3649 5621
rect 120 5443 138 5461
rect 4795 5589 4813 5607
rect 5174 5583 5192 5601
rect 1284 5429 1304 5449
rect 1387 5433 1407 5453
rect 1497 5429 1517 5449
rect 1600 5433 1620 5453
rect 1705 5429 1725 5449
rect 1808 5433 1828 5453
rect 1916 5433 1936 5453
rect 2019 5429 2039 5449
rect 7950 5642 7970 5662
rect 8053 5638 8073 5658
rect 8161 5638 8181 5658
rect 8264 5642 8284 5662
rect 8369 5638 8389 5658
rect 8472 5642 8492 5662
rect 8582 5638 8602 5658
rect 8685 5642 8705 5662
rect 4797 5490 4815 5508
rect 5176 5484 5194 5502
rect 9851 5630 9869 5648
rect 6340 5470 6360 5490
rect 6443 5474 6463 5494
rect 6553 5470 6573 5490
rect 6656 5474 6676 5494
rect 6761 5470 6781 5490
rect 6864 5474 6884 5494
rect 6972 5474 6992 5494
rect 7075 5470 7095 5490
rect 9853 5531 9871 5549
rect 118 5312 136 5330
rect 120 5213 138 5231
rect 3832 5357 3852 5377
rect 3935 5353 3955 5373
rect 4043 5353 4063 5373
rect 4146 5357 4166 5377
rect 4251 5353 4271 5373
rect 4354 5357 4374 5377
rect 4464 5353 4484 5373
rect 4567 5357 4587 5377
rect 4795 5360 4813 5378
rect 5174 5353 5192 5371
rect 4797 5261 4815 5279
rect 5176 5254 5194 5272
rect 8888 5398 8908 5418
rect 8991 5394 9011 5414
rect 9099 5394 9119 5414
rect 9202 5398 9222 5418
rect 9307 5394 9327 5414
rect 9410 5398 9430 5418
rect 9520 5394 9540 5414
rect 9623 5398 9643 5418
rect 9851 5401 9869 5419
rect 4795 5173 4813 5191
rect 9853 5302 9871 5320
rect 9851 5214 9869 5232
rect 345 5119 365 5139
rect 448 5123 468 5143
rect 558 5119 578 5139
rect 661 5123 681 5143
rect 766 5119 786 5139
rect 869 5123 889 5143
rect 977 5123 997 5143
rect 1080 5119 1100 5139
rect 5401 5160 5421 5180
rect 2785 5071 2805 5091
rect 2888 5067 2908 5087
rect 2996 5067 3016 5087
rect 3099 5071 3119 5091
rect 3204 5067 3224 5087
rect 3307 5071 3327 5091
rect 3417 5067 3437 5087
rect 3520 5071 3540 5091
rect 5504 5164 5524 5184
rect 5614 5160 5634 5180
rect 5717 5164 5737 5184
rect 5822 5160 5842 5180
rect 5925 5164 5945 5184
rect 6033 5164 6053 5184
rect 6136 5160 6156 5180
rect 4797 5074 4815 5092
rect 7841 5112 7861 5132
rect 7944 5108 7964 5128
rect 8052 5108 8072 5128
rect 8155 5112 8175 5132
rect 8260 5108 8280 5128
rect 8363 5112 8383 5132
rect 8473 5108 8493 5128
rect 8576 5112 8596 5132
rect 9853 5115 9871 5133
rect 118 4855 136 4873
rect 1393 4856 1413 4876
rect 1496 4860 1516 4880
rect 1606 4856 1626 4876
rect 1709 4860 1729 4880
rect 1814 4856 1834 4876
rect 1917 4860 1937 4880
rect 2025 4860 2045 4880
rect 2128 4856 2148 4876
rect 5174 4896 5192 4914
rect 3833 4808 3853 4828
rect 3936 4804 3956 4824
rect 4044 4804 4064 4824
rect 4147 4808 4167 4828
rect 4252 4804 4272 4824
rect 4355 4808 4375 4828
rect 4465 4804 4485 4824
rect 6449 4897 6469 4917
rect 6552 4901 6572 4921
rect 6662 4897 6682 4917
rect 6765 4901 6785 4921
rect 6870 4897 6890 4917
rect 6973 4901 6993 4921
rect 7081 4901 7101 4921
rect 7184 4897 7204 4917
rect 4568 4808 4588 4828
rect 8889 4849 8909 4869
rect 8992 4845 9012 4865
rect 9100 4845 9120 4865
rect 9203 4849 9223 4869
rect 9308 4845 9328 4865
rect 9411 4849 9431 4869
rect 9521 4845 9541 4865
rect 9624 4849 9644 4869
rect 120 4756 138 4774
rect 118 4668 136 4686
rect 5176 4797 5194 4815
rect 120 4569 138 4587
rect 346 4570 366 4590
rect 449 4574 469 4594
rect 559 4570 579 4590
rect 662 4574 682 4594
rect 767 4570 787 4590
rect 870 4574 890 4594
rect 978 4574 998 4594
rect 1081 4570 1101 4590
rect 4795 4716 4813 4734
rect 5174 4709 5192 4727
rect 4797 4617 4815 4635
rect 5176 4610 5194 4628
rect 5402 4611 5422 4631
rect 5505 4615 5525 4635
rect 5615 4611 5635 4631
rect 5718 4615 5738 4635
rect 5823 4611 5843 4631
rect 5926 4615 5946 4635
rect 6034 4615 6054 4635
rect 6137 4611 6157 4631
rect 9851 4757 9869 4775
rect 9853 4658 9871 4676
rect 118 4439 136 4457
rect 2894 4498 2914 4518
rect 2997 4494 3017 4514
rect 3105 4494 3125 4514
rect 3208 4498 3228 4518
rect 3313 4494 3333 4514
rect 3416 4498 3436 4518
rect 3526 4494 3546 4514
rect 3629 4498 3649 4518
rect 120 4340 138 4358
rect 4795 4486 4813 4504
rect 5174 4480 5192 4498
rect 1284 4326 1304 4346
rect 1387 4330 1407 4350
rect 1497 4326 1517 4346
rect 1600 4330 1620 4350
rect 1705 4326 1725 4346
rect 1808 4330 1828 4350
rect 1916 4330 1936 4350
rect 2019 4326 2039 4346
rect 7950 4539 7970 4559
rect 8053 4535 8073 4555
rect 8161 4535 8181 4555
rect 8264 4539 8284 4559
rect 8369 4535 8389 4555
rect 8472 4539 8492 4559
rect 8582 4535 8602 4555
rect 8685 4539 8705 4559
rect 4797 4387 4815 4405
rect 5176 4381 5194 4399
rect 9851 4527 9869 4545
rect 6340 4367 6360 4387
rect 6443 4371 6463 4391
rect 6553 4367 6573 4387
rect 6656 4371 6676 4391
rect 6761 4367 6781 4387
rect 6864 4371 6884 4391
rect 6972 4371 6992 4391
rect 7075 4367 7095 4387
rect 9853 4428 9871 4446
rect 118 4209 136 4227
rect 120 4110 138 4128
rect 3832 4254 3852 4274
rect 3935 4250 3955 4270
rect 4043 4250 4063 4270
rect 4146 4254 4166 4274
rect 4251 4250 4271 4270
rect 4354 4254 4374 4274
rect 4464 4250 4484 4270
rect 4567 4254 4587 4274
rect 4795 4257 4813 4275
rect 5174 4250 5192 4268
rect 4797 4158 4815 4176
rect 5176 4151 5194 4169
rect 8888 4295 8908 4315
rect 8991 4291 9011 4311
rect 9099 4291 9119 4311
rect 9202 4295 9222 4315
rect 9307 4291 9327 4311
rect 9410 4295 9430 4315
rect 9520 4291 9540 4311
rect 9623 4295 9643 4315
rect 9851 4298 9869 4316
rect 4795 4070 4813 4088
rect 9853 4199 9871 4217
rect 9851 4111 9869 4129
rect 5401 4057 5421 4077
rect 345 4016 365 4036
rect 448 4020 468 4040
rect 558 4016 578 4036
rect 661 4020 681 4040
rect 766 4016 786 4036
rect 869 4020 889 4040
rect 977 4020 997 4040
rect 1080 4016 1100 4036
rect 2754 3987 2774 4007
rect 2857 3983 2877 4003
rect 2965 3983 2985 4003
rect 3068 3987 3088 4007
rect 3173 3983 3193 4003
rect 3276 3987 3296 4007
rect 3386 3983 3406 4003
rect 3489 3987 3509 4007
rect 5504 4061 5524 4081
rect 5614 4057 5634 4077
rect 5717 4061 5737 4081
rect 5822 4057 5842 4077
rect 5925 4061 5945 4081
rect 6033 4061 6053 4081
rect 6136 4057 6156 4077
rect 7810 4028 7830 4048
rect 7913 4024 7933 4044
rect 8021 4024 8041 4044
rect 8124 4028 8144 4048
rect 8229 4024 8249 4044
rect 8332 4028 8352 4048
rect 8442 4024 8462 4044
rect 8545 4028 8565 4048
rect 4797 3971 4815 3989
rect 119 3752 137 3770
rect 9853 4012 9871 4030
rect 5175 3793 5193 3811
rect 1425 3734 1445 3754
rect 1528 3738 1548 3758
rect 1638 3734 1658 3754
rect 1741 3738 1761 3758
rect 1846 3734 1866 3754
rect 1949 3738 1969 3758
rect 2057 3738 2077 3758
rect 2160 3734 2180 3754
rect 3834 3705 3854 3725
rect 3937 3701 3957 3721
rect 4045 3701 4065 3721
rect 4148 3705 4168 3725
rect 4253 3701 4273 3721
rect 4356 3705 4376 3725
rect 4466 3701 4486 3721
rect 6481 3775 6501 3795
rect 6584 3779 6604 3799
rect 6694 3775 6714 3795
rect 6797 3779 6817 3799
rect 6902 3775 6922 3795
rect 7005 3779 7025 3799
rect 7113 3779 7133 3799
rect 7216 3775 7236 3795
rect 8890 3746 8910 3766
rect 8993 3742 9013 3762
rect 9101 3742 9121 3762
rect 9204 3746 9224 3766
rect 9309 3742 9329 3762
rect 9412 3746 9432 3766
rect 9522 3742 9542 3762
rect 9625 3746 9645 3766
rect 4569 3705 4589 3725
rect 121 3653 139 3671
rect 119 3565 137 3583
rect 5177 3694 5195 3712
rect 121 3466 139 3484
rect 347 3467 367 3487
rect 450 3471 470 3491
rect 560 3467 580 3487
rect 663 3471 683 3491
rect 768 3467 788 3487
rect 871 3471 891 3491
rect 979 3471 999 3491
rect 1082 3467 1102 3487
rect 4796 3613 4814 3631
rect 5175 3606 5193 3624
rect 4798 3514 4816 3532
rect 5177 3507 5195 3525
rect 5403 3508 5423 3528
rect 5506 3512 5526 3532
rect 5616 3508 5636 3528
rect 5719 3512 5739 3532
rect 5824 3508 5844 3528
rect 5927 3512 5947 3532
rect 6035 3512 6055 3532
rect 6138 3508 6158 3528
rect 9852 3654 9870 3672
rect 9854 3555 9872 3573
rect 119 3336 137 3354
rect 2895 3395 2915 3415
rect 2998 3391 3018 3411
rect 3106 3391 3126 3411
rect 3209 3395 3229 3415
rect 3314 3391 3334 3411
rect 3417 3395 3437 3415
rect 3527 3391 3547 3411
rect 3630 3395 3650 3415
rect 121 3237 139 3255
rect 4796 3383 4814 3401
rect 5175 3377 5193 3395
rect 1285 3223 1305 3243
rect 1388 3227 1408 3247
rect 1498 3223 1518 3243
rect 1601 3227 1621 3247
rect 1706 3223 1726 3243
rect 1809 3227 1829 3247
rect 1917 3227 1937 3247
rect 2020 3223 2040 3243
rect 7951 3436 7971 3456
rect 8054 3432 8074 3452
rect 8162 3432 8182 3452
rect 8265 3436 8285 3456
rect 8370 3432 8390 3452
rect 8473 3436 8493 3456
rect 8583 3432 8603 3452
rect 8686 3436 8706 3456
rect 4798 3284 4816 3302
rect 5177 3278 5195 3296
rect 9852 3424 9870 3442
rect 6341 3264 6361 3284
rect 6444 3268 6464 3288
rect 6554 3264 6574 3284
rect 6657 3268 6677 3288
rect 6762 3264 6782 3284
rect 6865 3268 6885 3288
rect 6973 3268 6993 3288
rect 7076 3264 7096 3284
rect 9854 3325 9872 3343
rect 119 3106 137 3124
rect 121 3007 139 3025
rect 3833 3151 3853 3171
rect 3936 3147 3956 3167
rect 4044 3147 4064 3167
rect 4147 3151 4167 3171
rect 4252 3147 4272 3167
rect 4355 3151 4375 3171
rect 4465 3147 4485 3167
rect 4568 3151 4588 3171
rect 4796 3154 4814 3172
rect 5175 3147 5193 3165
rect 4798 3055 4816 3073
rect 5177 3048 5195 3066
rect 8889 3192 8909 3212
rect 8992 3188 9012 3208
rect 9100 3188 9120 3208
rect 9203 3192 9223 3212
rect 9308 3188 9328 3208
rect 9411 3192 9431 3212
rect 9521 3188 9541 3208
rect 9624 3192 9644 3212
rect 9852 3195 9870 3213
rect 4796 2967 4814 2985
rect 9854 3096 9872 3114
rect 9852 3008 9870 3026
rect 5402 2954 5422 2974
rect 346 2913 366 2933
rect 449 2917 469 2937
rect 559 2913 579 2933
rect 662 2917 682 2937
rect 767 2913 787 2933
rect 870 2917 890 2937
rect 978 2917 998 2937
rect 1081 2913 1101 2933
rect 2785 2871 2805 2891
rect 2888 2867 2908 2887
rect 2996 2867 3016 2887
rect 3099 2871 3119 2891
rect 3204 2867 3224 2887
rect 3307 2871 3327 2891
rect 3417 2867 3437 2887
rect 3520 2871 3540 2891
rect 5505 2958 5525 2978
rect 5615 2954 5635 2974
rect 5718 2958 5738 2978
rect 5823 2954 5843 2974
rect 5926 2958 5946 2978
rect 6034 2958 6054 2978
rect 6137 2954 6157 2974
rect 7841 2912 7861 2932
rect 4798 2868 4816 2886
rect 7944 2908 7964 2928
rect 8052 2908 8072 2928
rect 8155 2912 8175 2932
rect 8260 2908 8280 2928
rect 8363 2912 8383 2932
rect 8473 2908 8493 2928
rect 8576 2912 8596 2932
rect 9854 2909 9872 2927
rect 119 2649 137 2667
rect 1395 2644 1415 2664
rect 1498 2648 1518 2668
rect 1608 2644 1628 2664
rect 1711 2648 1731 2668
rect 1816 2644 1836 2664
rect 1919 2648 1939 2668
rect 2027 2648 2047 2668
rect 5175 2690 5193 2708
rect 2130 2644 2150 2664
rect 3834 2602 3854 2622
rect 3937 2598 3957 2618
rect 4045 2598 4065 2618
rect 4148 2602 4168 2622
rect 4253 2598 4273 2618
rect 4356 2602 4376 2622
rect 4466 2598 4486 2618
rect 6451 2685 6471 2705
rect 6554 2689 6574 2709
rect 6664 2685 6684 2705
rect 6767 2689 6787 2709
rect 6872 2685 6892 2705
rect 6975 2689 6995 2709
rect 7083 2689 7103 2709
rect 7186 2685 7206 2705
rect 8890 2643 8910 2663
rect 8993 2639 9013 2659
rect 9101 2639 9121 2659
rect 9204 2643 9224 2663
rect 9309 2639 9329 2659
rect 9412 2643 9432 2663
rect 9522 2639 9542 2659
rect 9625 2643 9645 2663
rect 4569 2602 4589 2622
rect 121 2550 139 2568
rect 119 2462 137 2480
rect 5177 2591 5195 2609
rect 121 2363 139 2381
rect 347 2364 367 2384
rect 450 2368 470 2388
rect 560 2364 580 2384
rect 663 2368 683 2388
rect 768 2364 788 2384
rect 871 2368 891 2388
rect 979 2368 999 2388
rect 1082 2364 1102 2384
rect 4796 2510 4814 2528
rect 5175 2503 5193 2521
rect 4798 2411 4816 2429
rect 5177 2404 5195 2422
rect 5403 2405 5423 2425
rect 5506 2409 5526 2429
rect 5616 2405 5636 2425
rect 5719 2409 5739 2429
rect 5824 2405 5844 2425
rect 5927 2409 5947 2429
rect 6035 2409 6055 2429
rect 6138 2405 6158 2425
rect 9852 2551 9870 2569
rect 9854 2452 9872 2470
rect 119 2233 137 2251
rect 2895 2292 2915 2312
rect 2998 2288 3018 2308
rect 3106 2288 3126 2308
rect 3209 2292 3229 2312
rect 3314 2288 3334 2308
rect 3417 2292 3437 2312
rect 3527 2288 3547 2308
rect 3630 2292 3650 2312
rect 121 2134 139 2152
rect 4796 2280 4814 2298
rect 5175 2274 5193 2292
rect 1285 2120 1305 2140
rect 1388 2124 1408 2144
rect 1498 2120 1518 2140
rect 1601 2124 1621 2144
rect 1706 2120 1726 2140
rect 1809 2124 1829 2144
rect 1917 2124 1937 2144
rect 2020 2120 2040 2140
rect 7951 2333 7971 2353
rect 8054 2329 8074 2349
rect 8162 2329 8182 2349
rect 8265 2333 8285 2353
rect 8370 2329 8390 2349
rect 8473 2333 8493 2353
rect 8583 2329 8603 2349
rect 8686 2333 8706 2353
rect 4798 2181 4816 2199
rect 5177 2175 5195 2193
rect 9852 2321 9870 2339
rect 6341 2161 6361 2181
rect 6444 2165 6464 2185
rect 6554 2161 6574 2181
rect 6657 2165 6677 2185
rect 6762 2161 6782 2181
rect 6865 2165 6885 2185
rect 6973 2165 6993 2185
rect 7076 2161 7096 2181
rect 9854 2222 9872 2240
rect 119 2003 137 2021
rect 121 1904 139 1922
rect 3833 2048 3853 2068
rect 3936 2044 3956 2064
rect 4044 2044 4064 2064
rect 4147 2048 4167 2068
rect 4252 2044 4272 2064
rect 4355 2048 4375 2068
rect 4465 2044 4485 2064
rect 4568 2048 4588 2068
rect 4796 2051 4814 2069
rect 5175 2044 5193 2062
rect 4798 1952 4816 1970
rect 5177 1945 5195 1963
rect 8889 2089 8909 2109
rect 8992 2085 9012 2105
rect 9100 2085 9120 2105
rect 9203 2089 9223 2109
rect 9308 2085 9328 2105
rect 9411 2089 9431 2109
rect 9521 2085 9541 2105
rect 9624 2089 9644 2109
rect 9852 2092 9870 2110
rect 4796 1864 4814 1882
rect 9854 1993 9872 2011
rect 9852 1905 9870 1923
rect 5402 1851 5422 1871
rect 346 1810 366 1830
rect 449 1814 469 1834
rect 559 1810 579 1830
rect 662 1814 682 1834
rect 767 1810 787 1830
rect 870 1814 890 1834
rect 978 1814 998 1834
rect 1081 1810 1101 1830
rect 2755 1781 2775 1801
rect 2858 1777 2878 1797
rect 2966 1777 2986 1797
rect 3069 1781 3089 1801
rect 3174 1777 3194 1797
rect 3277 1781 3297 1801
rect 3387 1777 3407 1797
rect 3490 1781 3510 1801
rect 5505 1855 5525 1875
rect 5615 1851 5635 1871
rect 5718 1855 5738 1875
rect 5823 1851 5843 1871
rect 5926 1855 5946 1875
rect 6034 1855 6054 1875
rect 6137 1851 6157 1871
rect 7811 1822 7831 1842
rect 7914 1818 7934 1838
rect 8022 1818 8042 1838
rect 8125 1822 8145 1842
rect 8230 1818 8250 1838
rect 8333 1822 8353 1842
rect 8443 1818 8463 1838
rect 8546 1822 8566 1842
rect 4798 1765 4816 1783
rect 120 1546 138 1564
rect 9854 1806 9872 1824
rect 5176 1587 5194 1605
rect 1426 1528 1446 1548
rect 1529 1532 1549 1552
rect 1639 1528 1659 1548
rect 1742 1532 1762 1552
rect 1847 1528 1867 1548
rect 1950 1532 1970 1552
rect 2058 1532 2078 1552
rect 2161 1528 2181 1548
rect 3835 1499 3855 1519
rect 3938 1495 3958 1515
rect 4046 1495 4066 1515
rect 4149 1499 4169 1519
rect 4254 1495 4274 1515
rect 4357 1499 4377 1519
rect 4467 1495 4487 1515
rect 6482 1569 6502 1589
rect 6585 1573 6605 1593
rect 6695 1569 6715 1589
rect 6798 1573 6818 1593
rect 6903 1569 6923 1589
rect 7006 1573 7026 1593
rect 7114 1573 7134 1593
rect 7217 1569 7237 1589
rect 8891 1540 8911 1560
rect 8994 1536 9014 1556
rect 9102 1536 9122 1556
rect 9205 1540 9225 1560
rect 9310 1536 9330 1556
rect 9413 1540 9433 1560
rect 9523 1536 9543 1556
rect 9626 1540 9646 1560
rect 4570 1499 4590 1519
rect 122 1447 140 1465
rect 120 1359 138 1377
rect 5178 1488 5196 1506
rect 122 1260 140 1278
rect 348 1261 368 1281
rect 451 1265 471 1285
rect 561 1261 581 1281
rect 664 1265 684 1285
rect 769 1261 789 1281
rect 872 1265 892 1285
rect 980 1265 1000 1285
rect 1083 1261 1103 1281
rect 4797 1407 4815 1425
rect 5176 1400 5194 1418
rect 4799 1308 4817 1326
rect 5178 1301 5196 1319
rect 5404 1302 5424 1322
rect 5507 1306 5527 1326
rect 5617 1302 5637 1322
rect 5720 1306 5740 1326
rect 5825 1302 5845 1322
rect 5928 1306 5948 1326
rect 6036 1306 6056 1326
rect 6139 1302 6159 1322
rect 9853 1448 9871 1466
rect 9855 1349 9873 1367
rect 120 1130 138 1148
rect 2896 1189 2916 1209
rect 2999 1185 3019 1205
rect 3107 1185 3127 1205
rect 3210 1189 3230 1209
rect 3315 1185 3335 1205
rect 3418 1189 3438 1209
rect 3528 1185 3548 1205
rect 3631 1189 3651 1209
rect 122 1031 140 1049
rect 4797 1177 4815 1195
rect 5176 1171 5194 1189
rect 1286 1017 1306 1037
rect 1389 1021 1409 1041
rect 1499 1017 1519 1037
rect 1602 1021 1622 1041
rect 1707 1017 1727 1037
rect 1810 1021 1830 1041
rect 1918 1021 1938 1041
rect 2021 1017 2041 1037
rect 7952 1230 7972 1250
rect 8055 1226 8075 1246
rect 8163 1226 8183 1246
rect 8266 1230 8286 1250
rect 8371 1226 8391 1246
rect 8474 1230 8494 1250
rect 8584 1226 8604 1246
rect 8687 1230 8707 1250
rect 4799 1078 4817 1096
rect 5178 1072 5196 1090
rect 9853 1218 9871 1236
rect 6342 1058 6362 1078
rect 6445 1062 6465 1082
rect 6555 1058 6575 1078
rect 6658 1062 6678 1082
rect 6763 1058 6783 1078
rect 6866 1062 6886 1082
rect 6974 1062 6994 1082
rect 7077 1058 7097 1078
rect 9855 1119 9873 1137
rect 120 900 138 918
rect 122 801 140 819
rect 3834 945 3854 965
rect 3937 941 3957 961
rect 4045 941 4065 961
rect 4148 945 4168 965
rect 4253 941 4273 961
rect 4356 945 4376 965
rect 4466 941 4486 961
rect 4569 945 4589 965
rect 4797 948 4815 966
rect 5176 941 5194 959
rect 4799 849 4817 867
rect 5178 842 5196 860
rect 8890 986 8910 1006
rect 8993 982 9013 1002
rect 9101 982 9121 1002
rect 9204 986 9224 1006
rect 9309 982 9329 1002
rect 9412 986 9432 1006
rect 9522 982 9542 1002
rect 9625 986 9645 1006
rect 9853 989 9871 1007
rect 4797 761 4815 779
rect 9855 890 9873 908
rect 9853 802 9871 820
rect 5403 748 5423 768
rect 347 707 367 727
rect 450 711 470 731
rect 560 707 580 727
rect 663 711 683 731
rect 768 707 788 727
rect 871 711 891 731
rect 979 711 999 731
rect 1082 707 1102 727
rect 5506 752 5526 772
rect 5616 748 5636 768
rect 5719 752 5739 772
rect 5824 748 5844 768
rect 5927 752 5947 772
rect 6035 752 6055 772
rect 6138 748 6158 768
rect 9855 703 9873 721
rect 4799 662 4817 680
rect 1594 148 1614 168
rect 1697 152 1717 172
rect 1807 148 1827 168
rect 1910 152 1930 172
rect 2015 148 2035 168
rect 2118 152 2138 172
rect 2226 152 2246 172
rect 2329 148 2349 168
rect 6650 189 6670 209
rect 6753 193 6773 213
rect 6863 189 6883 209
rect 6966 193 6986 213
rect 7071 189 7091 209
rect 7174 193 7194 213
rect 7282 193 7302 213
rect 7385 189 7405 209
rect 4544 128 4564 148
rect 4647 132 4667 152
rect 4757 128 4777 148
rect 4860 132 4880 152
rect 4965 128 4985 148
rect 5068 132 5088 152
rect 5176 132 5196 152
rect 5279 128 5299 148
<< pdiffc >>
rect 350 9131 370 9151
rect 446 9131 466 9151
rect 563 9131 583 9151
rect 659 9131 679 9151
rect 771 9131 791 9151
rect 867 9131 887 9151
rect 977 9131 997 9151
rect 1073 9131 1093 9151
rect 5406 9172 5426 9192
rect 3837 9071 3857 9091
rect 3933 9071 3953 9091
rect 4043 9071 4063 9091
rect 4139 9071 4159 9091
rect 4251 9071 4271 9091
rect 4347 9071 4367 9091
rect 4464 9071 4484 9091
rect 5502 9172 5522 9192
rect 5619 9172 5639 9192
rect 5715 9172 5735 9192
rect 5827 9172 5847 9192
rect 5923 9172 5943 9192
rect 6033 9172 6053 9192
rect 6129 9172 6149 9192
rect 4560 9071 4580 9091
rect 8893 9112 8913 9132
rect 8989 9112 9009 9132
rect 9099 9112 9119 9132
rect 9195 9112 9215 9132
rect 9307 9112 9327 9132
rect 9403 9112 9423 9132
rect 9520 9112 9540 9132
rect 9616 9112 9636 9132
rect 1288 8887 1308 8907
rect 1384 8887 1404 8907
rect 1501 8887 1521 8907
rect 1597 8887 1617 8907
rect 1709 8887 1729 8907
rect 1805 8887 1825 8907
rect 1915 8887 1935 8907
rect 2011 8887 2031 8907
rect 6344 8928 6364 8948
rect 2898 8761 2918 8781
rect 2994 8761 3014 8781
rect 3104 8761 3124 8781
rect 3200 8761 3220 8781
rect 3312 8761 3332 8781
rect 3408 8761 3428 8781
rect 3525 8761 3545 8781
rect 6440 8928 6460 8948
rect 6557 8928 6577 8948
rect 6653 8928 6673 8948
rect 6765 8928 6785 8948
rect 6861 8928 6881 8948
rect 6971 8928 6991 8948
rect 7067 8928 7087 8948
rect 3621 8761 3641 8781
rect 7954 8802 7974 8822
rect 8050 8802 8070 8822
rect 8160 8802 8180 8822
rect 8256 8802 8276 8822
rect 8368 8802 8388 8822
rect 8464 8802 8484 8822
rect 8581 8802 8601 8822
rect 8677 8802 8697 8822
rect 349 8577 369 8597
rect 445 8577 465 8597
rect 562 8577 582 8597
rect 658 8577 678 8597
rect 770 8577 790 8597
rect 866 8577 886 8597
rect 976 8577 996 8597
rect 1072 8577 1092 8597
rect 5405 8618 5425 8638
rect 3836 8517 3856 8537
rect 3932 8517 3952 8537
rect 4042 8517 4062 8537
rect 4138 8517 4158 8537
rect 4250 8517 4270 8537
rect 4346 8517 4366 8537
rect 4463 8517 4483 8537
rect 5501 8618 5521 8638
rect 5618 8618 5638 8638
rect 5714 8618 5734 8638
rect 5826 8618 5846 8638
rect 5922 8618 5942 8638
rect 6032 8618 6052 8638
rect 6128 8618 6148 8638
rect 4559 8517 4579 8537
rect 8892 8558 8912 8578
rect 8988 8558 9008 8578
rect 9098 8558 9118 8578
rect 9194 8558 9214 8578
rect 9306 8558 9326 8578
rect 9402 8558 9422 8578
rect 9519 8558 9539 8578
rect 9615 8558 9635 8578
rect 1429 8295 1449 8315
rect 1525 8295 1545 8315
rect 1642 8295 1662 8315
rect 1738 8295 1758 8315
rect 1850 8295 1870 8315
rect 1946 8295 1966 8315
rect 2056 8295 2076 8315
rect 2152 8295 2172 8315
rect 6485 8336 6505 8356
rect 2758 8250 2778 8270
rect 2854 8250 2874 8270
rect 2964 8250 2984 8270
rect 3060 8250 3080 8270
rect 3172 8250 3192 8270
rect 3268 8250 3288 8270
rect 3385 8250 3405 8270
rect 6581 8336 6601 8356
rect 6698 8336 6718 8356
rect 6794 8336 6814 8356
rect 6906 8336 6926 8356
rect 7002 8336 7022 8356
rect 7112 8336 7132 8356
rect 7208 8336 7228 8356
rect 3481 8250 3501 8270
rect 7814 8291 7834 8311
rect 7910 8291 7930 8311
rect 8020 8291 8040 8311
rect 8116 8291 8136 8311
rect 8228 8291 8248 8311
rect 8324 8291 8344 8311
rect 8441 8291 8461 8311
rect 8537 8291 8557 8311
rect 351 8028 371 8048
rect 447 8028 467 8048
rect 564 8028 584 8048
rect 660 8028 680 8048
rect 772 8028 792 8048
rect 868 8028 888 8048
rect 978 8028 998 8048
rect 1074 8028 1094 8048
rect 5407 8069 5427 8089
rect 3838 7968 3858 7988
rect 3934 7968 3954 7988
rect 4044 7968 4064 7988
rect 4140 7968 4160 7988
rect 4252 7968 4272 7988
rect 4348 7968 4368 7988
rect 4465 7968 4485 7988
rect 5503 8069 5523 8089
rect 5620 8069 5640 8089
rect 5716 8069 5736 8089
rect 5828 8069 5848 8089
rect 5924 8069 5944 8089
rect 6034 8069 6054 8089
rect 6130 8069 6150 8089
rect 4561 7968 4581 7988
rect 8894 8009 8914 8029
rect 8990 8009 9010 8029
rect 9100 8009 9120 8029
rect 9196 8009 9216 8029
rect 9308 8009 9328 8029
rect 9404 8009 9424 8029
rect 9521 8009 9541 8029
rect 9617 8009 9637 8029
rect 1289 7784 1309 7804
rect 1385 7784 1405 7804
rect 1502 7784 1522 7804
rect 1598 7784 1618 7804
rect 1710 7784 1730 7804
rect 1806 7784 1826 7804
rect 1916 7784 1936 7804
rect 2012 7784 2032 7804
rect 6345 7825 6365 7845
rect 2899 7658 2919 7678
rect 2995 7658 3015 7678
rect 3105 7658 3125 7678
rect 3201 7658 3221 7678
rect 3313 7658 3333 7678
rect 3409 7658 3429 7678
rect 3526 7658 3546 7678
rect 6441 7825 6461 7845
rect 6558 7825 6578 7845
rect 6654 7825 6674 7845
rect 6766 7825 6786 7845
rect 6862 7825 6882 7845
rect 6972 7825 6992 7845
rect 7068 7825 7088 7845
rect 3622 7658 3642 7678
rect 7955 7699 7975 7719
rect 8051 7699 8071 7719
rect 8161 7699 8181 7719
rect 8257 7699 8277 7719
rect 8369 7699 8389 7719
rect 8465 7699 8485 7719
rect 8582 7699 8602 7719
rect 8678 7699 8698 7719
rect 350 7474 370 7494
rect 446 7474 466 7494
rect 563 7474 583 7494
rect 659 7474 679 7494
rect 771 7474 791 7494
rect 867 7474 887 7494
rect 977 7474 997 7494
rect 1073 7474 1093 7494
rect 5406 7515 5426 7535
rect 3837 7414 3857 7434
rect 3933 7414 3953 7434
rect 4043 7414 4063 7434
rect 4139 7414 4159 7434
rect 4251 7414 4271 7434
rect 4347 7414 4367 7434
rect 4464 7414 4484 7434
rect 5502 7515 5522 7535
rect 5619 7515 5639 7535
rect 5715 7515 5735 7535
rect 5827 7515 5847 7535
rect 5923 7515 5943 7535
rect 6033 7515 6053 7535
rect 6129 7515 6149 7535
rect 4560 7414 4580 7434
rect 8893 7455 8913 7475
rect 8989 7455 9009 7475
rect 9099 7455 9119 7475
rect 9195 7455 9215 7475
rect 9307 7455 9327 7475
rect 9403 7455 9423 7475
rect 9520 7455 9540 7475
rect 9616 7455 9636 7475
rect 1399 7205 1419 7225
rect 1495 7205 1515 7225
rect 1612 7205 1632 7225
rect 1708 7205 1728 7225
rect 1820 7205 1840 7225
rect 1916 7205 1936 7225
rect 2026 7205 2046 7225
rect 2122 7205 2142 7225
rect 6455 7246 6475 7266
rect 6551 7246 6571 7266
rect 6668 7246 6688 7266
rect 6764 7246 6784 7266
rect 6876 7246 6896 7266
rect 6972 7246 6992 7266
rect 7082 7246 7102 7266
rect 7178 7246 7198 7266
rect 2789 7134 2809 7154
rect 2885 7134 2905 7154
rect 2995 7134 3015 7154
rect 3091 7134 3111 7154
rect 3203 7134 3223 7154
rect 3299 7134 3319 7154
rect 3416 7134 3436 7154
rect 3512 7134 3532 7154
rect 7845 7175 7865 7195
rect 7941 7175 7961 7195
rect 8051 7175 8071 7195
rect 8147 7175 8167 7195
rect 8259 7175 8279 7195
rect 8355 7175 8375 7195
rect 8472 7175 8492 7195
rect 8568 7175 8588 7195
rect 351 6925 371 6945
rect 447 6925 467 6945
rect 564 6925 584 6945
rect 660 6925 680 6945
rect 772 6925 792 6945
rect 868 6925 888 6945
rect 978 6925 998 6945
rect 1074 6925 1094 6945
rect 5407 6966 5427 6986
rect 3838 6865 3858 6885
rect 3934 6865 3954 6885
rect 4044 6865 4064 6885
rect 4140 6865 4160 6885
rect 4252 6865 4272 6885
rect 4348 6865 4368 6885
rect 4465 6865 4485 6885
rect 5503 6966 5523 6986
rect 5620 6966 5640 6986
rect 5716 6966 5736 6986
rect 5828 6966 5848 6986
rect 5924 6966 5944 6986
rect 6034 6966 6054 6986
rect 6130 6966 6150 6986
rect 4561 6865 4581 6885
rect 8894 6906 8914 6926
rect 8990 6906 9010 6926
rect 9100 6906 9120 6926
rect 9196 6906 9216 6926
rect 9308 6906 9328 6926
rect 9404 6906 9424 6926
rect 9521 6906 9541 6926
rect 9617 6906 9637 6926
rect 1289 6681 1309 6701
rect 1385 6681 1405 6701
rect 1502 6681 1522 6701
rect 1598 6681 1618 6701
rect 1710 6681 1730 6701
rect 1806 6681 1826 6701
rect 1916 6681 1936 6701
rect 2012 6681 2032 6701
rect 6345 6722 6365 6742
rect 2899 6555 2919 6575
rect 2995 6555 3015 6575
rect 3105 6555 3125 6575
rect 3201 6555 3221 6575
rect 3313 6555 3333 6575
rect 3409 6555 3429 6575
rect 3526 6555 3546 6575
rect 6441 6722 6461 6742
rect 6558 6722 6578 6742
rect 6654 6722 6674 6742
rect 6766 6722 6786 6742
rect 6862 6722 6882 6742
rect 6972 6722 6992 6742
rect 7068 6722 7088 6742
rect 3622 6555 3642 6575
rect 7955 6596 7975 6616
rect 8051 6596 8071 6616
rect 8161 6596 8181 6616
rect 8257 6596 8277 6616
rect 8369 6596 8389 6616
rect 8465 6596 8485 6616
rect 8582 6596 8602 6616
rect 8678 6596 8698 6616
rect 350 6371 370 6391
rect 446 6371 466 6391
rect 563 6371 583 6391
rect 659 6371 679 6391
rect 771 6371 791 6391
rect 867 6371 887 6391
rect 977 6371 997 6391
rect 1073 6371 1093 6391
rect 5406 6412 5426 6432
rect 3837 6311 3857 6331
rect 3933 6311 3953 6331
rect 4043 6311 4063 6331
rect 4139 6311 4159 6331
rect 4251 6311 4271 6331
rect 4347 6311 4367 6331
rect 4464 6311 4484 6331
rect 5502 6412 5522 6432
rect 5619 6412 5639 6432
rect 5715 6412 5735 6432
rect 5827 6412 5847 6432
rect 5923 6412 5943 6432
rect 6033 6412 6053 6432
rect 6129 6412 6149 6432
rect 4560 6311 4580 6331
rect 8893 6352 8913 6372
rect 8989 6352 9009 6372
rect 9099 6352 9119 6372
rect 9195 6352 9215 6372
rect 9307 6352 9327 6372
rect 9403 6352 9423 6372
rect 9520 6352 9540 6372
rect 9616 6352 9636 6372
rect 1430 6089 1450 6109
rect 1526 6089 1546 6109
rect 1643 6089 1663 6109
rect 1739 6089 1759 6109
rect 1851 6089 1871 6109
rect 1947 6089 1967 6109
rect 2057 6089 2077 6109
rect 2153 6089 2173 6109
rect 6486 6130 6506 6150
rect 2759 6044 2779 6064
rect 2855 6044 2875 6064
rect 2965 6044 2985 6064
rect 3061 6044 3081 6064
rect 3173 6044 3193 6064
rect 3269 6044 3289 6064
rect 3386 6044 3406 6064
rect 6582 6130 6602 6150
rect 6699 6130 6719 6150
rect 6795 6130 6815 6150
rect 6907 6130 6927 6150
rect 7003 6130 7023 6150
rect 7113 6130 7133 6150
rect 7209 6130 7229 6150
rect 3482 6044 3502 6064
rect 7815 6085 7835 6105
rect 7911 6085 7931 6105
rect 8021 6085 8041 6105
rect 8117 6085 8137 6105
rect 8229 6085 8249 6105
rect 8325 6085 8345 6105
rect 8442 6085 8462 6105
rect 8538 6085 8558 6105
rect 352 5822 372 5842
rect 448 5822 468 5842
rect 565 5822 585 5842
rect 661 5822 681 5842
rect 773 5822 793 5842
rect 869 5822 889 5842
rect 979 5822 999 5842
rect 1075 5822 1095 5842
rect 5408 5863 5428 5883
rect 3839 5762 3859 5782
rect 3935 5762 3955 5782
rect 4045 5762 4065 5782
rect 4141 5762 4161 5782
rect 4253 5762 4273 5782
rect 4349 5762 4369 5782
rect 4466 5762 4486 5782
rect 5504 5863 5524 5883
rect 5621 5863 5641 5883
rect 5717 5863 5737 5883
rect 5829 5863 5849 5883
rect 5925 5863 5945 5883
rect 6035 5863 6055 5883
rect 6131 5863 6151 5883
rect 4562 5762 4582 5782
rect 8895 5803 8915 5823
rect 8991 5803 9011 5823
rect 9101 5803 9121 5823
rect 9197 5803 9217 5823
rect 9309 5803 9329 5823
rect 9405 5803 9425 5823
rect 9522 5803 9542 5823
rect 9618 5803 9638 5823
rect 1290 5578 1310 5598
rect 1386 5578 1406 5598
rect 1503 5578 1523 5598
rect 1599 5578 1619 5598
rect 1711 5578 1731 5598
rect 1807 5578 1827 5598
rect 1917 5578 1937 5598
rect 2013 5578 2033 5598
rect 6346 5619 6366 5639
rect 2900 5452 2920 5472
rect 2996 5452 3016 5472
rect 3106 5452 3126 5472
rect 3202 5452 3222 5472
rect 3314 5452 3334 5472
rect 3410 5452 3430 5472
rect 3527 5452 3547 5472
rect 6442 5619 6462 5639
rect 6559 5619 6579 5639
rect 6655 5619 6675 5639
rect 6767 5619 6787 5639
rect 6863 5619 6883 5639
rect 6973 5619 6993 5639
rect 7069 5619 7089 5639
rect 3623 5452 3643 5472
rect 7956 5493 7976 5513
rect 8052 5493 8072 5513
rect 8162 5493 8182 5513
rect 8258 5493 8278 5513
rect 8370 5493 8390 5513
rect 8466 5493 8486 5513
rect 8583 5493 8603 5513
rect 8679 5493 8699 5513
rect 351 5268 371 5288
rect 447 5268 467 5288
rect 564 5268 584 5288
rect 660 5268 680 5288
rect 772 5268 792 5288
rect 868 5268 888 5288
rect 978 5268 998 5288
rect 1074 5268 1094 5288
rect 5407 5309 5427 5329
rect 3838 5208 3858 5228
rect 3934 5208 3954 5228
rect 4044 5208 4064 5228
rect 4140 5208 4160 5228
rect 4252 5208 4272 5228
rect 4348 5208 4368 5228
rect 4465 5208 4485 5228
rect 5503 5309 5523 5329
rect 5620 5309 5640 5329
rect 5716 5309 5736 5329
rect 5828 5309 5848 5329
rect 5924 5309 5944 5329
rect 6034 5309 6054 5329
rect 6130 5309 6150 5329
rect 4561 5208 4581 5228
rect 8894 5249 8914 5269
rect 8990 5249 9010 5269
rect 9100 5249 9120 5269
rect 9196 5249 9216 5269
rect 9308 5249 9328 5269
rect 9404 5249 9424 5269
rect 9521 5249 9541 5269
rect 9617 5249 9637 5269
rect 1399 5005 1419 5025
rect 1495 5005 1515 5025
rect 1612 5005 1632 5025
rect 1708 5005 1728 5025
rect 1820 5005 1840 5025
rect 1916 5005 1936 5025
rect 2026 5005 2046 5025
rect 2122 5005 2142 5025
rect 6455 5046 6475 5066
rect 6551 5046 6571 5066
rect 6668 5046 6688 5066
rect 6764 5046 6784 5066
rect 6876 5046 6896 5066
rect 6972 5046 6992 5066
rect 7082 5046 7102 5066
rect 7178 5046 7198 5066
rect 2791 4922 2811 4942
rect 2887 4922 2907 4942
rect 2997 4922 3017 4942
rect 3093 4922 3113 4942
rect 3205 4922 3225 4942
rect 3301 4922 3321 4942
rect 3418 4922 3438 4942
rect 3514 4922 3534 4942
rect 7847 4963 7867 4983
rect 7943 4963 7963 4983
rect 8053 4963 8073 4983
rect 8149 4963 8169 4983
rect 8261 4963 8281 4983
rect 8357 4963 8377 4983
rect 8474 4963 8494 4983
rect 8570 4963 8590 4983
rect 352 4719 372 4739
rect 448 4719 468 4739
rect 565 4719 585 4739
rect 661 4719 681 4739
rect 773 4719 793 4739
rect 869 4719 889 4739
rect 979 4719 999 4739
rect 1075 4719 1095 4739
rect 5408 4760 5428 4780
rect 3839 4659 3859 4679
rect 3935 4659 3955 4679
rect 4045 4659 4065 4679
rect 4141 4659 4161 4679
rect 4253 4659 4273 4679
rect 4349 4659 4369 4679
rect 4466 4659 4486 4679
rect 5504 4760 5524 4780
rect 5621 4760 5641 4780
rect 5717 4760 5737 4780
rect 5829 4760 5849 4780
rect 5925 4760 5945 4780
rect 6035 4760 6055 4780
rect 6131 4760 6151 4780
rect 4562 4659 4582 4679
rect 8895 4700 8915 4720
rect 8991 4700 9011 4720
rect 9101 4700 9121 4720
rect 9197 4700 9217 4720
rect 9309 4700 9329 4720
rect 9405 4700 9425 4720
rect 9522 4700 9542 4720
rect 9618 4700 9638 4720
rect 1290 4475 1310 4495
rect 1386 4475 1406 4495
rect 1503 4475 1523 4495
rect 1599 4475 1619 4495
rect 1711 4475 1731 4495
rect 1807 4475 1827 4495
rect 1917 4475 1937 4495
rect 2013 4475 2033 4495
rect 6346 4516 6366 4536
rect 2900 4349 2920 4369
rect 2996 4349 3016 4369
rect 3106 4349 3126 4369
rect 3202 4349 3222 4369
rect 3314 4349 3334 4369
rect 3410 4349 3430 4369
rect 3527 4349 3547 4369
rect 6442 4516 6462 4536
rect 6559 4516 6579 4536
rect 6655 4516 6675 4536
rect 6767 4516 6787 4536
rect 6863 4516 6883 4536
rect 6973 4516 6993 4536
rect 7069 4516 7089 4536
rect 3623 4349 3643 4369
rect 7956 4390 7976 4410
rect 8052 4390 8072 4410
rect 8162 4390 8182 4410
rect 8258 4390 8278 4410
rect 8370 4390 8390 4410
rect 8466 4390 8486 4410
rect 8583 4390 8603 4410
rect 8679 4390 8699 4410
rect 351 4165 371 4185
rect 447 4165 467 4185
rect 564 4165 584 4185
rect 660 4165 680 4185
rect 772 4165 792 4185
rect 868 4165 888 4185
rect 978 4165 998 4185
rect 1074 4165 1094 4185
rect 5407 4206 5427 4226
rect 3838 4105 3858 4125
rect 3934 4105 3954 4125
rect 4044 4105 4064 4125
rect 4140 4105 4160 4125
rect 4252 4105 4272 4125
rect 4348 4105 4368 4125
rect 4465 4105 4485 4125
rect 5503 4206 5523 4226
rect 5620 4206 5640 4226
rect 5716 4206 5736 4226
rect 5828 4206 5848 4226
rect 5924 4206 5944 4226
rect 6034 4206 6054 4226
rect 6130 4206 6150 4226
rect 4561 4105 4581 4125
rect 8894 4146 8914 4166
rect 8990 4146 9010 4166
rect 9100 4146 9120 4166
rect 9196 4146 9216 4166
rect 9308 4146 9328 4166
rect 9404 4146 9424 4166
rect 9521 4146 9541 4166
rect 9617 4146 9637 4166
rect 1431 3883 1451 3903
rect 1527 3883 1547 3903
rect 1644 3883 1664 3903
rect 1740 3883 1760 3903
rect 1852 3883 1872 3903
rect 1948 3883 1968 3903
rect 2058 3883 2078 3903
rect 2154 3883 2174 3903
rect 6487 3924 6507 3944
rect 2760 3838 2780 3858
rect 2856 3838 2876 3858
rect 2966 3838 2986 3858
rect 3062 3838 3082 3858
rect 3174 3838 3194 3858
rect 3270 3838 3290 3858
rect 3387 3838 3407 3858
rect 6583 3924 6603 3944
rect 6700 3924 6720 3944
rect 6796 3924 6816 3944
rect 6908 3924 6928 3944
rect 7004 3924 7024 3944
rect 7114 3924 7134 3944
rect 7210 3924 7230 3944
rect 3483 3838 3503 3858
rect 7816 3879 7836 3899
rect 7912 3879 7932 3899
rect 8022 3879 8042 3899
rect 8118 3879 8138 3899
rect 8230 3879 8250 3899
rect 8326 3879 8346 3899
rect 8443 3879 8463 3899
rect 8539 3879 8559 3899
rect 353 3616 373 3636
rect 449 3616 469 3636
rect 566 3616 586 3636
rect 662 3616 682 3636
rect 774 3616 794 3636
rect 870 3616 890 3636
rect 980 3616 1000 3636
rect 1076 3616 1096 3636
rect 5409 3657 5429 3677
rect 3840 3556 3860 3576
rect 3936 3556 3956 3576
rect 4046 3556 4066 3576
rect 4142 3556 4162 3576
rect 4254 3556 4274 3576
rect 4350 3556 4370 3576
rect 4467 3556 4487 3576
rect 5505 3657 5525 3677
rect 5622 3657 5642 3677
rect 5718 3657 5738 3677
rect 5830 3657 5850 3677
rect 5926 3657 5946 3677
rect 6036 3657 6056 3677
rect 6132 3657 6152 3677
rect 4563 3556 4583 3576
rect 8896 3597 8916 3617
rect 8992 3597 9012 3617
rect 9102 3597 9122 3617
rect 9198 3597 9218 3617
rect 9310 3597 9330 3617
rect 9406 3597 9426 3617
rect 9523 3597 9543 3617
rect 9619 3597 9639 3617
rect 1291 3372 1311 3392
rect 1387 3372 1407 3392
rect 1504 3372 1524 3392
rect 1600 3372 1620 3392
rect 1712 3372 1732 3392
rect 1808 3372 1828 3392
rect 1918 3372 1938 3392
rect 2014 3372 2034 3392
rect 6347 3413 6367 3433
rect 2901 3246 2921 3266
rect 2997 3246 3017 3266
rect 3107 3246 3127 3266
rect 3203 3246 3223 3266
rect 3315 3246 3335 3266
rect 3411 3246 3431 3266
rect 3528 3246 3548 3266
rect 6443 3413 6463 3433
rect 6560 3413 6580 3433
rect 6656 3413 6676 3433
rect 6768 3413 6788 3433
rect 6864 3413 6884 3433
rect 6974 3413 6994 3433
rect 7070 3413 7090 3433
rect 3624 3246 3644 3266
rect 7957 3287 7977 3307
rect 8053 3287 8073 3307
rect 8163 3287 8183 3307
rect 8259 3287 8279 3307
rect 8371 3287 8391 3307
rect 8467 3287 8487 3307
rect 8584 3287 8604 3307
rect 8680 3287 8700 3307
rect 352 3062 372 3082
rect 448 3062 468 3082
rect 565 3062 585 3082
rect 661 3062 681 3082
rect 773 3062 793 3082
rect 869 3062 889 3082
rect 979 3062 999 3082
rect 1075 3062 1095 3082
rect 5408 3103 5428 3123
rect 3839 3002 3859 3022
rect 3935 3002 3955 3022
rect 4045 3002 4065 3022
rect 4141 3002 4161 3022
rect 4253 3002 4273 3022
rect 4349 3002 4369 3022
rect 4466 3002 4486 3022
rect 5504 3103 5524 3123
rect 5621 3103 5641 3123
rect 5717 3103 5737 3123
rect 5829 3103 5849 3123
rect 5925 3103 5945 3123
rect 6035 3103 6055 3123
rect 6131 3103 6151 3123
rect 4562 3002 4582 3022
rect 8895 3043 8915 3063
rect 8991 3043 9011 3063
rect 9101 3043 9121 3063
rect 9197 3043 9217 3063
rect 9309 3043 9329 3063
rect 9405 3043 9425 3063
rect 9522 3043 9542 3063
rect 9618 3043 9638 3063
rect 1401 2793 1421 2813
rect 1497 2793 1517 2813
rect 1614 2793 1634 2813
rect 1710 2793 1730 2813
rect 1822 2793 1842 2813
rect 1918 2793 1938 2813
rect 2028 2793 2048 2813
rect 2124 2793 2144 2813
rect 6457 2834 6477 2854
rect 6553 2834 6573 2854
rect 6670 2834 6690 2854
rect 6766 2834 6786 2854
rect 6878 2834 6898 2854
rect 6974 2834 6994 2854
rect 7084 2834 7104 2854
rect 7180 2834 7200 2854
rect 2791 2722 2811 2742
rect 2887 2722 2907 2742
rect 2997 2722 3017 2742
rect 3093 2722 3113 2742
rect 3205 2722 3225 2742
rect 3301 2722 3321 2742
rect 3418 2722 3438 2742
rect 3514 2722 3534 2742
rect 7847 2763 7867 2783
rect 7943 2763 7963 2783
rect 8053 2763 8073 2783
rect 8149 2763 8169 2783
rect 8261 2763 8281 2783
rect 8357 2763 8377 2783
rect 8474 2763 8494 2783
rect 8570 2763 8590 2783
rect 353 2513 373 2533
rect 449 2513 469 2533
rect 566 2513 586 2533
rect 662 2513 682 2533
rect 774 2513 794 2533
rect 870 2513 890 2533
rect 980 2513 1000 2533
rect 1076 2513 1096 2533
rect 5409 2554 5429 2574
rect 3840 2453 3860 2473
rect 3936 2453 3956 2473
rect 4046 2453 4066 2473
rect 4142 2453 4162 2473
rect 4254 2453 4274 2473
rect 4350 2453 4370 2473
rect 4467 2453 4487 2473
rect 5505 2554 5525 2574
rect 5622 2554 5642 2574
rect 5718 2554 5738 2574
rect 5830 2554 5850 2574
rect 5926 2554 5946 2574
rect 6036 2554 6056 2574
rect 6132 2554 6152 2574
rect 4563 2453 4583 2473
rect 8896 2494 8916 2514
rect 8992 2494 9012 2514
rect 9102 2494 9122 2514
rect 9198 2494 9218 2514
rect 9310 2494 9330 2514
rect 9406 2494 9426 2514
rect 9523 2494 9543 2514
rect 9619 2494 9639 2514
rect 1291 2269 1311 2289
rect 1387 2269 1407 2289
rect 1504 2269 1524 2289
rect 1600 2269 1620 2289
rect 1712 2269 1732 2289
rect 1808 2269 1828 2289
rect 1918 2269 1938 2289
rect 2014 2269 2034 2289
rect 6347 2310 6367 2330
rect 2901 2143 2921 2163
rect 2997 2143 3017 2163
rect 3107 2143 3127 2163
rect 3203 2143 3223 2163
rect 3315 2143 3335 2163
rect 3411 2143 3431 2163
rect 3528 2143 3548 2163
rect 6443 2310 6463 2330
rect 6560 2310 6580 2330
rect 6656 2310 6676 2330
rect 6768 2310 6788 2330
rect 6864 2310 6884 2330
rect 6974 2310 6994 2330
rect 7070 2310 7090 2330
rect 3624 2143 3644 2163
rect 7957 2184 7977 2204
rect 8053 2184 8073 2204
rect 8163 2184 8183 2204
rect 8259 2184 8279 2204
rect 8371 2184 8391 2204
rect 8467 2184 8487 2204
rect 8584 2184 8604 2204
rect 8680 2184 8700 2204
rect 352 1959 372 1979
rect 448 1959 468 1979
rect 565 1959 585 1979
rect 661 1959 681 1979
rect 773 1959 793 1979
rect 869 1959 889 1979
rect 979 1959 999 1979
rect 1075 1959 1095 1979
rect 5408 2000 5428 2020
rect 3839 1899 3859 1919
rect 3935 1899 3955 1919
rect 4045 1899 4065 1919
rect 4141 1899 4161 1919
rect 4253 1899 4273 1919
rect 4349 1899 4369 1919
rect 4466 1899 4486 1919
rect 5504 2000 5524 2020
rect 5621 2000 5641 2020
rect 5717 2000 5737 2020
rect 5829 2000 5849 2020
rect 5925 2000 5945 2020
rect 6035 2000 6055 2020
rect 6131 2000 6151 2020
rect 4562 1899 4582 1919
rect 8895 1940 8915 1960
rect 8991 1940 9011 1960
rect 9101 1940 9121 1960
rect 9197 1940 9217 1960
rect 9309 1940 9329 1960
rect 9405 1940 9425 1960
rect 9522 1940 9542 1960
rect 9618 1940 9638 1960
rect 1432 1677 1452 1697
rect 1528 1677 1548 1697
rect 1645 1677 1665 1697
rect 1741 1677 1761 1697
rect 1853 1677 1873 1697
rect 1949 1677 1969 1697
rect 2059 1677 2079 1697
rect 2155 1677 2175 1697
rect 6488 1718 6508 1738
rect 2761 1632 2781 1652
rect 2857 1632 2877 1652
rect 2967 1632 2987 1652
rect 3063 1632 3083 1652
rect 3175 1632 3195 1652
rect 3271 1632 3291 1652
rect 3388 1632 3408 1652
rect 6584 1718 6604 1738
rect 6701 1718 6721 1738
rect 6797 1718 6817 1738
rect 6909 1718 6929 1738
rect 7005 1718 7025 1738
rect 7115 1718 7135 1738
rect 7211 1718 7231 1738
rect 3484 1632 3504 1652
rect 7817 1673 7837 1693
rect 7913 1673 7933 1693
rect 8023 1673 8043 1693
rect 8119 1673 8139 1693
rect 8231 1673 8251 1693
rect 8327 1673 8347 1693
rect 8444 1673 8464 1693
rect 8540 1673 8560 1693
rect 354 1410 374 1430
rect 450 1410 470 1430
rect 567 1410 587 1430
rect 663 1410 683 1430
rect 775 1410 795 1430
rect 871 1410 891 1430
rect 981 1410 1001 1430
rect 1077 1410 1097 1430
rect 5410 1451 5430 1471
rect 3841 1350 3861 1370
rect 3937 1350 3957 1370
rect 4047 1350 4067 1370
rect 4143 1350 4163 1370
rect 4255 1350 4275 1370
rect 4351 1350 4371 1370
rect 4468 1350 4488 1370
rect 5506 1451 5526 1471
rect 5623 1451 5643 1471
rect 5719 1451 5739 1471
rect 5831 1451 5851 1471
rect 5927 1451 5947 1471
rect 6037 1451 6057 1471
rect 6133 1451 6153 1471
rect 4564 1350 4584 1370
rect 8897 1391 8917 1411
rect 8993 1391 9013 1411
rect 9103 1391 9123 1411
rect 9199 1391 9219 1411
rect 9311 1391 9331 1411
rect 9407 1391 9427 1411
rect 9524 1391 9544 1411
rect 9620 1391 9640 1411
rect 1292 1166 1312 1186
rect 1388 1166 1408 1186
rect 1505 1166 1525 1186
rect 1601 1166 1621 1186
rect 1713 1166 1733 1186
rect 1809 1166 1829 1186
rect 1919 1166 1939 1186
rect 2015 1166 2035 1186
rect 6348 1207 6368 1227
rect 2902 1040 2922 1060
rect 2998 1040 3018 1060
rect 3108 1040 3128 1060
rect 3204 1040 3224 1060
rect 3316 1040 3336 1060
rect 3412 1040 3432 1060
rect 3529 1040 3549 1060
rect 6444 1207 6464 1227
rect 6561 1207 6581 1227
rect 6657 1207 6677 1227
rect 6769 1207 6789 1227
rect 6865 1207 6885 1227
rect 6975 1207 6995 1227
rect 7071 1207 7091 1227
rect 3625 1040 3645 1060
rect 7958 1081 7978 1101
rect 8054 1081 8074 1101
rect 8164 1081 8184 1101
rect 8260 1081 8280 1101
rect 8372 1081 8392 1101
rect 8468 1081 8488 1101
rect 8585 1081 8605 1101
rect 8681 1081 8701 1101
rect 353 856 373 876
rect 449 856 469 876
rect 566 856 586 876
rect 662 856 682 876
rect 774 856 794 876
rect 870 856 890 876
rect 980 856 1000 876
rect 1076 856 1096 876
rect 5409 897 5429 917
rect 3840 796 3860 816
rect 3936 796 3956 816
rect 4046 796 4066 816
rect 4142 796 4162 816
rect 4254 796 4274 816
rect 4350 796 4370 816
rect 4467 796 4487 816
rect 5505 897 5525 917
rect 5622 897 5642 917
rect 5718 897 5738 917
rect 5830 897 5850 917
rect 5926 897 5946 917
rect 6036 897 6056 917
rect 6132 897 6152 917
rect 4563 796 4583 816
rect 8896 837 8916 857
rect 8992 837 9012 857
rect 9102 837 9122 857
rect 9198 837 9218 857
rect 9310 837 9330 857
rect 9406 837 9426 857
rect 9523 837 9543 857
rect 9619 837 9639 857
rect 1600 297 1620 317
rect 1696 297 1716 317
rect 1813 297 1833 317
rect 1909 297 1929 317
rect 2021 297 2041 317
rect 2117 297 2137 317
rect 2227 297 2247 317
rect 6656 338 6676 358
rect 2323 297 2343 317
rect 4550 277 4570 297
rect 4646 277 4666 297
rect 4763 277 4783 297
rect 4859 277 4879 297
rect 4971 277 4991 297
rect 5067 277 5087 297
rect 5177 277 5197 297
rect 5273 277 5293 297
rect 6752 338 6772 358
rect 6869 338 6889 358
rect 6965 338 6985 358
rect 7077 338 7097 358
rect 7173 338 7193 358
rect 7283 338 7303 358
rect 7379 338 7399 358
<< psubdiff >>
rect 9457 9378 9568 9393
rect 4401 9337 4512 9352
rect 9457 9348 9499 9378
rect 9527 9348 9568 9378
rect 4401 9307 4443 9337
rect 4471 9307 4512 9337
rect 9457 9334 9568 9348
rect 4401 9293 4512 9307
rect 3462 9027 3573 9042
rect 3462 8997 3504 9027
rect 3532 8997 3573 9027
rect 3462 8983 3573 8997
rect 8518 9068 8629 9083
rect 8518 9038 8560 9068
rect 8588 9038 8629 9068
rect 8518 9024 8629 9038
rect 418 8915 529 8929
rect 418 8885 459 8915
rect 487 8885 529 8915
rect 418 8870 529 8885
rect 5474 8956 5585 8970
rect 5474 8926 5515 8956
rect 5543 8926 5585 8956
rect 5474 8911 5585 8926
rect 4400 8783 4511 8798
rect 4400 8753 4442 8783
rect 4470 8753 4511 8783
rect 4400 8739 4511 8753
rect 9456 8824 9567 8839
rect 9456 8794 9498 8824
rect 9526 8794 9567 8824
rect 9456 8780 9567 8794
rect 1356 8671 1467 8685
rect 1356 8641 1397 8671
rect 1425 8641 1467 8671
rect 1356 8626 1467 8641
rect 6412 8712 6523 8726
rect 6412 8682 6453 8712
rect 6481 8682 6523 8712
rect 3322 8516 3433 8531
rect 3322 8486 3364 8516
rect 3392 8486 3433 8516
rect 3322 8472 3433 8486
rect 6412 8667 6523 8682
rect 8378 8557 8489 8572
rect 8378 8527 8420 8557
rect 8448 8527 8489 8557
rect 8378 8513 8489 8527
rect 417 8361 528 8375
rect 417 8331 458 8361
rect 486 8331 528 8361
rect 417 8316 528 8331
rect 5473 8402 5584 8416
rect 5473 8372 5514 8402
rect 5542 8372 5584 8402
rect 5473 8357 5584 8372
rect 4402 8234 4513 8249
rect 4402 8204 4444 8234
rect 4472 8204 4513 8234
rect 4402 8190 4513 8204
rect 9458 8275 9569 8290
rect 9458 8245 9500 8275
rect 9528 8245 9569 8275
rect 9458 8231 9569 8245
rect 1497 8079 1608 8093
rect 1497 8049 1538 8079
rect 1566 8049 1608 8079
rect 1497 8034 1608 8049
rect 3463 7924 3574 7939
rect 6553 8120 6664 8134
rect 6553 8090 6594 8120
rect 6622 8090 6664 8120
rect 6553 8075 6664 8090
rect 3463 7894 3505 7924
rect 3533 7894 3574 7924
rect 3463 7880 3574 7894
rect 8519 7965 8630 7980
rect 8519 7935 8561 7965
rect 8589 7935 8630 7965
rect 8519 7921 8630 7935
rect 419 7812 530 7826
rect 419 7782 460 7812
rect 488 7782 530 7812
rect 419 7767 530 7782
rect 5475 7853 5586 7867
rect 5475 7823 5516 7853
rect 5544 7823 5586 7853
rect 5475 7808 5586 7823
rect 4401 7680 4512 7695
rect 4401 7650 4443 7680
rect 4471 7650 4512 7680
rect 4401 7636 4512 7650
rect 9457 7721 9568 7736
rect 9457 7691 9499 7721
rect 9527 7691 9568 7721
rect 9457 7677 9568 7691
rect 1357 7568 1468 7582
rect 1357 7538 1398 7568
rect 1426 7538 1468 7568
rect 1357 7523 1468 7538
rect 6413 7609 6524 7623
rect 6413 7579 6454 7609
rect 6482 7579 6524 7609
rect 3353 7400 3464 7415
rect 3353 7370 3395 7400
rect 3423 7370 3464 7400
rect 6413 7564 6524 7579
rect 8409 7441 8520 7456
rect 8409 7411 8451 7441
rect 8479 7411 8520 7441
rect 8409 7397 8520 7411
rect 3353 7356 3464 7370
rect 418 7258 529 7272
rect 5474 7299 5585 7313
rect 418 7228 459 7258
rect 487 7228 529 7258
rect 418 7214 529 7228
rect 5474 7269 5515 7299
rect 5543 7269 5585 7299
rect 5474 7255 5585 7269
rect 4402 7131 4513 7145
rect 4402 7101 4444 7131
rect 4472 7101 4513 7131
rect 9458 7172 9569 7186
rect 9458 7142 9500 7172
rect 9528 7142 9569 7172
rect 4402 7087 4513 7101
rect 9458 7128 9569 7142
rect 6523 7030 6634 7044
rect 1467 6989 1578 7003
rect 1467 6959 1508 6989
rect 1536 6959 1578 6989
rect 1467 6944 1578 6959
rect 3463 6821 3574 6836
rect 6523 7000 6564 7030
rect 6592 7000 6634 7030
rect 6523 6985 6634 7000
rect 3463 6791 3505 6821
rect 3533 6791 3574 6821
rect 3463 6777 3574 6791
rect 8519 6862 8630 6877
rect 8519 6832 8561 6862
rect 8589 6832 8630 6862
rect 8519 6818 8630 6832
rect 419 6709 530 6723
rect 419 6679 460 6709
rect 488 6679 530 6709
rect 419 6664 530 6679
rect 5475 6750 5586 6764
rect 5475 6720 5516 6750
rect 5544 6720 5586 6750
rect 5475 6705 5586 6720
rect 4401 6577 4512 6592
rect 4401 6547 4443 6577
rect 4471 6547 4512 6577
rect 4401 6533 4512 6547
rect 9457 6618 9568 6633
rect 9457 6588 9499 6618
rect 9527 6588 9568 6618
rect 9457 6574 9568 6588
rect 1357 6465 1468 6479
rect 1357 6435 1398 6465
rect 1426 6435 1468 6465
rect 1357 6420 1468 6435
rect 6413 6506 6524 6520
rect 6413 6476 6454 6506
rect 6482 6476 6524 6506
rect 3323 6310 3434 6325
rect 3323 6280 3365 6310
rect 3393 6280 3434 6310
rect 3323 6266 3434 6280
rect 6413 6461 6524 6476
rect 8379 6351 8490 6366
rect 8379 6321 8421 6351
rect 8449 6321 8490 6351
rect 8379 6307 8490 6321
rect 418 6155 529 6169
rect 418 6125 459 6155
rect 487 6125 529 6155
rect 418 6110 529 6125
rect 5474 6196 5585 6210
rect 5474 6166 5515 6196
rect 5543 6166 5585 6196
rect 5474 6151 5585 6166
rect 4403 6028 4514 6043
rect 4403 5998 4445 6028
rect 4473 5998 4514 6028
rect 4403 5984 4514 5998
rect 9459 6069 9570 6084
rect 9459 6039 9501 6069
rect 9529 6039 9570 6069
rect 9459 6025 9570 6039
rect 1498 5873 1609 5887
rect 1498 5843 1539 5873
rect 1567 5843 1609 5873
rect 1498 5828 1609 5843
rect 3464 5718 3575 5733
rect 6554 5914 6665 5928
rect 6554 5884 6595 5914
rect 6623 5884 6665 5914
rect 6554 5869 6665 5884
rect 3464 5688 3506 5718
rect 3534 5688 3575 5718
rect 3464 5674 3575 5688
rect 8520 5759 8631 5774
rect 8520 5729 8562 5759
rect 8590 5729 8631 5759
rect 8520 5715 8631 5729
rect 420 5606 531 5620
rect 420 5576 461 5606
rect 489 5576 531 5606
rect 420 5561 531 5576
rect 5476 5647 5587 5661
rect 5476 5617 5517 5647
rect 5545 5617 5587 5647
rect 5476 5602 5587 5617
rect 4402 5474 4513 5489
rect 4402 5444 4444 5474
rect 4472 5444 4513 5474
rect 4402 5430 4513 5444
rect 9458 5515 9569 5530
rect 9458 5485 9500 5515
rect 9528 5485 9569 5515
rect 9458 5471 9569 5485
rect 1358 5362 1469 5376
rect 1358 5332 1399 5362
rect 1427 5332 1469 5362
rect 1358 5317 1469 5332
rect 6414 5403 6525 5417
rect 6414 5373 6455 5403
rect 6483 5373 6525 5403
rect 3355 5188 3466 5203
rect 3355 5158 3397 5188
rect 3425 5158 3466 5188
rect 6414 5358 6525 5373
rect 8411 5229 8522 5244
rect 8411 5199 8453 5229
rect 8481 5199 8522 5229
rect 3355 5144 3466 5158
rect 419 5052 530 5066
rect 419 5022 460 5052
rect 488 5022 530 5052
rect 419 5007 530 5022
rect 8411 5185 8522 5199
rect 5475 5093 5586 5107
rect 5475 5063 5516 5093
rect 5544 5063 5586 5093
rect 5475 5048 5586 5063
rect 4403 4925 4514 4940
rect 4403 4895 4445 4925
rect 4473 4895 4514 4925
rect 4403 4881 4514 4895
rect 1467 4789 1578 4803
rect 9459 4966 9570 4981
rect 9459 4936 9501 4966
rect 9529 4936 9570 4966
rect 9459 4922 9570 4936
rect 6523 4830 6634 4844
rect 1467 4759 1508 4789
rect 1536 4759 1578 4789
rect 1467 4744 1578 4759
rect 3464 4615 3575 4630
rect 6523 4800 6564 4830
rect 6592 4800 6634 4830
rect 6523 4785 6634 4800
rect 3464 4585 3506 4615
rect 3534 4585 3575 4615
rect 3464 4571 3575 4585
rect 8520 4656 8631 4671
rect 8520 4626 8562 4656
rect 8590 4626 8631 4656
rect 8520 4612 8631 4626
rect 420 4503 531 4517
rect 420 4473 461 4503
rect 489 4473 531 4503
rect 420 4458 531 4473
rect 5476 4544 5587 4558
rect 5476 4514 5517 4544
rect 5545 4514 5587 4544
rect 5476 4499 5587 4514
rect 4402 4371 4513 4386
rect 4402 4341 4444 4371
rect 4472 4341 4513 4371
rect 4402 4327 4513 4341
rect 9458 4412 9569 4427
rect 9458 4382 9500 4412
rect 9528 4382 9569 4412
rect 9458 4368 9569 4382
rect 1358 4259 1469 4273
rect 1358 4229 1399 4259
rect 1427 4229 1469 4259
rect 1358 4214 1469 4229
rect 6414 4300 6525 4314
rect 6414 4270 6455 4300
rect 6483 4270 6525 4300
rect 3324 4104 3435 4119
rect 3324 4074 3366 4104
rect 3394 4074 3435 4104
rect 3324 4060 3435 4074
rect 6414 4255 6525 4270
rect 8380 4145 8491 4160
rect 8380 4115 8422 4145
rect 8450 4115 8491 4145
rect 8380 4101 8491 4115
rect 419 3949 530 3963
rect 419 3919 460 3949
rect 488 3919 530 3949
rect 419 3904 530 3919
rect 5475 3990 5586 4004
rect 5475 3960 5516 3990
rect 5544 3960 5586 3990
rect 5475 3945 5586 3960
rect 4404 3822 4515 3837
rect 4404 3792 4446 3822
rect 4474 3792 4515 3822
rect 4404 3778 4515 3792
rect 9460 3863 9571 3878
rect 9460 3833 9502 3863
rect 9530 3833 9571 3863
rect 9460 3819 9571 3833
rect 1499 3667 1610 3681
rect 1499 3637 1540 3667
rect 1568 3637 1610 3667
rect 1499 3622 1610 3637
rect 3465 3512 3576 3527
rect 6555 3708 6666 3722
rect 6555 3678 6596 3708
rect 6624 3678 6666 3708
rect 6555 3663 6666 3678
rect 3465 3482 3507 3512
rect 3535 3482 3576 3512
rect 3465 3468 3576 3482
rect 8521 3553 8632 3568
rect 8521 3523 8563 3553
rect 8591 3523 8632 3553
rect 8521 3509 8632 3523
rect 421 3400 532 3414
rect 421 3370 462 3400
rect 490 3370 532 3400
rect 421 3355 532 3370
rect 5477 3441 5588 3455
rect 5477 3411 5518 3441
rect 5546 3411 5588 3441
rect 5477 3396 5588 3411
rect 4403 3268 4514 3283
rect 4403 3238 4445 3268
rect 4473 3238 4514 3268
rect 4403 3224 4514 3238
rect 9459 3309 9570 3324
rect 9459 3279 9501 3309
rect 9529 3279 9570 3309
rect 9459 3265 9570 3279
rect 1359 3156 1470 3170
rect 1359 3126 1400 3156
rect 1428 3126 1470 3156
rect 1359 3111 1470 3126
rect 6415 3197 6526 3211
rect 6415 3167 6456 3197
rect 6484 3167 6526 3197
rect 3355 2988 3466 3003
rect 3355 2958 3397 2988
rect 3425 2958 3466 2988
rect 6415 3152 6526 3167
rect 8411 3029 8522 3044
rect 8411 2999 8453 3029
rect 8481 2999 8522 3029
rect 8411 2985 8522 2999
rect 3355 2944 3466 2958
rect 420 2846 531 2860
rect 5476 2887 5587 2901
rect 420 2816 461 2846
rect 489 2816 531 2846
rect 420 2802 531 2816
rect 5476 2857 5517 2887
rect 5545 2857 5587 2887
rect 5476 2843 5587 2857
rect 4404 2719 4515 2733
rect 4404 2689 4446 2719
rect 4474 2689 4515 2719
rect 9460 2760 9571 2774
rect 9460 2730 9502 2760
rect 9530 2730 9571 2760
rect 4404 2675 4515 2689
rect 9460 2716 9571 2730
rect 6525 2618 6636 2632
rect 1469 2577 1580 2591
rect 1469 2547 1510 2577
rect 1538 2547 1580 2577
rect 1469 2532 1580 2547
rect 3465 2409 3576 2424
rect 6525 2588 6566 2618
rect 6594 2588 6636 2618
rect 6525 2573 6636 2588
rect 3465 2379 3507 2409
rect 3535 2379 3576 2409
rect 3465 2365 3576 2379
rect 8521 2450 8632 2465
rect 8521 2420 8563 2450
rect 8591 2420 8632 2450
rect 8521 2406 8632 2420
rect 421 2297 532 2311
rect 421 2267 462 2297
rect 490 2267 532 2297
rect 421 2252 532 2267
rect 5477 2338 5588 2352
rect 5477 2308 5518 2338
rect 5546 2308 5588 2338
rect 5477 2293 5588 2308
rect 4403 2165 4514 2180
rect 4403 2135 4445 2165
rect 4473 2135 4514 2165
rect 4403 2121 4514 2135
rect 9459 2206 9570 2221
rect 9459 2176 9501 2206
rect 9529 2176 9570 2206
rect 9459 2162 9570 2176
rect 1359 2053 1470 2067
rect 1359 2023 1400 2053
rect 1428 2023 1470 2053
rect 1359 2008 1470 2023
rect 6415 2094 6526 2108
rect 6415 2064 6456 2094
rect 6484 2064 6526 2094
rect 3325 1898 3436 1913
rect 3325 1868 3367 1898
rect 3395 1868 3436 1898
rect 3325 1854 3436 1868
rect 6415 2049 6526 2064
rect 8381 1939 8492 1954
rect 8381 1909 8423 1939
rect 8451 1909 8492 1939
rect 8381 1895 8492 1909
rect 420 1743 531 1757
rect 420 1713 461 1743
rect 489 1713 531 1743
rect 420 1698 531 1713
rect 5476 1784 5587 1798
rect 5476 1754 5517 1784
rect 5545 1754 5587 1784
rect 5476 1739 5587 1754
rect 4405 1616 4516 1631
rect 4405 1586 4447 1616
rect 4475 1586 4516 1616
rect 4405 1572 4516 1586
rect 9461 1657 9572 1672
rect 9461 1627 9503 1657
rect 9531 1627 9572 1657
rect 9461 1613 9572 1627
rect 1500 1461 1611 1475
rect 1500 1431 1541 1461
rect 1569 1431 1611 1461
rect 1500 1416 1611 1431
rect 3466 1306 3577 1321
rect 6556 1502 6667 1516
rect 6556 1472 6597 1502
rect 6625 1472 6667 1502
rect 6556 1457 6667 1472
rect 3466 1276 3508 1306
rect 3536 1276 3577 1306
rect 3466 1262 3577 1276
rect 8522 1347 8633 1362
rect 8522 1317 8564 1347
rect 8592 1317 8633 1347
rect 8522 1303 8633 1317
rect 422 1194 533 1208
rect 422 1164 463 1194
rect 491 1164 533 1194
rect 422 1149 533 1164
rect 5478 1235 5589 1249
rect 5478 1205 5519 1235
rect 5547 1205 5589 1235
rect 5478 1190 5589 1205
rect 4404 1062 4515 1077
rect 4404 1032 4446 1062
rect 4474 1032 4515 1062
rect 4404 1018 4515 1032
rect 9460 1103 9571 1118
rect 9460 1073 9502 1103
rect 9530 1073 9571 1103
rect 9460 1059 9571 1073
rect 1360 950 1471 964
rect 1360 920 1401 950
rect 1429 920 1471 950
rect 1360 905 1471 920
rect 6416 991 6527 1005
rect 6416 961 6457 991
rect 6485 961 6527 991
rect 6416 946 6527 961
rect 5477 681 5588 695
rect 421 640 532 654
rect 5477 651 5518 681
rect 5546 675 5588 681
rect 5546 651 5587 675
rect 421 610 462 640
rect 490 634 532 640
rect 5477 636 5587 651
rect 490 610 531 634
rect 421 595 531 610
rect 6724 122 6835 136
rect 1668 81 1779 95
rect 1668 51 1709 81
rect 1737 51 1779 81
rect 6724 92 6765 122
rect 6793 92 6835 122
rect 6724 77 6835 92
rect 1668 36 1779 51
rect 4618 61 4729 75
rect 4618 31 4659 61
rect 4687 31 4729 61
rect 4618 16 4729 31
<< nsubdiff >>
rect 5475 9303 5585 9317
rect 419 9262 529 9276
rect 419 9232 462 9262
rect 490 9232 529 9262
rect 419 9217 529 9232
rect 5475 9273 5518 9303
rect 5546 9273 5585 9303
rect 5475 9258 5585 9273
rect 1357 9018 1467 9032
rect 1357 8988 1400 9018
rect 1428 8988 1467 9018
rect 1357 8973 1467 8988
rect 6413 9059 6523 9073
rect 4401 8990 4511 9005
rect 6413 9029 6456 9059
rect 6484 9029 6523 9059
rect 6413 9014 6523 9029
rect 9457 9031 9567 9046
rect 9457 9001 9496 9031
rect 9524 9001 9567 9031
rect 4401 8960 4440 8990
rect 4468 8960 4511 8990
rect 4401 8946 4511 8960
rect 418 8708 528 8722
rect 9457 8987 9567 9001
rect 5474 8749 5584 8763
rect 5474 8719 5517 8749
rect 5545 8719 5584 8749
rect 418 8678 461 8708
rect 489 8678 528 8708
rect 418 8663 528 8678
rect 3462 8680 3572 8695
rect 3462 8650 3501 8680
rect 3529 8650 3572 8680
rect 5474 8704 5584 8719
rect 3462 8636 3572 8650
rect 8518 8721 8628 8736
rect 8518 8691 8557 8721
rect 8585 8691 8628 8721
rect 8518 8677 8628 8691
rect 1498 8426 1608 8440
rect 4400 8436 4510 8451
rect 1498 8396 1541 8426
rect 1569 8396 1608 8426
rect 1498 8381 1608 8396
rect 4400 8406 4439 8436
rect 4467 8406 4510 8436
rect 6554 8467 6664 8481
rect 9456 8477 9566 8492
rect 4400 8392 4510 8406
rect 6554 8437 6597 8467
rect 6625 8437 6664 8467
rect 6554 8422 6664 8437
rect 9456 8447 9495 8477
rect 9523 8447 9566 8477
rect 9456 8433 9566 8447
rect 420 8159 530 8173
rect 420 8129 463 8159
rect 491 8129 530 8159
rect 3322 8169 3432 8184
rect 3322 8139 3361 8169
rect 3389 8139 3432 8169
rect 5476 8200 5586 8214
rect 420 8114 530 8129
rect 3322 8125 3432 8139
rect 5476 8170 5519 8200
rect 5547 8170 5586 8200
rect 8378 8210 8488 8225
rect 8378 8180 8417 8210
rect 8445 8180 8488 8210
rect 5476 8155 5586 8170
rect 8378 8166 8488 8180
rect 1358 7915 1468 7929
rect 1358 7885 1401 7915
rect 1429 7885 1468 7915
rect 1358 7870 1468 7885
rect 6414 7956 6524 7970
rect 4402 7887 4512 7902
rect 6414 7926 6457 7956
rect 6485 7926 6524 7956
rect 6414 7911 6524 7926
rect 9458 7928 9568 7943
rect 9458 7898 9497 7928
rect 9525 7898 9568 7928
rect 4402 7857 4441 7887
rect 4469 7857 4512 7887
rect 4402 7843 4512 7857
rect 419 7605 529 7619
rect 9458 7884 9568 7898
rect 5475 7646 5585 7660
rect 5475 7616 5518 7646
rect 5546 7616 5585 7646
rect 419 7575 462 7605
rect 490 7575 529 7605
rect 419 7560 529 7575
rect 3463 7577 3573 7592
rect 3463 7547 3502 7577
rect 3530 7547 3573 7577
rect 5475 7601 5585 7616
rect 3463 7533 3573 7547
rect 8519 7618 8629 7633
rect 8519 7588 8558 7618
rect 8586 7588 8629 7618
rect 8519 7574 8629 7588
rect 1468 7336 1578 7350
rect 1468 7306 1511 7336
rect 1539 7306 1578 7336
rect 4401 7333 4511 7348
rect 1468 7291 1578 7306
rect 4401 7303 4440 7333
rect 4468 7303 4511 7333
rect 6524 7377 6634 7391
rect 6524 7347 6567 7377
rect 6595 7347 6634 7377
rect 9457 7374 9567 7389
rect 6524 7332 6634 7347
rect 4401 7289 4511 7303
rect 9457 7344 9496 7374
rect 9524 7344 9567 7374
rect 9457 7330 9567 7344
rect 420 7056 530 7070
rect 420 7026 463 7056
rect 491 7026 530 7056
rect 5476 7097 5586 7111
rect 3353 7053 3463 7068
rect 420 7011 530 7026
rect 3353 7023 3392 7053
rect 3420 7023 3463 7053
rect 3353 7009 3463 7023
rect 5476 7067 5519 7097
rect 5547 7067 5586 7097
rect 8409 7094 8519 7109
rect 5476 7052 5586 7067
rect 8409 7064 8448 7094
rect 8476 7064 8519 7094
rect 8409 7050 8519 7064
rect 1358 6812 1468 6826
rect 1358 6782 1401 6812
rect 1429 6782 1468 6812
rect 1358 6767 1468 6782
rect 6414 6853 6524 6867
rect 4402 6784 4512 6799
rect 6414 6823 6457 6853
rect 6485 6823 6524 6853
rect 6414 6808 6524 6823
rect 9458 6825 9568 6840
rect 9458 6795 9497 6825
rect 9525 6795 9568 6825
rect 4402 6754 4441 6784
rect 4469 6754 4512 6784
rect 4402 6740 4512 6754
rect 419 6502 529 6516
rect 9458 6781 9568 6795
rect 5475 6543 5585 6557
rect 5475 6513 5518 6543
rect 5546 6513 5585 6543
rect 419 6472 462 6502
rect 490 6472 529 6502
rect 419 6457 529 6472
rect 3463 6474 3573 6489
rect 3463 6444 3502 6474
rect 3530 6444 3573 6474
rect 5475 6498 5585 6513
rect 3463 6430 3573 6444
rect 8519 6515 8629 6530
rect 8519 6485 8558 6515
rect 8586 6485 8629 6515
rect 8519 6471 8629 6485
rect 1499 6220 1609 6234
rect 4401 6230 4511 6245
rect 1499 6190 1542 6220
rect 1570 6190 1609 6220
rect 1499 6175 1609 6190
rect 4401 6200 4440 6230
rect 4468 6200 4511 6230
rect 6555 6261 6665 6275
rect 9457 6271 9567 6286
rect 4401 6186 4511 6200
rect 6555 6231 6598 6261
rect 6626 6231 6665 6261
rect 6555 6216 6665 6231
rect 9457 6241 9496 6271
rect 9524 6241 9567 6271
rect 9457 6227 9567 6241
rect 421 5953 531 5967
rect 421 5923 464 5953
rect 492 5923 531 5953
rect 3323 5963 3433 5978
rect 3323 5933 3362 5963
rect 3390 5933 3433 5963
rect 5477 5994 5587 6008
rect 421 5908 531 5923
rect 3323 5919 3433 5933
rect 5477 5964 5520 5994
rect 5548 5964 5587 5994
rect 8379 6004 8489 6019
rect 8379 5974 8418 6004
rect 8446 5974 8489 6004
rect 5477 5949 5587 5964
rect 8379 5960 8489 5974
rect 1359 5709 1469 5723
rect 1359 5679 1402 5709
rect 1430 5679 1469 5709
rect 1359 5664 1469 5679
rect 6415 5750 6525 5764
rect 4403 5681 4513 5696
rect 6415 5720 6458 5750
rect 6486 5720 6525 5750
rect 6415 5705 6525 5720
rect 9459 5722 9569 5737
rect 9459 5692 9498 5722
rect 9526 5692 9569 5722
rect 4403 5651 4442 5681
rect 4470 5651 4513 5681
rect 4403 5637 4513 5651
rect 420 5399 530 5413
rect 9459 5678 9569 5692
rect 5476 5440 5586 5454
rect 5476 5410 5519 5440
rect 5547 5410 5586 5440
rect 420 5369 463 5399
rect 491 5369 530 5399
rect 420 5354 530 5369
rect 3464 5371 3574 5386
rect 3464 5341 3503 5371
rect 3531 5341 3574 5371
rect 5476 5395 5586 5410
rect 3464 5327 3574 5341
rect 8520 5412 8630 5427
rect 8520 5382 8559 5412
rect 8587 5382 8630 5412
rect 8520 5368 8630 5382
rect 1468 5136 1578 5150
rect 1468 5106 1511 5136
rect 1539 5106 1578 5136
rect 4402 5127 4512 5142
rect 1468 5091 1578 5106
rect 4402 5097 4441 5127
rect 4469 5097 4512 5127
rect 6524 5177 6634 5191
rect 6524 5147 6567 5177
rect 6595 5147 6634 5177
rect 9458 5168 9568 5183
rect 6524 5132 6634 5147
rect 4402 5083 4512 5097
rect 9458 5138 9497 5168
rect 9525 5138 9568 5168
rect 9458 5124 9568 5138
rect 421 4850 531 4864
rect 421 4820 464 4850
rect 492 4820 531 4850
rect 5477 4891 5587 4905
rect 3355 4841 3465 4856
rect 421 4805 531 4820
rect 3355 4811 3394 4841
rect 3422 4811 3465 4841
rect 3355 4797 3465 4811
rect 5477 4861 5520 4891
rect 5548 4861 5587 4891
rect 8411 4882 8521 4897
rect 5477 4846 5587 4861
rect 8411 4852 8450 4882
rect 8478 4852 8521 4882
rect 8411 4838 8521 4852
rect 1359 4606 1469 4620
rect 1359 4576 1402 4606
rect 1430 4576 1469 4606
rect 1359 4561 1469 4576
rect 6415 4647 6525 4661
rect 4403 4578 4513 4593
rect 6415 4617 6458 4647
rect 6486 4617 6525 4647
rect 6415 4602 6525 4617
rect 9459 4619 9569 4634
rect 9459 4589 9498 4619
rect 9526 4589 9569 4619
rect 4403 4548 4442 4578
rect 4470 4548 4513 4578
rect 4403 4534 4513 4548
rect 420 4296 530 4310
rect 9459 4575 9569 4589
rect 5476 4337 5586 4351
rect 5476 4307 5519 4337
rect 5547 4307 5586 4337
rect 420 4266 463 4296
rect 491 4266 530 4296
rect 420 4251 530 4266
rect 3464 4268 3574 4283
rect 3464 4238 3503 4268
rect 3531 4238 3574 4268
rect 5476 4292 5586 4307
rect 3464 4224 3574 4238
rect 8520 4309 8630 4324
rect 8520 4279 8559 4309
rect 8587 4279 8630 4309
rect 8520 4265 8630 4279
rect 1500 4014 1610 4028
rect 4402 4024 4512 4039
rect 1500 3984 1543 4014
rect 1571 3984 1610 4014
rect 1500 3969 1610 3984
rect 4402 3994 4441 4024
rect 4469 3994 4512 4024
rect 6556 4055 6666 4069
rect 9458 4065 9568 4080
rect 4402 3980 4512 3994
rect 6556 4025 6599 4055
rect 6627 4025 6666 4055
rect 6556 4010 6666 4025
rect 9458 4035 9497 4065
rect 9525 4035 9568 4065
rect 9458 4021 9568 4035
rect 422 3747 532 3761
rect 422 3717 465 3747
rect 493 3717 532 3747
rect 3324 3757 3434 3772
rect 3324 3727 3363 3757
rect 3391 3727 3434 3757
rect 5478 3788 5588 3802
rect 422 3702 532 3717
rect 3324 3713 3434 3727
rect 5478 3758 5521 3788
rect 5549 3758 5588 3788
rect 8380 3798 8490 3813
rect 8380 3768 8419 3798
rect 8447 3768 8490 3798
rect 5478 3743 5588 3758
rect 8380 3754 8490 3768
rect 1360 3503 1470 3517
rect 1360 3473 1403 3503
rect 1431 3473 1470 3503
rect 1360 3458 1470 3473
rect 6416 3544 6526 3558
rect 4404 3475 4514 3490
rect 6416 3514 6459 3544
rect 6487 3514 6526 3544
rect 6416 3499 6526 3514
rect 9460 3516 9570 3531
rect 9460 3486 9499 3516
rect 9527 3486 9570 3516
rect 4404 3445 4443 3475
rect 4471 3445 4514 3475
rect 4404 3431 4514 3445
rect 421 3193 531 3207
rect 9460 3472 9570 3486
rect 5477 3234 5587 3248
rect 5477 3204 5520 3234
rect 5548 3204 5587 3234
rect 421 3163 464 3193
rect 492 3163 531 3193
rect 421 3148 531 3163
rect 3465 3165 3575 3180
rect 3465 3135 3504 3165
rect 3532 3135 3575 3165
rect 5477 3189 5587 3204
rect 3465 3121 3575 3135
rect 8521 3206 8631 3221
rect 8521 3176 8560 3206
rect 8588 3176 8631 3206
rect 8521 3162 8631 3176
rect 1470 2924 1580 2938
rect 1470 2894 1513 2924
rect 1541 2894 1580 2924
rect 4403 2921 4513 2936
rect 1470 2879 1580 2894
rect 4403 2891 4442 2921
rect 4470 2891 4513 2921
rect 6526 2965 6636 2979
rect 6526 2935 6569 2965
rect 6597 2935 6636 2965
rect 9459 2962 9569 2977
rect 6526 2920 6636 2935
rect 4403 2877 4513 2891
rect 9459 2932 9498 2962
rect 9526 2932 9569 2962
rect 9459 2918 9569 2932
rect 422 2644 532 2658
rect 422 2614 465 2644
rect 493 2614 532 2644
rect 5478 2685 5588 2699
rect 3355 2641 3465 2656
rect 422 2599 532 2614
rect 3355 2611 3394 2641
rect 3422 2611 3465 2641
rect 3355 2597 3465 2611
rect 5478 2655 5521 2685
rect 5549 2655 5588 2685
rect 8411 2682 8521 2697
rect 5478 2640 5588 2655
rect 8411 2652 8450 2682
rect 8478 2652 8521 2682
rect 8411 2638 8521 2652
rect 1360 2400 1470 2414
rect 1360 2370 1403 2400
rect 1431 2370 1470 2400
rect 1360 2355 1470 2370
rect 6416 2441 6526 2455
rect 4404 2372 4514 2387
rect 6416 2411 6459 2441
rect 6487 2411 6526 2441
rect 6416 2396 6526 2411
rect 9460 2413 9570 2428
rect 9460 2383 9499 2413
rect 9527 2383 9570 2413
rect 4404 2342 4443 2372
rect 4471 2342 4514 2372
rect 4404 2328 4514 2342
rect 421 2090 531 2104
rect 9460 2369 9570 2383
rect 5477 2131 5587 2145
rect 5477 2101 5520 2131
rect 5548 2101 5587 2131
rect 421 2060 464 2090
rect 492 2060 531 2090
rect 421 2045 531 2060
rect 3465 2062 3575 2077
rect 3465 2032 3504 2062
rect 3532 2032 3575 2062
rect 5477 2086 5587 2101
rect 3465 2018 3575 2032
rect 8521 2103 8631 2118
rect 8521 2073 8560 2103
rect 8588 2073 8631 2103
rect 8521 2059 8631 2073
rect 1501 1808 1611 1822
rect 4403 1818 4513 1833
rect 1501 1778 1544 1808
rect 1572 1778 1611 1808
rect 1501 1763 1611 1778
rect 4403 1788 4442 1818
rect 4470 1788 4513 1818
rect 6557 1849 6667 1863
rect 9459 1859 9569 1874
rect 4403 1774 4513 1788
rect 6557 1819 6600 1849
rect 6628 1819 6667 1849
rect 6557 1804 6667 1819
rect 9459 1829 9498 1859
rect 9526 1829 9569 1859
rect 9459 1815 9569 1829
rect 423 1541 533 1555
rect 423 1511 466 1541
rect 494 1511 533 1541
rect 3325 1551 3435 1566
rect 3325 1521 3364 1551
rect 3392 1521 3435 1551
rect 5479 1582 5589 1596
rect 423 1496 533 1511
rect 3325 1507 3435 1521
rect 5479 1552 5522 1582
rect 5550 1552 5589 1582
rect 8381 1592 8491 1607
rect 8381 1562 8420 1592
rect 8448 1562 8491 1592
rect 5479 1537 5589 1552
rect 8381 1548 8491 1562
rect 1361 1297 1471 1311
rect 1361 1267 1404 1297
rect 1432 1267 1471 1297
rect 1361 1252 1471 1267
rect 6417 1338 6527 1352
rect 4405 1269 4515 1284
rect 6417 1308 6460 1338
rect 6488 1308 6527 1338
rect 6417 1293 6527 1308
rect 9461 1310 9571 1325
rect 9461 1280 9500 1310
rect 9528 1280 9571 1310
rect 4405 1239 4444 1269
rect 4472 1239 4515 1269
rect 4405 1225 4515 1239
rect 422 987 532 1001
rect 9461 1266 9571 1280
rect 5478 1028 5588 1042
rect 5478 998 5521 1028
rect 5549 998 5588 1028
rect 422 957 465 987
rect 493 957 532 987
rect 422 942 532 957
rect 3466 959 3576 974
rect 3466 929 3505 959
rect 3533 929 3576 959
rect 5478 983 5588 998
rect 3466 915 3576 929
rect 8522 1000 8632 1015
rect 8522 970 8561 1000
rect 8589 970 8632 1000
rect 8522 956 8632 970
rect 4404 715 4514 730
rect 4404 685 4443 715
rect 4471 685 4514 715
rect 9460 756 9570 771
rect 9460 726 9499 756
rect 9527 726 9570 756
rect 9460 712 9570 726
rect 4404 671 4514 685
rect 6725 469 6835 483
rect 1669 428 1779 442
rect 1669 398 1712 428
rect 1740 398 1779 428
rect 6725 439 6768 469
rect 6796 439 6835 469
rect 6725 424 6835 439
rect 1669 383 1779 398
rect 4619 408 4729 422
rect 4619 378 4662 408
rect 4690 378 4729 408
rect 4619 363 4729 378
<< psubdiffcont >>
rect 9499 9348 9527 9378
rect 4443 9307 4471 9337
rect 3504 8997 3532 9027
rect 8560 9038 8588 9068
rect 459 8885 487 8915
rect 5515 8926 5543 8956
rect 4442 8753 4470 8783
rect 9498 8794 9526 8824
rect 1397 8641 1425 8671
rect 6453 8682 6481 8712
rect 3364 8486 3392 8516
rect 8420 8527 8448 8557
rect 458 8331 486 8361
rect 5514 8372 5542 8402
rect 4444 8204 4472 8234
rect 9500 8245 9528 8275
rect 1538 8049 1566 8079
rect 6594 8090 6622 8120
rect 3505 7894 3533 7924
rect 8561 7935 8589 7965
rect 460 7782 488 7812
rect 5516 7823 5544 7853
rect 4443 7650 4471 7680
rect 9499 7691 9527 7721
rect 1398 7538 1426 7568
rect 6454 7579 6482 7609
rect 3395 7370 3423 7400
rect 8451 7411 8479 7441
rect 459 7228 487 7258
rect 5515 7269 5543 7299
rect 4444 7101 4472 7131
rect 9500 7142 9528 7172
rect 1508 6959 1536 6989
rect 6564 7000 6592 7030
rect 3505 6791 3533 6821
rect 8561 6832 8589 6862
rect 460 6679 488 6709
rect 5516 6720 5544 6750
rect 4443 6547 4471 6577
rect 9499 6588 9527 6618
rect 1398 6435 1426 6465
rect 6454 6476 6482 6506
rect 3365 6280 3393 6310
rect 8421 6321 8449 6351
rect 459 6125 487 6155
rect 5515 6166 5543 6196
rect 4445 5998 4473 6028
rect 9501 6039 9529 6069
rect 1539 5843 1567 5873
rect 6595 5884 6623 5914
rect 3506 5688 3534 5718
rect 8562 5729 8590 5759
rect 461 5576 489 5606
rect 5517 5617 5545 5647
rect 4444 5444 4472 5474
rect 9500 5485 9528 5515
rect 1399 5332 1427 5362
rect 6455 5373 6483 5403
rect 3397 5158 3425 5188
rect 8453 5199 8481 5229
rect 460 5022 488 5052
rect 5516 5063 5544 5093
rect 4445 4895 4473 4925
rect 9501 4936 9529 4966
rect 1508 4759 1536 4789
rect 6564 4800 6592 4830
rect 3506 4585 3534 4615
rect 8562 4626 8590 4656
rect 461 4473 489 4503
rect 5517 4514 5545 4544
rect 4444 4341 4472 4371
rect 9500 4382 9528 4412
rect 1399 4229 1427 4259
rect 6455 4270 6483 4300
rect 3366 4074 3394 4104
rect 8422 4115 8450 4145
rect 460 3919 488 3949
rect 5516 3960 5544 3990
rect 4446 3792 4474 3822
rect 9502 3833 9530 3863
rect 1540 3637 1568 3667
rect 6596 3678 6624 3708
rect 3507 3482 3535 3512
rect 8563 3523 8591 3553
rect 462 3370 490 3400
rect 5518 3411 5546 3441
rect 4445 3238 4473 3268
rect 9501 3279 9529 3309
rect 1400 3126 1428 3156
rect 6456 3167 6484 3197
rect 3397 2958 3425 2988
rect 8453 2999 8481 3029
rect 461 2816 489 2846
rect 5517 2857 5545 2887
rect 4446 2689 4474 2719
rect 9502 2730 9530 2760
rect 1510 2547 1538 2577
rect 6566 2588 6594 2618
rect 3507 2379 3535 2409
rect 8563 2420 8591 2450
rect 462 2267 490 2297
rect 5518 2308 5546 2338
rect 4445 2135 4473 2165
rect 9501 2176 9529 2206
rect 1400 2023 1428 2053
rect 6456 2064 6484 2094
rect 3367 1868 3395 1898
rect 8423 1909 8451 1939
rect 461 1713 489 1743
rect 5517 1754 5545 1784
rect 4447 1586 4475 1616
rect 9503 1627 9531 1657
rect 1541 1431 1569 1461
rect 6597 1472 6625 1502
rect 3508 1276 3536 1306
rect 8564 1317 8592 1347
rect 463 1164 491 1194
rect 5519 1205 5547 1235
rect 4446 1032 4474 1062
rect 9502 1073 9530 1103
rect 1401 920 1429 950
rect 6457 961 6485 991
rect 5518 651 5546 681
rect 462 610 490 640
rect 1709 51 1737 81
rect 6765 92 6793 122
rect 4659 31 4687 61
<< nsubdiffcont >>
rect 462 9232 490 9262
rect 5518 9273 5546 9303
rect 1400 8988 1428 9018
rect 6456 9029 6484 9059
rect 9496 9001 9524 9031
rect 4440 8960 4468 8990
rect 5517 8719 5545 8749
rect 461 8678 489 8708
rect 3501 8650 3529 8680
rect 8557 8691 8585 8721
rect 1541 8396 1569 8426
rect 4439 8406 4467 8436
rect 6597 8437 6625 8467
rect 9495 8447 9523 8477
rect 463 8129 491 8159
rect 3361 8139 3389 8169
rect 5519 8170 5547 8200
rect 8417 8180 8445 8210
rect 1401 7885 1429 7915
rect 6457 7926 6485 7956
rect 9497 7898 9525 7928
rect 4441 7857 4469 7887
rect 5518 7616 5546 7646
rect 462 7575 490 7605
rect 3502 7547 3530 7577
rect 8558 7588 8586 7618
rect 1511 7306 1539 7336
rect 4440 7303 4468 7333
rect 6567 7347 6595 7377
rect 9496 7344 9524 7374
rect 463 7026 491 7056
rect 3392 7023 3420 7053
rect 5519 7067 5547 7097
rect 8448 7064 8476 7094
rect 1401 6782 1429 6812
rect 6457 6823 6485 6853
rect 9497 6795 9525 6825
rect 4441 6754 4469 6784
rect 5518 6513 5546 6543
rect 462 6472 490 6502
rect 3502 6444 3530 6474
rect 8558 6485 8586 6515
rect 1542 6190 1570 6220
rect 4440 6200 4468 6230
rect 6598 6231 6626 6261
rect 9496 6241 9524 6271
rect 464 5923 492 5953
rect 3362 5933 3390 5963
rect 5520 5964 5548 5994
rect 8418 5974 8446 6004
rect 1402 5679 1430 5709
rect 6458 5720 6486 5750
rect 9498 5692 9526 5722
rect 4442 5651 4470 5681
rect 5519 5410 5547 5440
rect 463 5369 491 5399
rect 3503 5341 3531 5371
rect 8559 5382 8587 5412
rect 1511 5106 1539 5136
rect 4441 5097 4469 5127
rect 6567 5147 6595 5177
rect 9497 5138 9525 5168
rect 464 4820 492 4850
rect 3394 4811 3422 4841
rect 5520 4861 5548 4891
rect 8450 4852 8478 4882
rect 1402 4576 1430 4606
rect 6458 4617 6486 4647
rect 9498 4589 9526 4619
rect 4442 4548 4470 4578
rect 5519 4307 5547 4337
rect 463 4266 491 4296
rect 3503 4238 3531 4268
rect 8559 4279 8587 4309
rect 1543 3984 1571 4014
rect 4441 3994 4469 4024
rect 6599 4025 6627 4055
rect 9497 4035 9525 4065
rect 465 3717 493 3747
rect 3363 3727 3391 3757
rect 5521 3758 5549 3788
rect 8419 3768 8447 3798
rect 1403 3473 1431 3503
rect 6459 3514 6487 3544
rect 9499 3486 9527 3516
rect 4443 3445 4471 3475
rect 5520 3204 5548 3234
rect 464 3163 492 3193
rect 3504 3135 3532 3165
rect 8560 3176 8588 3206
rect 1513 2894 1541 2924
rect 4442 2891 4470 2921
rect 6569 2935 6597 2965
rect 9498 2932 9526 2962
rect 465 2614 493 2644
rect 3394 2611 3422 2641
rect 5521 2655 5549 2685
rect 8450 2652 8478 2682
rect 1403 2370 1431 2400
rect 6459 2411 6487 2441
rect 9499 2383 9527 2413
rect 4443 2342 4471 2372
rect 5520 2101 5548 2131
rect 464 2060 492 2090
rect 3504 2032 3532 2062
rect 8560 2073 8588 2103
rect 1544 1778 1572 1808
rect 4442 1788 4470 1818
rect 6600 1819 6628 1849
rect 9498 1829 9526 1859
rect 466 1511 494 1541
rect 3364 1521 3392 1551
rect 5522 1552 5550 1582
rect 8420 1562 8448 1592
rect 1404 1267 1432 1297
rect 6460 1308 6488 1338
rect 9500 1280 9528 1310
rect 4444 1239 4472 1269
rect 5521 998 5549 1028
rect 465 957 493 987
rect 3505 929 3533 959
rect 8561 970 8589 1000
rect 4443 685 4471 715
rect 9499 726 9527 756
rect 1712 398 1740 428
rect 6768 439 6796 469
rect 4662 378 4690 408
<< poly >>
rect 3869 9252 3919 9268
rect 4077 9252 4127 9268
rect 4285 9252 4335 9268
rect 4498 9252 4548 9268
rect 8925 9293 8975 9309
rect 9133 9293 9183 9309
rect 9341 9293 9391 9309
rect 9554 9293 9604 9309
rect 5438 9230 5488 9243
rect 5651 9230 5701 9243
rect 5859 9230 5909 9243
rect 6067 9230 6117 9243
rect 382 9189 432 9202
rect 595 9189 645 9202
rect 803 9189 853 9202
rect 1011 9189 1061 9202
rect 3869 9185 3919 9210
rect 3869 9159 3875 9185
rect 3901 9159 3919 9185
rect 3869 9133 3919 9159
rect 4077 9181 4127 9210
rect 4077 9157 4091 9181
rect 4115 9157 4127 9181
rect 4077 9133 4127 9157
rect 4285 9186 4335 9210
rect 4285 9162 4300 9186
rect 4324 9162 4335 9186
rect 4285 9133 4335 9162
rect 4498 9181 4548 9210
rect 4498 9161 4515 9181
rect 4535 9161 4548 9181
rect 4498 9133 4548 9161
rect 382 9061 432 9089
rect 382 9041 395 9061
rect 415 9041 432 9061
rect 382 9012 432 9041
rect 595 9060 645 9089
rect 595 9036 606 9060
rect 630 9036 645 9060
rect 595 9012 645 9036
rect 803 9065 853 9089
rect 803 9041 815 9065
rect 839 9041 853 9065
rect 803 9012 853 9041
rect 1011 9063 1061 9089
rect 1011 9037 1029 9063
rect 1055 9037 1061 9063
rect 1011 9012 1061 9037
rect 8925 9226 8975 9251
rect 8925 9200 8931 9226
rect 8957 9200 8975 9226
rect 8925 9174 8975 9200
rect 9133 9222 9183 9251
rect 9133 9198 9147 9222
rect 9171 9198 9183 9222
rect 9133 9174 9183 9198
rect 9341 9227 9391 9251
rect 9341 9203 9356 9227
rect 9380 9203 9391 9227
rect 9341 9174 9391 9203
rect 9554 9222 9604 9251
rect 9554 9202 9571 9222
rect 9591 9202 9604 9222
rect 9554 9174 9604 9202
rect 5438 9102 5488 9130
rect 5438 9082 5451 9102
rect 5471 9082 5488 9102
rect 3869 9020 3919 9033
rect 4077 9020 4127 9033
rect 4285 9020 4335 9033
rect 4498 9020 4548 9033
rect 5438 9053 5488 9082
rect 5651 9101 5701 9130
rect 5651 9077 5662 9101
rect 5686 9077 5701 9101
rect 5651 9053 5701 9077
rect 5859 9106 5909 9130
rect 5859 9082 5871 9106
rect 5895 9082 5909 9106
rect 5859 9053 5909 9082
rect 6067 9104 6117 9130
rect 6067 9078 6085 9104
rect 6111 9078 6117 9104
rect 6067 9053 6117 9078
rect 8925 9061 8975 9074
rect 9133 9061 9183 9074
rect 9341 9061 9391 9074
rect 9554 9061 9604 9074
rect 5438 8995 5488 9011
rect 5651 8995 5701 9011
rect 5859 8995 5909 9011
rect 6067 8995 6117 9011
rect 382 8954 432 8970
rect 595 8954 645 8970
rect 803 8954 853 8970
rect 1011 8954 1061 8970
rect 6376 8986 6426 8999
rect 6589 8986 6639 8999
rect 6797 8986 6847 8999
rect 7005 8986 7055 8999
rect 1320 8945 1370 8958
rect 1533 8945 1583 8958
rect 1741 8945 1791 8958
rect 1949 8945 1999 8958
rect 2930 8942 2980 8958
rect 3138 8942 3188 8958
rect 3346 8942 3396 8958
rect 3559 8942 3609 8958
rect 2930 8875 2980 8900
rect 2930 8849 2936 8875
rect 2962 8849 2980 8875
rect 1320 8817 1370 8845
rect 1320 8797 1333 8817
rect 1353 8797 1370 8817
rect 1320 8768 1370 8797
rect 1533 8816 1583 8845
rect 1533 8792 1544 8816
rect 1568 8792 1583 8816
rect 1533 8768 1583 8792
rect 1741 8821 1791 8845
rect 1741 8797 1753 8821
rect 1777 8797 1791 8821
rect 1741 8768 1791 8797
rect 1949 8819 1999 8845
rect 2930 8823 2980 8849
rect 3138 8871 3188 8900
rect 3138 8847 3152 8871
rect 3176 8847 3188 8871
rect 3138 8823 3188 8847
rect 3346 8876 3396 8900
rect 3346 8852 3361 8876
rect 3385 8852 3396 8876
rect 3346 8823 3396 8852
rect 3559 8871 3609 8900
rect 3559 8851 3576 8871
rect 3596 8851 3609 8871
rect 3559 8823 3609 8851
rect 1949 8793 1967 8819
rect 1993 8793 1999 8819
rect 1949 8768 1999 8793
rect 1320 8710 1370 8726
rect 1533 8710 1583 8726
rect 1741 8710 1791 8726
rect 1949 8710 1999 8726
rect 7986 8983 8036 8999
rect 8194 8983 8244 8999
rect 8402 8983 8452 8999
rect 8615 8983 8665 8999
rect 7986 8916 8036 8941
rect 7986 8890 7992 8916
rect 8018 8890 8036 8916
rect 6376 8858 6426 8886
rect 6376 8838 6389 8858
rect 6409 8838 6426 8858
rect 6376 8809 6426 8838
rect 6589 8857 6639 8886
rect 6589 8833 6600 8857
rect 6624 8833 6639 8857
rect 6589 8809 6639 8833
rect 6797 8862 6847 8886
rect 6797 8838 6809 8862
rect 6833 8838 6847 8862
rect 6797 8809 6847 8838
rect 7005 8860 7055 8886
rect 7986 8864 8036 8890
rect 8194 8912 8244 8941
rect 8194 8888 8208 8912
rect 8232 8888 8244 8912
rect 8194 8864 8244 8888
rect 8402 8917 8452 8941
rect 8402 8893 8417 8917
rect 8441 8893 8452 8917
rect 8402 8864 8452 8893
rect 8615 8912 8665 8941
rect 8615 8892 8632 8912
rect 8652 8892 8665 8912
rect 8615 8864 8665 8892
rect 7005 8834 7023 8860
rect 7049 8834 7055 8860
rect 7005 8809 7055 8834
rect 6376 8751 6426 8767
rect 6589 8751 6639 8767
rect 6797 8751 6847 8767
rect 7005 8751 7055 8767
rect 7986 8751 8036 8764
rect 8194 8751 8244 8764
rect 8402 8751 8452 8764
rect 8615 8751 8665 8764
rect 2930 8710 2980 8723
rect 3138 8710 3188 8723
rect 3346 8710 3396 8723
rect 3559 8710 3609 8723
rect 8924 8739 8974 8755
rect 9132 8739 9182 8755
rect 9340 8739 9390 8755
rect 9553 8739 9603 8755
rect 3868 8698 3918 8714
rect 4076 8698 4126 8714
rect 4284 8698 4334 8714
rect 4497 8698 4547 8714
rect 381 8635 431 8648
rect 594 8635 644 8648
rect 802 8635 852 8648
rect 1010 8635 1060 8648
rect 3868 8631 3918 8656
rect 3868 8605 3874 8631
rect 3900 8605 3918 8631
rect 3868 8579 3918 8605
rect 4076 8627 4126 8656
rect 4076 8603 4090 8627
rect 4114 8603 4126 8627
rect 4076 8579 4126 8603
rect 4284 8632 4334 8656
rect 4284 8608 4299 8632
rect 4323 8608 4334 8632
rect 4284 8579 4334 8608
rect 4497 8627 4547 8656
rect 5437 8676 5487 8689
rect 5650 8676 5700 8689
rect 5858 8676 5908 8689
rect 6066 8676 6116 8689
rect 4497 8607 4514 8627
rect 4534 8607 4547 8627
rect 4497 8579 4547 8607
rect 381 8507 431 8535
rect 381 8487 394 8507
rect 414 8487 431 8507
rect 381 8458 431 8487
rect 594 8506 644 8535
rect 594 8482 605 8506
rect 629 8482 644 8506
rect 594 8458 644 8482
rect 802 8511 852 8535
rect 802 8487 814 8511
rect 838 8487 852 8511
rect 802 8458 852 8487
rect 1010 8509 1060 8535
rect 1010 8483 1028 8509
rect 1054 8483 1060 8509
rect 1010 8458 1060 8483
rect 8924 8672 8974 8697
rect 8924 8646 8930 8672
rect 8956 8646 8974 8672
rect 8924 8620 8974 8646
rect 9132 8668 9182 8697
rect 9132 8644 9146 8668
rect 9170 8644 9182 8668
rect 9132 8620 9182 8644
rect 9340 8673 9390 8697
rect 9340 8649 9355 8673
rect 9379 8649 9390 8673
rect 9340 8620 9390 8649
rect 9553 8668 9603 8697
rect 9553 8648 9570 8668
rect 9590 8648 9603 8668
rect 9553 8620 9603 8648
rect 5437 8548 5487 8576
rect 5437 8528 5450 8548
rect 5470 8528 5487 8548
rect 5437 8499 5487 8528
rect 5650 8547 5700 8576
rect 5650 8523 5661 8547
rect 5685 8523 5700 8547
rect 5650 8499 5700 8523
rect 5858 8552 5908 8576
rect 5858 8528 5870 8552
rect 5894 8528 5908 8552
rect 5858 8499 5908 8528
rect 6066 8550 6116 8576
rect 6066 8524 6084 8550
rect 6110 8524 6116 8550
rect 6066 8499 6116 8524
rect 8924 8507 8974 8520
rect 9132 8507 9182 8520
rect 9340 8507 9390 8520
rect 9553 8507 9603 8520
rect 3868 8466 3918 8479
rect 4076 8466 4126 8479
rect 4284 8466 4334 8479
rect 4497 8466 4547 8479
rect 2790 8431 2840 8447
rect 2998 8431 3048 8447
rect 3206 8431 3256 8447
rect 3419 8431 3469 8447
rect 381 8400 431 8416
rect 594 8400 644 8416
rect 802 8400 852 8416
rect 1010 8400 1060 8416
rect 7846 8472 7896 8488
rect 8054 8472 8104 8488
rect 8262 8472 8312 8488
rect 8475 8472 8525 8488
rect 5437 8441 5487 8457
rect 5650 8441 5700 8457
rect 5858 8441 5908 8457
rect 6066 8441 6116 8457
rect 1461 8353 1511 8366
rect 1674 8353 1724 8366
rect 1882 8353 1932 8366
rect 2090 8353 2140 8366
rect 2790 8364 2840 8389
rect 2790 8338 2796 8364
rect 2822 8338 2840 8364
rect 2790 8312 2840 8338
rect 2998 8360 3048 8389
rect 2998 8336 3012 8360
rect 3036 8336 3048 8360
rect 2998 8312 3048 8336
rect 3206 8365 3256 8389
rect 3206 8341 3221 8365
rect 3245 8341 3256 8365
rect 3206 8312 3256 8341
rect 3419 8360 3469 8389
rect 6517 8394 6567 8407
rect 6730 8394 6780 8407
rect 6938 8394 6988 8407
rect 7146 8394 7196 8407
rect 7846 8405 7896 8430
rect 3419 8340 3436 8360
rect 3456 8340 3469 8360
rect 3419 8312 3469 8340
rect 1461 8225 1511 8253
rect 1461 8205 1474 8225
rect 1494 8205 1511 8225
rect 1461 8176 1511 8205
rect 1674 8224 1724 8253
rect 1674 8200 1685 8224
rect 1709 8200 1724 8224
rect 1674 8176 1724 8200
rect 1882 8229 1932 8253
rect 1882 8205 1894 8229
rect 1918 8205 1932 8229
rect 1882 8176 1932 8205
rect 2090 8227 2140 8253
rect 2090 8201 2108 8227
rect 2134 8201 2140 8227
rect 7846 8379 7852 8405
rect 7878 8379 7896 8405
rect 7846 8353 7896 8379
rect 8054 8401 8104 8430
rect 8054 8377 8068 8401
rect 8092 8377 8104 8401
rect 8054 8353 8104 8377
rect 8262 8406 8312 8430
rect 8262 8382 8277 8406
rect 8301 8382 8312 8406
rect 8262 8353 8312 8382
rect 8475 8401 8525 8430
rect 8475 8381 8492 8401
rect 8512 8381 8525 8401
rect 8475 8353 8525 8381
rect 6517 8266 6567 8294
rect 6517 8246 6530 8266
rect 6550 8246 6567 8266
rect 2090 8176 2140 8201
rect 2790 8199 2840 8212
rect 2998 8199 3048 8212
rect 3206 8199 3256 8212
rect 3419 8199 3469 8212
rect 6517 8217 6567 8246
rect 6730 8265 6780 8294
rect 6730 8241 6741 8265
rect 6765 8241 6780 8265
rect 6730 8217 6780 8241
rect 6938 8270 6988 8294
rect 6938 8246 6950 8270
rect 6974 8246 6988 8270
rect 6938 8217 6988 8246
rect 7146 8268 7196 8294
rect 7146 8242 7164 8268
rect 7190 8242 7196 8268
rect 7146 8217 7196 8242
rect 7846 8240 7896 8253
rect 8054 8240 8104 8253
rect 8262 8240 8312 8253
rect 8475 8240 8525 8253
rect 3870 8149 3920 8165
rect 4078 8149 4128 8165
rect 4286 8149 4336 8165
rect 4499 8149 4549 8165
rect 1461 8118 1511 8134
rect 1674 8118 1724 8134
rect 1882 8118 1932 8134
rect 2090 8118 2140 8134
rect 8926 8190 8976 8206
rect 9134 8190 9184 8206
rect 9342 8190 9392 8206
rect 9555 8190 9605 8206
rect 6517 8159 6567 8175
rect 6730 8159 6780 8175
rect 6938 8159 6988 8175
rect 7146 8159 7196 8175
rect 5439 8127 5489 8140
rect 5652 8127 5702 8140
rect 5860 8127 5910 8140
rect 6068 8127 6118 8140
rect 383 8086 433 8099
rect 596 8086 646 8099
rect 804 8086 854 8099
rect 1012 8086 1062 8099
rect 3870 8082 3920 8107
rect 3870 8056 3876 8082
rect 3902 8056 3920 8082
rect 3870 8030 3920 8056
rect 4078 8078 4128 8107
rect 4078 8054 4092 8078
rect 4116 8054 4128 8078
rect 4078 8030 4128 8054
rect 4286 8083 4336 8107
rect 4286 8059 4301 8083
rect 4325 8059 4336 8083
rect 4286 8030 4336 8059
rect 4499 8078 4549 8107
rect 4499 8058 4516 8078
rect 4536 8058 4549 8078
rect 4499 8030 4549 8058
rect 383 7958 433 7986
rect 383 7938 396 7958
rect 416 7938 433 7958
rect 383 7909 433 7938
rect 596 7957 646 7986
rect 596 7933 607 7957
rect 631 7933 646 7957
rect 596 7909 646 7933
rect 804 7962 854 7986
rect 804 7938 816 7962
rect 840 7938 854 7962
rect 804 7909 854 7938
rect 1012 7960 1062 7986
rect 1012 7934 1030 7960
rect 1056 7934 1062 7960
rect 1012 7909 1062 7934
rect 8926 8123 8976 8148
rect 8926 8097 8932 8123
rect 8958 8097 8976 8123
rect 8926 8071 8976 8097
rect 9134 8119 9184 8148
rect 9134 8095 9148 8119
rect 9172 8095 9184 8119
rect 9134 8071 9184 8095
rect 9342 8124 9392 8148
rect 9342 8100 9357 8124
rect 9381 8100 9392 8124
rect 9342 8071 9392 8100
rect 9555 8119 9605 8148
rect 9555 8099 9572 8119
rect 9592 8099 9605 8119
rect 9555 8071 9605 8099
rect 5439 7999 5489 8027
rect 5439 7979 5452 7999
rect 5472 7979 5489 7999
rect 3870 7917 3920 7930
rect 4078 7917 4128 7930
rect 4286 7917 4336 7930
rect 4499 7917 4549 7930
rect 5439 7950 5489 7979
rect 5652 7998 5702 8027
rect 5652 7974 5663 7998
rect 5687 7974 5702 7998
rect 5652 7950 5702 7974
rect 5860 8003 5910 8027
rect 5860 7979 5872 8003
rect 5896 7979 5910 8003
rect 5860 7950 5910 7979
rect 6068 8001 6118 8027
rect 6068 7975 6086 8001
rect 6112 7975 6118 8001
rect 6068 7950 6118 7975
rect 8926 7958 8976 7971
rect 9134 7958 9184 7971
rect 9342 7958 9392 7971
rect 9555 7958 9605 7971
rect 5439 7892 5489 7908
rect 5652 7892 5702 7908
rect 5860 7892 5910 7908
rect 6068 7892 6118 7908
rect 383 7851 433 7867
rect 596 7851 646 7867
rect 804 7851 854 7867
rect 1012 7851 1062 7867
rect 6377 7883 6427 7896
rect 6590 7883 6640 7896
rect 6798 7883 6848 7896
rect 7006 7883 7056 7896
rect 1321 7842 1371 7855
rect 1534 7842 1584 7855
rect 1742 7842 1792 7855
rect 1950 7842 2000 7855
rect 2931 7839 2981 7855
rect 3139 7839 3189 7855
rect 3347 7839 3397 7855
rect 3560 7839 3610 7855
rect 2931 7772 2981 7797
rect 2931 7746 2937 7772
rect 2963 7746 2981 7772
rect 1321 7714 1371 7742
rect 1321 7694 1334 7714
rect 1354 7694 1371 7714
rect 1321 7665 1371 7694
rect 1534 7713 1584 7742
rect 1534 7689 1545 7713
rect 1569 7689 1584 7713
rect 1534 7665 1584 7689
rect 1742 7718 1792 7742
rect 1742 7694 1754 7718
rect 1778 7694 1792 7718
rect 1742 7665 1792 7694
rect 1950 7716 2000 7742
rect 2931 7720 2981 7746
rect 3139 7768 3189 7797
rect 3139 7744 3153 7768
rect 3177 7744 3189 7768
rect 3139 7720 3189 7744
rect 3347 7773 3397 7797
rect 3347 7749 3362 7773
rect 3386 7749 3397 7773
rect 3347 7720 3397 7749
rect 3560 7768 3610 7797
rect 3560 7748 3577 7768
rect 3597 7748 3610 7768
rect 3560 7720 3610 7748
rect 1950 7690 1968 7716
rect 1994 7690 2000 7716
rect 1950 7665 2000 7690
rect 1321 7607 1371 7623
rect 1534 7607 1584 7623
rect 1742 7607 1792 7623
rect 1950 7607 2000 7623
rect 7987 7880 8037 7896
rect 8195 7880 8245 7896
rect 8403 7880 8453 7896
rect 8616 7880 8666 7896
rect 7987 7813 8037 7838
rect 7987 7787 7993 7813
rect 8019 7787 8037 7813
rect 6377 7755 6427 7783
rect 6377 7735 6390 7755
rect 6410 7735 6427 7755
rect 6377 7706 6427 7735
rect 6590 7754 6640 7783
rect 6590 7730 6601 7754
rect 6625 7730 6640 7754
rect 6590 7706 6640 7730
rect 6798 7759 6848 7783
rect 6798 7735 6810 7759
rect 6834 7735 6848 7759
rect 6798 7706 6848 7735
rect 7006 7757 7056 7783
rect 7987 7761 8037 7787
rect 8195 7809 8245 7838
rect 8195 7785 8209 7809
rect 8233 7785 8245 7809
rect 8195 7761 8245 7785
rect 8403 7814 8453 7838
rect 8403 7790 8418 7814
rect 8442 7790 8453 7814
rect 8403 7761 8453 7790
rect 8616 7809 8666 7838
rect 8616 7789 8633 7809
rect 8653 7789 8666 7809
rect 8616 7761 8666 7789
rect 7006 7731 7024 7757
rect 7050 7731 7056 7757
rect 7006 7706 7056 7731
rect 6377 7648 6427 7664
rect 6590 7648 6640 7664
rect 6798 7648 6848 7664
rect 7006 7648 7056 7664
rect 7987 7648 8037 7661
rect 8195 7648 8245 7661
rect 8403 7648 8453 7661
rect 8616 7648 8666 7661
rect 2931 7607 2981 7620
rect 3139 7607 3189 7620
rect 3347 7607 3397 7620
rect 3560 7607 3610 7620
rect 8925 7636 8975 7652
rect 9133 7636 9183 7652
rect 9341 7636 9391 7652
rect 9554 7636 9604 7652
rect 3869 7595 3919 7611
rect 4077 7595 4127 7611
rect 4285 7595 4335 7611
rect 4498 7595 4548 7611
rect 382 7532 432 7545
rect 595 7532 645 7545
rect 803 7532 853 7545
rect 1011 7532 1061 7545
rect 3869 7528 3919 7553
rect 3869 7502 3875 7528
rect 3901 7502 3919 7528
rect 3869 7476 3919 7502
rect 4077 7524 4127 7553
rect 4077 7500 4091 7524
rect 4115 7500 4127 7524
rect 4077 7476 4127 7500
rect 4285 7529 4335 7553
rect 4285 7505 4300 7529
rect 4324 7505 4335 7529
rect 4285 7476 4335 7505
rect 4498 7524 4548 7553
rect 5438 7573 5488 7586
rect 5651 7573 5701 7586
rect 5859 7573 5909 7586
rect 6067 7573 6117 7586
rect 4498 7504 4515 7524
rect 4535 7504 4548 7524
rect 4498 7476 4548 7504
rect 382 7404 432 7432
rect 382 7384 395 7404
rect 415 7384 432 7404
rect 382 7355 432 7384
rect 595 7403 645 7432
rect 595 7379 606 7403
rect 630 7379 645 7403
rect 595 7355 645 7379
rect 803 7408 853 7432
rect 803 7384 815 7408
rect 839 7384 853 7408
rect 803 7355 853 7384
rect 1011 7406 1061 7432
rect 1011 7380 1029 7406
rect 1055 7380 1061 7406
rect 1011 7355 1061 7380
rect 8925 7569 8975 7594
rect 8925 7543 8931 7569
rect 8957 7543 8975 7569
rect 8925 7517 8975 7543
rect 9133 7565 9183 7594
rect 9133 7541 9147 7565
rect 9171 7541 9183 7565
rect 9133 7517 9183 7541
rect 9341 7570 9391 7594
rect 9341 7546 9356 7570
rect 9380 7546 9391 7570
rect 9341 7517 9391 7546
rect 9554 7565 9604 7594
rect 9554 7545 9571 7565
rect 9591 7545 9604 7565
rect 9554 7517 9604 7545
rect 5438 7445 5488 7473
rect 5438 7425 5451 7445
rect 5471 7425 5488 7445
rect 5438 7396 5488 7425
rect 5651 7444 5701 7473
rect 5651 7420 5662 7444
rect 5686 7420 5701 7444
rect 5651 7396 5701 7420
rect 5859 7449 5909 7473
rect 5859 7425 5871 7449
rect 5895 7425 5909 7449
rect 5859 7396 5909 7425
rect 6067 7447 6117 7473
rect 6067 7421 6085 7447
rect 6111 7421 6117 7447
rect 6067 7396 6117 7421
rect 8925 7404 8975 7417
rect 9133 7404 9183 7417
rect 9341 7404 9391 7417
rect 9554 7404 9604 7417
rect 3869 7363 3919 7376
rect 4077 7363 4127 7376
rect 4285 7363 4335 7376
rect 4498 7363 4548 7376
rect 382 7297 432 7313
rect 595 7297 645 7313
rect 803 7297 853 7313
rect 1011 7297 1061 7313
rect 2821 7315 2871 7331
rect 3029 7315 3079 7331
rect 3237 7315 3287 7331
rect 3450 7315 3500 7331
rect 1431 7263 1481 7276
rect 1644 7263 1694 7276
rect 1852 7263 1902 7276
rect 2060 7263 2110 7276
rect 5438 7338 5488 7354
rect 5651 7338 5701 7354
rect 5859 7338 5909 7354
rect 6067 7338 6117 7354
rect 7877 7356 7927 7372
rect 8085 7356 8135 7372
rect 8293 7356 8343 7372
rect 8506 7356 8556 7372
rect 6487 7304 6537 7317
rect 6700 7304 6750 7317
rect 6908 7304 6958 7317
rect 7116 7304 7166 7317
rect 2821 7248 2871 7273
rect 2821 7222 2827 7248
rect 2853 7222 2871 7248
rect 2821 7196 2871 7222
rect 3029 7244 3079 7273
rect 3029 7220 3043 7244
rect 3067 7220 3079 7244
rect 3029 7196 3079 7220
rect 3237 7249 3287 7273
rect 3237 7225 3252 7249
rect 3276 7225 3287 7249
rect 3237 7196 3287 7225
rect 3450 7244 3500 7273
rect 3450 7224 3467 7244
rect 3487 7224 3500 7244
rect 3450 7196 3500 7224
rect 7877 7289 7927 7314
rect 7877 7263 7883 7289
rect 7909 7263 7927 7289
rect 7877 7237 7927 7263
rect 8085 7285 8135 7314
rect 8085 7261 8099 7285
rect 8123 7261 8135 7285
rect 8085 7237 8135 7261
rect 8293 7290 8343 7314
rect 8293 7266 8308 7290
rect 8332 7266 8343 7290
rect 8293 7237 8343 7266
rect 8506 7285 8556 7314
rect 8506 7265 8523 7285
rect 8543 7265 8556 7285
rect 8506 7237 8556 7265
rect 1431 7135 1481 7163
rect 1431 7115 1444 7135
rect 1464 7115 1481 7135
rect 1431 7086 1481 7115
rect 1644 7134 1694 7163
rect 1644 7110 1655 7134
rect 1679 7110 1694 7134
rect 1644 7086 1694 7110
rect 1852 7139 1902 7163
rect 1852 7115 1864 7139
rect 1888 7115 1902 7139
rect 1852 7086 1902 7115
rect 2060 7137 2110 7163
rect 2060 7111 2078 7137
rect 2104 7111 2110 7137
rect 2060 7086 2110 7111
rect 6487 7176 6537 7204
rect 6487 7156 6500 7176
rect 6520 7156 6537 7176
rect 6487 7127 6537 7156
rect 6700 7175 6750 7204
rect 6700 7151 6711 7175
rect 6735 7151 6750 7175
rect 6700 7127 6750 7151
rect 6908 7180 6958 7204
rect 6908 7156 6920 7180
rect 6944 7156 6958 7180
rect 6908 7127 6958 7156
rect 7116 7178 7166 7204
rect 7116 7152 7134 7178
rect 7160 7152 7166 7178
rect 7116 7127 7166 7152
rect 2821 7083 2871 7096
rect 3029 7083 3079 7096
rect 3237 7083 3287 7096
rect 3450 7083 3500 7096
rect 1431 7028 1481 7044
rect 1644 7028 1694 7044
rect 1852 7028 1902 7044
rect 2060 7028 2110 7044
rect 3870 7046 3920 7062
rect 4078 7046 4128 7062
rect 4286 7046 4336 7062
rect 4499 7046 4549 7062
rect 7877 7124 7927 7137
rect 8085 7124 8135 7137
rect 8293 7124 8343 7137
rect 8506 7124 8556 7137
rect 6487 7069 6537 7085
rect 6700 7069 6750 7085
rect 6908 7069 6958 7085
rect 7116 7069 7166 7085
rect 8926 7087 8976 7103
rect 9134 7087 9184 7103
rect 9342 7087 9392 7103
rect 9555 7087 9605 7103
rect 5439 7024 5489 7037
rect 5652 7024 5702 7037
rect 5860 7024 5910 7037
rect 6068 7024 6118 7037
rect 383 6983 433 6996
rect 596 6983 646 6996
rect 804 6983 854 6996
rect 1012 6983 1062 6996
rect 3870 6979 3920 7004
rect 3870 6953 3876 6979
rect 3902 6953 3920 6979
rect 3870 6927 3920 6953
rect 4078 6975 4128 7004
rect 4078 6951 4092 6975
rect 4116 6951 4128 6975
rect 4078 6927 4128 6951
rect 4286 6980 4336 7004
rect 4286 6956 4301 6980
rect 4325 6956 4336 6980
rect 4286 6927 4336 6956
rect 4499 6975 4549 7004
rect 4499 6955 4516 6975
rect 4536 6955 4549 6975
rect 4499 6927 4549 6955
rect 383 6855 433 6883
rect 383 6835 396 6855
rect 416 6835 433 6855
rect 383 6806 433 6835
rect 596 6854 646 6883
rect 596 6830 607 6854
rect 631 6830 646 6854
rect 596 6806 646 6830
rect 804 6859 854 6883
rect 804 6835 816 6859
rect 840 6835 854 6859
rect 804 6806 854 6835
rect 1012 6857 1062 6883
rect 1012 6831 1030 6857
rect 1056 6831 1062 6857
rect 1012 6806 1062 6831
rect 8926 7020 8976 7045
rect 8926 6994 8932 7020
rect 8958 6994 8976 7020
rect 8926 6968 8976 6994
rect 9134 7016 9184 7045
rect 9134 6992 9148 7016
rect 9172 6992 9184 7016
rect 9134 6968 9184 6992
rect 9342 7021 9392 7045
rect 9342 6997 9357 7021
rect 9381 6997 9392 7021
rect 9342 6968 9392 6997
rect 9555 7016 9605 7045
rect 9555 6996 9572 7016
rect 9592 6996 9605 7016
rect 9555 6968 9605 6996
rect 5439 6896 5489 6924
rect 5439 6876 5452 6896
rect 5472 6876 5489 6896
rect 3870 6814 3920 6827
rect 4078 6814 4128 6827
rect 4286 6814 4336 6827
rect 4499 6814 4549 6827
rect 5439 6847 5489 6876
rect 5652 6895 5702 6924
rect 5652 6871 5663 6895
rect 5687 6871 5702 6895
rect 5652 6847 5702 6871
rect 5860 6900 5910 6924
rect 5860 6876 5872 6900
rect 5896 6876 5910 6900
rect 5860 6847 5910 6876
rect 6068 6898 6118 6924
rect 6068 6872 6086 6898
rect 6112 6872 6118 6898
rect 6068 6847 6118 6872
rect 8926 6855 8976 6868
rect 9134 6855 9184 6868
rect 9342 6855 9392 6868
rect 9555 6855 9605 6868
rect 5439 6789 5489 6805
rect 5652 6789 5702 6805
rect 5860 6789 5910 6805
rect 6068 6789 6118 6805
rect 383 6748 433 6764
rect 596 6748 646 6764
rect 804 6748 854 6764
rect 1012 6748 1062 6764
rect 6377 6780 6427 6793
rect 6590 6780 6640 6793
rect 6798 6780 6848 6793
rect 7006 6780 7056 6793
rect 1321 6739 1371 6752
rect 1534 6739 1584 6752
rect 1742 6739 1792 6752
rect 1950 6739 2000 6752
rect 2931 6736 2981 6752
rect 3139 6736 3189 6752
rect 3347 6736 3397 6752
rect 3560 6736 3610 6752
rect 2931 6669 2981 6694
rect 2931 6643 2937 6669
rect 2963 6643 2981 6669
rect 1321 6611 1371 6639
rect 1321 6591 1334 6611
rect 1354 6591 1371 6611
rect 1321 6562 1371 6591
rect 1534 6610 1584 6639
rect 1534 6586 1545 6610
rect 1569 6586 1584 6610
rect 1534 6562 1584 6586
rect 1742 6615 1792 6639
rect 1742 6591 1754 6615
rect 1778 6591 1792 6615
rect 1742 6562 1792 6591
rect 1950 6613 2000 6639
rect 2931 6617 2981 6643
rect 3139 6665 3189 6694
rect 3139 6641 3153 6665
rect 3177 6641 3189 6665
rect 3139 6617 3189 6641
rect 3347 6670 3397 6694
rect 3347 6646 3362 6670
rect 3386 6646 3397 6670
rect 3347 6617 3397 6646
rect 3560 6665 3610 6694
rect 3560 6645 3577 6665
rect 3597 6645 3610 6665
rect 3560 6617 3610 6645
rect 1950 6587 1968 6613
rect 1994 6587 2000 6613
rect 1950 6562 2000 6587
rect 1321 6504 1371 6520
rect 1534 6504 1584 6520
rect 1742 6504 1792 6520
rect 1950 6504 2000 6520
rect 7987 6777 8037 6793
rect 8195 6777 8245 6793
rect 8403 6777 8453 6793
rect 8616 6777 8666 6793
rect 7987 6710 8037 6735
rect 7987 6684 7993 6710
rect 8019 6684 8037 6710
rect 6377 6652 6427 6680
rect 6377 6632 6390 6652
rect 6410 6632 6427 6652
rect 6377 6603 6427 6632
rect 6590 6651 6640 6680
rect 6590 6627 6601 6651
rect 6625 6627 6640 6651
rect 6590 6603 6640 6627
rect 6798 6656 6848 6680
rect 6798 6632 6810 6656
rect 6834 6632 6848 6656
rect 6798 6603 6848 6632
rect 7006 6654 7056 6680
rect 7987 6658 8037 6684
rect 8195 6706 8245 6735
rect 8195 6682 8209 6706
rect 8233 6682 8245 6706
rect 8195 6658 8245 6682
rect 8403 6711 8453 6735
rect 8403 6687 8418 6711
rect 8442 6687 8453 6711
rect 8403 6658 8453 6687
rect 8616 6706 8666 6735
rect 8616 6686 8633 6706
rect 8653 6686 8666 6706
rect 8616 6658 8666 6686
rect 7006 6628 7024 6654
rect 7050 6628 7056 6654
rect 7006 6603 7056 6628
rect 6377 6545 6427 6561
rect 6590 6545 6640 6561
rect 6798 6545 6848 6561
rect 7006 6545 7056 6561
rect 7987 6545 8037 6558
rect 8195 6545 8245 6558
rect 8403 6545 8453 6558
rect 8616 6545 8666 6558
rect 2931 6504 2981 6517
rect 3139 6504 3189 6517
rect 3347 6504 3397 6517
rect 3560 6504 3610 6517
rect 8925 6533 8975 6549
rect 9133 6533 9183 6549
rect 9341 6533 9391 6549
rect 9554 6533 9604 6549
rect 3869 6492 3919 6508
rect 4077 6492 4127 6508
rect 4285 6492 4335 6508
rect 4498 6492 4548 6508
rect 382 6429 432 6442
rect 595 6429 645 6442
rect 803 6429 853 6442
rect 1011 6429 1061 6442
rect 3869 6425 3919 6450
rect 3869 6399 3875 6425
rect 3901 6399 3919 6425
rect 3869 6373 3919 6399
rect 4077 6421 4127 6450
rect 4077 6397 4091 6421
rect 4115 6397 4127 6421
rect 4077 6373 4127 6397
rect 4285 6426 4335 6450
rect 4285 6402 4300 6426
rect 4324 6402 4335 6426
rect 4285 6373 4335 6402
rect 4498 6421 4548 6450
rect 5438 6470 5488 6483
rect 5651 6470 5701 6483
rect 5859 6470 5909 6483
rect 6067 6470 6117 6483
rect 4498 6401 4515 6421
rect 4535 6401 4548 6421
rect 4498 6373 4548 6401
rect 382 6301 432 6329
rect 382 6281 395 6301
rect 415 6281 432 6301
rect 382 6252 432 6281
rect 595 6300 645 6329
rect 595 6276 606 6300
rect 630 6276 645 6300
rect 595 6252 645 6276
rect 803 6305 853 6329
rect 803 6281 815 6305
rect 839 6281 853 6305
rect 803 6252 853 6281
rect 1011 6303 1061 6329
rect 1011 6277 1029 6303
rect 1055 6277 1061 6303
rect 1011 6252 1061 6277
rect 8925 6466 8975 6491
rect 8925 6440 8931 6466
rect 8957 6440 8975 6466
rect 8925 6414 8975 6440
rect 9133 6462 9183 6491
rect 9133 6438 9147 6462
rect 9171 6438 9183 6462
rect 9133 6414 9183 6438
rect 9341 6467 9391 6491
rect 9341 6443 9356 6467
rect 9380 6443 9391 6467
rect 9341 6414 9391 6443
rect 9554 6462 9604 6491
rect 9554 6442 9571 6462
rect 9591 6442 9604 6462
rect 9554 6414 9604 6442
rect 5438 6342 5488 6370
rect 5438 6322 5451 6342
rect 5471 6322 5488 6342
rect 5438 6293 5488 6322
rect 5651 6341 5701 6370
rect 5651 6317 5662 6341
rect 5686 6317 5701 6341
rect 5651 6293 5701 6317
rect 5859 6346 5909 6370
rect 5859 6322 5871 6346
rect 5895 6322 5909 6346
rect 5859 6293 5909 6322
rect 6067 6344 6117 6370
rect 6067 6318 6085 6344
rect 6111 6318 6117 6344
rect 6067 6293 6117 6318
rect 8925 6301 8975 6314
rect 9133 6301 9183 6314
rect 9341 6301 9391 6314
rect 9554 6301 9604 6314
rect 3869 6260 3919 6273
rect 4077 6260 4127 6273
rect 4285 6260 4335 6273
rect 4498 6260 4548 6273
rect 2791 6225 2841 6241
rect 2999 6225 3049 6241
rect 3207 6225 3257 6241
rect 3420 6225 3470 6241
rect 382 6194 432 6210
rect 595 6194 645 6210
rect 803 6194 853 6210
rect 1011 6194 1061 6210
rect 7847 6266 7897 6282
rect 8055 6266 8105 6282
rect 8263 6266 8313 6282
rect 8476 6266 8526 6282
rect 5438 6235 5488 6251
rect 5651 6235 5701 6251
rect 5859 6235 5909 6251
rect 6067 6235 6117 6251
rect 1462 6147 1512 6160
rect 1675 6147 1725 6160
rect 1883 6147 1933 6160
rect 2091 6147 2141 6160
rect 2791 6158 2841 6183
rect 2791 6132 2797 6158
rect 2823 6132 2841 6158
rect 2791 6106 2841 6132
rect 2999 6154 3049 6183
rect 2999 6130 3013 6154
rect 3037 6130 3049 6154
rect 2999 6106 3049 6130
rect 3207 6159 3257 6183
rect 3207 6135 3222 6159
rect 3246 6135 3257 6159
rect 3207 6106 3257 6135
rect 3420 6154 3470 6183
rect 6518 6188 6568 6201
rect 6731 6188 6781 6201
rect 6939 6188 6989 6201
rect 7147 6188 7197 6201
rect 7847 6199 7897 6224
rect 3420 6134 3437 6154
rect 3457 6134 3470 6154
rect 3420 6106 3470 6134
rect 1462 6019 1512 6047
rect 1462 5999 1475 6019
rect 1495 5999 1512 6019
rect 1462 5970 1512 5999
rect 1675 6018 1725 6047
rect 1675 5994 1686 6018
rect 1710 5994 1725 6018
rect 1675 5970 1725 5994
rect 1883 6023 1933 6047
rect 1883 5999 1895 6023
rect 1919 5999 1933 6023
rect 1883 5970 1933 5999
rect 2091 6021 2141 6047
rect 2091 5995 2109 6021
rect 2135 5995 2141 6021
rect 7847 6173 7853 6199
rect 7879 6173 7897 6199
rect 7847 6147 7897 6173
rect 8055 6195 8105 6224
rect 8055 6171 8069 6195
rect 8093 6171 8105 6195
rect 8055 6147 8105 6171
rect 8263 6200 8313 6224
rect 8263 6176 8278 6200
rect 8302 6176 8313 6200
rect 8263 6147 8313 6176
rect 8476 6195 8526 6224
rect 8476 6175 8493 6195
rect 8513 6175 8526 6195
rect 8476 6147 8526 6175
rect 6518 6060 6568 6088
rect 6518 6040 6531 6060
rect 6551 6040 6568 6060
rect 2091 5970 2141 5995
rect 2791 5993 2841 6006
rect 2999 5993 3049 6006
rect 3207 5993 3257 6006
rect 3420 5993 3470 6006
rect 6518 6011 6568 6040
rect 6731 6059 6781 6088
rect 6731 6035 6742 6059
rect 6766 6035 6781 6059
rect 6731 6011 6781 6035
rect 6939 6064 6989 6088
rect 6939 6040 6951 6064
rect 6975 6040 6989 6064
rect 6939 6011 6989 6040
rect 7147 6062 7197 6088
rect 7147 6036 7165 6062
rect 7191 6036 7197 6062
rect 7147 6011 7197 6036
rect 7847 6034 7897 6047
rect 8055 6034 8105 6047
rect 8263 6034 8313 6047
rect 8476 6034 8526 6047
rect 3871 5943 3921 5959
rect 4079 5943 4129 5959
rect 4287 5943 4337 5959
rect 4500 5943 4550 5959
rect 1462 5912 1512 5928
rect 1675 5912 1725 5928
rect 1883 5912 1933 5928
rect 2091 5912 2141 5928
rect 8927 5984 8977 6000
rect 9135 5984 9185 6000
rect 9343 5984 9393 6000
rect 9556 5984 9606 6000
rect 6518 5953 6568 5969
rect 6731 5953 6781 5969
rect 6939 5953 6989 5969
rect 7147 5953 7197 5969
rect 5440 5921 5490 5934
rect 5653 5921 5703 5934
rect 5861 5921 5911 5934
rect 6069 5921 6119 5934
rect 384 5880 434 5893
rect 597 5880 647 5893
rect 805 5880 855 5893
rect 1013 5880 1063 5893
rect 3871 5876 3921 5901
rect 3871 5850 3877 5876
rect 3903 5850 3921 5876
rect 3871 5824 3921 5850
rect 4079 5872 4129 5901
rect 4079 5848 4093 5872
rect 4117 5848 4129 5872
rect 4079 5824 4129 5848
rect 4287 5877 4337 5901
rect 4287 5853 4302 5877
rect 4326 5853 4337 5877
rect 4287 5824 4337 5853
rect 4500 5872 4550 5901
rect 4500 5852 4517 5872
rect 4537 5852 4550 5872
rect 4500 5824 4550 5852
rect 384 5752 434 5780
rect 384 5732 397 5752
rect 417 5732 434 5752
rect 384 5703 434 5732
rect 597 5751 647 5780
rect 597 5727 608 5751
rect 632 5727 647 5751
rect 597 5703 647 5727
rect 805 5756 855 5780
rect 805 5732 817 5756
rect 841 5732 855 5756
rect 805 5703 855 5732
rect 1013 5754 1063 5780
rect 1013 5728 1031 5754
rect 1057 5728 1063 5754
rect 1013 5703 1063 5728
rect 8927 5917 8977 5942
rect 8927 5891 8933 5917
rect 8959 5891 8977 5917
rect 8927 5865 8977 5891
rect 9135 5913 9185 5942
rect 9135 5889 9149 5913
rect 9173 5889 9185 5913
rect 9135 5865 9185 5889
rect 9343 5918 9393 5942
rect 9343 5894 9358 5918
rect 9382 5894 9393 5918
rect 9343 5865 9393 5894
rect 9556 5913 9606 5942
rect 9556 5893 9573 5913
rect 9593 5893 9606 5913
rect 9556 5865 9606 5893
rect 5440 5793 5490 5821
rect 5440 5773 5453 5793
rect 5473 5773 5490 5793
rect 3871 5711 3921 5724
rect 4079 5711 4129 5724
rect 4287 5711 4337 5724
rect 4500 5711 4550 5724
rect 5440 5744 5490 5773
rect 5653 5792 5703 5821
rect 5653 5768 5664 5792
rect 5688 5768 5703 5792
rect 5653 5744 5703 5768
rect 5861 5797 5911 5821
rect 5861 5773 5873 5797
rect 5897 5773 5911 5797
rect 5861 5744 5911 5773
rect 6069 5795 6119 5821
rect 6069 5769 6087 5795
rect 6113 5769 6119 5795
rect 6069 5744 6119 5769
rect 8927 5752 8977 5765
rect 9135 5752 9185 5765
rect 9343 5752 9393 5765
rect 9556 5752 9606 5765
rect 5440 5686 5490 5702
rect 5653 5686 5703 5702
rect 5861 5686 5911 5702
rect 6069 5686 6119 5702
rect 384 5645 434 5661
rect 597 5645 647 5661
rect 805 5645 855 5661
rect 1013 5645 1063 5661
rect 6378 5677 6428 5690
rect 6591 5677 6641 5690
rect 6799 5677 6849 5690
rect 7007 5677 7057 5690
rect 1322 5636 1372 5649
rect 1535 5636 1585 5649
rect 1743 5636 1793 5649
rect 1951 5636 2001 5649
rect 2932 5633 2982 5649
rect 3140 5633 3190 5649
rect 3348 5633 3398 5649
rect 3561 5633 3611 5649
rect 2932 5566 2982 5591
rect 2932 5540 2938 5566
rect 2964 5540 2982 5566
rect 1322 5508 1372 5536
rect 1322 5488 1335 5508
rect 1355 5488 1372 5508
rect 1322 5459 1372 5488
rect 1535 5507 1585 5536
rect 1535 5483 1546 5507
rect 1570 5483 1585 5507
rect 1535 5459 1585 5483
rect 1743 5512 1793 5536
rect 1743 5488 1755 5512
rect 1779 5488 1793 5512
rect 1743 5459 1793 5488
rect 1951 5510 2001 5536
rect 2932 5514 2982 5540
rect 3140 5562 3190 5591
rect 3140 5538 3154 5562
rect 3178 5538 3190 5562
rect 3140 5514 3190 5538
rect 3348 5567 3398 5591
rect 3348 5543 3363 5567
rect 3387 5543 3398 5567
rect 3348 5514 3398 5543
rect 3561 5562 3611 5591
rect 3561 5542 3578 5562
rect 3598 5542 3611 5562
rect 3561 5514 3611 5542
rect 1951 5484 1969 5510
rect 1995 5484 2001 5510
rect 1951 5459 2001 5484
rect 1322 5401 1372 5417
rect 1535 5401 1585 5417
rect 1743 5401 1793 5417
rect 1951 5401 2001 5417
rect 7988 5674 8038 5690
rect 8196 5674 8246 5690
rect 8404 5674 8454 5690
rect 8617 5674 8667 5690
rect 7988 5607 8038 5632
rect 7988 5581 7994 5607
rect 8020 5581 8038 5607
rect 6378 5549 6428 5577
rect 6378 5529 6391 5549
rect 6411 5529 6428 5549
rect 6378 5500 6428 5529
rect 6591 5548 6641 5577
rect 6591 5524 6602 5548
rect 6626 5524 6641 5548
rect 6591 5500 6641 5524
rect 6799 5553 6849 5577
rect 6799 5529 6811 5553
rect 6835 5529 6849 5553
rect 6799 5500 6849 5529
rect 7007 5551 7057 5577
rect 7988 5555 8038 5581
rect 8196 5603 8246 5632
rect 8196 5579 8210 5603
rect 8234 5579 8246 5603
rect 8196 5555 8246 5579
rect 8404 5608 8454 5632
rect 8404 5584 8419 5608
rect 8443 5584 8454 5608
rect 8404 5555 8454 5584
rect 8617 5603 8667 5632
rect 8617 5583 8634 5603
rect 8654 5583 8667 5603
rect 8617 5555 8667 5583
rect 7007 5525 7025 5551
rect 7051 5525 7057 5551
rect 7007 5500 7057 5525
rect 6378 5442 6428 5458
rect 6591 5442 6641 5458
rect 6799 5442 6849 5458
rect 7007 5442 7057 5458
rect 7988 5442 8038 5455
rect 8196 5442 8246 5455
rect 8404 5442 8454 5455
rect 8617 5442 8667 5455
rect 2932 5401 2982 5414
rect 3140 5401 3190 5414
rect 3348 5401 3398 5414
rect 3561 5401 3611 5414
rect 8926 5430 8976 5446
rect 9134 5430 9184 5446
rect 9342 5430 9392 5446
rect 9555 5430 9605 5446
rect 3870 5389 3920 5405
rect 4078 5389 4128 5405
rect 4286 5389 4336 5405
rect 4499 5389 4549 5405
rect 383 5326 433 5339
rect 596 5326 646 5339
rect 804 5326 854 5339
rect 1012 5326 1062 5339
rect 3870 5322 3920 5347
rect 3870 5296 3876 5322
rect 3902 5296 3920 5322
rect 3870 5270 3920 5296
rect 4078 5318 4128 5347
rect 4078 5294 4092 5318
rect 4116 5294 4128 5318
rect 4078 5270 4128 5294
rect 4286 5323 4336 5347
rect 4286 5299 4301 5323
rect 4325 5299 4336 5323
rect 4286 5270 4336 5299
rect 4499 5318 4549 5347
rect 5439 5367 5489 5380
rect 5652 5367 5702 5380
rect 5860 5367 5910 5380
rect 6068 5367 6118 5380
rect 4499 5298 4516 5318
rect 4536 5298 4549 5318
rect 4499 5270 4549 5298
rect 383 5198 433 5226
rect 383 5178 396 5198
rect 416 5178 433 5198
rect 383 5149 433 5178
rect 596 5197 646 5226
rect 596 5173 607 5197
rect 631 5173 646 5197
rect 596 5149 646 5173
rect 804 5202 854 5226
rect 804 5178 816 5202
rect 840 5178 854 5202
rect 804 5149 854 5178
rect 1012 5200 1062 5226
rect 1012 5174 1030 5200
rect 1056 5174 1062 5200
rect 1012 5149 1062 5174
rect 8926 5363 8976 5388
rect 8926 5337 8932 5363
rect 8958 5337 8976 5363
rect 8926 5311 8976 5337
rect 9134 5359 9184 5388
rect 9134 5335 9148 5359
rect 9172 5335 9184 5359
rect 9134 5311 9184 5335
rect 9342 5364 9392 5388
rect 9342 5340 9357 5364
rect 9381 5340 9392 5364
rect 9342 5311 9392 5340
rect 9555 5359 9605 5388
rect 9555 5339 9572 5359
rect 9592 5339 9605 5359
rect 9555 5311 9605 5339
rect 5439 5239 5489 5267
rect 5439 5219 5452 5239
rect 5472 5219 5489 5239
rect 5439 5190 5489 5219
rect 5652 5238 5702 5267
rect 5652 5214 5663 5238
rect 5687 5214 5702 5238
rect 5652 5190 5702 5214
rect 5860 5243 5910 5267
rect 5860 5219 5872 5243
rect 5896 5219 5910 5243
rect 5860 5190 5910 5219
rect 6068 5241 6118 5267
rect 6068 5215 6086 5241
rect 6112 5215 6118 5241
rect 6068 5190 6118 5215
rect 3870 5157 3920 5170
rect 4078 5157 4128 5170
rect 4286 5157 4336 5170
rect 4499 5157 4549 5170
rect 383 5091 433 5107
rect 596 5091 646 5107
rect 804 5091 854 5107
rect 1012 5091 1062 5107
rect 2823 5103 2873 5119
rect 3031 5103 3081 5119
rect 3239 5103 3289 5119
rect 3452 5103 3502 5119
rect 1431 5063 1481 5076
rect 1644 5063 1694 5076
rect 1852 5063 1902 5076
rect 2060 5063 2110 5076
rect 8926 5198 8976 5211
rect 9134 5198 9184 5211
rect 9342 5198 9392 5211
rect 9555 5198 9605 5211
rect 5439 5132 5489 5148
rect 5652 5132 5702 5148
rect 5860 5132 5910 5148
rect 6068 5132 6118 5148
rect 7879 5144 7929 5160
rect 8087 5144 8137 5160
rect 8295 5144 8345 5160
rect 8508 5144 8558 5160
rect 6487 5104 6537 5117
rect 6700 5104 6750 5117
rect 6908 5104 6958 5117
rect 7116 5104 7166 5117
rect 2823 5036 2873 5061
rect 2823 5010 2829 5036
rect 2855 5010 2873 5036
rect 2823 4984 2873 5010
rect 3031 5032 3081 5061
rect 3031 5008 3045 5032
rect 3069 5008 3081 5032
rect 3031 4984 3081 5008
rect 3239 5037 3289 5061
rect 3239 5013 3254 5037
rect 3278 5013 3289 5037
rect 3239 4984 3289 5013
rect 3452 5032 3502 5061
rect 3452 5012 3469 5032
rect 3489 5012 3502 5032
rect 3452 4984 3502 5012
rect 7879 5077 7929 5102
rect 7879 5051 7885 5077
rect 7911 5051 7929 5077
rect 7879 5025 7929 5051
rect 8087 5073 8137 5102
rect 8087 5049 8101 5073
rect 8125 5049 8137 5073
rect 8087 5025 8137 5049
rect 8295 5078 8345 5102
rect 8295 5054 8310 5078
rect 8334 5054 8345 5078
rect 8295 5025 8345 5054
rect 8508 5073 8558 5102
rect 8508 5053 8525 5073
rect 8545 5053 8558 5073
rect 8508 5025 8558 5053
rect 1431 4935 1481 4963
rect 1431 4915 1444 4935
rect 1464 4915 1481 4935
rect 1431 4886 1481 4915
rect 1644 4934 1694 4963
rect 1644 4910 1655 4934
rect 1679 4910 1694 4934
rect 1644 4886 1694 4910
rect 1852 4939 1902 4963
rect 1852 4915 1864 4939
rect 1888 4915 1902 4939
rect 1852 4886 1902 4915
rect 2060 4937 2110 4963
rect 2060 4911 2078 4937
rect 2104 4911 2110 4937
rect 2060 4886 2110 4911
rect 6487 4976 6537 5004
rect 6487 4956 6500 4976
rect 6520 4956 6537 4976
rect 6487 4927 6537 4956
rect 6700 4975 6750 5004
rect 6700 4951 6711 4975
rect 6735 4951 6750 4975
rect 6700 4927 6750 4951
rect 6908 4980 6958 5004
rect 6908 4956 6920 4980
rect 6944 4956 6958 4980
rect 6908 4927 6958 4956
rect 7116 4978 7166 5004
rect 7116 4952 7134 4978
rect 7160 4952 7166 4978
rect 7116 4927 7166 4952
rect 2823 4871 2873 4884
rect 3031 4871 3081 4884
rect 3239 4871 3289 4884
rect 3452 4871 3502 4884
rect 1431 4828 1481 4844
rect 1644 4828 1694 4844
rect 1852 4828 1902 4844
rect 2060 4828 2110 4844
rect 3871 4840 3921 4856
rect 4079 4840 4129 4856
rect 4287 4840 4337 4856
rect 4500 4840 4550 4856
rect 384 4777 434 4790
rect 597 4777 647 4790
rect 805 4777 855 4790
rect 1013 4777 1063 4790
rect 7879 4912 7929 4925
rect 8087 4912 8137 4925
rect 8295 4912 8345 4925
rect 8508 4912 8558 4925
rect 6487 4869 6537 4885
rect 6700 4869 6750 4885
rect 6908 4869 6958 4885
rect 7116 4869 7166 4885
rect 8927 4881 8977 4897
rect 9135 4881 9185 4897
rect 9343 4881 9393 4897
rect 9556 4881 9606 4897
rect 5440 4818 5490 4831
rect 5653 4818 5703 4831
rect 5861 4818 5911 4831
rect 6069 4818 6119 4831
rect 3871 4773 3921 4798
rect 3871 4747 3877 4773
rect 3903 4747 3921 4773
rect 3871 4721 3921 4747
rect 4079 4769 4129 4798
rect 4079 4745 4093 4769
rect 4117 4745 4129 4769
rect 4079 4721 4129 4745
rect 4287 4774 4337 4798
rect 4287 4750 4302 4774
rect 4326 4750 4337 4774
rect 4287 4721 4337 4750
rect 4500 4769 4550 4798
rect 4500 4749 4517 4769
rect 4537 4749 4550 4769
rect 4500 4721 4550 4749
rect 384 4649 434 4677
rect 384 4629 397 4649
rect 417 4629 434 4649
rect 384 4600 434 4629
rect 597 4648 647 4677
rect 597 4624 608 4648
rect 632 4624 647 4648
rect 597 4600 647 4624
rect 805 4653 855 4677
rect 805 4629 817 4653
rect 841 4629 855 4653
rect 805 4600 855 4629
rect 1013 4651 1063 4677
rect 1013 4625 1031 4651
rect 1057 4625 1063 4651
rect 1013 4600 1063 4625
rect 8927 4814 8977 4839
rect 8927 4788 8933 4814
rect 8959 4788 8977 4814
rect 8927 4762 8977 4788
rect 9135 4810 9185 4839
rect 9135 4786 9149 4810
rect 9173 4786 9185 4810
rect 9135 4762 9185 4786
rect 9343 4815 9393 4839
rect 9343 4791 9358 4815
rect 9382 4791 9393 4815
rect 9343 4762 9393 4791
rect 9556 4810 9606 4839
rect 9556 4790 9573 4810
rect 9593 4790 9606 4810
rect 9556 4762 9606 4790
rect 5440 4690 5490 4718
rect 5440 4670 5453 4690
rect 5473 4670 5490 4690
rect 3871 4608 3921 4621
rect 4079 4608 4129 4621
rect 4287 4608 4337 4621
rect 4500 4608 4550 4621
rect 5440 4641 5490 4670
rect 5653 4689 5703 4718
rect 5653 4665 5664 4689
rect 5688 4665 5703 4689
rect 5653 4641 5703 4665
rect 5861 4694 5911 4718
rect 5861 4670 5873 4694
rect 5897 4670 5911 4694
rect 5861 4641 5911 4670
rect 6069 4692 6119 4718
rect 6069 4666 6087 4692
rect 6113 4666 6119 4692
rect 6069 4641 6119 4666
rect 8927 4649 8977 4662
rect 9135 4649 9185 4662
rect 9343 4649 9393 4662
rect 9556 4649 9606 4662
rect 5440 4583 5490 4599
rect 5653 4583 5703 4599
rect 5861 4583 5911 4599
rect 6069 4583 6119 4599
rect 384 4542 434 4558
rect 597 4542 647 4558
rect 805 4542 855 4558
rect 1013 4542 1063 4558
rect 6378 4574 6428 4587
rect 6591 4574 6641 4587
rect 6799 4574 6849 4587
rect 7007 4574 7057 4587
rect 1322 4533 1372 4546
rect 1535 4533 1585 4546
rect 1743 4533 1793 4546
rect 1951 4533 2001 4546
rect 2932 4530 2982 4546
rect 3140 4530 3190 4546
rect 3348 4530 3398 4546
rect 3561 4530 3611 4546
rect 2932 4463 2982 4488
rect 2932 4437 2938 4463
rect 2964 4437 2982 4463
rect 1322 4405 1372 4433
rect 1322 4385 1335 4405
rect 1355 4385 1372 4405
rect 1322 4356 1372 4385
rect 1535 4404 1585 4433
rect 1535 4380 1546 4404
rect 1570 4380 1585 4404
rect 1535 4356 1585 4380
rect 1743 4409 1793 4433
rect 1743 4385 1755 4409
rect 1779 4385 1793 4409
rect 1743 4356 1793 4385
rect 1951 4407 2001 4433
rect 2932 4411 2982 4437
rect 3140 4459 3190 4488
rect 3140 4435 3154 4459
rect 3178 4435 3190 4459
rect 3140 4411 3190 4435
rect 3348 4464 3398 4488
rect 3348 4440 3363 4464
rect 3387 4440 3398 4464
rect 3348 4411 3398 4440
rect 3561 4459 3611 4488
rect 3561 4439 3578 4459
rect 3598 4439 3611 4459
rect 3561 4411 3611 4439
rect 1951 4381 1969 4407
rect 1995 4381 2001 4407
rect 1951 4356 2001 4381
rect 1322 4298 1372 4314
rect 1535 4298 1585 4314
rect 1743 4298 1793 4314
rect 1951 4298 2001 4314
rect 7988 4571 8038 4587
rect 8196 4571 8246 4587
rect 8404 4571 8454 4587
rect 8617 4571 8667 4587
rect 7988 4504 8038 4529
rect 7988 4478 7994 4504
rect 8020 4478 8038 4504
rect 6378 4446 6428 4474
rect 6378 4426 6391 4446
rect 6411 4426 6428 4446
rect 6378 4397 6428 4426
rect 6591 4445 6641 4474
rect 6591 4421 6602 4445
rect 6626 4421 6641 4445
rect 6591 4397 6641 4421
rect 6799 4450 6849 4474
rect 6799 4426 6811 4450
rect 6835 4426 6849 4450
rect 6799 4397 6849 4426
rect 7007 4448 7057 4474
rect 7988 4452 8038 4478
rect 8196 4500 8246 4529
rect 8196 4476 8210 4500
rect 8234 4476 8246 4500
rect 8196 4452 8246 4476
rect 8404 4505 8454 4529
rect 8404 4481 8419 4505
rect 8443 4481 8454 4505
rect 8404 4452 8454 4481
rect 8617 4500 8667 4529
rect 8617 4480 8634 4500
rect 8654 4480 8667 4500
rect 8617 4452 8667 4480
rect 7007 4422 7025 4448
rect 7051 4422 7057 4448
rect 7007 4397 7057 4422
rect 6378 4339 6428 4355
rect 6591 4339 6641 4355
rect 6799 4339 6849 4355
rect 7007 4339 7057 4355
rect 7988 4339 8038 4352
rect 8196 4339 8246 4352
rect 8404 4339 8454 4352
rect 8617 4339 8667 4352
rect 2932 4298 2982 4311
rect 3140 4298 3190 4311
rect 3348 4298 3398 4311
rect 3561 4298 3611 4311
rect 8926 4327 8976 4343
rect 9134 4327 9184 4343
rect 9342 4327 9392 4343
rect 9555 4327 9605 4343
rect 3870 4286 3920 4302
rect 4078 4286 4128 4302
rect 4286 4286 4336 4302
rect 4499 4286 4549 4302
rect 383 4223 433 4236
rect 596 4223 646 4236
rect 804 4223 854 4236
rect 1012 4223 1062 4236
rect 3870 4219 3920 4244
rect 3870 4193 3876 4219
rect 3902 4193 3920 4219
rect 3870 4167 3920 4193
rect 4078 4215 4128 4244
rect 4078 4191 4092 4215
rect 4116 4191 4128 4215
rect 4078 4167 4128 4191
rect 4286 4220 4336 4244
rect 4286 4196 4301 4220
rect 4325 4196 4336 4220
rect 4286 4167 4336 4196
rect 4499 4215 4549 4244
rect 5439 4264 5489 4277
rect 5652 4264 5702 4277
rect 5860 4264 5910 4277
rect 6068 4264 6118 4277
rect 4499 4195 4516 4215
rect 4536 4195 4549 4215
rect 4499 4167 4549 4195
rect 383 4095 433 4123
rect 383 4075 396 4095
rect 416 4075 433 4095
rect 383 4046 433 4075
rect 596 4094 646 4123
rect 596 4070 607 4094
rect 631 4070 646 4094
rect 596 4046 646 4070
rect 804 4099 854 4123
rect 804 4075 816 4099
rect 840 4075 854 4099
rect 804 4046 854 4075
rect 1012 4097 1062 4123
rect 1012 4071 1030 4097
rect 1056 4071 1062 4097
rect 1012 4046 1062 4071
rect 8926 4260 8976 4285
rect 8926 4234 8932 4260
rect 8958 4234 8976 4260
rect 8926 4208 8976 4234
rect 9134 4256 9184 4285
rect 9134 4232 9148 4256
rect 9172 4232 9184 4256
rect 9134 4208 9184 4232
rect 9342 4261 9392 4285
rect 9342 4237 9357 4261
rect 9381 4237 9392 4261
rect 9342 4208 9392 4237
rect 9555 4256 9605 4285
rect 9555 4236 9572 4256
rect 9592 4236 9605 4256
rect 9555 4208 9605 4236
rect 5439 4136 5489 4164
rect 5439 4116 5452 4136
rect 5472 4116 5489 4136
rect 5439 4087 5489 4116
rect 5652 4135 5702 4164
rect 5652 4111 5663 4135
rect 5687 4111 5702 4135
rect 5652 4087 5702 4111
rect 5860 4140 5910 4164
rect 5860 4116 5872 4140
rect 5896 4116 5910 4140
rect 5860 4087 5910 4116
rect 6068 4138 6118 4164
rect 6068 4112 6086 4138
rect 6112 4112 6118 4138
rect 6068 4087 6118 4112
rect 8926 4095 8976 4108
rect 9134 4095 9184 4108
rect 9342 4095 9392 4108
rect 9555 4095 9605 4108
rect 3870 4054 3920 4067
rect 4078 4054 4128 4067
rect 4286 4054 4336 4067
rect 4499 4054 4549 4067
rect 2792 4019 2842 4035
rect 3000 4019 3050 4035
rect 3208 4019 3258 4035
rect 3421 4019 3471 4035
rect 383 3988 433 4004
rect 596 3988 646 4004
rect 804 3988 854 4004
rect 1012 3988 1062 4004
rect 7848 4060 7898 4076
rect 8056 4060 8106 4076
rect 8264 4060 8314 4076
rect 8477 4060 8527 4076
rect 5439 4029 5489 4045
rect 5652 4029 5702 4045
rect 5860 4029 5910 4045
rect 6068 4029 6118 4045
rect 1463 3941 1513 3954
rect 1676 3941 1726 3954
rect 1884 3941 1934 3954
rect 2092 3941 2142 3954
rect 2792 3952 2842 3977
rect 2792 3926 2798 3952
rect 2824 3926 2842 3952
rect 2792 3900 2842 3926
rect 3000 3948 3050 3977
rect 3000 3924 3014 3948
rect 3038 3924 3050 3948
rect 3000 3900 3050 3924
rect 3208 3953 3258 3977
rect 3208 3929 3223 3953
rect 3247 3929 3258 3953
rect 3208 3900 3258 3929
rect 3421 3948 3471 3977
rect 6519 3982 6569 3995
rect 6732 3982 6782 3995
rect 6940 3982 6990 3995
rect 7148 3982 7198 3995
rect 7848 3993 7898 4018
rect 3421 3928 3438 3948
rect 3458 3928 3471 3948
rect 3421 3900 3471 3928
rect 1463 3813 1513 3841
rect 1463 3793 1476 3813
rect 1496 3793 1513 3813
rect 1463 3764 1513 3793
rect 1676 3812 1726 3841
rect 1676 3788 1687 3812
rect 1711 3788 1726 3812
rect 1676 3764 1726 3788
rect 1884 3817 1934 3841
rect 1884 3793 1896 3817
rect 1920 3793 1934 3817
rect 1884 3764 1934 3793
rect 2092 3815 2142 3841
rect 2092 3789 2110 3815
rect 2136 3789 2142 3815
rect 7848 3967 7854 3993
rect 7880 3967 7898 3993
rect 7848 3941 7898 3967
rect 8056 3989 8106 4018
rect 8056 3965 8070 3989
rect 8094 3965 8106 3989
rect 8056 3941 8106 3965
rect 8264 3994 8314 4018
rect 8264 3970 8279 3994
rect 8303 3970 8314 3994
rect 8264 3941 8314 3970
rect 8477 3989 8527 4018
rect 8477 3969 8494 3989
rect 8514 3969 8527 3989
rect 8477 3941 8527 3969
rect 6519 3854 6569 3882
rect 6519 3834 6532 3854
rect 6552 3834 6569 3854
rect 2092 3764 2142 3789
rect 2792 3787 2842 3800
rect 3000 3787 3050 3800
rect 3208 3787 3258 3800
rect 3421 3787 3471 3800
rect 6519 3805 6569 3834
rect 6732 3853 6782 3882
rect 6732 3829 6743 3853
rect 6767 3829 6782 3853
rect 6732 3805 6782 3829
rect 6940 3858 6990 3882
rect 6940 3834 6952 3858
rect 6976 3834 6990 3858
rect 6940 3805 6990 3834
rect 7148 3856 7198 3882
rect 7148 3830 7166 3856
rect 7192 3830 7198 3856
rect 7148 3805 7198 3830
rect 7848 3828 7898 3841
rect 8056 3828 8106 3841
rect 8264 3828 8314 3841
rect 8477 3828 8527 3841
rect 3872 3737 3922 3753
rect 4080 3737 4130 3753
rect 4288 3737 4338 3753
rect 4501 3737 4551 3753
rect 1463 3706 1513 3722
rect 1676 3706 1726 3722
rect 1884 3706 1934 3722
rect 2092 3706 2142 3722
rect 8928 3778 8978 3794
rect 9136 3778 9186 3794
rect 9344 3778 9394 3794
rect 9557 3778 9607 3794
rect 6519 3747 6569 3763
rect 6732 3747 6782 3763
rect 6940 3747 6990 3763
rect 7148 3747 7198 3763
rect 5441 3715 5491 3728
rect 5654 3715 5704 3728
rect 5862 3715 5912 3728
rect 6070 3715 6120 3728
rect 385 3674 435 3687
rect 598 3674 648 3687
rect 806 3674 856 3687
rect 1014 3674 1064 3687
rect 3872 3670 3922 3695
rect 3872 3644 3878 3670
rect 3904 3644 3922 3670
rect 3872 3618 3922 3644
rect 4080 3666 4130 3695
rect 4080 3642 4094 3666
rect 4118 3642 4130 3666
rect 4080 3618 4130 3642
rect 4288 3671 4338 3695
rect 4288 3647 4303 3671
rect 4327 3647 4338 3671
rect 4288 3618 4338 3647
rect 4501 3666 4551 3695
rect 4501 3646 4518 3666
rect 4538 3646 4551 3666
rect 4501 3618 4551 3646
rect 385 3546 435 3574
rect 385 3526 398 3546
rect 418 3526 435 3546
rect 385 3497 435 3526
rect 598 3545 648 3574
rect 598 3521 609 3545
rect 633 3521 648 3545
rect 598 3497 648 3521
rect 806 3550 856 3574
rect 806 3526 818 3550
rect 842 3526 856 3550
rect 806 3497 856 3526
rect 1014 3548 1064 3574
rect 1014 3522 1032 3548
rect 1058 3522 1064 3548
rect 1014 3497 1064 3522
rect 8928 3711 8978 3736
rect 8928 3685 8934 3711
rect 8960 3685 8978 3711
rect 8928 3659 8978 3685
rect 9136 3707 9186 3736
rect 9136 3683 9150 3707
rect 9174 3683 9186 3707
rect 9136 3659 9186 3683
rect 9344 3712 9394 3736
rect 9344 3688 9359 3712
rect 9383 3688 9394 3712
rect 9344 3659 9394 3688
rect 9557 3707 9607 3736
rect 9557 3687 9574 3707
rect 9594 3687 9607 3707
rect 9557 3659 9607 3687
rect 5441 3587 5491 3615
rect 5441 3567 5454 3587
rect 5474 3567 5491 3587
rect 3872 3505 3922 3518
rect 4080 3505 4130 3518
rect 4288 3505 4338 3518
rect 4501 3505 4551 3518
rect 5441 3538 5491 3567
rect 5654 3586 5704 3615
rect 5654 3562 5665 3586
rect 5689 3562 5704 3586
rect 5654 3538 5704 3562
rect 5862 3591 5912 3615
rect 5862 3567 5874 3591
rect 5898 3567 5912 3591
rect 5862 3538 5912 3567
rect 6070 3589 6120 3615
rect 6070 3563 6088 3589
rect 6114 3563 6120 3589
rect 6070 3538 6120 3563
rect 8928 3546 8978 3559
rect 9136 3546 9186 3559
rect 9344 3546 9394 3559
rect 9557 3546 9607 3559
rect 5441 3480 5491 3496
rect 5654 3480 5704 3496
rect 5862 3480 5912 3496
rect 6070 3480 6120 3496
rect 385 3439 435 3455
rect 598 3439 648 3455
rect 806 3439 856 3455
rect 1014 3439 1064 3455
rect 6379 3471 6429 3484
rect 6592 3471 6642 3484
rect 6800 3471 6850 3484
rect 7008 3471 7058 3484
rect 1323 3430 1373 3443
rect 1536 3430 1586 3443
rect 1744 3430 1794 3443
rect 1952 3430 2002 3443
rect 2933 3427 2983 3443
rect 3141 3427 3191 3443
rect 3349 3427 3399 3443
rect 3562 3427 3612 3443
rect 2933 3360 2983 3385
rect 2933 3334 2939 3360
rect 2965 3334 2983 3360
rect 1323 3302 1373 3330
rect 1323 3282 1336 3302
rect 1356 3282 1373 3302
rect 1323 3253 1373 3282
rect 1536 3301 1586 3330
rect 1536 3277 1547 3301
rect 1571 3277 1586 3301
rect 1536 3253 1586 3277
rect 1744 3306 1794 3330
rect 1744 3282 1756 3306
rect 1780 3282 1794 3306
rect 1744 3253 1794 3282
rect 1952 3304 2002 3330
rect 2933 3308 2983 3334
rect 3141 3356 3191 3385
rect 3141 3332 3155 3356
rect 3179 3332 3191 3356
rect 3141 3308 3191 3332
rect 3349 3361 3399 3385
rect 3349 3337 3364 3361
rect 3388 3337 3399 3361
rect 3349 3308 3399 3337
rect 3562 3356 3612 3385
rect 3562 3336 3579 3356
rect 3599 3336 3612 3356
rect 3562 3308 3612 3336
rect 1952 3278 1970 3304
rect 1996 3278 2002 3304
rect 1952 3253 2002 3278
rect 1323 3195 1373 3211
rect 1536 3195 1586 3211
rect 1744 3195 1794 3211
rect 1952 3195 2002 3211
rect 7989 3468 8039 3484
rect 8197 3468 8247 3484
rect 8405 3468 8455 3484
rect 8618 3468 8668 3484
rect 7989 3401 8039 3426
rect 7989 3375 7995 3401
rect 8021 3375 8039 3401
rect 6379 3343 6429 3371
rect 6379 3323 6392 3343
rect 6412 3323 6429 3343
rect 6379 3294 6429 3323
rect 6592 3342 6642 3371
rect 6592 3318 6603 3342
rect 6627 3318 6642 3342
rect 6592 3294 6642 3318
rect 6800 3347 6850 3371
rect 6800 3323 6812 3347
rect 6836 3323 6850 3347
rect 6800 3294 6850 3323
rect 7008 3345 7058 3371
rect 7989 3349 8039 3375
rect 8197 3397 8247 3426
rect 8197 3373 8211 3397
rect 8235 3373 8247 3397
rect 8197 3349 8247 3373
rect 8405 3402 8455 3426
rect 8405 3378 8420 3402
rect 8444 3378 8455 3402
rect 8405 3349 8455 3378
rect 8618 3397 8668 3426
rect 8618 3377 8635 3397
rect 8655 3377 8668 3397
rect 8618 3349 8668 3377
rect 7008 3319 7026 3345
rect 7052 3319 7058 3345
rect 7008 3294 7058 3319
rect 6379 3236 6429 3252
rect 6592 3236 6642 3252
rect 6800 3236 6850 3252
rect 7008 3236 7058 3252
rect 7989 3236 8039 3249
rect 8197 3236 8247 3249
rect 8405 3236 8455 3249
rect 8618 3236 8668 3249
rect 2933 3195 2983 3208
rect 3141 3195 3191 3208
rect 3349 3195 3399 3208
rect 3562 3195 3612 3208
rect 8927 3224 8977 3240
rect 9135 3224 9185 3240
rect 9343 3224 9393 3240
rect 9556 3224 9606 3240
rect 3871 3183 3921 3199
rect 4079 3183 4129 3199
rect 4287 3183 4337 3199
rect 4500 3183 4550 3199
rect 384 3120 434 3133
rect 597 3120 647 3133
rect 805 3120 855 3133
rect 1013 3120 1063 3133
rect 3871 3116 3921 3141
rect 3871 3090 3877 3116
rect 3903 3090 3921 3116
rect 3871 3064 3921 3090
rect 4079 3112 4129 3141
rect 4079 3088 4093 3112
rect 4117 3088 4129 3112
rect 4079 3064 4129 3088
rect 4287 3117 4337 3141
rect 4287 3093 4302 3117
rect 4326 3093 4337 3117
rect 4287 3064 4337 3093
rect 4500 3112 4550 3141
rect 5440 3161 5490 3174
rect 5653 3161 5703 3174
rect 5861 3161 5911 3174
rect 6069 3161 6119 3174
rect 4500 3092 4517 3112
rect 4537 3092 4550 3112
rect 4500 3064 4550 3092
rect 384 2992 434 3020
rect 384 2972 397 2992
rect 417 2972 434 2992
rect 384 2943 434 2972
rect 597 2991 647 3020
rect 597 2967 608 2991
rect 632 2967 647 2991
rect 597 2943 647 2967
rect 805 2996 855 3020
rect 805 2972 817 2996
rect 841 2972 855 2996
rect 805 2943 855 2972
rect 1013 2994 1063 3020
rect 1013 2968 1031 2994
rect 1057 2968 1063 2994
rect 1013 2943 1063 2968
rect 8927 3157 8977 3182
rect 8927 3131 8933 3157
rect 8959 3131 8977 3157
rect 8927 3105 8977 3131
rect 9135 3153 9185 3182
rect 9135 3129 9149 3153
rect 9173 3129 9185 3153
rect 9135 3105 9185 3129
rect 9343 3158 9393 3182
rect 9343 3134 9358 3158
rect 9382 3134 9393 3158
rect 9343 3105 9393 3134
rect 9556 3153 9606 3182
rect 9556 3133 9573 3153
rect 9593 3133 9606 3153
rect 9556 3105 9606 3133
rect 5440 3033 5490 3061
rect 5440 3013 5453 3033
rect 5473 3013 5490 3033
rect 5440 2984 5490 3013
rect 5653 3032 5703 3061
rect 5653 3008 5664 3032
rect 5688 3008 5703 3032
rect 5653 2984 5703 3008
rect 5861 3037 5911 3061
rect 5861 3013 5873 3037
rect 5897 3013 5911 3037
rect 5861 2984 5911 3013
rect 6069 3035 6119 3061
rect 6069 3009 6087 3035
rect 6113 3009 6119 3035
rect 6069 2984 6119 3009
rect 8927 2992 8977 3005
rect 9135 2992 9185 3005
rect 9343 2992 9393 3005
rect 9556 2992 9606 3005
rect 3871 2951 3921 2964
rect 4079 2951 4129 2964
rect 4287 2951 4337 2964
rect 4500 2951 4550 2964
rect 384 2885 434 2901
rect 597 2885 647 2901
rect 805 2885 855 2901
rect 1013 2885 1063 2901
rect 2823 2903 2873 2919
rect 3031 2903 3081 2919
rect 3239 2903 3289 2919
rect 3452 2903 3502 2919
rect 1433 2851 1483 2864
rect 1646 2851 1696 2864
rect 1854 2851 1904 2864
rect 2062 2851 2112 2864
rect 5440 2926 5490 2942
rect 5653 2926 5703 2942
rect 5861 2926 5911 2942
rect 6069 2926 6119 2942
rect 7879 2944 7929 2960
rect 8087 2944 8137 2960
rect 8295 2944 8345 2960
rect 8508 2944 8558 2960
rect 6489 2892 6539 2905
rect 6702 2892 6752 2905
rect 6910 2892 6960 2905
rect 7118 2892 7168 2905
rect 2823 2836 2873 2861
rect 2823 2810 2829 2836
rect 2855 2810 2873 2836
rect 2823 2784 2873 2810
rect 3031 2832 3081 2861
rect 3031 2808 3045 2832
rect 3069 2808 3081 2832
rect 3031 2784 3081 2808
rect 3239 2837 3289 2861
rect 3239 2813 3254 2837
rect 3278 2813 3289 2837
rect 3239 2784 3289 2813
rect 3452 2832 3502 2861
rect 3452 2812 3469 2832
rect 3489 2812 3502 2832
rect 3452 2784 3502 2812
rect 7879 2877 7929 2902
rect 7879 2851 7885 2877
rect 7911 2851 7929 2877
rect 7879 2825 7929 2851
rect 8087 2873 8137 2902
rect 8087 2849 8101 2873
rect 8125 2849 8137 2873
rect 8087 2825 8137 2849
rect 8295 2878 8345 2902
rect 8295 2854 8310 2878
rect 8334 2854 8345 2878
rect 8295 2825 8345 2854
rect 8508 2873 8558 2902
rect 8508 2853 8525 2873
rect 8545 2853 8558 2873
rect 8508 2825 8558 2853
rect 1433 2723 1483 2751
rect 1433 2703 1446 2723
rect 1466 2703 1483 2723
rect 1433 2674 1483 2703
rect 1646 2722 1696 2751
rect 1646 2698 1657 2722
rect 1681 2698 1696 2722
rect 1646 2674 1696 2698
rect 1854 2727 1904 2751
rect 1854 2703 1866 2727
rect 1890 2703 1904 2727
rect 1854 2674 1904 2703
rect 2062 2725 2112 2751
rect 2062 2699 2080 2725
rect 2106 2699 2112 2725
rect 2062 2674 2112 2699
rect 6489 2764 6539 2792
rect 6489 2744 6502 2764
rect 6522 2744 6539 2764
rect 6489 2715 6539 2744
rect 6702 2763 6752 2792
rect 6702 2739 6713 2763
rect 6737 2739 6752 2763
rect 6702 2715 6752 2739
rect 6910 2768 6960 2792
rect 6910 2744 6922 2768
rect 6946 2744 6960 2768
rect 6910 2715 6960 2744
rect 7118 2766 7168 2792
rect 7118 2740 7136 2766
rect 7162 2740 7168 2766
rect 7118 2715 7168 2740
rect 2823 2671 2873 2684
rect 3031 2671 3081 2684
rect 3239 2671 3289 2684
rect 3452 2671 3502 2684
rect 1433 2616 1483 2632
rect 1646 2616 1696 2632
rect 1854 2616 1904 2632
rect 2062 2616 2112 2632
rect 3872 2634 3922 2650
rect 4080 2634 4130 2650
rect 4288 2634 4338 2650
rect 4501 2634 4551 2650
rect 7879 2712 7929 2725
rect 8087 2712 8137 2725
rect 8295 2712 8345 2725
rect 8508 2712 8558 2725
rect 6489 2657 6539 2673
rect 6702 2657 6752 2673
rect 6910 2657 6960 2673
rect 7118 2657 7168 2673
rect 8928 2675 8978 2691
rect 9136 2675 9186 2691
rect 9344 2675 9394 2691
rect 9557 2675 9607 2691
rect 5441 2612 5491 2625
rect 5654 2612 5704 2625
rect 5862 2612 5912 2625
rect 6070 2612 6120 2625
rect 385 2571 435 2584
rect 598 2571 648 2584
rect 806 2571 856 2584
rect 1014 2571 1064 2584
rect 3872 2567 3922 2592
rect 3872 2541 3878 2567
rect 3904 2541 3922 2567
rect 3872 2515 3922 2541
rect 4080 2563 4130 2592
rect 4080 2539 4094 2563
rect 4118 2539 4130 2563
rect 4080 2515 4130 2539
rect 4288 2568 4338 2592
rect 4288 2544 4303 2568
rect 4327 2544 4338 2568
rect 4288 2515 4338 2544
rect 4501 2563 4551 2592
rect 4501 2543 4518 2563
rect 4538 2543 4551 2563
rect 4501 2515 4551 2543
rect 385 2443 435 2471
rect 385 2423 398 2443
rect 418 2423 435 2443
rect 385 2394 435 2423
rect 598 2442 648 2471
rect 598 2418 609 2442
rect 633 2418 648 2442
rect 598 2394 648 2418
rect 806 2447 856 2471
rect 806 2423 818 2447
rect 842 2423 856 2447
rect 806 2394 856 2423
rect 1014 2445 1064 2471
rect 1014 2419 1032 2445
rect 1058 2419 1064 2445
rect 1014 2394 1064 2419
rect 8928 2608 8978 2633
rect 8928 2582 8934 2608
rect 8960 2582 8978 2608
rect 8928 2556 8978 2582
rect 9136 2604 9186 2633
rect 9136 2580 9150 2604
rect 9174 2580 9186 2604
rect 9136 2556 9186 2580
rect 9344 2609 9394 2633
rect 9344 2585 9359 2609
rect 9383 2585 9394 2609
rect 9344 2556 9394 2585
rect 9557 2604 9607 2633
rect 9557 2584 9574 2604
rect 9594 2584 9607 2604
rect 9557 2556 9607 2584
rect 5441 2484 5491 2512
rect 5441 2464 5454 2484
rect 5474 2464 5491 2484
rect 3872 2402 3922 2415
rect 4080 2402 4130 2415
rect 4288 2402 4338 2415
rect 4501 2402 4551 2415
rect 5441 2435 5491 2464
rect 5654 2483 5704 2512
rect 5654 2459 5665 2483
rect 5689 2459 5704 2483
rect 5654 2435 5704 2459
rect 5862 2488 5912 2512
rect 5862 2464 5874 2488
rect 5898 2464 5912 2488
rect 5862 2435 5912 2464
rect 6070 2486 6120 2512
rect 6070 2460 6088 2486
rect 6114 2460 6120 2486
rect 6070 2435 6120 2460
rect 8928 2443 8978 2456
rect 9136 2443 9186 2456
rect 9344 2443 9394 2456
rect 9557 2443 9607 2456
rect 5441 2377 5491 2393
rect 5654 2377 5704 2393
rect 5862 2377 5912 2393
rect 6070 2377 6120 2393
rect 385 2336 435 2352
rect 598 2336 648 2352
rect 806 2336 856 2352
rect 1014 2336 1064 2352
rect 6379 2368 6429 2381
rect 6592 2368 6642 2381
rect 6800 2368 6850 2381
rect 7008 2368 7058 2381
rect 1323 2327 1373 2340
rect 1536 2327 1586 2340
rect 1744 2327 1794 2340
rect 1952 2327 2002 2340
rect 2933 2324 2983 2340
rect 3141 2324 3191 2340
rect 3349 2324 3399 2340
rect 3562 2324 3612 2340
rect 2933 2257 2983 2282
rect 2933 2231 2939 2257
rect 2965 2231 2983 2257
rect 1323 2199 1373 2227
rect 1323 2179 1336 2199
rect 1356 2179 1373 2199
rect 1323 2150 1373 2179
rect 1536 2198 1586 2227
rect 1536 2174 1547 2198
rect 1571 2174 1586 2198
rect 1536 2150 1586 2174
rect 1744 2203 1794 2227
rect 1744 2179 1756 2203
rect 1780 2179 1794 2203
rect 1744 2150 1794 2179
rect 1952 2201 2002 2227
rect 2933 2205 2983 2231
rect 3141 2253 3191 2282
rect 3141 2229 3155 2253
rect 3179 2229 3191 2253
rect 3141 2205 3191 2229
rect 3349 2258 3399 2282
rect 3349 2234 3364 2258
rect 3388 2234 3399 2258
rect 3349 2205 3399 2234
rect 3562 2253 3612 2282
rect 3562 2233 3579 2253
rect 3599 2233 3612 2253
rect 3562 2205 3612 2233
rect 1952 2175 1970 2201
rect 1996 2175 2002 2201
rect 1952 2150 2002 2175
rect 1323 2092 1373 2108
rect 1536 2092 1586 2108
rect 1744 2092 1794 2108
rect 1952 2092 2002 2108
rect 7989 2365 8039 2381
rect 8197 2365 8247 2381
rect 8405 2365 8455 2381
rect 8618 2365 8668 2381
rect 7989 2298 8039 2323
rect 7989 2272 7995 2298
rect 8021 2272 8039 2298
rect 6379 2240 6429 2268
rect 6379 2220 6392 2240
rect 6412 2220 6429 2240
rect 6379 2191 6429 2220
rect 6592 2239 6642 2268
rect 6592 2215 6603 2239
rect 6627 2215 6642 2239
rect 6592 2191 6642 2215
rect 6800 2244 6850 2268
rect 6800 2220 6812 2244
rect 6836 2220 6850 2244
rect 6800 2191 6850 2220
rect 7008 2242 7058 2268
rect 7989 2246 8039 2272
rect 8197 2294 8247 2323
rect 8197 2270 8211 2294
rect 8235 2270 8247 2294
rect 8197 2246 8247 2270
rect 8405 2299 8455 2323
rect 8405 2275 8420 2299
rect 8444 2275 8455 2299
rect 8405 2246 8455 2275
rect 8618 2294 8668 2323
rect 8618 2274 8635 2294
rect 8655 2274 8668 2294
rect 8618 2246 8668 2274
rect 7008 2216 7026 2242
rect 7052 2216 7058 2242
rect 7008 2191 7058 2216
rect 6379 2133 6429 2149
rect 6592 2133 6642 2149
rect 6800 2133 6850 2149
rect 7008 2133 7058 2149
rect 7989 2133 8039 2146
rect 8197 2133 8247 2146
rect 8405 2133 8455 2146
rect 8618 2133 8668 2146
rect 2933 2092 2983 2105
rect 3141 2092 3191 2105
rect 3349 2092 3399 2105
rect 3562 2092 3612 2105
rect 8927 2121 8977 2137
rect 9135 2121 9185 2137
rect 9343 2121 9393 2137
rect 9556 2121 9606 2137
rect 3871 2080 3921 2096
rect 4079 2080 4129 2096
rect 4287 2080 4337 2096
rect 4500 2080 4550 2096
rect 384 2017 434 2030
rect 597 2017 647 2030
rect 805 2017 855 2030
rect 1013 2017 1063 2030
rect 3871 2013 3921 2038
rect 3871 1987 3877 2013
rect 3903 1987 3921 2013
rect 3871 1961 3921 1987
rect 4079 2009 4129 2038
rect 4079 1985 4093 2009
rect 4117 1985 4129 2009
rect 4079 1961 4129 1985
rect 4287 2014 4337 2038
rect 4287 1990 4302 2014
rect 4326 1990 4337 2014
rect 4287 1961 4337 1990
rect 4500 2009 4550 2038
rect 5440 2058 5490 2071
rect 5653 2058 5703 2071
rect 5861 2058 5911 2071
rect 6069 2058 6119 2071
rect 4500 1989 4517 2009
rect 4537 1989 4550 2009
rect 4500 1961 4550 1989
rect 384 1889 434 1917
rect 384 1869 397 1889
rect 417 1869 434 1889
rect 384 1840 434 1869
rect 597 1888 647 1917
rect 597 1864 608 1888
rect 632 1864 647 1888
rect 597 1840 647 1864
rect 805 1893 855 1917
rect 805 1869 817 1893
rect 841 1869 855 1893
rect 805 1840 855 1869
rect 1013 1891 1063 1917
rect 1013 1865 1031 1891
rect 1057 1865 1063 1891
rect 1013 1840 1063 1865
rect 8927 2054 8977 2079
rect 8927 2028 8933 2054
rect 8959 2028 8977 2054
rect 8927 2002 8977 2028
rect 9135 2050 9185 2079
rect 9135 2026 9149 2050
rect 9173 2026 9185 2050
rect 9135 2002 9185 2026
rect 9343 2055 9393 2079
rect 9343 2031 9358 2055
rect 9382 2031 9393 2055
rect 9343 2002 9393 2031
rect 9556 2050 9606 2079
rect 9556 2030 9573 2050
rect 9593 2030 9606 2050
rect 9556 2002 9606 2030
rect 5440 1930 5490 1958
rect 5440 1910 5453 1930
rect 5473 1910 5490 1930
rect 5440 1881 5490 1910
rect 5653 1929 5703 1958
rect 5653 1905 5664 1929
rect 5688 1905 5703 1929
rect 5653 1881 5703 1905
rect 5861 1934 5911 1958
rect 5861 1910 5873 1934
rect 5897 1910 5911 1934
rect 5861 1881 5911 1910
rect 6069 1932 6119 1958
rect 6069 1906 6087 1932
rect 6113 1906 6119 1932
rect 6069 1881 6119 1906
rect 8927 1889 8977 1902
rect 9135 1889 9185 1902
rect 9343 1889 9393 1902
rect 9556 1889 9606 1902
rect 3871 1848 3921 1861
rect 4079 1848 4129 1861
rect 4287 1848 4337 1861
rect 4500 1848 4550 1861
rect 2793 1813 2843 1829
rect 3001 1813 3051 1829
rect 3209 1813 3259 1829
rect 3422 1813 3472 1829
rect 384 1782 434 1798
rect 597 1782 647 1798
rect 805 1782 855 1798
rect 1013 1782 1063 1798
rect 7849 1854 7899 1870
rect 8057 1854 8107 1870
rect 8265 1854 8315 1870
rect 8478 1854 8528 1870
rect 5440 1823 5490 1839
rect 5653 1823 5703 1839
rect 5861 1823 5911 1839
rect 6069 1823 6119 1839
rect 1464 1735 1514 1748
rect 1677 1735 1727 1748
rect 1885 1735 1935 1748
rect 2093 1735 2143 1748
rect 2793 1746 2843 1771
rect 2793 1720 2799 1746
rect 2825 1720 2843 1746
rect 2793 1694 2843 1720
rect 3001 1742 3051 1771
rect 3001 1718 3015 1742
rect 3039 1718 3051 1742
rect 3001 1694 3051 1718
rect 3209 1747 3259 1771
rect 3209 1723 3224 1747
rect 3248 1723 3259 1747
rect 3209 1694 3259 1723
rect 3422 1742 3472 1771
rect 6520 1776 6570 1789
rect 6733 1776 6783 1789
rect 6941 1776 6991 1789
rect 7149 1776 7199 1789
rect 7849 1787 7899 1812
rect 3422 1722 3439 1742
rect 3459 1722 3472 1742
rect 3422 1694 3472 1722
rect 1464 1607 1514 1635
rect 1464 1587 1477 1607
rect 1497 1587 1514 1607
rect 1464 1558 1514 1587
rect 1677 1606 1727 1635
rect 1677 1582 1688 1606
rect 1712 1582 1727 1606
rect 1677 1558 1727 1582
rect 1885 1611 1935 1635
rect 1885 1587 1897 1611
rect 1921 1587 1935 1611
rect 1885 1558 1935 1587
rect 2093 1609 2143 1635
rect 2093 1583 2111 1609
rect 2137 1583 2143 1609
rect 7849 1761 7855 1787
rect 7881 1761 7899 1787
rect 7849 1735 7899 1761
rect 8057 1783 8107 1812
rect 8057 1759 8071 1783
rect 8095 1759 8107 1783
rect 8057 1735 8107 1759
rect 8265 1788 8315 1812
rect 8265 1764 8280 1788
rect 8304 1764 8315 1788
rect 8265 1735 8315 1764
rect 8478 1783 8528 1812
rect 8478 1763 8495 1783
rect 8515 1763 8528 1783
rect 8478 1735 8528 1763
rect 6520 1648 6570 1676
rect 6520 1628 6533 1648
rect 6553 1628 6570 1648
rect 2093 1558 2143 1583
rect 2793 1581 2843 1594
rect 3001 1581 3051 1594
rect 3209 1581 3259 1594
rect 3422 1581 3472 1594
rect 6520 1599 6570 1628
rect 6733 1647 6783 1676
rect 6733 1623 6744 1647
rect 6768 1623 6783 1647
rect 6733 1599 6783 1623
rect 6941 1652 6991 1676
rect 6941 1628 6953 1652
rect 6977 1628 6991 1652
rect 6941 1599 6991 1628
rect 7149 1650 7199 1676
rect 7149 1624 7167 1650
rect 7193 1624 7199 1650
rect 7149 1599 7199 1624
rect 7849 1622 7899 1635
rect 8057 1622 8107 1635
rect 8265 1622 8315 1635
rect 8478 1622 8528 1635
rect 3873 1531 3923 1547
rect 4081 1531 4131 1547
rect 4289 1531 4339 1547
rect 4502 1531 4552 1547
rect 1464 1500 1514 1516
rect 1677 1500 1727 1516
rect 1885 1500 1935 1516
rect 2093 1500 2143 1516
rect 8929 1572 8979 1588
rect 9137 1572 9187 1588
rect 9345 1572 9395 1588
rect 9558 1572 9608 1588
rect 6520 1541 6570 1557
rect 6733 1541 6783 1557
rect 6941 1541 6991 1557
rect 7149 1541 7199 1557
rect 5442 1509 5492 1522
rect 5655 1509 5705 1522
rect 5863 1509 5913 1522
rect 6071 1509 6121 1522
rect 386 1468 436 1481
rect 599 1468 649 1481
rect 807 1468 857 1481
rect 1015 1468 1065 1481
rect 3873 1464 3923 1489
rect 3873 1438 3879 1464
rect 3905 1438 3923 1464
rect 3873 1412 3923 1438
rect 4081 1460 4131 1489
rect 4081 1436 4095 1460
rect 4119 1436 4131 1460
rect 4081 1412 4131 1436
rect 4289 1465 4339 1489
rect 4289 1441 4304 1465
rect 4328 1441 4339 1465
rect 4289 1412 4339 1441
rect 4502 1460 4552 1489
rect 4502 1440 4519 1460
rect 4539 1440 4552 1460
rect 4502 1412 4552 1440
rect 386 1340 436 1368
rect 386 1320 399 1340
rect 419 1320 436 1340
rect 386 1291 436 1320
rect 599 1339 649 1368
rect 599 1315 610 1339
rect 634 1315 649 1339
rect 599 1291 649 1315
rect 807 1344 857 1368
rect 807 1320 819 1344
rect 843 1320 857 1344
rect 807 1291 857 1320
rect 1015 1342 1065 1368
rect 1015 1316 1033 1342
rect 1059 1316 1065 1342
rect 1015 1291 1065 1316
rect 8929 1505 8979 1530
rect 8929 1479 8935 1505
rect 8961 1479 8979 1505
rect 8929 1453 8979 1479
rect 9137 1501 9187 1530
rect 9137 1477 9151 1501
rect 9175 1477 9187 1501
rect 9137 1453 9187 1477
rect 9345 1506 9395 1530
rect 9345 1482 9360 1506
rect 9384 1482 9395 1506
rect 9345 1453 9395 1482
rect 9558 1501 9608 1530
rect 9558 1481 9575 1501
rect 9595 1481 9608 1501
rect 9558 1453 9608 1481
rect 5442 1381 5492 1409
rect 5442 1361 5455 1381
rect 5475 1361 5492 1381
rect 3873 1299 3923 1312
rect 4081 1299 4131 1312
rect 4289 1299 4339 1312
rect 4502 1299 4552 1312
rect 5442 1332 5492 1361
rect 5655 1380 5705 1409
rect 5655 1356 5666 1380
rect 5690 1356 5705 1380
rect 5655 1332 5705 1356
rect 5863 1385 5913 1409
rect 5863 1361 5875 1385
rect 5899 1361 5913 1385
rect 5863 1332 5913 1361
rect 6071 1383 6121 1409
rect 6071 1357 6089 1383
rect 6115 1357 6121 1383
rect 6071 1332 6121 1357
rect 8929 1340 8979 1353
rect 9137 1340 9187 1353
rect 9345 1340 9395 1353
rect 9558 1340 9608 1353
rect 5442 1274 5492 1290
rect 5655 1274 5705 1290
rect 5863 1274 5913 1290
rect 6071 1274 6121 1290
rect 386 1233 436 1249
rect 599 1233 649 1249
rect 807 1233 857 1249
rect 1015 1233 1065 1249
rect 6380 1265 6430 1278
rect 6593 1265 6643 1278
rect 6801 1265 6851 1278
rect 7009 1265 7059 1278
rect 1324 1224 1374 1237
rect 1537 1224 1587 1237
rect 1745 1224 1795 1237
rect 1953 1224 2003 1237
rect 2934 1221 2984 1237
rect 3142 1221 3192 1237
rect 3350 1221 3400 1237
rect 3563 1221 3613 1237
rect 2934 1154 2984 1179
rect 2934 1128 2940 1154
rect 2966 1128 2984 1154
rect 1324 1096 1374 1124
rect 1324 1076 1337 1096
rect 1357 1076 1374 1096
rect 1324 1047 1374 1076
rect 1537 1095 1587 1124
rect 1537 1071 1548 1095
rect 1572 1071 1587 1095
rect 1537 1047 1587 1071
rect 1745 1100 1795 1124
rect 1745 1076 1757 1100
rect 1781 1076 1795 1100
rect 1745 1047 1795 1076
rect 1953 1098 2003 1124
rect 2934 1102 2984 1128
rect 3142 1150 3192 1179
rect 3142 1126 3156 1150
rect 3180 1126 3192 1150
rect 3142 1102 3192 1126
rect 3350 1155 3400 1179
rect 3350 1131 3365 1155
rect 3389 1131 3400 1155
rect 3350 1102 3400 1131
rect 3563 1150 3613 1179
rect 3563 1130 3580 1150
rect 3600 1130 3613 1150
rect 3563 1102 3613 1130
rect 1953 1072 1971 1098
rect 1997 1072 2003 1098
rect 1953 1047 2003 1072
rect 1324 989 1374 1005
rect 1537 989 1587 1005
rect 1745 989 1795 1005
rect 1953 989 2003 1005
rect 7990 1262 8040 1278
rect 8198 1262 8248 1278
rect 8406 1262 8456 1278
rect 8619 1262 8669 1278
rect 7990 1195 8040 1220
rect 7990 1169 7996 1195
rect 8022 1169 8040 1195
rect 6380 1137 6430 1165
rect 6380 1117 6393 1137
rect 6413 1117 6430 1137
rect 6380 1088 6430 1117
rect 6593 1136 6643 1165
rect 6593 1112 6604 1136
rect 6628 1112 6643 1136
rect 6593 1088 6643 1112
rect 6801 1141 6851 1165
rect 6801 1117 6813 1141
rect 6837 1117 6851 1141
rect 6801 1088 6851 1117
rect 7009 1139 7059 1165
rect 7990 1143 8040 1169
rect 8198 1191 8248 1220
rect 8198 1167 8212 1191
rect 8236 1167 8248 1191
rect 8198 1143 8248 1167
rect 8406 1196 8456 1220
rect 8406 1172 8421 1196
rect 8445 1172 8456 1196
rect 8406 1143 8456 1172
rect 8619 1191 8669 1220
rect 8619 1171 8636 1191
rect 8656 1171 8669 1191
rect 8619 1143 8669 1171
rect 7009 1113 7027 1139
rect 7053 1113 7059 1139
rect 7009 1088 7059 1113
rect 6380 1030 6430 1046
rect 6593 1030 6643 1046
rect 6801 1030 6851 1046
rect 7009 1030 7059 1046
rect 7990 1030 8040 1043
rect 8198 1030 8248 1043
rect 8406 1030 8456 1043
rect 8619 1030 8669 1043
rect 2934 989 2984 1002
rect 3142 989 3192 1002
rect 3350 989 3400 1002
rect 3563 989 3613 1002
rect 8928 1018 8978 1034
rect 9136 1018 9186 1034
rect 9344 1018 9394 1034
rect 9557 1018 9607 1034
rect 3872 977 3922 993
rect 4080 977 4130 993
rect 4288 977 4338 993
rect 4501 977 4551 993
rect 385 914 435 927
rect 598 914 648 927
rect 806 914 856 927
rect 1014 914 1064 927
rect 3872 910 3922 935
rect 3872 884 3878 910
rect 3904 884 3922 910
rect 3872 858 3922 884
rect 4080 906 4130 935
rect 4080 882 4094 906
rect 4118 882 4130 906
rect 4080 858 4130 882
rect 4288 911 4338 935
rect 4288 887 4303 911
rect 4327 887 4338 911
rect 4288 858 4338 887
rect 4501 906 4551 935
rect 5441 955 5491 968
rect 5654 955 5704 968
rect 5862 955 5912 968
rect 6070 955 6120 968
rect 4501 886 4518 906
rect 4538 886 4551 906
rect 4501 858 4551 886
rect 385 786 435 814
rect 385 766 398 786
rect 418 766 435 786
rect 385 737 435 766
rect 598 785 648 814
rect 598 761 609 785
rect 633 761 648 785
rect 598 737 648 761
rect 806 790 856 814
rect 806 766 818 790
rect 842 766 856 790
rect 806 737 856 766
rect 1014 788 1064 814
rect 1014 762 1032 788
rect 1058 762 1064 788
rect 1014 737 1064 762
rect 8928 951 8978 976
rect 8928 925 8934 951
rect 8960 925 8978 951
rect 8928 899 8978 925
rect 9136 947 9186 976
rect 9136 923 9150 947
rect 9174 923 9186 947
rect 9136 899 9186 923
rect 9344 952 9394 976
rect 9344 928 9359 952
rect 9383 928 9394 952
rect 9344 899 9394 928
rect 9557 947 9607 976
rect 9557 927 9574 947
rect 9594 927 9607 947
rect 9557 899 9607 927
rect 5441 827 5491 855
rect 5441 807 5454 827
rect 5474 807 5491 827
rect 5441 778 5491 807
rect 5654 826 5704 855
rect 5654 802 5665 826
rect 5689 802 5704 826
rect 5654 778 5704 802
rect 5862 831 5912 855
rect 5862 807 5874 831
rect 5898 807 5912 831
rect 5862 778 5912 807
rect 6070 829 6120 855
rect 6070 803 6088 829
rect 6114 803 6120 829
rect 6070 778 6120 803
rect 8928 786 8978 799
rect 9136 786 9186 799
rect 9344 786 9394 799
rect 9557 786 9607 799
rect 3872 745 3922 758
rect 4080 745 4130 758
rect 4288 745 4338 758
rect 4501 745 4551 758
rect 385 679 435 695
rect 598 679 648 695
rect 806 679 856 695
rect 1014 679 1064 695
rect 5441 720 5491 736
rect 5654 720 5704 736
rect 5862 720 5912 736
rect 6070 720 6120 736
rect 6688 396 6738 409
rect 6901 396 6951 409
rect 7109 396 7159 409
rect 7317 396 7367 409
rect 1632 355 1682 368
rect 1845 355 1895 368
rect 2053 355 2103 368
rect 2261 355 2311 368
rect 4582 335 4632 348
rect 4795 335 4845 348
rect 5003 335 5053 348
rect 5211 335 5261 348
rect 1632 227 1682 255
rect 1632 207 1645 227
rect 1665 207 1682 227
rect 1632 178 1682 207
rect 1845 226 1895 255
rect 1845 202 1856 226
rect 1880 202 1895 226
rect 1845 178 1895 202
rect 2053 231 2103 255
rect 2053 207 2065 231
rect 2089 207 2103 231
rect 2053 178 2103 207
rect 2261 229 2311 255
rect 6688 268 6738 296
rect 6688 248 6701 268
rect 6721 248 6738 268
rect 2261 203 2279 229
rect 2305 203 2311 229
rect 2261 178 2311 203
rect 4582 207 4632 235
rect 4582 187 4595 207
rect 4615 187 4632 207
rect 4582 158 4632 187
rect 4795 206 4845 235
rect 4795 182 4806 206
rect 4830 182 4845 206
rect 4795 158 4845 182
rect 5003 211 5053 235
rect 5003 187 5015 211
rect 5039 187 5053 211
rect 5003 158 5053 187
rect 5211 209 5261 235
rect 6688 219 6738 248
rect 6901 267 6951 296
rect 6901 243 6912 267
rect 6936 243 6951 267
rect 6901 219 6951 243
rect 7109 272 7159 296
rect 7109 248 7121 272
rect 7145 248 7159 272
rect 7109 219 7159 248
rect 7317 270 7367 296
rect 7317 244 7335 270
rect 7361 244 7367 270
rect 7317 219 7367 244
rect 5211 183 5229 209
rect 5255 183 5261 209
rect 5211 158 5261 183
rect 6688 161 6738 177
rect 6901 161 6951 177
rect 7109 161 7159 177
rect 7317 161 7367 177
rect 1632 120 1682 136
rect 1845 120 1895 136
rect 2053 120 2103 136
rect 2261 120 2311 136
rect 4582 100 4632 116
rect 4795 100 4845 116
rect 5003 100 5053 116
rect 5211 100 5261 116
<< polycont >>
rect 3875 9159 3901 9185
rect 4091 9157 4115 9181
rect 4300 9162 4324 9186
rect 4515 9161 4535 9181
rect 395 9041 415 9061
rect 606 9036 630 9060
rect 815 9041 839 9065
rect 1029 9037 1055 9063
rect 8931 9200 8957 9226
rect 9147 9198 9171 9222
rect 9356 9203 9380 9227
rect 9571 9202 9591 9222
rect 5451 9082 5471 9102
rect 5662 9077 5686 9101
rect 5871 9082 5895 9106
rect 6085 9078 6111 9104
rect 2936 8849 2962 8875
rect 1333 8797 1353 8817
rect 1544 8792 1568 8816
rect 1753 8797 1777 8821
rect 3152 8847 3176 8871
rect 3361 8852 3385 8876
rect 3576 8851 3596 8871
rect 1967 8793 1993 8819
rect 7992 8890 8018 8916
rect 6389 8838 6409 8858
rect 6600 8833 6624 8857
rect 6809 8838 6833 8862
rect 8208 8888 8232 8912
rect 8417 8893 8441 8917
rect 8632 8892 8652 8912
rect 7023 8834 7049 8860
rect 3874 8605 3900 8631
rect 4090 8603 4114 8627
rect 4299 8608 4323 8632
rect 4514 8607 4534 8627
rect 394 8487 414 8507
rect 605 8482 629 8506
rect 814 8487 838 8511
rect 1028 8483 1054 8509
rect 8930 8646 8956 8672
rect 9146 8644 9170 8668
rect 9355 8649 9379 8673
rect 9570 8648 9590 8668
rect 5450 8528 5470 8548
rect 5661 8523 5685 8547
rect 5870 8528 5894 8552
rect 6084 8524 6110 8550
rect 2796 8338 2822 8364
rect 3012 8336 3036 8360
rect 3221 8341 3245 8365
rect 3436 8340 3456 8360
rect 1474 8205 1494 8225
rect 1685 8200 1709 8224
rect 1894 8205 1918 8229
rect 2108 8201 2134 8227
rect 7852 8379 7878 8405
rect 8068 8377 8092 8401
rect 8277 8382 8301 8406
rect 8492 8381 8512 8401
rect 6530 8246 6550 8266
rect 6741 8241 6765 8265
rect 6950 8246 6974 8270
rect 7164 8242 7190 8268
rect 3876 8056 3902 8082
rect 4092 8054 4116 8078
rect 4301 8059 4325 8083
rect 4516 8058 4536 8078
rect 396 7938 416 7958
rect 607 7933 631 7957
rect 816 7938 840 7962
rect 1030 7934 1056 7960
rect 8932 8097 8958 8123
rect 9148 8095 9172 8119
rect 9357 8100 9381 8124
rect 9572 8099 9592 8119
rect 5452 7979 5472 7999
rect 5663 7974 5687 7998
rect 5872 7979 5896 8003
rect 6086 7975 6112 8001
rect 2937 7746 2963 7772
rect 1334 7694 1354 7714
rect 1545 7689 1569 7713
rect 1754 7694 1778 7718
rect 3153 7744 3177 7768
rect 3362 7749 3386 7773
rect 3577 7748 3597 7768
rect 1968 7690 1994 7716
rect 7993 7787 8019 7813
rect 6390 7735 6410 7755
rect 6601 7730 6625 7754
rect 6810 7735 6834 7759
rect 8209 7785 8233 7809
rect 8418 7790 8442 7814
rect 8633 7789 8653 7809
rect 7024 7731 7050 7757
rect 3875 7502 3901 7528
rect 4091 7500 4115 7524
rect 4300 7505 4324 7529
rect 4515 7504 4535 7524
rect 395 7384 415 7404
rect 606 7379 630 7403
rect 815 7384 839 7408
rect 1029 7380 1055 7406
rect 8931 7543 8957 7569
rect 9147 7541 9171 7565
rect 9356 7546 9380 7570
rect 9571 7545 9591 7565
rect 5451 7425 5471 7445
rect 5662 7420 5686 7444
rect 5871 7425 5895 7449
rect 6085 7421 6111 7447
rect 2827 7222 2853 7248
rect 3043 7220 3067 7244
rect 3252 7225 3276 7249
rect 3467 7224 3487 7244
rect 7883 7263 7909 7289
rect 8099 7261 8123 7285
rect 8308 7266 8332 7290
rect 8523 7265 8543 7285
rect 1444 7115 1464 7135
rect 1655 7110 1679 7134
rect 1864 7115 1888 7139
rect 2078 7111 2104 7137
rect 6500 7156 6520 7176
rect 6711 7151 6735 7175
rect 6920 7156 6944 7180
rect 7134 7152 7160 7178
rect 3876 6953 3902 6979
rect 4092 6951 4116 6975
rect 4301 6956 4325 6980
rect 4516 6955 4536 6975
rect 396 6835 416 6855
rect 607 6830 631 6854
rect 816 6835 840 6859
rect 1030 6831 1056 6857
rect 8932 6994 8958 7020
rect 9148 6992 9172 7016
rect 9357 6997 9381 7021
rect 9572 6996 9592 7016
rect 5452 6876 5472 6896
rect 5663 6871 5687 6895
rect 5872 6876 5896 6900
rect 6086 6872 6112 6898
rect 2937 6643 2963 6669
rect 1334 6591 1354 6611
rect 1545 6586 1569 6610
rect 1754 6591 1778 6615
rect 3153 6641 3177 6665
rect 3362 6646 3386 6670
rect 3577 6645 3597 6665
rect 1968 6587 1994 6613
rect 7993 6684 8019 6710
rect 6390 6632 6410 6652
rect 6601 6627 6625 6651
rect 6810 6632 6834 6656
rect 8209 6682 8233 6706
rect 8418 6687 8442 6711
rect 8633 6686 8653 6706
rect 7024 6628 7050 6654
rect 3875 6399 3901 6425
rect 4091 6397 4115 6421
rect 4300 6402 4324 6426
rect 4515 6401 4535 6421
rect 395 6281 415 6301
rect 606 6276 630 6300
rect 815 6281 839 6305
rect 1029 6277 1055 6303
rect 8931 6440 8957 6466
rect 9147 6438 9171 6462
rect 9356 6443 9380 6467
rect 9571 6442 9591 6462
rect 5451 6322 5471 6342
rect 5662 6317 5686 6341
rect 5871 6322 5895 6346
rect 6085 6318 6111 6344
rect 2797 6132 2823 6158
rect 3013 6130 3037 6154
rect 3222 6135 3246 6159
rect 3437 6134 3457 6154
rect 1475 5999 1495 6019
rect 1686 5994 1710 6018
rect 1895 5999 1919 6023
rect 2109 5995 2135 6021
rect 7853 6173 7879 6199
rect 8069 6171 8093 6195
rect 8278 6176 8302 6200
rect 8493 6175 8513 6195
rect 6531 6040 6551 6060
rect 6742 6035 6766 6059
rect 6951 6040 6975 6064
rect 7165 6036 7191 6062
rect 3877 5850 3903 5876
rect 4093 5848 4117 5872
rect 4302 5853 4326 5877
rect 4517 5852 4537 5872
rect 397 5732 417 5752
rect 608 5727 632 5751
rect 817 5732 841 5756
rect 1031 5728 1057 5754
rect 8933 5891 8959 5917
rect 9149 5889 9173 5913
rect 9358 5894 9382 5918
rect 9573 5893 9593 5913
rect 5453 5773 5473 5793
rect 5664 5768 5688 5792
rect 5873 5773 5897 5797
rect 6087 5769 6113 5795
rect 2938 5540 2964 5566
rect 1335 5488 1355 5508
rect 1546 5483 1570 5507
rect 1755 5488 1779 5512
rect 3154 5538 3178 5562
rect 3363 5543 3387 5567
rect 3578 5542 3598 5562
rect 1969 5484 1995 5510
rect 7994 5581 8020 5607
rect 6391 5529 6411 5549
rect 6602 5524 6626 5548
rect 6811 5529 6835 5553
rect 8210 5579 8234 5603
rect 8419 5584 8443 5608
rect 8634 5583 8654 5603
rect 7025 5525 7051 5551
rect 3876 5296 3902 5322
rect 4092 5294 4116 5318
rect 4301 5299 4325 5323
rect 4516 5298 4536 5318
rect 396 5178 416 5198
rect 607 5173 631 5197
rect 816 5178 840 5202
rect 1030 5174 1056 5200
rect 8932 5337 8958 5363
rect 9148 5335 9172 5359
rect 9357 5340 9381 5364
rect 9572 5339 9592 5359
rect 5452 5219 5472 5239
rect 5663 5214 5687 5238
rect 5872 5219 5896 5243
rect 6086 5215 6112 5241
rect 2829 5010 2855 5036
rect 3045 5008 3069 5032
rect 3254 5013 3278 5037
rect 3469 5012 3489 5032
rect 7885 5051 7911 5077
rect 8101 5049 8125 5073
rect 8310 5054 8334 5078
rect 8525 5053 8545 5073
rect 1444 4915 1464 4935
rect 1655 4910 1679 4934
rect 1864 4915 1888 4939
rect 2078 4911 2104 4937
rect 6500 4956 6520 4976
rect 6711 4951 6735 4975
rect 6920 4956 6944 4980
rect 7134 4952 7160 4978
rect 3877 4747 3903 4773
rect 4093 4745 4117 4769
rect 4302 4750 4326 4774
rect 4517 4749 4537 4769
rect 397 4629 417 4649
rect 608 4624 632 4648
rect 817 4629 841 4653
rect 1031 4625 1057 4651
rect 8933 4788 8959 4814
rect 9149 4786 9173 4810
rect 9358 4791 9382 4815
rect 9573 4790 9593 4810
rect 5453 4670 5473 4690
rect 5664 4665 5688 4689
rect 5873 4670 5897 4694
rect 6087 4666 6113 4692
rect 2938 4437 2964 4463
rect 1335 4385 1355 4405
rect 1546 4380 1570 4404
rect 1755 4385 1779 4409
rect 3154 4435 3178 4459
rect 3363 4440 3387 4464
rect 3578 4439 3598 4459
rect 1969 4381 1995 4407
rect 7994 4478 8020 4504
rect 6391 4426 6411 4446
rect 6602 4421 6626 4445
rect 6811 4426 6835 4450
rect 8210 4476 8234 4500
rect 8419 4481 8443 4505
rect 8634 4480 8654 4500
rect 7025 4422 7051 4448
rect 3876 4193 3902 4219
rect 4092 4191 4116 4215
rect 4301 4196 4325 4220
rect 4516 4195 4536 4215
rect 396 4075 416 4095
rect 607 4070 631 4094
rect 816 4075 840 4099
rect 1030 4071 1056 4097
rect 8932 4234 8958 4260
rect 9148 4232 9172 4256
rect 9357 4237 9381 4261
rect 9572 4236 9592 4256
rect 5452 4116 5472 4136
rect 5663 4111 5687 4135
rect 5872 4116 5896 4140
rect 6086 4112 6112 4138
rect 2798 3926 2824 3952
rect 3014 3924 3038 3948
rect 3223 3929 3247 3953
rect 3438 3928 3458 3948
rect 1476 3793 1496 3813
rect 1687 3788 1711 3812
rect 1896 3793 1920 3817
rect 2110 3789 2136 3815
rect 7854 3967 7880 3993
rect 8070 3965 8094 3989
rect 8279 3970 8303 3994
rect 8494 3969 8514 3989
rect 6532 3834 6552 3854
rect 6743 3829 6767 3853
rect 6952 3834 6976 3858
rect 7166 3830 7192 3856
rect 3878 3644 3904 3670
rect 4094 3642 4118 3666
rect 4303 3647 4327 3671
rect 4518 3646 4538 3666
rect 398 3526 418 3546
rect 609 3521 633 3545
rect 818 3526 842 3550
rect 1032 3522 1058 3548
rect 8934 3685 8960 3711
rect 9150 3683 9174 3707
rect 9359 3688 9383 3712
rect 9574 3687 9594 3707
rect 5454 3567 5474 3587
rect 5665 3562 5689 3586
rect 5874 3567 5898 3591
rect 6088 3563 6114 3589
rect 2939 3334 2965 3360
rect 1336 3282 1356 3302
rect 1547 3277 1571 3301
rect 1756 3282 1780 3306
rect 3155 3332 3179 3356
rect 3364 3337 3388 3361
rect 3579 3336 3599 3356
rect 1970 3278 1996 3304
rect 7995 3375 8021 3401
rect 6392 3323 6412 3343
rect 6603 3318 6627 3342
rect 6812 3323 6836 3347
rect 8211 3373 8235 3397
rect 8420 3378 8444 3402
rect 8635 3377 8655 3397
rect 7026 3319 7052 3345
rect 3877 3090 3903 3116
rect 4093 3088 4117 3112
rect 4302 3093 4326 3117
rect 4517 3092 4537 3112
rect 397 2972 417 2992
rect 608 2967 632 2991
rect 817 2972 841 2996
rect 1031 2968 1057 2994
rect 8933 3131 8959 3157
rect 9149 3129 9173 3153
rect 9358 3134 9382 3158
rect 9573 3133 9593 3153
rect 5453 3013 5473 3033
rect 5664 3008 5688 3032
rect 5873 3013 5897 3037
rect 6087 3009 6113 3035
rect 2829 2810 2855 2836
rect 3045 2808 3069 2832
rect 3254 2813 3278 2837
rect 3469 2812 3489 2832
rect 7885 2851 7911 2877
rect 8101 2849 8125 2873
rect 8310 2854 8334 2878
rect 8525 2853 8545 2873
rect 1446 2703 1466 2723
rect 1657 2698 1681 2722
rect 1866 2703 1890 2727
rect 2080 2699 2106 2725
rect 6502 2744 6522 2764
rect 6713 2739 6737 2763
rect 6922 2744 6946 2768
rect 7136 2740 7162 2766
rect 3878 2541 3904 2567
rect 4094 2539 4118 2563
rect 4303 2544 4327 2568
rect 4518 2543 4538 2563
rect 398 2423 418 2443
rect 609 2418 633 2442
rect 818 2423 842 2447
rect 1032 2419 1058 2445
rect 8934 2582 8960 2608
rect 9150 2580 9174 2604
rect 9359 2585 9383 2609
rect 9574 2584 9594 2604
rect 5454 2464 5474 2484
rect 5665 2459 5689 2483
rect 5874 2464 5898 2488
rect 6088 2460 6114 2486
rect 2939 2231 2965 2257
rect 1336 2179 1356 2199
rect 1547 2174 1571 2198
rect 1756 2179 1780 2203
rect 3155 2229 3179 2253
rect 3364 2234 3388 2258
rect 3579 2233 3599 2253
rect 1970 2175 1996 2201
rect 7995 2272 8021 2298
rect 6392 2220 6412 2240
rect 6603 2215 6627 2239
rect 6812 2220 6836 2244
rect 8211 2270 8235 2294
rect 8420 2275 8444 2299
rect 8635 2274 8655 2294
rect 7026 2216 7052 2242
rect 3877 1987 3903 2013
rect 4093 1985 4117 2009
rect 4302 1990 4326 2014
rect 4517 1989 4537 2009
rect 397 1869 417 1889
rect 608 1864 632 1888
rect 817 1869 841 1893
rect 1031 1865 1057 1891
rect 8933 2028 8959 2054
rect 9149 2026 9173 2050
rect 9358 2031 9382 2055
rect 9573 2030 9593 2050
rect 5453 1910 5473 1930
rect 5664 1905 5688 1929
rect 5873 1910 5897 1934
rect 6087 1906 6113 1932
rect 2799 1720 2825 1746
rect 3015 1718 3039 1742
rect 3224 1723 3248 1747
rect 3439 1722 3459 1742
rect 1477 1587 1497 1607
rect 1688 1582 1712 1606
rect 1897 1587 1921 1611
rect 2111 1583 2137 1609
rect 7855 1761 7881 1787
rect 8071 1759 8095 1783
rect 8280 1764 8304 1788
rect 8495 1763 8515 1783
rect 6533 1628 6553 1648
rect 6744 1623 6768 1647
rect 6953 1628 6977 1652
rect 7167 1624 7193 1650
rect 3879 1438 3905 1464
rect 4095 1436 4119 1460
rect 4304 1441 4328 1465
rect 4519 1440 4539 1460
rect 399 1320 419 1340
rect 610 1315 634 1339
rect 819 1320 843 1344
rect 1033 1316 1059 1342
rect 8935 1479 8961 1505
rect 9151 1477 9175 1501
rect 9360 1482 9384 1506
rect 9575 1481 9595 1501
rect 5455 1361 5475 1381
rect 5666 1356 5690 1380
rect 5875 1361 5899 1385
rect 6089 1357 6115 1383
rect 2940 1128 2966 1154
rect 1337 1076 1357 1096
rect 1548 1071 1572 1095
rect 1757 1076 1781 1100
rect 3156 1126 3180 1150
rect 3365 1131 3389 1155
rect 3580 1130 3600 1150
rect 1971 1072 1997 1098
rect 7996 1169 8022 1195
rect 6393 1117 6413 1137
rect 6604 1112 6628 1136
rect 6813 1117 6837 1141
rect 8212 1167 8236 1191
rect 8421 1172 8445 1196
rect 8636 1171 8656 1191
rect 7027 1113 7053 1139
rect 3878 884 3904 910
rect 4094 882 4118 906
rect 4303 887 4327 911
rect 4518 886 4538 906
rect 398 766 418 786
rect 609 761 633 785
rect 818 766 842 790
rect 1032 762 1058 788
rect 8934 925 8960 951
rect 9150 923 9174 947
rect 9359 928 9383 952
rect 9574 927 9594 947
rect 5454 807 5474 827
rect 5665 802 5689 826
rect 5874 807 5898 831
rect 6088 803 6114 829
rect 1645 207 1665 227
rect 1856 202 1880 226
rect 2065 207 2089 231
rect 6701 248 6721 268
rect 2279 203 2305 229
rect 4595 187 4615 207
rect 4806 182 4830 206
rect 5015 187 5039 211
rect 6912 243 6936 267
rect 7121 248 7145 272
rect 7335 244 7361 270
rect 5229 183 5255 209
<< ndiffres >>
rect 5151 9326 5208 9345
rect 5151 9323 5172 9326
rect 95 9285 152 9304
rect 5057 9308 5172 9323
rect 5190 9308 5208 9326
rect 95 9282 116 9285
rect 1 9267 116 9282
rect 134 9267 152 9285
rect 5057 9285 5208 9308
rect 1 9244 152 9267
rect 1 9208 43 9244
rect 5057 9249 5099 9285
rect 5056 9248 5156 9249
rect 5056 9227 5212 9248
rect 0 9207 100 9208
rect 0 9186 156 9207
rect 0 9168 118 9186
rect 136 9168 156 9186
rect 0 9164 156 9168
rect 95 9148 156 9164
rect 95 9098 152 9117
rect 95 9095 116 9098
rect 1 9080 116 9095
rect 134 9080 152 9098
rect 5056 9209 5174 9227
rect 5192 9209 5212 9227
rect 5056 9205 5212 9209
rect 5151 9189 5212 9205
rect 4773 9150 4834 9166
rect 4773 9146 4929 9150
rect 1 9057 152 9080
rect 1 9021 43 9057
rect 0 9020 100 9021
rect 0 8999 156 9020
rect 0 8981 118 8999
rect 136 8981 156 8999
rect 0 8977 156 8981
rect 95 8961 156 8977
rect 4773 9128 4793 9146
rect 4811 9128 4929 9146
rect 5151 9139 5208 9158
rect 5151 9136 5172 9139
rect 4773 9107 4929 9128
rect 4829 9106 4929 9107
rect 5057 9121 5172 9136
rect 5190 9121 5208 9139
rect 9829 9191 9890 9207
rect 9829 9187 9985 9191
rect 4886 9070 4928 9106
rect 4777 9047 4928 9070
rect 5057 9098 5208 9121
rect 5057 9062 5099 9098
rect 4777 9029 4795 9047
rect 4813 9032 4928 9047
rect 5056 9061 5156 9062
rect 5056 9040 5212 9061
rect 4813 9029 4834 9032
rect 4777 9010 4834 9029
rect 5056 9022 5174 9040
rect 5192 9022 5212 9040
rect 5056 9018 5212 9022
rect 5151 9002 5212 9018
rect 9829 9169 9849 9187
rect 9867 9169 9985 9187
rect 9829 9148 9985 9169
rect 9885 9147 9985 9148
rect 9942 9111 9984 9147
rect 9833 9088 9984 9111
rect 9833 9070 9851 9088
rect 9869 9073 9984 9088
rect 9869 9070 9890 9073
rect 9833 9051 9890 9070
rect 95 8869 152 8888
rect 95 8866 116 8869
rect 1 8851 116 8866
rect 134 8851 152 8869
rect 1 8828 152 8851
rect 4773 8920 4834 8936
rect 4773 8916 4929 8920
rect 1 8792 43 8828
rect 0 8791 100 8792
rect 0 8770 156 8791
rect 0 8752 118 8770
rect 136 8752 156 8770
rect 4773 8898 4793 8916
rect 4811 8898 4929 8916
rect 5151 8910 5208 8929
rect 5151 8907 5172 8910
rect 4773 8877 4929 8898
rect 4829 8876 4929 8877
rect 5057 8892 5172 8907
rect 5190 8892 5208 8910
rect 4886 8840 4928 8876
rect 0 8748 156 8752
rect 95 8732 156 8748
rect 4777 8817 4928 8840
rect 5057 8869 5208 8892
rect 9829 8961 9890 8977
rect 9829 8957 9985 8961
rect 5057 8833 5099 8869
rect 4777 8799 4795 8817
rect 4813 8802 4928 8817
rect 5056 8832 5156 8833
rect 5056 8811 5212 8832
rect 4813 8799 4834 8802
rect 4777 8780 4834 8799
rect 5056 8793 5174 8811
rect 5192 8793 5212 8811
rect 9829 8939 9849 8957
rect 9867 8939 9985 8957
rect 9829 8918 9985 8939
rect 9885 8917 9985 8918
rect 9942 8881 9984 8917
rect 5056 8789 5212 8793
rect 5151 8773 5212 8789
rect 9833 8858 9984 8881
rect 9833 8840 9851 8858
rect 9869 8843 9984 8858
rect 9869 8840 9890 8843
rect 9833 8821 9890 8840
rect 95 8639 152 8658
rect 95 8636 116 8639
rect 1 8621 116 8636
rect 134 8621 152 8639
rect 1 8598 152 8621
rect 1 8562 43 8598
rect 0 8561 100 8562
rect 0 8540 156 8561
rect 0 8522 118 8540
rect 136 8522 156 8540
rect 4773 8691 4834 8707
rect 4773 8687 4929 8691
rect 4773 8669 4793 8687
rect 4811 8669 4929 8687
rect 5151 8680 5208 8699
rect 5151 8677 5172 8680
rect 4773 8648 4929 8669
rect 4829 8647 4929 8648
rect 5057 8662 5172 8677
rect 5190 8662 5208 8680
rect 4886 8611 4928 8647
rect 4777 8588 4928 8611
rect 5057 8639 5208 8662
rect 5057 8603 5099 8639
rect 0 8518 156 8522
rect 95 8502 156 8518
rect 4777 8570 4795 8588
rect 4813 8573 4928 8588
rect 5056 8602 5156 8603
rect 5056 8581 5212 8602
rect 4813 8570 4834 8573
rect 4777 8551 4834 8570
rect 5056 8563 5174 8581
rect 5192 8563 5212 8581
rect 9829 8732 9890 8748
rect 9829 8728 9985 8732
rect 9829 8710 9849 8728
rect 9867 8710 9985 8728
rect 9829 8689 9985 8710
rect 9885 8688 9985 8689
rect 9942 8652 9984 8688
rect 9833 8629 9984 8652
rect 5056 8559 5212 8563
rect 5151 8543 5212 8559
rect 4773 8504 4834 8520
rect 4773 8500 4929 8504
rect 4773 8482 4793 8500
rect 4811 8482 4929 8500
rect 9833 8611 9851 8629
rect 9869 8614 9984 8629
rect 9869 8611 9890 8614
rect 9833 8592 9890 8611
rect 9829 8545 9890 8561
rect 9829 8541 9985 8545
rect 9829 8523 9849 8541
rect 9867 8523 9985 8541
rect 9829 8502 9985 8523
rect 9885 8501 9985 8502
rect 4773 8461 4929 8482
rect 4829 8460 4929 8461
rect 4886 8424 4928 8460
rect 4777 8401 4928 8424
rect 9942 8465 9984 8501
rect 9833 8442 9984 8465
rect 4777 8383 4795 8401
rect 4813 8386 4928 8401
rect 4813 8383 4834 8386
rect 4777 8364 4834 8383
rect 96 8182 153 8201
rect 96 8179 117 8182
rect 2 8164 117 8179
rect 135 8164 153 8182
rect 9833 8424 9851 8442
rect 9869 8427 9984 8442
rect 9869 8424 9890 8427
rect 9833 8405 9890 8424
rect 5152 8223 5209 8242
rect 5152 8220 5173 8223
rect 5058 8205 5173 8220
rect 5191 8205 5209 8223
rect 2 8141 153 8164
rect 2 8105 44 8141
rect 5058 8182 5209 8205
rect 5058 8146 5100 8182
rect 5057 8145 5157 8146
rect 5057 8124 5213 8145
rect 1 8104 101 8105
rect 1 8083 157 8104
rect 1 8065 119 8083
rect 137 8065 157 8083
rect 1 8061 157 8065
rect 96 8045 157 8061
rect 96 7995 153 8014
rect 96 7992 117 7995
rect 2 7977 117 7992
rect 135 7977 153 7995
rect 5057 8106 5175 8124
rect 5193 8106 5213 8124
rect 5057 8102 5213 8106
rect 5152 8086 5213 8102
rect 4774 8047 4835 8063
rect 4774 8043 4930 8047
rect 2 7954 153 7977
rect 2 7918 44 7954
rect 1 7917 101 7918
rect 1 7896 157 7917
rect 1 7878 119 7896
rect 137 7878 157 7896
rect 1 7874 157 7878
rect 96 7858 157 7874
rect 4774 8025 4794 8043
rect 4812 8025 4930 8043
rect 5152 8036 5209 8055
rect 5152 8033 5173 8036
rect 4774 8004 4930 8025
rect 4830 8003 4930 8004
rect 5058 8018 5173 8033
rect 5191 8018 5209 8036
rect 9830 8088 9891 8104
rect 9830 8084 9986 8088
rect 4887 7967 4929 8003
rect 4778 7944 4929 7967
rect 5058 7995 5209 8018
rect 5058 7959 5100 7995
rect 4778 7926 4796 7944
rect 4814 7929 4929 7944
rect 5057 7958 5157 7959
rect 5057 7937 5213 7958
rect 4814 7926 4835 7929
rect 4778 7907 4835 7926
rect 5057 7919 5175 7937
rect 5193 7919 5213 7937
rect 5057 7915 5213 7919
rect 5152 7899 5213 7915
rect 9830 8066 9850 8084
rect 9868 8066 9986 8084
rect 9830 8045 9986 8066
rect 9886 8044 9986 8045
rect 9943 8008 9985 8044
rect 9834 7985 9985 8008
rect 9834 7967 9852 7985
rect 9870 7970 9985 7985
rect 9870 7967 9891 7970
rect 9834 7948 9891 7967
rect 96 7766 153 7785
rect 96 7763 117 7766
rect 2 7748 117 7763
rect 135 7748 153 7766
rect 2 7725 153 7748
rect 4774 7817 4835 7833
rect 4774 7813 4930 7817
rect 2 7689 44 7725
rect 1 7688 101 7689
rect 1 7667 157 7688
rect 1 7649 119 7667
rect 137 7649 157 7667
rect 4774 7795 4794 7813
rect 4812 7795 4930 7813
rect 5152 7807 5209 7826
rect 5152 7804 5173 7807
rect 4774 7774 4930 7795
rect 4830 7773 4930 7774
rect 5058 7789 5173 7804
rect 5191 7789 5209 7807
rect 4887 7737 4929 7773
rect 1 7645 157 7649
rect 96 7629 157 7645
rect 4778 7714 4929 7737
rect 5058 7766 5209 7789
rect 9830 7858 9891 7874
rect 9830 7854 9986 7858
rect 5058 7730 5100 7766
rect 4778 7696 4796 7714
rect 4814 7699 4929 7714
rect 5057 7729 5157 7730
rect 5057 7708 5213 7729
rect 4814 7696 4835 7699
rect 4778 7677 4835 7696
rect 5057 7690 5175 7708
rect 5193 7690 5213 7708
rect 9830 7836 9850 7854
rect 9868 7836 9986 7854
rect 9830 7815 9986 7836
rect 9886 7814 9986 7815
rect 9943 7778 9985 7814
rect 5057 7686 5213 7690
rect 5152 7670 5213 7686
rect 9834 7755 9985 7778
rect 9834 7737 9852 7755
rect 9870 7740 9985 7755
rect 9870 7737 9891 7740
rect 9834 7718 9891 7737
rect 96 7536 153 7555
rect 96 7533 117 7536
rect 2 7518 117 7533
rect 135 7518 153 7536
rect 2 7495 153 7518
rect 2 7459 44 7495
rect 1 7458 101 7459
rect 1 7437 157 7458
rect 1 7419 119 7437
rect 137 7419 157 7437
rect 4774 7588 4835 7604
rect 4774 7584 4930 7588
rect 4774 7566 4794 7584
rect 4812 7566 4930 7584
rect 5152 7577 5209 7596
rect 5152 7574 5173 7577
rect 4774 7545 4930 7566
rect 4830 7544 4930 7545
rect 5058 7559 5173 7574
rect 5191 7559 5209 7577
rect 4887 7508 4929 7544
rect 4778 7485 4929 7508
rect 5058 7536 5209 7559
rect 5058 7500 5100 7536
rect 1 7415 157 7419
rect 96 7399 157 7415
rect 4778 7467 4796 7485
rect 4814 7470 4929 7485
rect 5057 7499 5157 7500
rect 5057 7478 5213 7499
rect 4814 7467 4835 7470
rect 4778 7448 4835 7467
rect 5057 7460 5175 7478
rect 5193 7460 5213 7478
rect 9830 7629 9891 7645
rect 9830 7625 9986 7629
rect 9830 7607 9850 7625
rect 9868 7607 9986 7625
rect 9830 7586 9986 7607
rect 9886 7585 9986 7586
rect 9943 7549 9985 7585
rect 9834 7526 9985 7549
rect 5057 7456 5213 7460
rect 5152 7440 5213 7456
rect 4774 7401 4835 7417
rect 4774 7397 4930 7401
rect 4774 7379 4794 7397
rect 4812 7379 4930 7397
rect 9834 7508 9852 7526
rect 9870 7511 9985 7526
rect 9870 7508 9891 7511
rect 9834 7489 9891 7508
rect 9830 7442 9891 7458
rect 9830 7438 9986 7442
rect 9830 7420 9850 7438
rect 9868 7420 9986 7438
rect 9830 7399 9986 7420
rect 9886 7398 9986 7399
rect 4774 7358 4930 7379
rect 4830 7357 4930 7358
rect 4887 7321 4929 7357
rect 4778 7298 4929 7321
rect 4778 7280 4796 7298
rect 4814 7283 4929 7298
rect 9943 7362 9985 7398
rect 9834 7339 9985 7362
rect 9834 7321 9852 7339
rect 9870 7324 9985 7339
rect 9870 7321 9891 7324
rect 4814 7280 4835 7283
rect 4778 7261 4835 7280
rect 9834 7302 9891 7321
rect 96 7079 153 7098
rect 5152 7120 5209 7139
rect 5152 7117 5173 7120
rect 96 7076 117 7079
rect 2 7061 117 7076
rect 135 7061 153 7079
rect 2 7038 153 7061
rect 2 7002 44 7038
rect 5058 7102 5173 7117
rect 5191 7102 5209 7120
rect 5058 7079 5209 7102
rect 5058 7043 5100 7079
rect 5057 7042 5157 7043
rect 5057 7021 5213 7042
rect 1 7001 101 7002
rect 1 6980 157 7001
rect 1 6962 119 6980
rect 137 6962 157 6980
rect 1 6958 157 6962
rect 96 6942 157 6958
rect 96 6892 153 6911
rect 96 6889 117 6892
rect 2 6874 117 6889
rect 135 6874 153 6892
rect 5057 7003 5175 7021
rect 5193 7003 5213 7021
rect 5057 6999 5213 7003
rect 5152 6983 5213 6999
rect 4774 6944 4835 6960
rect 4774 6940 4930 6944
rect 2 6851 153 6874
rect 2 6815 44 6851
rect 1 6814 101 6815
rect 1 6793 157 6814
rect 1 6775 119 6793
rect 137 6775 157 6793
rect 1 6771 157 6775
rect 96 6755 157 6771
rect 4774 6922 4794 6940
rect 4812 6922 4930 6940
rect 5152 6933 5209 6952
rect 5152 6930 5173 6933
rect 4774 6901 4930 6922
rect 4830 6900 4930 6901
rect 5058 6915 5173 6930
rect 5191 6915 5209 6933
rect 9830 6985 9891 7001
rect 9830 6981 9986 6985
rect 4887 6864 4929 6900
rect 4778 6841 4929 6864
rect 5058 6892 5209 6915
rect 5058 6856 5100 6892
rect 4778 6823 4796 6841
rect 4814 6826 4929 6841
rect 5057 6855 5157 6856
rect 5057 6834 5213 6855
rect 4814 6823 4835 6826
rect 4778 6804 4835 6823
rect 5057 6816 5175 6834
rect 5193 6816 5213 6834
rect 5057 6812 5213 6816
rect 5152 6796 5213 6812
rect 9830 6963 9850 6981
rect 9868 6963 9986 6981
rect 9830 6942 9986 6963
rect 9886 6941 9986 6942
rect 9943 6905 9985 6941
rect 9834 6882 9985 6905
rect 9834 6864 9852 6882
rect 9870 6867 9985 6882
rect 9870 6864 9891 6867
rect 9834 6845 9891 6864
rect 96 6663 153 6682
rect 96 6660 117 6663
rect 2 6645 117 6660
rect 135 6645 153 6663
rect 2 6622 153 6645
rect 4774 6714 4835 6730
rect 4774 6710 4930 6714
rect 2 6586 44 6622
rect 1 6585 101 6586
rect 1 6564 157 6585
rect 1 6546 119 6564
rect 137 6546 157 6564
rect 4774 6692 4794 6710
rect 4812 6692 4930 6710
rect 5152 6704 5209 6723
rect 5152 6701 5173 6704
rect 4774 6671 4930 6692
rect 4830 6670 4930 6671
rect 5058 6686 5173 6701
rect 5191 6686 5209 6704
rect 4887 6634 4929 6670
rect 1 6542 157 6546
rect 96 6526 157 6542
rect 4778 6611 4929 6634
rect 5058 6663 5209 6686
rect 9830 6755 9891 6771
rect 9830 6751 9986 6755
rect 5058 6627 5100 6663
rect 4778 6593 4796 6611
rect 4814 6596 4929 6611
rect 5057 6626 5157 6627
rect 5057 6605 5213 6626
rect 4814 6593 4835 6596
rect 4778 6574 4835 6593
rect 5057 6587 5175 6605
rect 5193 6587 5213 6605
rect 9830 6733 9850 6751
rect 9868 6733 9986 6751
rect 9830 6712 9986 6733
rect 9886 6711 9986 6712
rect 9943 6675 9985 6711
rect 5057 6583 5213 6587
rect 5152 6567 5213 6583
rect 9834 6652 9985 6675
rect 9834 6634 9852 6652
rect 9870 6637 9985 6652
rect 9870 6634 9891 6637
rect 9834 6615 9891 6634
rect 96 6433 153 6452
rect 96 6430 117 6433
rect 2 6415 117 6430
rect 135 6415 153 6433
rect 2 6392 153 6415
rect 2 6356 44 6392
rect 1 6355 101 6356
rect 1 6334 157 6355
rect 1 6316 119 6334
rect 137 6316 157 6334
rect 4774 6485 4835 6501
rect 4774 6481 4930 6485
rect 4774 6463 4794 6481
rect 4812 6463 4930 6481
rect 5152 6474 5209 6493
rect 5152 6471 5173 6474
rect 4774 6442 4930 6463
rect 4830 6441 4930 6442
rect 5058 6456 5173 6471
rect 5191 6456 5209 6474
rect 4887 6405 4929 6441
rect 4778 6382 4929 6405
rect 5058 6433 5209 6456
rect 5058 6397 5100 6433
rect 1 6312 157 6316
rect 96 6296 157 6312
rect 4778 6364 4796 6382
rect 4814 6367 4929 6382
rect 5057 6396 5157 6397
rect 5057 6375 5213 6396
rect 4814 6364 4835 6367
rect 4778 6345 4835 6364
rect 5057 6357 5175 6375
rect 5193 6357 5213 6375
rect 9830 6526 9891 6542
rect 9830 6522 9986 6526
rect 9830 6504 9850 6522
rect 9868 6504 9986 6522
rect 9830 6483 9986 6504
rect 9886 6482 9986 6483
rect 9943 6446 9985 6482
rect 9834 6423 9985 6446
rect 5057 6353 5213 6357
rect 5152 6337 5213 6353
rect 4774 6298 4835 6314
rect 4774 6294 4930 6298
rect 4774 6276 4794 6294
rect 4812 6276 4930 6294
rect 9834 6405 9852 6423
rect 9870 6408 9985 6423
rect 9870 6405 9891 6408
rect 9834 6386 9891 6405
rect 9830 6339 9891 6355
rect 9830 6335 9986 6339
rect 9830 6317 9850 6335
rect 9868 6317 9986 6335
rect 9830 6296 9986 6317
rect 9886 6295 9986 6296
rect 4774 6255 4930 6276
rect 4830 6254 4930 6255
rect 4887 6218 4929 6254
rect 4778 6195 4929 6218
rect 9943 6259 9985 6295
rect 9834 6236 9985 6259
rect 4778 6177 4796 6195
rect 4814 6180 4929 6195
rect 4814 6177 4835 6180
rect 4778 6158 4835 6177
rect 97 5976 154 5995
rect 97 5973 118 5976
rect 3 5958 118 5973
rect 136 5958 154 5976
rect 9834 6218 9852 6236
rect 9870 6221 9985 6236
rect 9870 6218 9891 6221
rect 9834 6199 9891 6218
rect 5153 6017 5210 6036
rect 5153 6014 5174 6017
rect 5059 5999 5174 6014
rect 5192 5999 5210 6017
rect 3 5935 154 5958
rect 3 5899 45 5935
rect 5059 5976 5210 5999
rect 5059 5940 5101 5976
rect 5058 5939 5158 5940
rect 5058 5918 5214 5939
rect 2 5898 102 5899
rect 2 5877 158 5898
rect 2 5859 120 5877
rect 138 5859 158 5877
rect 2 5855 158 5859
rect 97 5839 158 5855
rect 97 5789 154 5808
rect 97 5786 118 5789
rect 3 5771 118 5786
rect 136 5771 154 5789
rect 5058 5900 5176 5918
rect 5194 5900 5214 5918
rect 5058 5896 5214 5900
rect 5153 5880 5214 5896
rect 4775 5841 4836 5857
rect 4775 5837 4931 5841
rect 3 5748 154 5771
rect 3 5712 45 5748
rect 2 5711 102 5712
rect 2 5690 158 5711
rect 2 5672 120 5690
rect 138 5672 158 5690
rect 2 5668 158 5672
rect 97 5652 158 5668
rect 4775 5819 4795 5837
rect 4813 5819 4931 5837
rect 5153 5830 5210 5849
rect 5153 5827 5174 5830
rect 4775 5798 4931 5819
rect 4831 5797 4931 5798
rect 5059 5812 5174 5827
rect 5192 5812 5210 5830
rect 9831 5882 9892 5898
rect 9831 5878 9987 5882
rect 4888 5761 4930 5797
rect 4779 5738 4930 5761
rect 5059 5789 5210 5812
rect 5059 5753 5101 5789
rect 4779 5720 4797 5738
rect 4815 5723 4930 5738
rect 5058 5752 5158 5753
rect 5058 5731 5214 5752
rect 4815 5720 4836 5723
rect 4779 5701 4836 5720
rect 5058 5713 5176 5731
rect 5194 5713 5214 5731
rect 5058 5709 5214 5713
rect 5153 5693 5214 5709
rect 9831 5860 9851 5878
rect 9869 5860 9987 5878
rect 9831 5839 9987 5860
rect 9887 5838 9987 5839
rect 9944 5802 9986 5838
rect 9835 5779 9986 5802
rect 9835 5761 9853 5779
rect 9871 5764 9986 5779
rect 9871 5761 9892 5764
rect 9835 5742 9892 5761
rect 97 5560 154 5579
rect 97 5557 118 5560
rect 3 5542 118 5557
rect 136 5542 154 5560
rect 3 5519 154 5542
rect 4775 5611 4836 5627
rect 4775 5607 4931 5611
rect 3 5483 45 5519
rect 2 5482 102 5483
rect 2 5461 158 5482
rect 2 5443 120 5461
rect 138 5443 158 5461
rect 4775 5589 4795 5607
rect 4813 5589 4931 5607
rect 5153 5601 5210 5620
rect 5153 5598 5174 5601
rect 4775 5568 4931 5589
rect 4831 5567 4931 5568
rect 5059 5583 5174 5598
rect 5192 5583 5210 5601
rect 4888 5531 4930 5567
rect 2 5439 158 5443
rect 97 5423 158 5439
rect 4779 5508 4930 5531
rect 5059 5560 5210 5583
rect 9831 5652 9892 5668
rect 9831 5648 9987 5652
rect 5059 5524 5101 5560
rect 4779 5490 4797 5508
rect 4815 5493 4930 5508
rect 5058 5523 5158 5524
rect 5058 5502 5214 5523
rect 4815 5490 4836 5493
rect 4779 5471 4836 5490
rect 5058 5484 5176 5502
rect 5194 5484 5214 5502
rect 9831 5630 9851 5648
rect 9869 5630 9987 5648
rect 9831 5609 9987 5630
rect 9887 5608 9987 5609
rect 9944 5572 9986 5608
rect 5058 5480 5214 5484
rect 5153 5464 5214 5480
rect 9835 5549 9986 5572
rect 9835 5531 9853 5549
rect 9871 5534 9986 5549
rect 9871 5531 9892 5534
rect 9835 5512 9892 5531
rect 97 5330 154 5349
rect 97 5327 118 5330
rect 3 5312 118 5327
rect 136 5312 154 5330
rect 3 5289 154 5312
rect 3 5253 45 5289
rect 2 5252 102 5253
rect 2 5231 158 5252
rect 2 5213 120 5231
rect 138 5213 158 5231
rect 4775 5382 4836 5398
rect 4775 5378 4931 5382
rect 4775 5360 4795 5378
rect 4813 5360 4931 5378
rect 5153 5371 5210 5390
rect 5153 5368 5174 5371
rect 4775 5339 4931 5360
rect 4831 5338 4931 5339
rect 5059 5353 5174 5368
rect 5192 5353 5210 5371
rect 4888 5302 4930 5338
rect 4779 5279 4930 5302
rect 5059 5330 5210 5353
rect 5059 5294 5101 5330
rect 2 5209 158 5213
rect 97 5193 158 5209
rect 4779 5261 4797 5279
rect 4815 5264 4930 5279
rect 5058 5293 5158 5294
rect 5058 5272 5214 5293
rect 4815 5261 4836 5264
rect 4779 5242 4836 5261
rect 5058 5254 5176 5272
rect 5194 5254 5214 5272
rect 9831 5423 9892 5439
rect 9831 5419 9987 5423
rect 9831 5401 9851 5419
rect 9869 5401 9987 5419
rect 9831 5380 9987 5401
rect 9887 5379 9987 5380
rect 9944 5343 9986 5379
rect 9835 5320 9986 5343
rect 5058 5250 5214 5254
rect 5153 5234 5214 5250
rect 4775 5195 4836 5211
rect 4775 5191 4931 5195
rect 4775 5173 4795 5191
rect 4813 5173 4931 5191
rect 9835 5302 9853 5320
rect 9871 5305 9986 5320
rect 9871 5302 9892 5305
rect 9835 5283 9892 5302
rect 9831 5236 9892 5252
rect 9831 5232 9987 5236
rect 9831 5214 9851 5232
rect 9869 5214 9987 5232
rect 4775 5152 4931 5173
rect 4831 5151 4931 5152
rect 4888 5115 4930 5151
rect 9831 5193 9987 5214
rect 9887 5192 9987 5193
rect 4779 5092 4930 5115
rect 4779 5074 4797 5092
rect 4815 5077 4930 5092
rect 4815 5074 4836 5077
rect 4779 5055 4836 5074
rect 9944 5156 9986 5192
rect 9835 5133 9986 5156
rect 9835 5115 9853 5133
rect 9871 5118 9986 5133
rect 9871 5115 9892 5118
rect 9835 5096 9892 5115
rect 97 4873 154 4892
rect 97 4870 118 4873
rect 3 4855 118 4870
rect 136 4855 154 4873
rect 3 4832 154 4855
rect 3 4796 45 4832
rect 5153 4914 5210 4933
rect 5153 4911 5174 4914
rect 5059 4896 5174 4911
rect 5192 4896 5210 4914
rect 5059 4873 5210 4896
rect 2 4795 102 4796
rect 2 4774 158 4795
rect 5059 4837 5101 4873
rect 5058 4836 5158 4837
rect 5058 4815 5214 4836
rect 2 4756 120 4774
rect 138 4756 158 4774
rect 2 4752 158 4756
rect 97 4736 158 4752
rect 97 4686 154 4705
rect 97 4683 118 4686
rect 3 4668 118 4683
rect 136 4668 154 4686
rect 5058 4797 5176 4815
rect 5194 4797 5214 4815
rect 5058 4793 5214 4797
rect 5153 4777 5214 4793
rect 4775 4738 4836 4754
rect 4775 4734 4931 4738
rect 3 4645 154 4668
rect 3 4609 45 4645
rect 2 4608 102 4609
rect 2 4587 158 4608
rect 2 4569 120 4587
rect 138 4569 158 4587
rect 2 4565 158 4569
rect 97 4549 158 4565
rect 4775 4716 4795 4734
rect 4813 4716 4931 4734
rect 5153 4727 5210 4746
rect 5153 4724 5174 4727
rect 4775 4695 4931 4716
rect 4831 4694 4931 4695
rect 5059 4709 5174 4724
rect 5192 4709 5210 4727
rect 9831 4779 9892 4795
rect 9831 4775 9987 4779
rect 4888 4658 4930 4694
rect 4779 4635 4930 4658
rect 5059 4686 5210 4709
rect 5059 4650 5101 4686
rect 4779 4617 4797 4635
rect 4815 4620 4930 4635
rect 5058 4649 5158 4650
rect 5058 4628 5214 4649
rect 4815 4617 4836 4620
rect 4779 4598 4836 4617
rect 5058 4610 5176 4628
rect 5194 4610 5214 4628
rect 5058 4606 5214 4610
rect 5153 4590 5214 4606
rect 9831 4757 9851 4775
rect 9869 4757 9987 4775
rect 9831 4736 9987 4757
rect 9887 4735 9987 4736
rect 9944 4699 9986 4735
rect 9835 4676 9986 4699
rect 9835 4658 9853 4676
rect 9871 4661 9986 4676
rect 9871 4658 9892 4661
rect 9835 4639 9892 4658
rect 97 4457 154 4476
rect 97 4454 118 4457
rect 3 4439 118 4454
rect 136 4439 154 4457
rect 3 4416 154 4439
rect 4775 4508 4836 4524
rect 4775 4504 4931 4508
rect 3 4380 45 4416
rect 2 4379 102 4380
rect 2 4358 158 4379
rect 2 4340 120 4358
rect 138 4340 158 4358
rect 4775 4486 4795 4504
rect 4813 4486 4931 4504
rect 5153 4498 5210 4517
rect 5153 4495 5174 4498
rect 4775 4465 4931 4486
rect 4831 4464 4931 4465
rect 5059 4480 5174 4495
rect 5192 4480 5210 4498
rect 4888 4428 4930 4464
rect 2 4336 158 4340
rect 97 4320 158 4336
rect 4779 4405 4930 4428
rect 5059 4457 5210 4480
rect 9831 4549 9892 4565
rect 9831 4545 9987 4549
rect 5059 4421 5101 4457
rect 4779 4387 4797 4405
rect 4815 4390 4930 4405
rect 5058 4420 5158 4421
rect 5058 4399 5214 4420
rect 4815 4387 4836 4390
rect 4779 4368 4836 4387
rect 5058 4381 5176 4399
rect 5194 4381 5214 4399
rect 9831 4527 9851 4545
rect 9869 4527 9987 4545
rect 9831 4506 9987 4527
rect 9887 4505 9987 4506
rect 9944 4469 9986 4505
rect 5058 4377 5214 4381
rect 5153 4361 5214 4377
rect 9835 4446 9986 4469
rect 9835 4428 9853 4446
rect 9871 4431 9986 4446
rect 9871 4428 9892 4431
rect 9835 4409 9892 4428
rect 97 4227 154 4246
rect 97 4224 118 4227
rect 3 4209 118 4224
rect 136 4209 154 4227
rect 3 4186 154 4209
rect 3 4150 45 4186
rect 2 4149 102 4150
rect 2 4128 158 4149
rect 2 4110 120 4128
rect 138 4110 158 4128
rect 4775 4279 4836 4295
rect 4775 4275 4931 4279
rect 4775 4257 4795 4275
rect 4813 4257 4931 4275
rect 5153 4268 5210 4287
rect 5153 4265 5174 4268
rect 4775 4236 4931 4257
rect 4831 4235 4931 4236
rect 5059 4250 5174 4265
rect 5192 4250 5210 4268
rect 4888 4199 4930 4235
rect 4779 4176 4930 4199
rect 5059 4227 5210 4250
rect 5059 4191 5101 4227
rect 2 4106 158 4110
rect 97 4090 158 4106
rect 4779 4158 4797 4176
rect 4815 4161 4930 4176
rect 5058 4190 5158 4191
rect 5058 4169 5214 4190
rect 4815 4158 4836 4161
rect 4779 4139 4836 4158
rect 5058 4151 5176 4169
rect 5194 4151 5214 4169
rect 9831 4320 9892 4336
rect 9831 4316 9987 4320
rect 9831 4298 9851 4316
rect 9869 4298 9987 4316
rect 9831 4277 9987 4298
rect 9887 4276 9987 4277
rect 9944 4240 9986 4276
rect 9835 4217 9986 4240
rect 5058 4147 5214 4151
rect 5153 4131 5214 4147
rect 4775 4092 4836 4108
rect 4775 4088 4931 4092
rect 4775 4070 4795 4088
rect 4813 4070 4931 4088
rect 9835 4199 9853 4217
rect 9871 4202 9986 4217
rect 9871 4199 9892 4202
rect 9835 4180 9892 4199
rect 9831 4133 9892 4149
rect 9831 4129 9987 4133
rect 9831 4111 9851 4129
rect 9869 4111 9987 4129
rect 9831 4090 9987 4111
rect 9887 4089 9987 4090
rect 4775 4049 4931 4070
rect 4831 4048 4931 4049
rect 4888 4012 4930 4048
rect 4779 3989 4930 4012
rect 9944 4053 9986 4089
rect 9835 4030 9986 4053
rect 4779 3971 4797 3989
rect 4815 3974 4930 3989
rect 4815 3971 4836 3974
rect 4779 3952 4836 3971
rect 98 3770 155 3789
rect 98 3767 119 3770
rect 4 3752 119 3767
rect 137 3752 155 3770
rect 9835 4012 9853 4030
rect 9871 4015 9986 4030
rect 9871 4012 9892 4015
rect 9835 3993 9892 4012
rect 5154 3811 5211 3830
rect 5154 3808 5175 3811
rect 5060 3793 5175 3808
rect 5193 3793 5211 3811
rect 4 3729 155 3752
rect 4 3693 46 3729
rect 5060 3770 5211 3793
rect 5060 3734 5102 3770
rect 5059 3733 5159 3734
rect 5059 3712 5215 3733
rect 3 3692 103 3693
rect 3 3671 159 3692
rect 3 3653 121 3671
rect 139 3653 159 3671
rect 3 3649 159 3653
rect 98 3633 159 3649
rect 98 3583 155 3602
rect 98 3580 119 3583
rect 4 3565 119 3580
rect 137 3565 155 3583
rect 5059 3694 5177 3712
rect 5195 3694 5215 3712
rect 5059 3690 5215 3694
rect 5154 3674 5215 3690
rect 4776 3635 4837 3651
rect 4776 3631 4932 3635
rect 4 3542 155 3565
rect 4 3506 46 3542
rect 3 3505 103 3506
rect 3 3484 159 3505
rect 3 3466 121 3484
rect 139 3466 159 3484
rect 3 3462 159 3466
rect 98 3446 159 3462
rect 4776 3613 4796 3631
rect 4814 3613 4932 3631
rect 5154 3624 5211 3643
rect 5154 3621 5175 3624
rect 4776 3592 4932 3613
rect 4832 3591 4932 3592
rect 5060 3606 5175 3621
rect 5193 3606 5211 3624
rect 9832 3676 9893 3692
rect 9832 3672 9988 3676
rect 4889 3555 4931 3591
rect 4780 3532 4931 3555
rect 5060 3583 5211 3606
rect 5060 3547 5102 3583
rect 4780 3514 4798 3532
rect 4816 3517 4931 3532
rect 5059 3546 5159 3547
rect 5059 3525 5215 3546
rect 4816 3514 4837 3517
rect 4780 3495 4837 3514
rect 5059 3507 5177 3525
rect 5195 3507 5215 3525
rect 5059 3503 5215 3507
rect 5154 3487 5215 3503
rect 9832 3654 9852 3672
rect 9870 3654 9988 3672
rect 9832 3633 9988 3654
rect 9888 3632 9988 3633
rect 9945 3596 9987 3632
rect 9836 3573 9987 3596
rect 9836 3555 9854 3573
rect 9872 3558 9987 3573
rect 9872 3555 9893 3558
rect 9836 3536 9893 3555
rect 98 3354 155 3373
rect 98 3351 119 3354
rect 4 3336 119 3351
rect 137 3336 155 3354
rect 4 3313 155 3336
rect 4776 3405 4837 3421
rect 4776 3401 4932 3405
rect 4 3277 46 3313
rect 3 3276 103 3277
rect 3 3255 159 3276
rect 3 3237 121 3255
rect 139 3237 159 3255
rect 4776 3383 4796 3401
rect 4814 3383 4932 3401
rect 5154 3395 5211 3414
rect 5154 3392 5175 3395
rect 4776 3362 4932 3383
rect 4832 3361 4932 3362
rect 5060 3377 5175 3392
rect 5193 3377 5211 3395
rect 4889 3325 4931 3361
rect 3 3233 159 3237
rect 98 3217 159 3233
rect 4780 3302 4931 3325
rect 5060 3354 5211 3377
rect 9832 3446 9893 3462
rect 9832 3442 9988 3446
rect 5060 3318 5102 3354
rect 4780 3284 4798 3302
rect 4816 3287 4931 3302
rect 5059 3317 5159 3318
rect 5059 3296 5215 3317
rect 4816 3284 4837 3287
rect 4780 3265 4837 3284
rect 5059 3278 5177 3296
rect 5195 3278 5215 3296
rect 9832 3424 9852 3442
rect 9870 3424 9988 3442
rect 9832 3403 9988 3424
rect 9888 3402 9988 3403
rect 9945 3366 9987 3402
rect 5059 3274 5215 3278
rect 5154 3258 5215 3274
rect 9836 3343 9987 3366
rect 9836 3325 9854 3343
rect 9872 3328 9987 3343
rect 9872 3325 9893 3328
rect 9836 3306 9893 3325
rect 98 3124 155 3143
rect 98 3121 119 3124
rect 4 3106 119 3121
rect 137 3106 155 3124
rect 4 3083 155 3106
rect 4 3047 46 3083
rect 3 3046 103 3047
rect 3 3025 159 3046
rect 3 3007 121 3025
rect 139 3007 159 3025
rect 4776 3176 4837 3192
rect 4776 3172 4932 3176
rect 4776 3154 4796 3172
rect 4814 3154 4932 3172
rect 5154 3165 5211 3184
rect 5154 3162 5175 3165
rect 4776 3133 4932 3154
rect 4832 3132 4932 3133
rect 5060 3147 5175 3162
rect 5193 3147 5211 3165
rect 4889 3096 4931 3132
rect 4780 3073 4931 3096
rect 5060 3124 5211 3147
rect 5060 3088 5102 3124
rect 3 3003 159 3007
rect 98 2987 159 3003
rect 4780 3055 4798 3073
rect 4816 3058 4931 3073
rect 5059 3087 5159 3088
rect 5059 3066 5215 3087
rect 4816 3055 4837 3058
rect 4780 3036 4837 3055
rect 5059 3048 5177 3066
rect 5195 3048 5215 3066
rect 9832 3217 9893 3233
rect 9832 3213 9988 3217
rect 9832 3195 9852 3213
rect 9870 3195 9988 3213
rect 9832 3174 9988 3195
rect 9888 3173 9988 3174
rect 9945 3137 9987 3173
rect 9836 3114 9987 3137
rect 5059 3044 5215 3048
rect 5154 3028 5215 3044
rect 4776 2989 4837 3005
rect 4776 2985 4932 2989
rect 4776 2967 4796 2985
rect 4814 2967 4932 2985
rect 9836 3096 9854 3114
rect 9872 3099 9987 3114
rect 9872 3096 9893 3099
rect 9836 3077 9893 3096
rect 9832 3030 9893 3046
rect 9832 3026 9988 3030
rect 9832 3008 9852 3026
rect 9870 3008 9988 3026
rect 9832 2987 9988 3008
rect 9888 2986 9988 2987
rect 4776 2946 4932 2967
rect 4832 2945 4932 2946
rect 4889 2909 4931 2945
rect 4780 2886 4931 2909
rect 4780 2868 4798 2886
rect 4816 2871 4931 2886
rect 9945 2950 9987 2986
rect 9836 2927 9987 2950
rect 9836 2909 9854 2927
rect 9872 2912 9987 2927
rect 9872 2909 9893 2912
rect 4816 2868 4837 2871
rect 4780 2849 4837 2868
rect 9836 2890 9893 2909
rect 98 2667 155 2686
rect 5154 2708 5211 2727
rect 5154 2705 5175 2708
rect 98 2664 119 2667
rect 4 2649 119 2664
rect 137 2649 155 2667
rect 4 2626 155 2649
rect 4 2590 46 2626
rect 5060 2690 5175 2705
rect 5193 2690 5211 2708
rect 5060 2667 5211 2690
rect 5060 2631 5102 2667
rect 5059 2630 5159 2631
rect 5059 2609 5215 2630
rect 3 2589 103 2590
rect 3 2568 159 2589
rect 3 2550 121 2568
rect 139 2550 159 2568
rect 3 2546 159 2550
rect 98 2530 159 2546
rect 98 2480 155 2499
rect 98 2477 119 2480
rect 4 2462 119 2477
rect 137 2462 155 2480
rect 5059 2591 5177 2609
rect 5195 2591 5215 2609
rect 5059 2587 5215 2591
rect 5154 2571 5215 2587
rect 4776 2532 4837 2548
rect 4776 2528 4932 2532
rect 4 2439 155 2462
rect 4 2403 46 2439
rect 3 2402 103 2403
rect 3 2381 159 2402
rect 3 2363 121 2381
rect 139 2363 159 2381
rect 3 2359 159 2363
rect 98 2343 159 2359
rect 4776 2510 4796 2528
rect 4814 2510 4932 2528
rect 5154 2521 5211 2540
rect 5154 2518 5175 2521
rect 4776 2489 4932 2510
rect 4832 2488 4932 2489
rect 5060 2503 5175 2518
rect 5193 2503 5211 2521
rect 9832 2573 9893 2589
rect 9832 2569 9988 2573
rect 4889 2452 4931 2488
rect 4780 2429 4931 2452
rect 5060 2480 5211 2503
rect 5060 2444 5102 2480
rect 4780 2411 4798 2429
rect 4816 2414 4931 2429
rect 5059 2443 5159 2444
rect 5059 2422 5215 2443
rect 4816 2411 4837 2414
rect 4780 2392 4837 2411
rect 5059 2404 5177 2422
rect 5195 2404 5215 2422
rect 5059 2400 5215 2404
rect 5154 2384 5215 2400
rect 9832 2551 9852 2569
rect 9870 2551 9988 2569
rect 9832 2530 9988 2551
rect 9888 2529 9988 2530
rect 9945 2493 9987 2529
rect 9836 2470 9987 2493
rect 9836 2452 9854 2470
rect 9872 2455 9987 2470
rect 9872 2452 9893 2455
rect 9836 2433 9893 2452
rect 98 2251 155 2270
rect 98 2248 119 2251
rect 4 2233 119 2248
rect 137 2233 155 2251
rect 4 2210 155 2233
rect 4776 2302 4837 2318
rect 4776 2298 4932 2302
rect 4 2174 46 2210
rect 3 2173 103 2174
rect 3 2152 159 2173
rect 3 2134 121 2152
rect 139 2134 159 2152
rect 4776 2280 4796 2298
rect 4814 2280 4932 2298
rect 5154 2292 5211 2311
rect 5154 2289 5175 2292
rect 4776 2259 4932 2280
rect 4832 2258 4932 2259
rect 5060 2274 5175 2289
rect 5193 2274 5211 2292
rect 4889 2222 4931 2258
rect 3 2130 159 2134
rect 98 2114 159 2130
rect 4780 2199 4931 2222
rect 5060 2251 5211 2274
rect 9832 2343 9893 2359
rect 9832 2339 9988 2343
rect 5060 2215 5102 2251
rect 4780 2181 4798 2199
rect 4816 2184 4931 2199
rect 5059 2214 5159 2215
rect 5059 2193 5215 2214
rect 4816 2181 4837 2184
rect 4780 2162 4837 2181
rect 5059 2175 5177 2193
rect 5195 2175 5215 2193
rect 9832 2321 9852 2339
rect 9870 2321 9988 2339
rect 9832 2300 9988 2321
rect 9888 2299 9988 2300
rect 9945 2263 9987 2299
rect 5059 2171 5215 2175
rect 5154 2155 5215 2171
rect 9836 2240 9987 2263
rect 9836 2222 9854 2240
rect 9872 2225 9987 2240
rect 9872 2222 9893 2225
rect 9836 2203 9893 2222
rect 98 2021 155 2040
rect 98 2018 119 2021
rect 4 2003 119 2018
rect 137 2003 155 2021
rect 4 1980 155 2003
rect 4 1944 46 1980
rect 3 1943 103 1944
rect 3 1922 159 1943
rect 3 1904 121 1922
rect 139 1904 159 1922
rect 4776 2073 4837 2089
rect 4776 2069 4932 2073
rect 4776 2051 4796 2069
rect 4814 2051 4932 2069
rect 5154 2062 5211 2081
rect 5154 2059 5175 2062
rect 4776 2030 4932 2051
rect 4832 2029 4932 2030
rect 5060 2044 5175 2059
rect 5193 2044 5211 2062
rect 4889 1993 4931 2029
rect 4780 1970 4931 1993
rect 5060 2021 5211 2044
rect 5060 1985 5102 2021
rect 3 1900 159 1904
rect 98 1884 159 1900
rect 4780 1952 4798 1970
rect 4816 1955 4931 1970
rect 5059 1984 5159 1985
rect 5059 1963 5215 1984
rect 4816 1952 4837 1955
rect 4780 1933 4837 1952
rect 5059 1945 5177 1963
rect 5195 1945 5215 1963
rect 9832 2114 9893 2130
rect 9832 2110 9988 2114
rect 9832 2092 9852 2110
rect 9870 2092 9988 2110
rect 9832 2071 9988 2092
rect 9888 2070 9988 2071
rect 9945 2034 9987 2070
rect 9836 2011 9987 2034
rect 5059 1941 5215 1945
rect 5154 1925 5215 1941
rect 4776 1886 4837 1902
rect 4776 1882 4932 1886
rect 4776 1864 4796 1882
rect 4814 1864 4932 1882
rect 9836 1993 9854 2011
rect 9872 1996 9987 2011
rect 9872 1993 9893 1996
rect 9836 1974 9893 1993
rect 9832 1927 9893 1943
rect 9832 1923 9988 1927
rect 9832 1905 9852 1923
rect 9870 1905 9988 1923
rect 9832 1884 9988 1905
rect 9888 1883 9988 1884
rect 4776 1843 4932 1864
rect 4832 1842 4932 1843
rect 4889 1806 4931 1842
rect 4780 1783 4931 1806
rect 9945 1847 9987 1883
rect 9836 1824 9987 1847
rect 4780 1765 4798 1783
rect 4816 1768 4931 1783
rect 4816 1765 4837 1768
rect 4780 1746 4837 1765
rect 99 1564 156 1583
rect 99 1561 120 1564
rect 5 1546 120 1561
rect 138 1546 156 1564
rect 9836 1806 9854 1824
rect 9872 1809 9987 1824
rect 9872 1806 9893 1809
rect 9836 1787 9893 1806
rect 5155 1605 5212 1624
rect 5155 1602 5176 1605
rect 5061 1587 5176 1602
rect 5194 1587 5212 1605
rect 5 1523 156 1546
rect 5 1487 47 1523
rect 5061 1564 5212 1587
rect 5061 1528 5103 1564
rect 5060 1527 5160 1528
rect 5060 1506 5216 1527
rect 4 1486 104 1487
rect 4 1465 160 1486
rect 4 1447 122 1465
rect 140 1447 160 1465
rect 4 1443 160 1447
rect 99 1427 160 1443
rect 99 1377 156 1396
rect 99 1374 120 1377
rect 5 1359 120 1374
rect 138 1359 156 1377
rect 5060 1488 5178 1506
rect 5196 1488 5216 1506
rect 5060 1484 5216 1488
rect 5155 1468 5216 1484
rect 4777 1429 4838 1445
rect 4777 1425 4933 1429
rect 5 1336 156 1359
rect 5 1300 47 1336
rect 4 1299 104 1300
rect 4 1278 160 1299
rect 4 1260 122 1278
rect 140 1260 160 1278
rect 4 1256 160 1260
rect 99 1240 160 1256
rect 4777 1407 4797 1425
rect 4815 1407 4933 1425
rect 5155 1418 5212 1437
rect 5155 1415 5176 1418
rect 4777 1386 4933 1407
rect 4833 1385 4933 1386
rect 5061 1400 5176 1415
rect 5194 1400 5212 1418
rect 9833 1470 9894 1486
rect 9833 1466 9989 1470
rect 4890 1349 4932 1385
rect 4781 1326 4932 1349
rect 5061 1377 5212 1400
rect 5061 1341 5103 1377
rect 4781 1308 4799 1326
rect 4817 1311 4932 1326
rect 5060 1340 5160 1341
rect 5060 1319 5216 1340
rect 4817 1308 4838 1311
rect 4781 1289 4838 1308
rect 5060 1301 5178 1319
rect 5196 1301 5216 1319
rect 5060 1297 5216 1301
rect 5155 1281 5216 1297
rect 9833 1448 9853 1466
rect 9871 1448 9989 1466
rect 9833 1427 9989 1448
rect 9889 1426 9989 1427
rect 9946 1390 9988 1426
rect 9837 1367 9988 1390
rect 9837 1349 9855 1367
rect 9873 1352 9988 1367
rect 9873 1349 9894 1352
rect 9837 1330 9894 1349
rect 99 1148 156 1167
rect 99 1145 120 1148
rect 5 1130 120 1145
rect 138 1130 156 1148
rect 5 1107 156 1130
rect 4777 1199 4838 1215
rect 4777 1195 4933 1199
rect 5 1071 47 1107
rect 4 1070 104 1071
rect 4 1049 160 1070
rect 4 1031 122 1049
rect 140 1031 160 1049
rect 4777 1177 4797 1195
rect 4815 1177 4933 1195
rect 5155 1189 5212 1208
rect 5155 1186 5176 1189
rect 4777 1156 4933 1177
rect 4833 1155 4933 1156
rect 5061 1171 5176 1186
rect 5194 1171 5212 1189
rect 4890 1119 4932 1155
rect 4 1027 160 1031
rect 99 1011 160 1027
rect 4781 1096 4932 1119
rect 5061 1148 5212 1171
rect 9833 1240 9894 1256
rect 9833 1236 9989 1240
rect 5061 1112 5103 1148
rect 4781 1078 4799 1096
rect 4817 1081 4932 1096
rect 5060 1111 5160 1112
rect 5060 1090 5216 1111
rect 4817 1078 4838 1081
rect 4781 1059 4838 1078
rect 5060 1072 5178 1090
rect 5196 1072 5216 1090
rect 9833 1218 9853 1236
rect 9871 1218 9989 1236
rect 9833 1197 9989 1218
rect 9889 1196 9989 1197
rect 9946 1160 9988 1196
rect 5060 1068 5216 1072
rect 5155 1052 5216 1068
rect 9837 1137 9988 1160
rect 9837 1119 9855 1137
rect 9873 1122 9988 1137
rect 9873 1119 9894 1122
rect 9837 1100 9894 1119
rect 99 918 156 937
rect 99 915 120 918
rect 5 900 120 915
rect 138 900 156 918
rect 5 877 156 900
rect 5 841 47 877
rect 4 840 104 841
rect 4 819 160 840
rect 4 801 122 819
rect 140 801 160 819
rect 4777 970 4838 986
rect 4777 966 4933 970
rect 4777 948 4797 966
rect 4815 948 4933 966
rect 5155 959 5212 978
rect 5155 956 5176 959
rect 4777 927 4933 948
rect 4833 926 4933 927
rect 5061 941 5176 956
rect 5194 941 5212 959
rect 4890 890 4932 926
rect 4781 867 4932 890
rect 5061 918 5212 941
rect 5061 882 5103 918
rect 4 797 160 801
rect 99 781 160 797
rect 4781 849 4799 867
rect 4817 852 4932 867
rect 5060 881 5160 882
rect 5060 860 5216 881
rect 4817 849 4838 852
rect 4781 830 4838 849
rect 5060 842 5178 860
rect 5196 842 5216 860
rect 9833 1011 9894 1027
rect 9833 1007 9989 1011
rect 9833 989 9853 1007
rect 9871 989 9989 1007
rect 9833 968 9989 989
rect 9889 967 9989 968
rect 9946 931 9988 967
rect 9837 908 9988 931
rect 5060 838 5216 842
rect 5155 822 5216 838
rect 4777 783 4838 799
rect 4777 779 4933 783
rect 4777 761 4797 779
rect 4815 761 4933 779
rect 9837 890 9855 908
rect 9873 893 9988 908
rect 9873 890 9894 893
rect 9837 871 9894 890
rect 9833 824 9894 840
rect 9833 820 9989 824
rect 9833 802 9853 820
rect 9871 802 9989 820
rect 9833 781 9989 802
rect 9889 780 9989 781
rect 4777 740 4933 761
rect 4833 739 4933 740
rect 4890 703 4932 739
rect 9946 744 9988 780
rect 9837 721 9988 744
rect 4781 680 4932 703
rect 9837 703 9855 721
rect 9873 706 9988 721
rect 9873 703 9894 706
rect 4781 662 4799 680
rect 4817 665 4932 680
rect 9837 684 9894 703
rect 4817 662 4838 665
rect 4781 643 4838 662
<< locali >>
rect 9193 9468 9231 9470
rect 9193 9435 9879 9468
rect 4137 9427 4175 9429
rect 4780 9427 5205 9429
rect 4137 9396 5214 9427
rect 4137 9394 4386 9396
rect 4542 9394 5214 9396
rect 105 9287 144 9344
rect 3729 9306 3897 9307
rect 4137 9306 4175 9394
rect 4780 9393 5215 9394
rect 4783 9370 4823 9393
rect 5135 9389 5215 9393
rect 4400 9337 4512 9355
rect 4400 9336 4443 9337
rect 105 9285 153 9287
rect 105 9267 116 9285
rect 134 9267 153 9285
rect 3729 9283 4175 9306
rect 4401 9335 4443 9336
rect 4401 9315 4408 9335
rect 4427 9315 4443 9335
rect 4401 9307 4443 9315
rect 4471 9335 4512 9337
rect 4471 9315 4485 9335
rect 4504 9315 4512 9335
rect 4784 9326 4823 9370
rect 5157 9345 5215 9389
rect 5159 9331 5215 9345
rect 4471 9307 4512 9315
rect 4401 9301 4512 9307
rect 3729 9280 4173 9283
rect 3729 9278 3897 9280
rect 105 9258 153 9267
rect 106 9257 153 9258
rect 419 9262 529 9276
rect 419 9259 462 9262
rect 419 9254 423 9259
rect 341 9232 423 9254
rect 452 9232 462 9259
rect 490 9235 497 9262
rect 526 9254 529 9262
rect 526 9235 591 9254
rect 490 9232 591 9235
rect 341 9230 591 9232
rect 109 9194 146 9195
rect 105 9191 146 9194
rect 105 9186 147 9191
rect 105 9168 118 9186
rect 136 9168 147 9186
rect 105 9154 147 9168
rect 185 9154 232 9158
rect 105 9148 232 9154
rect 105 9119 193 9148
rect 222 9119 232 9148
rect 341 9151 378 9230
rect 419 9217 529 9230
rect 493 9161 524 9162
rect 341 9131 350 9151
rect 370 9131 378 9151
rect 341 9121 378 9131
rect 437 9151 524 9161
rect 437 9131 446 9151
rect 466 9131 524 9151
rect 437 9122 524 9131
rect 437 9121 474 9122
rect 105 9115 232 9119
rect 105 9098 144 9115
rect 185 9114 232 9115
rect 105 9080 116 9098
rect 134 9080 144 9098
rect 105 9071 144 9080
rect 106 9070 143 9071
rect 493 9069 524 9122
rect 554 9151 591 9230
rect 762 9227 1155 9247
rect 1175 9227 1178 9247
rect 762 9222 1178 9227
rect 762 9221 1103 9222
rect 706 9161 737 9162
rect 554 9131 563 9151
rect 583 9131 591 9151
rect 554 9121 591 9131
rect 650 9154 737 9161
rect 650 9151 711 9154
rect 650 9131 659 9151
rect 679 9134 711 9151
rect 732 9134 737 9154
rect 679 9131 737 9134
rect 650 9124 737 9131
rect 762 9151 799 9221
rect 1065 9220 1102 9221
rect 914 9161 950 9162
rect 762 9131 771 9151
rect 791 9131 799 9151
rect 650 9122 706 9124
rect 650 9121 687 9122
rect 762 9121 799 9131
rect 858 9151 1006 9161
rect 1106 9158 1202 9160
rect 858 9131 867 9151
rect 887 9131 977 9151
rect 997 9131 1006 9151
rect 858 9122 1006 9131
rect 1064 9151 1202 9158
rect 1064 9131 1073 9151
rect 1093 9131 1202 9151
rect 1064 9122 1202 9131
rect 858 9121 895 9122
rect 914 9070 950 9122
rect 969 9121 1006 9122
rect 1065 9121 1102 9122
rect 385 9068 426 9069
rect 277 9061 426 9068
rect 277 9041 395 9061
rect 415 9041 426 9061
rect 277 9033 426 9041
rect 493 9065 852 9069
rect 493 9060 815 9065
rect 493 9036 606 9060
rect 630 9041 815 9060
rect 839 9041 852 9065
rect 630 9036 852 9041
rect 493 9033 852 9036
rect 914 9033 949 9070
rect 1017 9067 1117 9070
rect 1017 9063 1084 9067
rect 1017 9037 1029 9063
rect 1055 9041 1084 9063
rect 1110 9041 1117 9067
rect 1055 9037 1117 9041
rect 1017 9033 1117 9037
rect 493 9012 524 9033
rect 914 9012 950 9033
rect 336 9011 373 9012
rect 110 9008 144 9009
rect 109 8999 146 9008
rect 109 8981 118 8999
rect 136 8981 146 8999
rect 109 8971 146 8981
rect 335 9002 373 9011
rect 335 8982 344 9002
rect 364 8982 373 9002
rect 335 8974 373 8982
rect 439 9006 524 9012
rect 549 9011 586 9012
rect 439 8986 447 9006
rect 467 8986 524 9006
rect 439 8978 524 8986
rect 548 9002 586 9011
rect 548 8982 557 9002
rect 577 8982 586 9002
rect 439 8977 475 8978
rect 548 8974 586 8982
rect 652 9006 737 9012
rect 757 9011 794 9012
rect 652 8986 660 9006
rect 680 9005 737 9006
rect 680 8986 709 9005
rect 652 8985 709 8986
rect 730 8985 737 9005
rect 652 8978 737 8985
rect 756 9002 794 9011
rect 756 8982 765 9002
rect 785 8982 794 9002
rect 652 8977 688 8978
rect 756 8974 794 8982
rect 860 9006 1004 9012
rect 860 8986 868 9006
rect 888 9005 976 9006
rect 888 8986 919 9005
rect 860 8985 919 8986
rect 944 8986 976 9005
rect 996 8986 1004 9006
rect 944 8985 1004 8986
rect 860 8978 1004 8985
rect 860 8977 896 8978
rect 968 8977 1004 8978
rect 1070 9011 1107 9012
rect 1070 9010 1108 9011
rect 1070 9002 1134 9010
rect 1070 8982 1079 9002
rect 1099 8988 1134 9002
rect 1154 8988 1157 9008
rect 1099 8983 1157 8988
rect 1099 8982 1134 8983
rect 110 8943 144 8971
rect 336 8945 373 8974
rect 337 8943 373 8945
rect 549 8943 586 8974
rect 110 8942 282 8943
rect 110 8910 296 8942
rect 337 8921 586 8943
rect 757 8942 794 8974
rect 1070 8970 1134 8982
rect 1174 8944 1201 9122
rect 3729 9100 3756 9278
rect 3796 9240 3860 9252
rect 4136 9248 4173 9280
rect 4344 9279 4593 9301
rect 4344 9248 4381 9279
rect 4557 9277 4593 9279
rect 4557 9248 4594 9277
rect 3796 9239 3831 9240
rect 3773 9234 3831 9239
rect 3773 9214 3776 9234
rect 3796 9220 3831 9234
rect 3851 9220 3860 9240
rect 3796 9212 3860 9220
rect 3822 9211 3860 9212
rect 3823 9210 3860 9211
rect 3926 9244 3962 9245
rect 4034 9244 4070 9245
rect 3926 9239 4070 9244
rect 3926 9236 3988 9239
rect 3926 9216 3934 9236
rect 3954 9219 3988 9236
rect 4011 9236 4070 9239
rect 4011 9219 4042 9236
rect 3954 9216 4042 9219
rect 4062 9216 4070 9236
rect 3926 9210 4070 9216
rect 4136 9240 4174 9248
rect 4242 9244 4278 9245
rect 4136 9220 4145 9240
rect 4165 9220 4174 9240
rect 4136 9211 4174 9220
rect 4193 9237 4278 9244
rect 4193 9217 4200 9237
rect 4221 9236 4278 9237
rect 4221 9217 4250 9236
rect 4193 9216 4250 9217
rect 4270 9216 4278 9236
rect 4136 9210 4173 9211
rect 4193 9210 4278 9216
rect 4344 9240 4382 9248
rect 4455 9244 4491 9245
rect 4344 9220 4353 9240
rect 4373 9220 4382 9240
rect 4344 9211 4382 9220
rect 4406 9236 4491 9244
rect 4406 9216 4463 9236
rect 4483 9216 4491 9236
rect 4344 9210 4381 9211
rect 4406 9210 4491 9216
rect 4557 9240 4595 9248
rect 4557 9220 4566 9240
rect 4586 9220 4595 9240
rect 4557 9211 4595 9220
rect 4557 9210 4594 9211
rect 3980 9189 4016 9210
rect 4406 9189 4437 9210
rect 3813 9185 3913 9189
rect 3813 9181 3875 9185
rect 3813 9155 3820 9181
rect 3846 9159 3875 9181
rect 3901 9159 3913 9185
rect 3846 9155 3913 9159
rect 3813 9152 3913 9155
rect 3981 9152 4016 9189
rect 4078 9186 4437 9189
rect 4078 9181 4300 9186
rect 4078 9157 4091 9181
rect 4115 9162 4300 9181
rect 4324 9162 4437 9186
rect 4115 9157 4437 9162
rect 4078 9153 4437 9157
rect 4504 9181 4653 9189
rect 4504 9161 4515 9181
rect 4535 9161 4653 9181
rect 4504 9154 4653 9161
rect 4504 9153 4545 9154
rect 3828 9100 3865 9101
rect 3924 9100 3961 9101
rect 3980 9100 4016 9152
rect 4035 9100 4072 9101
rect 3728 9091 3866 9100
rect 3728 9071 3837 9091
rect 3857 9071 3866 9091
rect 3728 9064 3866 9071
rect 3924 9091 4072 9100
rect 3924 9071 3933 9091
rect 3953 9071 4043 9091
rect 4063 9071 4072 9091
rect 3728 9062 3824 9064
rect 3924 9061 4072 9071
rect 4131 9091 4168 9101
rect 4243 9100 4280 9101
rect 4224 9098 4280 9100
rect 4131 9071 4139 9091
rect 4159 9071 4168 9091
rect 3980 9060 4016 9061
rect 1357 9018 1467 9032
rect 1357 9015 1400 9018
rect 1357 9010 1361 9015
rect 1033 8942 1201 8944
rect 757 8936 1201 8942
rect 110 8878 144 8910
rect 106 8869 144 8878
rect 106 8851 116 8869
rect 134 8851 144 8869
rect 106 8845 144 8851
rect 262 8847 296 8910
rect 418 8915 529 8921
rect 418 8907 459 8915
rect 418 8887 426 8907
rect 445 8887 459 8907
rect 418 8885 459 8887
rect 487 8907 529 8915
rect 487 8887 503 8907
rect 522 8887 529 8907
rect 487 8885 529 8887
rect 418 8870 529 8885
rect 756 8916 1201 8936
rect 756 8847 794 8916
rect 1033 8915 1201 8916
rect 1279 8988 1361 9010
rect 1390 8988 1400 9015
rect 1428 8991 1435 9018
rect 1464 9010 1467 9018
rect 3462 9027 3573 9042
rect 3462 9025 3504 9027
rect 1464 8991 1529 9010
rect 1428 8988 1529 8991
rect 1279 8986 1529 8988
rect 1279 8907 1316 8986
rect 1357 8973 1467 8986
rect 1431 8917 1462 8918
rect 1279 8887 1288 8907
rect 1308 8887 1316 8907
rect 1279 8877 1316 8887
rect 1375 8907 1462 8917
rect 1375 8887 1384 8907
rect 1404 8887 1462 8907
rect 1375 8878 1462 8887
rect 1375 8877 1412 8878
rect 106 8841 143 8845
rect 262 8836 794 8847
rect 261 8820 794 8836
rect 1431 8825 1462 8878
rect 1492 8907 1529 8986
rect 1700 8983 2093 9003
rect 2113 8983 2116 9003
rect 3195 8998 3236 9007
rect 1700 8978 2116 8983
rect 2790 8996 2958 8997
rect 3195 8996 3204 8998
rect 1700 8977 2041 8978
rect 1644 8917 1675 8918
rect 1492 8887 1501 8907
rect 1521 8887 1529 8907
rect 1492 8877 1529 8887
rect 1588 8910 1675 8917
rect 1588 8907 1649 8910
rect 1588 8887 1597 8907
rect 1617 8890 1649 8907
rect 1670 8890 1675 8910
rect 1617 8887 1675 8890
rect 1588 8880 1675 8887
rect 1700 8907 1737 8977
rect 2003 8976 2040 8977
rect 2790 8976 3204 8996
rect 3230 8976 3236 8998
rect 3462 9005 3469 9025
rect 3488 9005 3504 9025
rect 3462 8997 3504 9005
rect 3532 9025 3573 9027
rect 3532 9005 3546 9025
rect 3565 9005 3573 9025
rect 3532 8997 3573 9005
rect 3828 9001 3865 9002
rect 4131 9001 4168 9071
rect 4193 9091 4280 9098
rect 4193 9088 4251 9091
rect 4193 9068 4198 9088
rect 4219 9071 4251 9088
rect 4271 9071 4280 9091
rect 4219 9068 4280 9071
rect 4193 9061 4280 9068
rect 4339 9091 4376 9101
rect 4339 9071 4347 9091
rect 4367 9071 4376 9091
rect 4193 9060 4224 9061
rect 3827 9000 4168 9001
rect 3462 8991 3573 8997
rect 3752 8995 4168 9000
rect 2790 8970 3236 8976
rect 2790 8968 2958 8970
rect 1852 8917 1888 8918
rect 1700 8887 1709 8907
rect 1729 8887 1737 8907
rect 1588 8878 1644 8880
rect 1588 8877 1625 8878
rect 1700 8877 1737 8887
rect 1796 8907 1944 8917
rect 2044 8914 2140 8916
rect 1796 8887 1805 8907
rect 1825 8887 1915 8907
rect 1935 8887 1944 8907
rect 1796 8878 1944 8887
rect 2002 8907 2140 8914
rect 2002 8887 2011 8907
rect 2031 8887 2140 8907
rect 2002 8878 2140 8887
rect 1796 8877 1833 8878
rect 1852 8826 1888 8878
rect 1907 8877 1944 8878
rect 2003 8877 2040 8878
rect 1323 8824 1364 8825
rect 261 8819 775 8820
rect 1215 8817 1364 8824
rect 1215 8797 1333 8817
rect 1353 8797 1364 8817
rect 1215 8789 1364 8797
rect 1431 8821 1790 8825
rect 1431 8816 1753 8821
rect 1431 8792 1544 8816
rect 1568 8797 1753 8816
rect 1777 8797 1790 8821
rect 1568 8792 1790 8797
rect 1431 8789 1790 8792
rect 1852 8789 1887 8826
rect 1955 8823 2055 8826
rect 1955 8819 2022 8823
rect 1955 8793 1967 8819
rect 1993 8797 2022 8819
rect 2048 8797 2055 8823
rect 1993 8793 2055 8797
rect 1955 8789 2055 8793
rect 109 8778 146 8779
rect 107 8770 147 8778
rect 107 8752 118 8770
rect 136 8752 147 8770
rect 1431 8768 1462 8789
rect 1852 8768 1888 8789
rect 1274 8767 1311 8768
rect 107 8704 147 8752
rect 1273 8758 1311 8767
rect 1273 8738 1282 8758
rect 1302 8738 1311 8758
rect 1273 8730 1311 8738
rect 1377 8762 1462 8768
rect 1487 8767 1524 8768
rect 1377 8742 1385 8762
rect 1405 8742 1462 8762
rect 1377 8734 1462 8742
rect 1486 8758 1524 8767
rect 1486 8738 1495 8758
rect 1515 8738 1524 8758
rect 1377 8733 1413 8734
rect 1486 8730 1524 8738
rect 1590 8762 1675 8768
rect 1695 8767 1732 8768
rect 1590 8742 1598 8762
rect 1618 8761 1675 8762
rect 1618 8742 1647 8761
rect 1590 8741 1647 8742
rect 1668 8741 1675 8761
rect 1590 8734 1675 8741
rect 1694 8758 1732 8767
rect 1694 8738 1703 8758
rect 1723 8738 1732 8758
rect 1590 8733 1626 8734
rect 1694 8730 1732 8738
rect 1798 8762 1942 8768
rect 1798 8742 1806 8762
rect 1826 8745 1862 8762
rect 1882 8745 1914 8762
rect 1826 8742 1914 8745
rect 1934 8742 1942 8762
rect 1798 8734 1942 8742
rect 1798 8733 1834 8734
rect 1906 8733 1942 8734
rect 2008 8767 2045 8768
rect 2008 8766 2046 8767
rect 2008 8758 2072 8766
rect 2008 8738 2017 8758
rect 2037 8744 2072 8758
rect 2092 8744 2095 8764
rect 2037 8739 2095 8744
rect 2037 8738 2072 8739
rect 418 8708 528 8722
rect 418 8705 461 8708
rect 107 8697 232 8704
rect 418 8700 422 8705
rect 107 8678 199 8697
rect 224 8678 232 8697
rect 107 8668 232 8678
rect 340 8678 422 8700
rect 451 8678 461 8705
rect 489 8681 496 8708
rect 525 8700 528 8708
rect 1274 8701 1311 8730
rect 525 8681 590 8700
rect 1275 8699 1311 8701
rect 1487 8699 1524 8730
rect 1695 8703 1732 8730
rect 2008 8726 2072 8738
rect 489 8678 590 8681
rect 340 8676 590 8678
rect 107 8648 147 8668
rect 106 8639 147 8648
rect 106 8621 116 8639
rect 134 8621 147 8639
rect 106 8612 147 8621
rect 106 8611 143 8612
rect 340 8597 377 8676
rect 418 8663 528 8676
rect 492 8607 523 8608
rect 340 8577 349 8597
rect 369 8577 377 8597
rect 340 8567 377 8577
rect 436 8597 523 8607
rect 436 8577 445 8597
rect 465 8577 523 8597
rect 436 8568 523 8577
rect 436 8567 473 8568
rect 109 8545 146 8549
rect 106 8540 146 8545
rect 106 8522 118 8540
rect 136 8522 146 8540
rect 106 8342 146 8522
rect 492 8515 523 8568
rect 553 8597 590 8676
rect 761 8673 1154 8693
rect 1174 8673 1177 8693
rect 1275 8677 1524 8699
rect 1693 8698 1734 8703
rect 2112 8700 2139 8878
rect 2790 8790 2817 8968
rect 3195 8965 3236 8970
rect 3405 8969 3654 8991
rect 3752 8975 3755 8995
rect 3775 8975 4168 8995
rect 4339 8992 4376 9071
rect 4406 9100 4437 9153
rect 4783 9146 4823 9326
rect 5161 9326 5215 9331
rect 5161 9308 5172 9326
rect 5190 9308 5215 9326
rect 8785 9347 8953 9348
rect 9193 9347 9231 9435
rect 9492 9417 9539 9435
rect 9456 9378 9568 9417
rect 9839 9411 9879 9435
rect 9456 9377 9499 9378
rect 8785 9324 9231 9347
rect 9457 9376 9499 9377
rect 9457 9356 9464 9376
rect 9483 9356 9499 9376
rect 9457 9348 9499 9356
rect 9527 9376 9568 9378
rect 9527 9356 9541 9376
rect 9560 9356 9568 9376
rect 9840 9367 9879 9411
rect 9527 9348 9568 9356
rect 9457 9342 9568 9348
rect 8785 9321 9229 9324
rect 8785 9319 8953 9321
rect 5161 9299 5215 9308
rect 5162 9298 5215 9299
rect 5475 9303 5585 9317
rect 5475 9300 5518 9303
rect 5475 9295 5479 9300
rect 5397 9273 5479 9295
rect 5508 9273 5518 9300
rect 5546 9276 5553 9303
rect 5582 9295 5585 9303
rect 5582 9276 5647 9295
rect 5546 9273 5647 9276
rect 5397 9271 5647 9273
rect 5165 9235 5202 9236
rect 4783 9128 4793 9146
rect 4811 9128 4823 9146
rect 4783 9123 4823 9128
rect 5161 9232 5202 9235
rect 5161 9227 5203 9232
rect 5161 9209 5174 9227
rect 5192 9209 5203 9227
rect 5161 9195 5203 9209
rect 5241 9195 5288 9199
rect 5161 9189 5288 9195
rect 5161 9160 5249 9189
rect 5278 9160 5288 9189
rect 5397 9192 5434 9271
rect 5475 9258 5585 9271
rect 5549 9202 5580 9203
rect 5397 9172 5406 9192
rect 5426 9172 5434 9192
rect 5397 9162 5434 9172
rect 5493 9192 5580 9202
rect 5493 9172 5502 9192
rect 5522 9172 5580 9192
rect 5493 9163 5580 9172
rect 5493 9162 5530 9163
rect 5161 9156 5288 9160
rect 5161 9139 5200 9156
rect 5241 9155 5288 9156
rect 4783 9119 4820 9123
rect 5161 9121 5172 9139
rect 5190 9121 5200 9139
rect 5161 9112 5200 9121
rect 5162 9111 5199 9112
rect 5549 9110 5580 9163
rect 5610 9192 5647 9271
rect 5818 9268 6211 9288
rect 6231 9268 6234 9288
rect 5818 9263 6234 9268
rect 5818 9262 6159 9263
rect 5762 9202 5793 9203
rect 5610 9172 5619 9192
rect 5639 9172 5647 9192
rect 5610 9162 5647 9172
rect 5706 9195 5793 9202
rect 5706 9192 5767 9195
rect 5706 9172 5715 9192
rect 5735 9175 5767 9192
rect 5788 9175 5793 9195
rect 5735 9172 5793 9175
rect 5706 9165 5793 9172
rect 5818 9192 5855 9262
rect 6121 9261 6158 9262
rect 5970 9202 6006 9203
rect 5818 9172 5827 9192
rect 5847 9172 5855 9192
rect 5706 9163 5762 9165
rect 5706 9162 5743 9163
rect 5818 9162 5855 9172
rect 5914 9192 6062 9202
rect 6162 9199 6258 9201
rect 5914 9172 5923 9192
rect 5943 9172 6033 9192
rect 6053 9172 6062 9192
rect 5914 9163 6062 9172
rect 6120 9192 6258 9199
rect 6120 9172 6129 9192
rect 6149 9172 6258 9192
rect 6120 9163 6258 9172
rect 5914 9162 5951 9163
rect 5970 9111 6006 9163
rect 6025 9162 6062 9163
rect 6121 9162 6158 9163
rect 5441 9109 5482 9110
rect 5333 9102 5482 9109
rect 4456 9100 4493 9101
rect 4406 9091 4493 9100
rect 4406 9071 4464 9091
rect 4484 9071 4493 9091
rect 4406 9061 4493 9071
rect 4552 9091 4589 9101
rect 4552 9071 4560 9091
rect 4580 9071 4589 9091
rect 5333 9082 5451 9102
rect 5471 9082 5482 9102
rect 5333 9074 5482 9082
rect 5549 9106 5908 9110
rect 5549 9101 5871 9106
rect 5549 9077 5662 9101
rect 5686 9082 5871 9101
rect 5895 9082 5908 9106
rect 5686 9077 5908 9082
rect 5549 9074 5908 9077
rect 5970 9074 6005 9111
rect 6073 9108 6173 9111
rect 6073 9104 6140 9108
rect 6073 9078 6085 9104
rect 6111 9082 6140 9104
rect 6166 9082 6173 9108
rect 6111 9078 6173 9082
rect 6073 9074 6173 9078
rect 4406 9060 4437 9061
rect 4401 8992 4511 9005
rect 4552 8992 4589 9071
rect 4786 9056 4823 9057
rect 4782 9047 4823 9056
rect 5549 9053 5580 9074
rect 5970 9053 6006 9074
rect 5392 9052 5429 9053
rect 5166 9049 5200 9050
rect 4782 9029 4795 9047
rect 4813 9029 4823 9047
rect 4782 9020 4823 9029
rect 5165 9040 5202 9049
rect 5165 9022 5174 9040
rect 5192 9022 5202 9040
rect 4782 9000 4822 9020
rect 5165 9012 5202 9022
rect 5391 9043 5429 9052
rect 5391 9023 5400 9043
rect 5420 9023 5429 9043
rect 5391 9015 5429 9023
rect 5495 9047 5580 9053
rect 5605 9052 5642 9053
rect 5495 9027 5503 9047
rect 5523 9027 5580 9047
rect 5495 9019 5580 9027
rect 5604 9043 5642 9052
rect 5604 9023 5613 9043
rect 5633 9023 5642 9043
rect 5495 9018 5531 9019
rect 5604 9015 5642 9023
rect 5708 9047 5793 9053
rect 5813 9052 5850 9053
rect 5708 9027 5716 9047
rect 5736 9046 5793 9047
rect 5736 9027 5765 9046
rect 5708 9026 5765 9027
rect 5786 9026 5793 9046
rect 5708 9019 5793 9026
rect 5812 9043 5850 9052
rect 5812 9023 5821 9043
rect 5841 9023 5850 9043
rect 5708 9018 5744 9019
rect 5812 9015 5850 9023
rect 5916 9047 6060 9053
rect 5916 9027 5924 9047
rect 5944 9046 6032 9047
rect 5944 9027 5975 9046
rect 5916 9026 5975 9027
rect 6000 9027 6032 9046
rect 6052 9027 6060 9047
rect 6000 9026 6060 9027
rect 5916 9019 6060 9026
rect 5916 9018 5952 9019
rect 6024 9018 6060 9019
rect 6126 9052 6163 9053
rect 6126 9051 6164 9052
rect 6126 9043 6190 9051
rect 6126 9023 6135 9043
rect 6155 9029 6190 9043
rect 6210 9029 6213 9049
rect 6155 9024 6213 9029
rect 6155 9023 6190 9024
rect 4339 8990 4589 8992
rect 4339 8987 4440 8990
rect 2857 8930 2921 8942
rect 3197 8938 3234 8965
rect 3405 8938 3442 8969
rect 3618 8967 3654 8969
rect 4339 8968 4404 8987
rect 3618 8938 3655 8967
rect 4401 8960 4404 8968
rect 4433 8960 4440 8987
rect 4468 8963 4478 8990
rect 4507 8968 4589 8990
rect 4697 8990 4822 9000
rect 4697 8971 4705 8990
rect 4730 8971 4822 8990
rect 4507 8963 4511 8968
rect 4697 8964 4822 8971
rect 4468 8960 4511 8963
rect 4401 8946 4511 8960
rect 2857 8929 2892 8930
rect 2834 8924 2892 8929
rect 2834 8904 2837 8924
rect 2857 8910 2892 8924
rect 2912 8910 2921 8930
rect 2857 8902 2921 8910
rect 2883 8901 2921 8902
rect 2884 8900 2921 8901
rect 2987 8934 3023 8935
rect 3095 8934 3131 8935
rect 2987 8926 3131 8934
rect 2987 8906 2995 8926
rect 3015 8906 3103 8926
rect 3123 8906 3131 8926
rect 2987 8900 3131 8906
rect 3197 8930 3235 8938
rect 3303 8934 3339 8935
rect 3197 8910 3206 8930
rect 3226 8910 3235 8930
rect 3197 8901 3235 8910
rect 3254 8927 3339 8934
rect 3254 8907 3261 8927
rect 3282 8926 3339 8927
rect 3282 8907 3311 8926
rect 3254 8906 3311 8907
rect 3331 8906 3339 8926
rect 3197 8900 3234 8901
rect 3254 8900 3339 8906
rect 3405 8930 3443 8938
rect 3516 8934 3552 8935
rect 3405 8910 3414 8930
rect 3434 8910 3443 8930
rect 3405 8901 3443 8910
rect 3467 8926 3552 8934
rect 3467 8906 3524 8926
rect 3544 8906 3552 8926
rect 3405 8900 3442 8901
rect 3467 8900 3552 8906
rect 3618 8930 3656 8938
rect 3618 8910 3627 8930
rect 3647 8910 3656 8930
rect 3618 8901 3656 8910
rect 4782 8916 4822 8964
rect 5166 8984 5200 9012
rect 5392 8986 5429 9015
rect 5393 8984 5429 8986
rect 5605 8984 5642 9015
rect 5166 8983 5338 8984
rect 5166 8951 5352 8983
rect 5393 8962 5642 8984
rect 5813 8983 5850 9015
rect 6126 9011 6190 9023
rect 6230 8985 6257 9163
rect 8785 9141 8812 9319
rect 8852 9281 8916 9293
rect 9192 9289 9229 9321
rect 9400 9320 9649 9342
rect 9400 9289 9437 9320
rect 9613 9318 9649 9320
rect 9613 9289 9650 9318
rect 8852 9280 8887 9281
rect 8829 9275 8887 9280
rect 8829 9255 8832 9275
rect 8852 9261 8887 9275
rect 8907 9261 8916 9281
rect 8852 9253 8916 9261
rect 8878 9252 8916 9253
rect 8879 9251 8916 9252
rect 8982 9285 9018 9286
rect 9090 9285 9126 9286
rect 8982 9280 9126 9285
rect 8982 9277 9044 9280
rect 8982 9257 8990 9277
rect 9010 9260 9044 9277
rect 9067 9277 9126 9280
rect 9067 9260 9098 9277
rect 9010 9257 9098 9260
rect 9118 9257 9126 9277
rect 8982 9251 9126 9257
rect 9192 9281 9230 9289
rect 9298 9285 9334 9286
rect 9192 9261 9201 9281
rect 9221 9261 9230 9281
rect 9192 9252 9230 9261
rect 9249 9278 9334 9285
rect 9249 9258 9256 9278
rect 9277 9277 9334 9278
rect 9277 9258 9306 9277
rect 9249 9257 9306 9258
rect 9326 9257 9334 9277
rect 9192 9251 9229 9252
rect 9249 9251 9334 9257
rect 9400 9281 9438 9289
rect 9511 9285 9547 9286
rect 9400 9261 9409 9281
rect 9429 9261 9438 9281
rect 9400 9252 9438 9261
rect 9462 9277 9547 9285
rect 9462 9257 9519 9277
rect 9539 9257 9547 9277
rect 9400 9251 9437 9252
rect 9462 9251 9547 9257
rect 9613 9281 9651 9289
rect 9613 9261 9622 9281
rect 9642 9261 9651 9281
rect 9613 9252 9651 9261
rect 9613 9251 9650 9252
rect 9036 9230 9072 9251
rect 9462 9230 9493 9251
rect 8869 9226 8969 9230
rect 8869 9222 8931 9226
rect 8869 9196 8876 9222
rect 8902 9200 8931 9222
rect 8957 9200 8969 9226
rect 8902 9196 8969 9200
rect 8869 9193 8969 9196
rect 9037 9193 9072 9230
rect 9134 9227 9493 9230
rect 9134 9222 9356 9227
rect 9134 9198 9147 9222
rect 9171 9203 9356 9222
rect 9380 9203 9493 9227
rect 9171 9198 9493 9203
rect 9134 9194 9493 9198
rect 9560 9222 9709 9230
rect 9560 9202 9571 9222
rect 9591 9202 9709 9222
rect 9560 9195 9709 9202
rect 9560 9194 9601 9195
rect 8884 9141 8921 9142
rect 8980 9141 9017 9142
rect 9036 9141 9072 9193
rect 9091 9141 9128 9142
rect 8784 9132 8922 9141
rect 8784 9112 8893 9132
rect 8913 9112 8922 9132
rect 8784 9105 8922 9112
rect 8980 9132 9128 9141
rect 8980 9112 8989 9132
rect 9009 9112 9099 9132
rect 9119 9112 9128 9132
rect 8784 9103 8880 9105
rect 8980 9102 9128 9112
rect 9187 9132 9224 9142
rect 9299 9141 9336 9142
rect 9280 9139 9336 9141
rect 9187 9112 9195 9132
rect 9215 9112 9224 9132
rect 9036 9101 9072 9102
rect 6413 9059 6523 9073
rect 6413 9056 6456 9059
rect 6413 9051 6417 9056
rect 6089 8983 6257 8985
rect 5813 8977 6257 8983
rect 5166 8919 5200 8951
rect 3618 8900 3655 8901
rect 3041 8879 3077 8900
rect 3467 8879 3498 8900
rect 4782 8898 4793 8916
rect 4811 8898 4822 8916
rect 4782 8890 4822 8898
rect 5162 8910 5200 8919
rect 5162 8892 5172 8910
rect 5190 8892 5200 8910
rect 4783 8889 4820 8890
rect 5162 8886 5200 8892
rect 5318 8888 5352 8951
rect 5474 8956 5585 8962
rect 5474 8948 5515 8956
rect 5474 8928 5482 8948
rect 5501 8928 5515 8948
rect 5474 8926 5515 8928
rect 5543 8948 5585 8956
rect 5543 8928 5559 8948
rect 5578 8928 5585 8948
rect 5543 8926 5585 8928
rect 5474 8911 5585 8926
rect 5812 8957 6257 8977
rect 5812 8888 5850 8957
rect 6089 8956 6257 8957
rect 6335 9029 6417 9051
rect 6446 9029 6456 9056
rect 6484 9032 6491 9059
rect 6520 9051 6523 9059
rect 8518 9068 8629 9083
rect 8518 9066 8560 9068
rect 6520 9032 6585 9051
rect 6484 9029 6585 9032
rect 6335 9027 6585 9029
rect 6335 8948 6372 9027
rect 6413 9014 6523 9027
rect 6487 8958 6518 8959
rect 6335 8928 6344 8948
rect 6364 8928 6372 8948
rect 6335 8918 6372 8928
rect 6431 8948 6518 8958
rect 6431 8928 6440 8948
rect 6460 8928 6518 8948
rect 6431 8919 6518 8928
rect 6431 8918 6468 8919
rect 5162 8882 5199 8886
rect 2874 8875 2974 8879
rect 2874 8871 2936 8875
rect 2874 8845 2881 8871
rect 2907 8849 2936 8871
rect 2962 8849 2974 8875
rect 2907 8845 2974 8849
rect 2874 8842 2974 8845
rect 3042 8842 3077 8879
rect 3139 8876 3498 8879
rect 3139 8871 3361 8876
rect 3139 8847 3152 8871
rect 3176 8852 3361 8871
rect 3385 8852 3498 8876
rect 3176 8847 3498 8852
rect 3139 8843 3498 8847
rect 3565 8871 3714 8879
rect 5318 8877 5850 8888
rect 3565 8851 3576 8871
rect 3596 8851 3714 8871
rect 5317 8861 5850 8877
rect 6487 8866 6518 8919
rect 6548 8948 6585 9027
rect 6756 9024 7149 9044
rect 7169 9024 7172 9044
rect 8251 9039 8292 9048
rect 6756 9019 7172 9024
rect 7846 9037 8014 9038
rect 8251 9037 8260 9039
rect 6756 9018 7097 9019
rect 6700 8958 6731 8959
rect 6548 8928 6557 8948
rect 6577 8928 6585 8948
rect 6548 8918 6585 8928
rect 6644 8951 6731 8958
rect 6644 8948 6705 8951
rect 6644 8928 6653 8948
rect 6673 8931 6705 8948
rect 6726 8931 6731 8951
rect 6673 8928 6731 8931
rect 6644 8921 6731 8928
rect 6756 8948 6793 9018
rect 7059 9017 7096 9018
rect 7846 9017 8260 9037
rect 8286 9017 8292 9039
rect 8518 9046 8525 9066
rect 8544 9046 8560 9066
rect 8518 9038 8560 9046
rect 8588 9066 8629 9068
rect 8588 9046 8602 9066
rect 8621 9046 8629 9066
rect 8588 9038 8629 9046
rect 8884 9042 8921 9043
rect 9187 9042 9224 9112
rect 9249 9132 9336 9139
rect 9249 9129 9307 9132
rect 9249 9109 9254 9129
rect 9275 9112 9307 9129
rect 9327 9112 9336 9132
rect 9275 9109 9336 9112
rect 9249 9102 9336 9109
rect 9395 9132 9432 9142
rect 9395 9112 9403 9132
rect 9423 9112 9432 9132
rect 9249 9101 9280 9102
rect 8883 9041 9224 9042
rect 8518 9032 8629 9038
rect 8808 9036 9224 9041
rect 7846 9011 8292 9017
rect 7846 9009 8014 9011
rect 6908 8958 6944 8959
rect 6756 8928 6765 8948
rect 6785 8928 6793 8948
rect 6644 8919 6700 8921
rect 6644 8918 6681 8919
rect 6756 8918 6793 8928
rect 6852 8948 7000 8958
rect 7100 8955 7196 8957
rect 6852 8928 6861 8948
rect 6881 8928 6971 8948
rect 6991 8928 7000 8948
rect 6852 8919 7000 8928
rect 7058 8948 7196 8955
rect 7058 8928 7067 8948
rect 7087 8928 7196 8948
rect 7058 8919 7196 8928
rect 6852 8918 6889 8919
rect 6908 8867 6944 8919
rect 6963 8918 7000 8919
rect 7059 8918 7096 8919
rect 6379 8865 6420 8866
rect 5317 8860 5831 8861
rect 3565 8844 3714 8851
rect 6271 8858 6420 8865
rect 4154 8848 4668 8849
rect 3565 8843 3606 8844
rect 3041 8807 3077 8842
rect 2889 8790 2926 8791
rect 2985 8790 3022 8791
rect 3041 8790 3048 8807
rect 2789 8781 2927 8790
rect 2789 8761 2898 8781
rect 2918 8761 2927 8781
rect 2789 8754 2927 8761
rect 2985 8781 3048 8790
rect 2985 8761 2994 8781
rect 3014 8766 3048 8781
rect 3069 8790 3077 8807
rect 3096 8790 3133 8791
rect 3069 8781 3133 8790
rect 3069 8766 3104 8781
rect 3014 8761 3104 8766
rect 3124 8761 3133 8781
rect 2789 8752 2885 8754
rect 2985 8751 3133 8761
rect 3192 8781 3229 8791
rect 3304 8790 3341 8791
rect 3285 8788 3341 8790
rect 3192 8761 3200 8781
rect 3220 8761 3229 8781
rect 3041 8750 3077 8751
rect 1971 8698 2139 8700
rect 1693 8692 2139 8698
rect 761 8668 1177 8673
rect 1356 8671 1467 8677
rect 761 8667 1102 8668
rect 705 8607 736 8608
rect 553 8577 562 8597
rect 582 8577 590 8597
rect 553 8567 590 8577
rect 649 8600 736 8607
rect 649 8597 710 8600
rect 649 8577 658 8597
rect 678 8580 710 8597
rect 731 8580 736 8600
rect 678 8577 736 8580
rect 649 8570 736 8577
rect 761 8597 798 8667
rect 1064 8666 1101 8667
rect 1356 8663 1397 8671
rect 1356 8643 1364 8663
rect 1383 8643 1397 8663
rect 1356 8641 1397 8643
rect 1425 8663 1467 8671
rect 1425 8643 1441 8663
rect 1460 8643 1467 8663
rect 1693 8670 1699 8692
rect 1725 8672 2139 8692
rect 2889 8691 2926 8692
rect 3192 8691 3229 8761
rect 3254 8781 3341 8788
rect 3254 8778 3312 8781
rect 3254 8758 3259 8778
rect 3280 8761 3312 8778
rect 3332 8761 3341 8781
rect 3280 8758 3341 8761
rect 3254 8751 3341 8758
rect 3400 8781 3437 8791
rect 3400 8761 3408 8781
rect 3428 8761 3437 8781
rect 3254 8750 3285 8751
rect 2888 8690 3229 8691
rect 1725 8670 1734 8672
rect 1971 8671 2139 8672
rect 2813 8689 3229 8690
rect 2813 8685 3189 8689
rect 1693 8661 1734 8670
rect 2813 8665 2816 8685
rect 2836 8672 3189 8685
rect 3221 8672 3229 8689
rect 2836 8665 3229 8672
rect 3400 8682 3437 8761
rect 3467 8790 3498 8843
rect 4135 8832 4668 8848
rect 6271 8838 6389 8858
rect 6409 8838 6420 8858
rect 4135 8821 4667 8832
rect 6271 8830 6420 8838
rect 6487 8862 6846 8866
rect 6487 8857 6809 8862
rect 6487 8833 6600 8857
rect 6624 8838 6809 8857
rect 6833 8838 6846 8862
rect 6624 8833 6846 8838
rect 6487 8830 6846 8833
rect 6908 8830 6943 8867
rect 7011 8864 7111 8867
rect 7011 8860 7078 8864
rect 7011 8834 7023 8860
rect 7049 8838 7078 8860
rect 7104 8838 7111 8864
rect 7049 8834 7111 8838
rect 7011 8830 7111 8834
rect 4786 8823 4823 8827
rect 3517 8790 3554 8791
rect 3467 8781 3554 8790
rect 3467 8761 3525 8781
rect 3545 8761 3554 8781
rect 3467 8751 3554 8761
rect 3613 8781 3650 8791
rect 3613 8761 3621 8781
rect 3641 8761 3650 8781
rect 3467 8750 3498 8751
rect 3462 8682 3572 8695
rect 3613 8682 3650 8761
rect 3400 8680 3650 8682
rect 3400 8677 3501 8680
rect 3400 8658 3465 8677
rect 1425 8641 1467 8643
rect 1356 8626 1467 8641
rect 3462 8650 3465 8658
rect 3494 8650 3501 8677
rect 3529 8653 3539 8680
rect 3568 8658 3650 8680
rect 3728 8752 3896 8753
rect 4135 8752 4173 8821
rect 3728 8732 4173 8752
rect 4400 8783 4511 8798
rect 4400 8781 4442 8783
rect 4400 8761 4407 8781
rect 4426 8761 4442 8781
rect 4400 8753 4442 8761
rect 4470 8781 4511 8783
rect 4470 8761 4484 8781
rect 4503 8761 4511 8781
rect 4470 8753 4511 8761
rect 4400 8747 4511 8753
rect 4633 8758 4667 8821
rect 4785 8817 4823 8823
rect 5165 8819 5202 8820
rect 4785 8799 4795 8817
rect 4813 8799 4823 8817
rect 4785 8790 4823 8799
rect 5163 8811 5203 8819
rect 5163 8793 5174 8811
rect 5192 8793 5203 8811
rect 6487 8809 6518 8830
rect 6908 8809 6944 8830
rect 6330 8808 6367 8809
rect 4785 8758 4819 8790
rect 3728 8726 4172 8732
rect 3728 8724 3896 8726
rect 3568 8653 3572 8658
rect 3529 8650 3572 8653
rect 3462 8636 3572 8650
rect 913 8607 949 8608
rect 761 8577 770 8597
rect 790 8577 798 8597
rect 649 8568 705 8570
rect 649 8567 686 8568
rect 761 8567 798 8577
rect 857 8597 1005 8607
rect 1105 8604 1201 8606
rect 857 8577 866 8597
rect 886 8577 976 8597
rect 996 8577 1005 8597
rect 857 8568 1005 8577
rect 1063 8597 1201 8604
rect 1063 8577 1072 8597
rect 1092 8577 1201 8597
rect 1063 8568 1201 8577
rect 857 8567 894 8568
rect 913 8516 949 8568
rect 968 8567 1005 8568
rect 1064 8567 1101 8568
rect 384 8514 425 8515
rect 276 8507 425 8514
rect 276 8487 394 8507
rect 414 8487 425 8507
rect 276 8479 425 8487
rect 492 8511 851 8515
rect 492 8506 814 8511
rect 492 8482 605 8506
rect 629 8487 814 8506
rect 838 8487 851 8511
rect 629 8482 851 8487
rect 492 8479 851 8482
rect 913 8479 948 8516
rect 1016 8513 1116 8516
rect 1016 8509 1083 8513
rect 1016 8483 1028 8509
rect 1054 8487 1083 8509
rect 1109 8487 1116 8513
rect 1054 8483 1116 8487
rect 1016 8479 1116 8483
rect 492 8458 523 8479
rect 913 8458 949 8479
rect 335 8457 372 8458
rect 334 8448 372 8457
rect 334 8428 343 8448
rect 363 8428 372 8448
rect 334 8420 372 8428
rect 438 8452 523 8458
rect 548 8457 585 8458
rect 438 8432 446 8452
rect 466 8432 523 8452
rect 438 8424 523 8432
rect 547 8448 585 8457
rect 547 8428 556 8448
rect 576 8428 585 8448
rect 438 8423 474 8424
rect 547 8420 585 8428
rect 651 8452 736 8458
rect 756 8457 793 8458
rect 651 8432 659 8452
rect 679 8451 736 8452
rect 679 8432 708 8451
rect 651 8431 708 8432
rect 729 8431 736 8451
rect 651 8424 736 8431
rect 755 8448 793 8457
rect 755 8428 764 8448
rect 784 8428 793 8448
rect 651 8423 687 8424
rect 755 8420 793 8428
rect 859 8452 1003 8458
rect 859 8432 867 8452
rect 887 8449 975 8452
rect 887 8432 918 8449
rect 859 8429 918 8432
rect 941 8432 975 8449
rect 995 8432 1003 8452
rect 941 8429 1003 8432
rect 859 8424 1003 8429
rect 859 8423 895 8424
rect 967 8423 1003 8424
rect 1069 8457 1106 8458
rect 1069 8456 1107 8457
rect 1069 8448 1133 8456
rect 1069 8428 1078 8448
rect 1098 8434 1133 8448
rect 1153 8434 1156 8454
rect 1098 8429 1156 8434
rect 1098 8428 1133 8429
rect 335 8391 372 8420
rect 336 8389 372 8391
rect 548 8389 585 8420
rect 336 8367 585 8389
rect 756 8388 793 8420
rect 1069 8416 1133 8428
rect 1173 8390 1200 8568
rect 3728 8546 3755 8724
rect 3795 8686 3859 8698
rect 4135 8694 4172 8726
rect 4343 8725 4592 8747
rect 4633 8726 4819 8758
rect 4647 8725 4819 8726
rect 4343 8694 4380 8725
rect 4556 8723 4592 8725
rect 4556 8694 4593 8723
rect 4785 8697 4819 8725
rect 5163 8745 5203 8793
rect 6329 8799 6367 8808
rect 6329 8779 6338 8799
rect 6358 8779 6367 8799
rect 6329 8771 6367 8779
rect 6433 8803 6518 8809
rect 6543 8808 6580 8809
rect 6433 8783 6441 8803
rect 6461 8783 6518 8803
rect 6433 8775 6518 8783
rect 6542 8799 6580 8808
rect 6542 8779 6551 8799
rect 6571 8779 6580 8799
rect 6433 8774 6469 8775
rect 6542 8771 6580 8779
rect 6646 8803 6731 8809
rect 6751 8808 6788 8809
rect 6646 8783 6654 8803
rect 6674 8802 6731 8803
rect 6674 8783 6703 8802
rect 6646 8782 6703 8783
rect 6724 8782 6731 8802
rect 6646 8775 6731 8782
rect 6750 8799 6788 8808
rect 6750 8779 6759 8799
rect 6779 8779 6788 8799
rect 6646 8774 6682 8775
rect 6750 8771 6788 8779
rect 6854 8803 6998 8809
rect 6854 8783 6862 8803
rect 6882 8786 6918 8803
rect 6938 8786 6970 8803
rect 6882 8783 6970 8786
rect 6990 8783 6998 8803
rect 6854 8775 6998 8783
rect 6854 8774 6890 8775
rect 6962 8774 6998 8775
rect 7064 8808 7101 8809
rect 7064 8807 7102 8808
rect 7064 8799 7128 8807
rect 7064 8779 7073 8799
rect 7093 8785 7128 8799
rect 7148 8785 7151 8805
rect 7093 8780 7151 8785
rect 7093 8779 7128 8780
rect 5474 8749 5584 8763
rect 5474 8746 5517 8749
rect 5163 8738 5288 8745
rect 5474 8741 5478 8746
rect 5163 8719 5255 8738
rect 5280 8719 5288 8738
rect 5163 8709 5288 8719
rect 5396 8719 5478 8741
rect 5507 8719 5517 8746
rect 5545 8722 5552 8749
rect 5581 8741 5584 8749
rect 6330 8742 6367 8771
rect 5581 8722 5646 8741
rect 6331 8740 6367 8742
rect 6543 8740 6580 8771
rect 6751 8744 6788 8771
rect 7064 8767 7128 8779
rect 5545 8719 5646 8722
rect 5396 8717 5646 8719
rect 3795 8685 3830 8686
rect 3772 8680 3830 8685
rect 3772 8660 3775 8680
rect 3795 8666 3830 8680
rect 3850 8666 3859 8686
rect 3795 8658 3859 8666
rect 3821 8657 3859 8658
rect 3822 8656 3859 8657
rect 3925 8690 3961 8691
rect 4033 8690 4069 8691
rect 3925 8683 4069 8690
rect 3925 8682 3985 8683
rect 3925 8662 3933 8682
rect 3953 8663 3985 8682
rect 4010 8682 4069 8683
rect 4010 8663 4041 8682
rect 3953 8662 4041 8663
rect 4061 8662 4069 8682
rect 3925 8656 4069 8662
rect 4135 8686 4173 8694
rect 4241 8690 4277 8691
rect 4135 8666 4144 8686
rect 4164 8666 4173 8686
rect 4135 8657 4173 8666
rect 4192 8683 4277 8690
rect 4192 8663 4199 8683
rect 4220 8682 4277 8683
rect 4220 8663 4249 8682
rect 4192 8662 4249 8663
rect 4269 8662 4277 8682
rect 4135 8656 4172 8657
rect 4192 8656 4277 8662
rect 4343 8686 4381 8694
rect 4454 8690 4490 8691
rect 4343 8666 4352 8686
rect 4372 8666 4381 8686
rect 4343 8657 4381 8666
rect 4405 8682 4490 8690
rect 4405 8662 4462 8682
rect 4482 8662 4490 8682
rect 4343 8656 4380 8657
rect 4405 8656 4490 8662
rect 4556 8686 4594 8694
rect 4556 8666 4565 8686
rect 4585 8666 4594 8686
rect 4556 8657 4594 8666
rect 4783 8687 4820 8697
rect 5163 8689 5203 8709
rect 4783 8669 4793 8687
rect 4811 8669 4820 8687
rect 4783 8660 4820 8669
rect 5162 8680 5203 8689
rect 5162 8662 5172 8680
rect 5190 8662 5203 8680
rect 4785 8659 4819 8660
rect 4556 8656 4593 8657
rect 3979 8635 4015 8656
rect 4405 8635 4436 8656
rect 5162 8653 5203 8662
rect 5162 8652 5199 8653
rect 5396 8638 5433 8717
rect 5474 8704 5584 8717
rect 5548 8648 5579 8649
rect 3812 8631 3912 8635
rect 3812 8627 3874 8631
rect 3812 8601 3819 8627
rect 3845 8605 3874 8627
rect 3900 8605 3912 8631
rect 3845 8601 3912 8605
rect 3812 8598 3912 8601
rect 3980 8598 4015 8635
rect 4077 8632 4436 8635
rect 4077 8627 4299 8632
rect 4077 8603 4090 8627
rect 4114 8608 4299 8627
rect 4323 8608 4436 8632
rect 4114 8603 4436 8608
rect 4077 8599 4436 8603
rect 4503 8627 4652 8635
rect 4503 8607 4514 8627
rect 4534 8607 4652 8627
rect 5396 8618 5405 8638
rect 5425 8618 5433 8638
rect 5396 8608 5433 8618
rect 5492 8638 5579 8648
rect 5492 8618 5501 8638
rect 5521 8618 5579 8638
rect 5492 8609 5579 8618
rect 5492 8608 5529 8609
rect 4503 8600 4652 8607
rect 4503 8599 4544 8600
rect 3827 8546 3864 8547
rect 3923 8546 3960 8547
rect 3979 8546 4015 8598
rect 4034 8546 4071 8547
rect 3727 8537 3865 8546
rect 3322 8516 3433 8531
rect 3322 8514 3364 8516
rect 2992 8493 3097 8495
rect 2648 8485 2818 8486
rect 2992 8485 3041 8493
rect 2648 8466 3041 8485
rect 3072 8466 3097 8493
rect 3322 8494 3329 8514
rect 3348 8494 3364 8514
rect 3322 8486 3364 8494
rect 3392 8514 3433 8516
rect 3392 8494 3406 8514
rect 3425 8494 3433 8514
rect 3727 8517 3836 8537
rect 3856 8517 3865 8537
rect 3727 8510 3865 8517
rect 3923 8537 4071 8546
rect 3923 8517 3932 8537
rect 3952 8517 4042 8537
rect 4062 8517 4071 8537
rect 3727 8508 3823 8510
rect 3923 8507 4071 8517
rect 4130 8537 4167 8547
rect 4242 8546 4279 8547
rect 4223 8544 4279 8546
rect 4130 8517 4138 8537
rect 4158 8517 4167 8537
rect 3979 8506 4015 8507
rect 3392 8486 3433 8494
rect 3322 8480 3433 8486
rect 2648 8459 3097 8466
rect 2648 8457 2818 8459
rect 1498 8426 1608 8440
rect 1498 8423 1541 8426
rect 1498 8418 1502 8423
rect 1032 8388 1200 8390
rect 756 8385 1200 8388
rect 417 8361 528 8367
rect 417 8353 458 8361
rect 106 8298 145 8342
rect 417 8333 425 8353
rect 444 8333 458 8353
rect 417 8331 458 8333
rect 486 8353 528 8361
rect 486 8333 502 8353
rect 521 8333 528 8353
rect 486 8331 528 8333
rect 417 8316 528 8331
rect 754 8362 1200 8385
rect 106 8274 146 8298
rect 446 8274 493 8276
rect 754 8274 792 8362
rect 1032 8361 1200 8362
rect 1420 8396 1502 8418
rect 1531 8396 1541 8423
rect 1569 8399 1576 8426
rect 1605 8418 1608 8426
rect 1605 8399 1670 8418
rect 1569 8396 1670 8399
rect 1420 8394 1670 8396
rect 1420 8315 1457 8394
rect 1498 8381 1608 8394
rect 1572 8325 1603 8326
rect 1420 8295 1429 8315
rect 1449 8295 1457 8315
rect 1420 8285 1457 8295
rect 1516 8315 1603 8325
rect 1516 8295 1525 8315
rect 1545 8295 1603 8315
rect 1516 8286 1603 8295
rect 1516 8285 1553 8286
rect 106 8241 792 8274
rect 106 8184 145 8241
rect 754 8239 792 8241
rect 1572 8233 1603 8286
rect 1633 8315 1670 8394
rect 1841 8407 2234 8411
rect 1841 8390 1860 8407
rect 1880 8391 2234 8407
rect 2254 8391 2257 8411
rect 1880 8390 2257 8391
rect 1841 8386 2257 8390
rect 1841 8385 2182 8386
rect 1785 8325 1816 8326
rect 1633 8295 1642 8315
rect 1662 8295 1670 8315
rect 1633 8285 1670 8295
rect 1729 8318 1816 8325
rect 1729 8315 1790 8318
rect 1729 8295 1738 8315
rect 1758 8298 1790 8315
rect 1811 8298 1816 8318
rect 1758 8295 1816 8298
rect 1729 8288 1816 8295
rect 1841 8315 1878 8385
rect 2144 8384 2181 8385
rect 1993 8325 2029 8326
rect 1841 8295 1850 8315
rect 1870 8295 1878 8315
rect 1729 8286 1785 8288
rect 1729 8285 1766 8286
rect 1841 8285 1878 8295
rect 1937 8315 2085 8325
rect 2185 8322 2281 8324
rect 1937 8295 1946 8315
rect 1966 8295 2056 8315
rect 2076 8295 2085 8315
rect 1937 8286 2085 8295
rect 2143 8315 2281 8322
rect 2143 8295 2152 8315
rect 2172 8295 2281 8315
rect 2143 8286 2281 8295
rect 1937 8285 1974 8286
rect 1993 8234 2029 8286
rect 2048 8285 2085 8286
rect 2144 8285 2181 8286
rect 1464 8232 1505 8233
rect 1356 8225 1505 8232
rect 1356 8205 1474 8225
rect 1494 8205 1505 8225
rect 1356 8197 1505 8205
rect 1572 8229 1931 8233
rect 1572 8224 1894 8229
rect 1572 8200 1685 8224
rect 1709 8205 1894 8224
rect 1918 8205 1931 8229
rect 1709 8200 1931 8205
rect 1572 8197 1931 8200
rect 1993 8197 2028 8234
rect 2096 8231 2196 8234
rect 2096 8227 2163 8231
rect 2096 8201 2108 8227
rect 2134 8205 2163 8227
rect 2189 8205 2196 8231
rect 2134 8201 2196 8205
rect 2096 8197 2196 8201
rect 106 8182 154 8184
rect 106 8164 117 8182
rect 135 8164 154 8182
rect 1572 8176 1603 8197
rect 1993 8176 2029 8197
rect 1415 8175 1452 8176
rect 106 8155 154 8164
rect 107 8154 154 8155
rect 420 8159 530 8173
rect 420 8156 463 8159
rect 420 8151 424 8156
rect 342 8129 424 8151
rect 453 8129 463 8156
rect 491 8132 498 8159
rect 527 8151 530 8159
rect 1414 8166 1452 8175
rect 527 8132 592 8151
rect 1414 8146 1423 8166
rect 1443 8146 1452 8166
rect 491 8129 592 8132
rect 342 8127 592 8129
rect 110 8091 147 8092
rect 106 8088 147 8091
rect 106 8083 148 8088
rect 106 8065 119 8083
rect 137 8065 148 8083
rect 106 8051 148 8065
rect 186 8051 233 8055
rect 106 8045 233 8051
rect 106 8016 194 8045
rect 223 8016 233 8045
rect 342 8048 379 8127
rect 420 8114 530 8127
rect 494 8058 525 8059
rect 342 8028 351 8048
rect 371 8028 379 8048
rect 342 8018 379 8028
rect 438 8048 525 8058
rect 438 8028 447 8048
rect 467 8028 525 8048
rect 438 8019 525 8028
rect 438 8018 475 8019
rect 106 8012 233 8016
rect 106 7995 145 8012
rect 186 8011 233 8012
rect 106 7977 117 7995
rect 135 7977 145 7995
rect 106 7968 145 7977
rect 107 7967 144 7968
rect 494 7966 525 8019
rect 555 8048 592 8127
rect 763 8124 1156 8144
rect 1176 8124 1179 8144
rect 1414 8138 1452 8146
rect 1518 8170 1603 8176
rect 1628 8175 1665 8176
rect 1518 8150 1526 8170
rect 1546 8150 1603 8170
rect 1518 8142 1603 8150
rect 1627 8166 1665 8175
rect 1627 8146 1636 8166
rect 1656 8146 1665 8166
rect 1518 8141 1554 8142
rect 1627 8138 1665 8146
rect 1731 8170 1816 8176
rect 1836 8175 1873 8176
rect 1731 8150 1739 8170
rect 1759 8169 1816 8170
rect 1759 8150 1788 8169
rect 1731 8149 1788 8150
rect 1809 8149 1816 8169
rect 1731 8142 1816 8149
rect 1835 8166 1873 8175
rect 1835 8146 1844 8166
rect 1864 8146 1873 8166
rect 1731 8141 1767 8142
rect 1835 8138 1873 8146
rect 1939 8170 2083 8176
rect 1939 8150 1947 8170
rect 1967 8168 2055 8170
rect 1967 8150 1996 8168
rect 1939 8147 1996 8150
rect 2023 8150 2055 8168
rect 2075 8150 2083 8170
rect 2023 8147 2083 8150
rect 1939 8142 2083 8147
rect 1939 8141 1975 8142
rect 2047 8141 2083 8142
rect 2149 8175 2186 8176
rect 2149 8174 2187 8175
rect 2149 8166 2213 8174
rect 2149 8146 2158 8166
rect 2178 8152 2213 8166
rect 2233 8152 2236 8172
rect 2178 8147 2236 8152
rect 2178 8146 2213 8147
rect 763 8119 1179 8124
rect 763 8118 1104 8119
rect 707 8058 738 8059
rect 555 8028 564 8048
rect 584 8028 592 8048
rect 555 8018 592 8028
rect 651 8051 738 8058
rect 651 8048 712 8051
rect 651 8028 660 8048
rect 680 8031 712 8048
rect 733 8031 738 8051
rect 680 8028 738 8031
rect 651 8021 738 8028
rect 763 8048 800 8118
rect 1066 8117 1103 8118
rect 1415 8109 1452 8138
rect 1416 8107 1452 8109
rect 1628 8107 1665 8138
rect 1416 8085 1665 8107
rect 1836 8106 1873 8138
rect 2149 8134 2213 8146
rect 2253 8108 2280 8286
rect 2648 8279 2677 8457
rect 2717 8419 2781 8431
rect 3057 8427 3094 8459
rect 3265 8458 3514 8480
rect 3265 8427 3302 8458
rect 3478 8456 3514 8458
rect 3478 8427 3515 8456
rect 3827 8447 3864 8448
rect 4130 8447 4167 8517
rect 4192 8537 4279 8544
rect 4192 8534 4250 8537
rect 4192 8514 4197 8534
rect 4218 8517 4250 8534
rect 4270 8517 4279 8537
rect 4218 8514 4279 8517
rect 4192 8507 4279 8514
rect 4338 8537 4375 8547
rect 4338 8517 4346 8537
rect 4366 8517 4375 8537
rect 4192 8506 4223 8507
rect 3826 8446 4167 8447
rect 3751 8441 4167 8446
rect 2717 8418 2752 8419
rect 2694 8413 2752 8418
rect 2694 8393 2697 8413
rect 2717 8399 2752 8413
rect 2772 8399 2781 8419
rect 2717 8391 2781 8399
rect 2743 8390 2781 8391
rect 2744 8389 2781 8390
rect 2847 8423 2883 8424
rect 2955 8423 2991 8424
rect 2847 8415 2991 8423
rect 2847 8395 2855 8415
rect 2875 8395 2963 8415
rect 2983 8395 2991 8415
rect 2847 8389 2991 8395
rect 3057 8419 3095 8427
rect 3163 8423 3199 8424
rect 3057 8399 3066 8419
rect 3086 8399 3095 8419
rect 3057 8390 3095 8399
rect 3114 8416 3199 8423
rect 3114 8396 3121 8416
rect 3142 8415 3199 8416
rect 3142 8396 3171 8415
rect 3114 8395 3171 8396
rect 3191 8395 3199 8415
rect 3057 8389 3094 8390
rect 3114 8389 3199 8395
rect 3265 8419 3303 8427
rect 3376 8423 3412 8424
rect 3265 8399 3274 8419
rect 3294 8399 3303 8419
rect 3265 8390 3303 8399
rect 3327 8415 3412 8423
rect 3327 8395 3384 8415
rect 3404 8395 3412 8415
rect 3265 8389 3302 8390
rect 3327 8389 3412 8395
rect 3478 8419 3516 8427
rect 3751 8421 3754 8441
rect 3774 8421 4167 8441
rect 4338 8438 4375 8517
rect 4405 8546 4436 8599
rect 4786 8597 4823 8598
rect 4785 8588 4824 8597
rect 4785 8570 4795 8588
rect 4813 8570 4824 8588
rect 5165 8586 5202 8590
rect 4697 8553 4744 8554
rect 4785 8553 4824 8570
rect 4697 8549 4824 8553
rect 4455 8546 4492 8547
rect 4405 8537 4492 8546
rect 4405 8517 4463 8537
rect 4483 8517 4492 8537
rect 4405 8507 4492 8517
rect 4551 8537 4588 8547
rect 4551 8517 4559 8537
rect 4579 8517 4588 8537
rect 4405 8506 4436 8507
rect 4400 8438 4510 8451
rect 4551 8438 4588 8517
rect 4697 8520 4707 8549
rect 4736 8520 4824 8549
rect 4697 8514 4824 8520
rect 4697 8510 4744 8514
rect 4782 8500 4824 8514
rect 4782 8482 4793 8500
rect 4811 8482 4824 8500
rect 4782 8477 4824 8482
rect 4783 8474 4824 8477
rect 5162 8581 5202 8586
rect 5162 8563 5174 8581
rect 5192 8563 5202 8581
rect 4783 8473 4820 8474
rect 4338 8436 4588 8438
rect 4338 8433 4439 8436
rect 3478 8399 3487 8419
rect 3507 8399 3516 8419
rect 4338 8414 4403 8433
rect 3478 8390 3516 8399
rect 4400 8406 4403 8414
rect 4432 8406 4439 8433
rect 4467 8409 4477 8436
rect 4506 8414 4588 8436
rect 4506 8409 4510 8414
rect 4467 8406 4510 8409
rect 4400 8392 4510 8406
rect 4776 8410 4823 8411
rect 4776 8401 4824 8410
rect 3478 8389 3515 8390
rect 2901 8368 2937 8389
rect 3327 8368 3358 8389
rect 4776 8383 4795 8401
rect 4813 8383 4824 8401
rect 4776 8381 4824 8383
rect 2734 8364 2834 8368
rect 2734 8360 2796 8364
rect 2734 8334 2741 8360
rect 2767 8338 2796 8360
rect 2822 8338 2834 8364
rect 2767 8334 2834 8338
rect 2734 8331 2834 8334
rect 2902 8331 2937 8368
rect 2999 8365 3358 8368
rect 2999 8360 3221 8365
rect 2999 8336 3012 8360
rect 3036 8341 3221 8360
rect 3245 8341 3358 8365
rect 3036 8336 3358 8341
rect 2999 8332 3358 8336
rect 3425 8360 3574 8368
rect 3425 8340 3436 8360
rect 3456 8340 3574 8360
rect 3425 8333 3574 8340
rect 3425 8332 3466 8333
rect 2901 8292 2937 8331
rect 2749 8279 2786 8280
rect 2845 8279 2882 8280
rect 2901 8279 2908 8292
rect 2648 8270 2787 8279
rect 2648 8250 2758 8270
rect 2778 8250 2787 8270
rect 2648 8243 2787 8250
rect 2845 8270 2908 8279
rect 2845 8250 2854 8270
rect 2874 8254 2908 8270
rect 2931 8279 2937 8292
rect 2956 8279 2993 8280
rect 2931 8270 2993 8279
rect 2931 8254 2964 8270
rect 2874 8250 2964 8254
rect 2984 8250 2993 8270
rect 2648 8241 2745 8243
rect 2648 8240 2677 8241
rect 2845 8240 2993 8250
rect 3052 8270 3089 8280
rect 3164 8279 3201 8280
rect 3145 8277 3201 8279
rect 3052 8250 3060 8270
rect 3080 8250 3089 8270
rect 2901 8239 2937 8240
rect 2749 8180 2786 8181
rect 3052 8180 3089 8250
rect 3114 8270 3201 8277
rect 3114 8267 3172 8270
rect 3114 8247 3119 8267
rect 3140 8250 3172 8267
rect 3192 8250 3201 8270
rect 3140 8247 3201 8250
rect 3114 8240 3201 8247
rect 3260 8270 3297 8280
rect 3260 8250 3268 8270
rect 3288 8250 3297 8270
rect 3114 8239 3145 8240
rect 2748 8179 3089 8180
rect 2673 8175 3089 8179
rect 2673 8174 3050 8175
rect 2673 8154 2676 8174
rect 2696 8158 3050 8174
rect 3070 8158 3089 8175
rect 2696 8154 3089 8158
rect 3260 8171 3297 8250
rect 3327 8279 3358 8332
rect 4138 8324 4176 8326
rect 4785 8324 4824 8381
rect 4138 8291 4824 8324
rect 3377 8279 3414 8280
rect 3327 8270 3414 8279
rect 3327 8250 3385 8270
rect 3405 8250 3414 8270
rect 3327 8240 3414 8250
rect 3473 8270 3510 8280
rect 3473 8250 3481 8270
rect 3501 8250 3510 8270
rect 3327 8239 3358 8240
rect 3322 8171 3432 8184
rect 3473 8171 3510 8250
rect 3260 8169 3510 8171
rect 3260 8166 3361 8169
rect 3260 8147 3325 8166
rect 3322 8139 3325 8147
rect 3354 8139 3361 8166
rect 3389 8142 3399 8169
rect 3428 8147 3510 8169
rect 3730 8203 3898 8204
rect 4138 8203 4176 8291
rect 4437 8289 4484 8291
rect 4784 8267 4824 8291
rect 3730 8180 4176 8203
rect 4402 8234 4513 8249
rect 4402 8232 4444 8234
rect 4402 8212 4409 8232
rect 4428 8212 4444 8232
rect 4402 8204 4444 8212
rect 4472 8232 4513 8234
rect 4472 8212 4486 8232
rect 4505 8212 4513 8232
rect 4785 8223 4824 8267
rect 4472 8204 4513 8212
rect 4402 8198 4513 8204
rect 3730 8177 4174 8180
rect 3730 8175 3898 8177
rect 3428 8142 3432 8147
rect 3389 8139 3432 8142
rect 3322 8125 3432 8139
rect 2112 8106 2280 8108
rect 1833 8099 2280 8106
rect 1497 8079 1608 8085
rect 1497 8071 1538 8079
rect 915 8058 951 8059
rect 763 8028 772 8048
rect 792 8028 800 8048
rect 651 8019 707 8021
rect 651 8018 688 8019
rect 763 8018 800 8028
rect 859 8048 1007 8058
rect 1107 8055 1203 8057
rect 859 8028 868 8048
rect 888 8028 978 8048
rect 998 8028 1007 8048
rect 859 8019 1007 8028
rect 1065 8048 1203 8055
rect 1065 8028 1074 8048
rect 1094 8028 1203 8048
rect 1497 8051 1505 8071
rect 1524 8051 1538 8071
rect 1497 8049 1538 8051
rect 1566 8071 1608 8079
rect 1566 8051 1582 8071
rect 1601 8051 1608 8071
rect 1833 8072 1858 8099
rect 1889 8080 2280 8099
rect 1889 8072 1938 8080
rect 2112 8079 2280 8080
rect 1833 8070 1938 8072
rect 1566 8049 1608 8051
rect 1497 8034 1608 8049
rect 1065 8019 1203 8028
rect 859 8018 896 8019
rect 915 7967 951 8019
rect 970 8018 1007 8019
rect 1066 8018 1103 8019
rect 386 7965 427 7966
rect 278 7958 427 7965
rect 278 7938 396 7958
rect 416 7938 427 7958
rect 278 7930 427 7938
rect 494 7962 853 7966
rect 494 7957 816 7962
rect 494 7933 607 7957
rect 631 7938 816 7957
rect 840 7938 853 7962
rect 631 7933 853 7938
rect 494 7930 853 7933
rect 915 7930 950 7967
rect 1018 7964 1118 7967
rect 1018 7960 1085 7964
rect 1018 7934 1030 7960
rect 1056 7938 1085 7960
rect 1111 7938 1118 7964
rect 1056 7934 1118 7938
rect 1018 7930 1118 7934
rect 494 7909 525 7930
rect 915 7909 951 7930
rect 337 7908 374 7909
rect 111 7905 145 7906
rect 110 7896 147 7905
rect 110 7878 119 7896
rect 137 7878 147 7896
rect 110 7868 147 7878
rect 336 7899 374 7908
rect 336 7879 345 7899
rect 365 7879 374 7899
rect 336 7871 374 7879
rect 440 7903 525 7909
rect 550 7908 587 7909
rect 440 7883 448 7903
rect 468 7883 525 7903
rect 440 7875 525 7883
rect 549 7899 587 7908
rect 549 7879 558 7899
rect 578 7879 587 7899
rect 440 7874 476 7875
rect 549 7871 587 7879
rect 653 7903 738 7909
rect 758 7908 795 7909
rect 653 7883 661 7903
rect 681 7902 738 7903
rect 681 7883 710 7902
rect 653 7882 710 7883
rect 731 7882 738 7902
rect 653 7875 738 7882
rect 757 7899 795 7908
rect 757 7879 766 7899
rect 786 7879 795 7899
rect 653 7874 689 7875
rect 757 7871 795 7879
rect 861 7903 1005 7909
rect 861 7883 869 7903
rect 889 7902 977 7903
rect 889 7883 920 7902
rect 861 7882 920 7883
rect 945 7883 977 7902
rect 997 7883 1005 7903
rect 945 7882 1005 7883
rect 861 7875 1005 7882
rect 861 7874 897 7875
rect 969 7874 1005 7875
rect 1071 7908 1108 7909
rect 1071 7907 1109 7908
rect 1071 7899 1135 7907
rect 1071 7879 1080 7899
rect 1100 7885 1135 7899
rect 1155 7885 1158 7905
rect 1100 7880 1158 7885
rect 1100 7879 1135 7880
rect 111 7840 145 7868
rect 337 7842 374 7871
rect 338 7840 374 7842
rect 550 7840 587 7871
rect 111 7839 283 7840
rect 111 7807 297 7839
rect 338 7818 587 7840
rect 758 7839 795 7871
rect 1071 7867 1135 7879
rect 1175 7841 1202 8019
rect 3730 7997 3757 8175
rect 3797 8137 3861 8149
rect 4137 8145 4174 8177
rect 4345 8176 4594 8198
rect 4345 8145 4382 8176
rect 4558 8174 4594 8176
rect 4558 8145 4595 8174
rect 3797 8136 3832 8137
rect 3774 8131 3832 8136
rect 3774 8111 3777 8131
rect 3797 8117 3832 8131
rect 3852 8117 3861 8137
rect 3797 8109 3861 8117
rect 3823 8108 3861 8109
rect 3824 8107 3861 8108
rect 3927 8141 3963 8142
rect 4035 8141 4071 8142
rect 3927 8136 4071 8141
rect 3927 8133 3989 8136
rect 3927 8113 3935 8133
rect 3955 8116 3989 8133
rect 4012 8133 4071 8136
rect 4012 8116 4043 8133
rect 3955 8113 4043 8116
rect 4063 8113 4071 8133
rect 3927 8107 4071 8113
rect 4137 8137 4175 8145
rect 4243 8141 4279 8142
rect 4137 8117 4146 8137
rect 4166 8117 4175 8137
rect 4137 8108 4175 8117
rect 4194 8134 4279 8141
rect 4194 8114 4201 8134
rect 4222 8133 4279 8134
rect 4222 8114 4251 8133
rect 4194 8113 4251 8114
rect 4271 8113 4279 8133
rect 4137 8107 4174 8108
rect 4194 8107 4279 8113
rect 4345 8137 4383 8145
rect 4456 8141 4492 8142
rect 4345 8117 4354 8137
rect 4374 8117 4383 8137
rect 4345 8108 4383 8117
rect 4407 8133 4492 8141
rect 4407 8113 4464 8133
rect 4484 8113 4492 8133
rect 4345 8107 4382 8108
rect 4407 8107 4492 8113
rect 4558 8137 4596 8145
rect 4558 8117 4567 8137
rect 4587 8117 4596 8137
rect 4558 8108 4596 8117
rect 4558 8107 4595 8108
rect 3981 8086 4017 8107
rect 4407 8086 4438 8107
rect 3814 8082 3914 8086
rect 3814 8078 3876 8082
rect 3814 8052 3821 8078
rect 3847 8056 3876 8078
rect 3902 8056 3914 8082
rect 3847 8052 3914 8056
rect 3814 8049 3914 8052
rect 3982 8049 4017 8086
rect 4079 8083 4438 8086
rect 4079 8078 4301 8083
rect 4079 8054 4092 8078
rect 4116 8059 4301 8078
rect 4325 8059 4438 8083
rect 4116 8054 4438 8059
rect 4079 8050 4438 8054
rect 4505 8078 4654 8086
rect 4505 8058 4516 8078
rect 4536 8058 4654 8078
rect 4505 8051 4654 8058
rect 4505 8050 4546 8051
rect 3829 7997 3866 7998
rect 3925 7997 3962 7998
rect 3981 7997 4017 8049
rect 4036 7997 4073 7998
rect 3729 7988 3867 7997
rect 3729 7968 3838 7988
rect 3858 7968 3867 7988
rect 3729 7961 3867 7968
rect 3925 7988 4073 7997
rect 3925 7968 3934 7988
rect 3954 7968 4044 7988
rect 4064 7968 4073 7988
rect 3729 7959 3825 7961
rect 3925 7958 4073 7968
rect 4132 7988 4169 7998
rect 4244 7997 4281 7998
rect 4225 7995 4281 7997
rect 4132 7968 4140 7988
rect 4160 7968 4169 7988
rect 3981 7957 4017 7958
rect 1358 7915 1468 7929
rect 1358 7912 1401 7915
rect 1358 7907 1362 7912
rect 1034 7839 1202 7841
rect 758 7833 1202 7839
rect 111 7775 145 7807
rect 107 7766 145 7775
rect 107 7748 117 7766
rect 135 7748 145 7766
rect 107 7742 145 7748
rect 263 7744 297 7807
rect 419 7812 530 7818
rect 419 7804 460 7812
rect 419 7784 427 7804
rect 446 7784 460 7804
rect 419 7782 460 7784
rect 488 7804 530 7812
rect 488 7784 504 7804
rect 523 7784 530 7804
rect 488 7782 530 7784
rect 419 7767 530 7782
rect 757 7813 1202 7833
rect 757 7744 795 7813
rect 1034 7812 1202 7813
rect 1280 7885 1362 7907
rect 1391 7885 1401 7912
rect 1429 7888 1436 7915
rect 1465 7907 1468 7915
rect 3463 7924 3574 7939
rect 3463 7922 3505 7924
rect 1465 7888 1530 7907
rect 1429 7885 1530 7888
rect 1280 7883 1530 7885
rect 1280 7804 1317 7883
rect 1358 7870 1468 7883
rect 1432 7814 1463 7815
rect 1280 7784 1289 7804
rect 1309 7784 1317 7804
rect 1280 7774 1317 7784
rect 1376 7804 1463 7814
rect 1376 7784 1385 7804
rect 1405 7784 1463 7804
rect 1376 7775 1463 7784
rect 1376 7774 1413 7775
rect 107 7738 144 7742
rect 263 7733 795 7744
rect 262 7717 795 7733
rect 1432 7722 1463 7775
rect 1493 7804 1530 7883
rect 1701 7893 2094 7900
rect 1701 7876 1709 7893
rect 1741 7880 2094 7893
rect 2114 7880 2117 7900
rect 3196 7895 3237 7904
rect 1741 7876 2117 7880
rect 1701 7875 2117 7876
rect 2791 7893 2959 7894
rect 3196 7893 3205 7895
rect 1701 7874 2042 7875
rect 1645 7814 1676 7815
rect 1493 7784 1502 7804
rect 1522 7784 1530 7804
rect 1493 7774 1530 7784
rect 1589 7807 1676 7814
rect 1589 7804 1650 7807
rect 1589 7784 1598 7804
rect 1618 7787 1650 7804
rect 1671 7787 1676 7807
rect 1618 7784 1676 7787
rect 1589 7777 1676 7784
rect 1701 7804 1738 7874
rect 2004 7873 2041 7874
rect 2791 7873 3205 7893
rect 3231 7873 3237 7895
rect 3463 7902 3470 7922
rect 3489 7902 3505 7922
rect 3463 7894 3505 7902
rect 3533 7922 3574 7924
rect 3533 7902 3547 7922
rect 3566 7902 3574 7922
rect 3533 7894 3574 7902
rect 3829 7898 3866 7899
rect 4132 7898 4169 7968
rect 4194 7988 4281 7995
rect 4194 7985 4252 7988
rect 4194 7965 4199 7985
rect 4220 7968 4252 7985
rect 4272 7968 4281 7988
rect 4220 7965 4281 7968
rect 4194 7958 4281 7965
rect 4340 7988 4377 7998
rect 4340 7968 4348 7988
rect 4368 7968 4377 7988
rect 4194 7957 4225 7958
rect 3828 7897 4169 7898
rect 3463 7888 3574 7894
rect 3753 7892 4169 7897
rect 2791 7867 3237 7873
rect 2791 7865 2959 7867
rect 1853 7814 1889 7815
rect 1701 7784 1710 7804
rect 1730 7784 1738 7804
rect 1589 7775 1645 7777
rect 1589 7774 1626 7775
rect 1701 7774 1738 7784
rect 1797 7804 1945 7814
rect 2045 7811 2141 7813
rect 1797 7784 1806 7804
rect 1826 7799 1916 7804
rect 1826 7784 1861 7799
rect 1797 7775 1861 7784
rect 1797 7774 1834 7775
rect 1853 7758 1861 7775
rect 1882 7784 1916 7799
rect 1936 7784 1945 7804
rect 1882 7775 1945 7784
rect 2003 7804 2141 7811
rect 2003 7784 2012 7804
rect 2032 7784 2141 7804
rect 2003 7775 2141 7784
rect 1882 7758 1889 7775
rect 1908 7774 1945 7775
rect 2004 7774 2041 7775
rect 1853 7723 1889 7758
rect 1324 7721 1365 7722
rect 262 7716 776 7717
rect 1216 7714 1365 7721
rect 1216 7694 1334 7714
rect 1354 7694 1365 7714
rect 1216 7686 1365 7694
rect 1432 7718 1791 7722
rect 1432 7713 1754 7718
rect 1432 7689 1545 7713
rect 1569 7694 1754 7713
rect 1778 7694 1791 7718
rect 1569 7689 1791 7694
rect 1432 7686 1791 7689
rect 1853 7686 1888 7723
rect 1956 7720 2056 7723
rect 1956 7716 2023 7720
rect 1956 7690 1968 7716
rect 1994 7694 2023 7716
rect 2049 7694 2056 7720
rect 1994 7690 2056 7694
rect 1956 7686 2056 7690
rect 110 7675 147 7676
rect 108 7667 148 7675
rect 108 7649 119 7667
rect 137 7649 148 7667
rect 1432 7665 1463 7686
rect 1853 7665 1889 7686
rect 1275 7664 1312 7665
rect 108 7601 148 7649
rect 1274 7655 1312 7664
rect 1274 7635 1283 7655
rect 1303 7635 1312 7655
rect 1274 7627 1312 7635
rect 1378 7659 1463 7665
rect 1488 7664 1525 7665
rect 1378 7639 1386 7659
rect 1406 7639 1463 7659
rect 1378 7631 1463 7639
rect 1487 7655 1525 7664
rect 1487 7635 1496 7655
rect 1516 7635 1525 7655
rect 1378 7630 1414 7631
rect 1487 7627 1525 7635
rect 1591 7659 1676 7665
rect 1696 7664 1733 7665
rect 1591 7639 1599 7659
rect 1619 7658 1676 7659
rect 1619 7639 1648 7658
rect 1591 7638 1648 7639
rect 1669 7638 1676 7658
rect 1591 7631 1676 7638
rect 1695 7655 1733 7664
rect 1695 7635 1704 7655
rect 1724 7635 1733 7655
rect 1591 7630 1627 7631
rect 1695 7627 1733 7635
rect 1799 7659 1943 7665
rect 1799 7639 1807 7659
rect 1827 7639 1915 7659
rect 1935 7639 1943 7659
rect 1799 7631 1943 7639
rect 1799 7630 1835 7631
rect 1907 7630 1943 7631
rect 2009 7664 2046 7665
rect 2009 7663 2047 7664
rect 2009 7655 2073 7663
rect 2009 7635 2018 7655
rect 2038 7641 2073 7655
rect 2093 7641 2096 7661
rect 2038 7636 2096 7641
rect 2038 7635 2073 7636
rect 419 7605 529 7619
rect 419 7602 462 7605
rect 108 7594 233 7601
rect 419 7597 423 7602
rect 108 7575 200 7594
rect 225 7575 233 7594
rect 108 7565 233 7575
rect 341 7575 423 7597
rect 452 7575 462 7602
rect 490 7578 497 7605
rect 526 7597 529 7605
rect 1275 7598 1312 7627
rect 526 7578 591 7597
rect 1276 7596 1312 7598
rect 1488 7596 1525 7627
rect 1696 7600 1733 7627
rect 2009 7623 2073 7635
rect 490 7575 591 7578
rect 341 7573 591 7575
rect 108 7545 148 7565
rect 107 7536 148 7545
rect 107 7518 117 7536
rect 135 7518 148 7536
rect 107 7509 148 7518
rect 107 7508 144 7509
rect 341 7494 378 7573
rect 419 7560 529 7573
rect 493 7504 524 7505
rect 341 7474 350 7494
rect 370 7474 378 7494
rect 341 7464 378 7474
rect 437 7494 524 7504
rect 437 7474 446 7494
rect 466 7474 524 7494
rect 437 7465 524 7474
rect 437 7464 474 7465
rect 110 7442 147 7446
rect 107 7437 147 7442
rect 107 7419 119 7437
rect 137 7419 147 7437
rect 107 7239 147 7419
rect 493 7412 524 7465
rect 554 7494 591 7573
rect 762 7570 1155 7590
rect 1175 7570 1178 7590
rect 1276 7574 1525 7596
rect 1694 7595 1735 7600
rect 2113 7597 2140 7775
rect 2791 7687 2818 7865
rect 3196 7862 3237 7867
rect 3406 7866 3655 7888
rect 3753 7872 3756 7892
rect 3776 7872 4169 7892
rect 4340 7889 4377 7968
rect 4407 7997 4438 8050
rect 4784 8043 4824 8223
rect 5162 8383 5202 8563
rect 5548 8556 5579 8609
rect 5609 8638 5646 8717
rect 5817 8714 6210 8734
rect 6230 8714 6233 8734
rect 6331 8718 6580 8740
rect 6749 8739 6790 8744
rect 7168 8741 7195 8919
rect 7846 8831 7873 9009
rect 8251 9006 8292 9011
rect 8461 9010 8710 9032
rect 8808 9016 8811 9036
rect 8831 9016 9224 9036
rect 9395 9033 9432 9112
rect 9462 9141 9493 9194
rect 9839 9187 9879 9367
rect 9839 9169 9849 9187
rect 9867 9169 9879 9187
rect 9839 9164 9879 9169
rect 9839 9160 9876 9164
rect 9512 9141 9549 9142
rect 9462 9132 9549 9141
rect 9462 9112 9520 9132
rect 9540 9112 9549 9132
rect 9462 9102 9549 9112
rect 9608 9132 9645 9142
rect 9608 9112 9616 9132
rect 9636 9112 9645 9132
rect 9462 9101 9493 9102
rect 9457 9033 9567 9046
rect 9608 9033 9645 9112
rect 9842 9097 9879 9098
rect 9838 9088 9879 9097
rect 9838 9070 9851 9088
rect 9869 9070 9879 9088
rect 9838 9061 9879 9070
rect 9838 9041 9878 9061
rect 9395 9031 9645 9033
rect 9395 9028 9496 9031
rect 7913 8971 7977 8983
rect 8253 8979 8290 9006
rect 8461 8979 8498 9010
rect 8674 9008 8710 9010
rect 9395 9009 9460 9028
rect 8674 8979 8711 9008
rect 9457 9001 9460 9009
rect 9489 9001 9496 9028
rect 9524 9004 9534 9031
rect 9563 9009 9645 9031
rect 9753 9031 9878 9041
rect 9753 9012 9761 9031
rect 9786 9012 9878 9031
rect 9563 9004 9567 9009
rect 9753 9005 9878 9012
rect 9524 9001 9567 9004
rect 9457 8987 9567 9001
rect 7913 8970 7948 8971
rect 7890 8965 7948 8970
rect 7890 8945 7893 8965
rect 7913 8951 7948 8965
rect 7968 8951 7977 8971
rect 7913 8943 7977 8951
rect 7939 8942 7977 8943
rect 7940 8941 7977 8942
rect 8043 8975 8079 8976
rect 8151 8975 8187 8976
rect 8043 8967 8187 8975
rect 8043 8947 8051 8967
rect 8071 8947 8159 8967
rect 8179 8947 8187 8967
rect 8043 8941 8187 8947
rect 8253 8971 8291 8979
rect 8359 8975 8395 8976
rect 8253 8951 8262 8971
rect 8282 8951 8291 8971
rect 8253 8942 8291 8951
rect 8310 8968 8395 8975
rect 8310 8948 8317 8968
rect 8338 8967 8395 8968
rect 8338 8948 8367 8967
rect 8310 8947 8367 8948
rect 8387 8947 8395 8967
rect 8253 8941 8290 8942
rect 8310 8941 8395 8947
rect 8461 8971 8499 8979
rect 8572 8975 8608 8976
rect 8461 8951 8470 8971
rect 8490 8951 8499 8971
rect 8461 8942 8499 8951
rect 8523 8967 8608 8975
rect 8523 8947 8580 8967
rect 8600 8947 8608 8967
rect 8461 8941 8498 8942
rect 8523 8941 8608 8947
rect 8674 8971 8712 8979
rect 8674 8951 8683 8971
rect 8703 8951 8712 8971
rect 8674 8942 8712 8951
rect 9838 8957 9878 9005
rect 8674 8941 8711 8942
rect 8097 8920 8133 8941
rect 8523 8920 8554 8941
rect 9838 8939 9849 8957
rect 9867 8939 9878 8957
rect 9838 8931 9878 8939
rect 9839 8930 9876 8931
rect 7930 8916 8030 8920
rect 7930 8912 7992 8916
rect 7930 8886 7937 8912
rect 7963 8890 7992 8912
rect 8018 8890 8030 8916
rect 7963 8886 8030 8890
rect 7930 8883 8030 8886
rect 8098 8883 8133 8920
rect 8195 8917 8554 8920
rect 8195 8912 8417 8917
rect 8195 8888 8208 8912
rect 8232 8893 8417 8912
rect 8441 8893 8554 8917
rect 8232 8888 8554 8893
rect 8195 8884 8554 8888
rect 8621 8912 8770 8920
rect 8621 8892 8632 8912
rect 8652 8892 8770 8912
rect 8621 8885 8770 8892
rect 9210 8889 9724 8890
rect 8621 8884 8662 8885
rect 8097 8848 8133 8883
rect 7945 8831 7982 8832
rect 8041 8831 8078 8832
rect 8097 8831 8104 8848
rect 7845 8822 7983 8831
rect 7845 8802 7954 8822
rect 7974 8802 7983 8822
rect 7845 8795 7983 8802
rect 8041 8822 8104 8831
rect 8041 8802 8050 8822
rect 8070 8807 8104 8822
rect 8125 8831 8133 8848
rect 8152 8831 8189 8832
rect 8125 8822 8189 8831
rect 8125 8807 8160 8822
rect 8070 8802 8160 8807
rect 8180 8802 8189 8822
rect 7845 8793 7941 8795
rect 8041 8792 8189 8802
rect 8248 8822 8285 8832
rect 8360 8831 8397 8832
rect 8341 8829 8397 8831
rect 8248 8802 8256 8822
rect 8276 8802 8285 8822
rect 8097 8791 8133 8792
rect 7027 8739 7195 8741
rect 6749 8733 7195 8739
rect 5817 8709 6233 8714
rect 6412 8712 6523 8718
rect 5817 8708 6158 8709
rect 5761 8648 5792 8649
rect 5609 8618 5618 8638
rect 5638 8618 5646 8638
rect 5609 8608 5646 8618
rect 5705 8641 5792 8648
rect 5705 8638 5766 8641
rect 5705 8618 5714 8638
rect 5734 8621 5766 8638
rect 5787 8621 5792 8641
rect 5734 8618 5792 8621
rect 5705 8611 5792 8618
rect 5817 8638 5854 8708
rect 6120 8707 6157 8708
rect 6412 8704 6453 8712
rect 6412 8684 6420 8704
rect 6439 8684 6453 8704
rect 6412 8682 6453 8684
rect 6481 8704 6523 8712
rect 6481 8684 6497 8704
rect 6516 8684 6523 8704
rect 6749 8711 6755 8733
rect 6781 8713 7195 8733
rect 7945 8732 7982 8733
rect 8248 8732 8285 8802
rect 8310 8822 8397 8829
rect 8310 8819 8368 8822
rect 8310 8799 8315 8819
rect 8336 8802 8368 8819
rect 8388 8802 8397 8822
rect 8336 8799 8397 8802
rect 8310 8792 8397 8799
rect 8456 8822 8493 8832
rect 8456 8802 8464 8822
rect 8484 8802 8493 8822
rect 8310 8791 8341 8792
rect 7944 8731 8285 8732
rect 6781 8711 6790 8713
rect 7027 8712 7195 8713
rect 7869 8730 8285 8731
rect 7869 8726 8245 8730
rect 6749 8702 6790 8711
rect 7869 8706 7872 8726
rect 7892 8713 8245 8726
rect 8277 8713 8285 8730
rect 7892 8706 8285 8713
rect 8456 8723 8493 8802
rect 8523 8831 8554 8884
rect 9191 8873 9724 8889
rect 9191 8862 9723 8873
rect 9842 8864 9879 8868
rect 8573 8831 8610 8832
rect 8523 8822 8610 8831
rect 8523 8802 8581 8822
rect 8601 8802 8610 8822
rect 8523 8792 8610 8802
rect 8669 8822 8706 8832
rect 8669 8802 8677 8822
rect 8697 8802 8706 8822
rect 8523 8791 8554 8792
rect 8518 8723 8628 8736
rect 8669 8723 8706 8802
rect 8456 8721 8706 8723
rect 8456 8718 8557 8721
rect 8456 8699 8521 8718
rect 6481 8682 6523 8684
rect 6412 8667 6523 8682
rect 8518 8691 8521 8699
rect 8550 8691 8557 8718
rect 8585 8694 8595 8721
rect 8624 8699 8706 8721
rect 8784 8793 8952 8794
rect 9191 8793 9229 8862
rect 8784 8773 9229 8793
rect 9456 8824 9567 8839
rect 9456 8822 9498 8824
rect 9456 8802 9463 8822
rect 9482 8802 9498 8822
rect 9456 8794 9498 8802
rect 9526 8822 9567 8824
rect 9526 8802 9540 8822
rect 9559 8802 9567 8822
rect 9526 8794 9567 8802
rect 9456 8788 9567 8794
rect 9689 8799 9723 8862
rect 9841 8858 9879 8864
rect 9841 8840 9851 8858
rect 9869 8840 9879 8858
rect 9841 8831 9879 8840
rect 9841 8799 9875 8831
rect 8784 8767 9228 8773
rect 8784 8765 8952 8767
rect 8624 8694 8628 8699
rect 8585 8691 8628 8694
rect 8518 8677 8628 8691
rect 5969 8648 6005 8649
rect 5817 8618 5826 8638
rect 5846 8618 5854 8638
rect 5705 8609 5761 8611
rect 5705 8608 5742 8609
rect 5817 8608 5854 8618
rect 5913 8638 6061 8648
rect 6161 8645 6257 8647
rect 5913 8618 5922 8638
rect 5942 8618 6032 8638
rect 6052 8618 6061 8638
rect 5913 8609 6061 8618
rect 6119 8638 6257 8645
rect 6119 8618 6128 8638
rect 6148 8618 6257 8638
rect 6119 8609 6257 8618
rect 5913 8608 5950 8609
rect 5969 8557 6005 8609
rect 6024 8608 6061 8609
rect 6120 8608 6157 8609
rect 5440 8555 5481 8556
rect 5332 8548 5481 8555
rect 5332 8528 5450 8548
rect 5470 8528 5481 8548
rect 5332 8520 5481 8528
rect 5548 8552 5907 8556
rect 5548 8547 5870 8552
rect 5548 8523 5661 8547
rect 5685 8528 5870 8547
rect 5894 8528 5907 8552
rect 5685 8523 5907 8528
rect 5548 8520 5907 8523
rect 5969 8520 6004 8557
rect 6072 8554 6172 8557
rect 6072 8550 6139 8554
rect 6072 8524 6084 8550
rect 6110 8528 6139 8550
rect 6165 8528 6172 8554
rect 6110 8524 6172 8528
rect 6072 8520 6172 8524
rect 5548 8499 5579 8520
rect 5969 8499 6005 8520
rect 5391 8498 5428 8499
rect 5390 8489 5428 8498
rect 5390 8469 5399 8489
rect 5419 8469 5428 8489
rect 5390 8461 5428 8469
rect 5494 8493 5579 8499
rect 5604 8498 5641 8499
rect 5494 8473 5502 8493
rect 5522 8473 5579 8493
rect 5494 8465 5579 8473
rect 5603 8489 5641 8498
rect 5603 8469 5612 8489
rect 5632 8469 5641 8489
rect 5494 8464 5530 8465
rect 5603 8461 5641 8469
rect 5707 8493 5792 8499
rect 5812 8498 5849 8499
rect 5707 8473 5715 8493
rect 5735 8492 5792 8493
rect 5735 8473 5764 8492
rect 5707 8472 5764 8473
rect 5785 8472 5792 8492
rect 5707 8465 5792 8472
rect 5811 8489 5849 8498
rect 5811 8469 5820 8489
rect 5840 8469 5849 8489
rect 5707 8464 5743 8465
rect 5811 8461 5849 8469
rect 5915 8493 6059 8499
rect 5915 8473 5923 8493
rect 5943 8490 6031 8493
rect 5943 8473 5974 8490
rect 5915 8470 5974 8473
rect 5997 8473 6031 8490
rect 6051 8473 6059 8493
rect 5997 8470 6059 8473
rect 5915 8465 6059 8470
rect 5915 8464 5951 8465
rect 6023 8464 6059 8465
rect 6125 8498 6162 8499
rect 6125 8497 6163 8498
rect 6125 8489 6189 8497
rect 6125 8469 6134 8489
rect 6154 8475 6189 8489
rect 6209 8475 6212 8495
rect 6154 8470 6212 8475
rect 6154 8469 6189 8470
rect 5391 8432 5428 8461
rect 5392 8430 5428 8432
rect 5604 8430 5641 8461
rect 5392 8408 5641 8430
rect 5812 8429 5849 8461
rect 6125 8457 6189 8469
rect 6229 8431 6256 8609
rect 8784 8587 8811 8765
rect 8851 8727 8915 8739
rect 9191 8735 9228 8767
rect 9399 8766 9648 8788
rect 9689 8767 9875 8799
rect 9703 8766 9875 8767
rect 9399 8735 9436 8766
rect 9612 8764 9648 8766
rect 9612 8735 9649 8764
rect 9841 8738 9875 8766
rect 8851 8726 8886 8727
rect 8828 8721 8886 8726
rect 8828 8701 8831 8721
rect 8851 8707 8886 8721
rect 8906 8707 8915 8727
rect 8851 8699 8915 8707
rect 8877 8698 8915 8699
rect 8878 8697 8915 8698
rect 8981 8731 9017 8732
rect 9089 8731 9125 8732
rect 8981 8724 9125 8731
rect 8981 8723 9041 8724
rect 8981 8703 8989 8723
rect 9009 8704 9041 8723
rect 9066 8723 9125 8724
rect 9066 8704 9097 8723
rect 9009 8703 9097 8704
rect 9117 8703 9125 8723
rect 8981 8697 9125 8703
rect 9191 8727 9229 8735
rect 9297 8731 9333 8732
rect 9191 8707 9200 8727
rect 9220 8707 9229 8727
rect 9191 8698 9229 8707
rect 9248 8724 9333 8731
rect 9248 8704 9255 8724
rect 9276 8723 9333 8724
rect 9276 8704 9305 8723
rect 9248 8703 9305 8704
rect 9325 8703 9333 8723
rect 9191 8697 9228 8698
rect 9248 8697 9333 8703
rect 9399 8727 9437 8735
rect 9510 8731 9546 8732
rect 9399 8707 9408 8727
rect 9428 8707 9437 8727
rect 9399 8698 9437 8707
rect 9461 8723 9546 8731
rect 9461 8703 9518 8723
rect 9538 8703 9546 8723
rect 9399 8697 9436 8698
rect 9461 8697 9546 8703
rect 9612 8727 9650 8735
rect 9612 8707 9621 8727
rect 9641 8707 9650 8727
rect 9612 8698 9650 8707
rect 9839 8728 9876 8738
rect 9839 8710 9849 8728
rect 9867 8710 9876 8728
rect 9839 8701 9876 8710
rect 9841 8700 9875 8701
rect 9612 8697 9649 8698
rect 9035 8676 9071 8697
rect 9461 8676 9492 8697
rect 8868 8672 8968 8676
rect 8868 8668 8930 8672
rect 8868 8642 8875 8668
rect 8901 8646 8930 8668
rect 8956 8646 8968 8672
rect 8901 8642 8968 8646
rect 8868 8639 8968 8642
rect 9036 8639 9071 8676
rect 9133 8673 9492 8676
rect 9133 8668 9355 8673
rect 9133 8644 9146 8668
rect 9170 8649 9355 8668
rect 9379 8649 9492 8673
rect 9170 8644 9492 8649
rect 9133 8640 9492 8644
rect 9559 8668 9708 8676
rect 9559 8648 9570 8668
rect 9590 8648 9708 8668
rect 9559 8641 9708 8648
rect 9559 8640 9600 8641
rect 8883 8587 8920 8588
rect 8979 8587 9016 8588
rect 9035 8587 9071 8639
rect 9090 8587 9127 8588
rect 8783 8578 8921 8587
rect 8378 8557 8489 8572
rect 8378 8555 8420 8557
rect 8048 8534 8153 8536
rect 7704 8526 7874 8527
rect 8048 8526 8097 8534
rect 7704 8507 8097 8526
rect 8128 8507 8153 8534
rect 8378 8535 8385 8555
rect 8404 8535 8420 8555
rect 8378 8527 8420 8535
rect 8448 8555 8489 8557
rect 8448 8535 8462 8555
rect 8481 8535 8489 8555
rect 8783 8558 8892 8578
rect 8912 8558 8921 8578
rect 8783 8551 8921 8558
rect 8979 8578 9127 8587
rect 8979 8558 8988 8578
rect 9008 8558 9098 8578
rect 9118 8558 9127 8578
rect 8783 8549 8879 8551
rect 8979 8548 9127 8558
rect 9186 8578 9223 8588
rect 9298 8587 9335 8588
rect 9279 8585 9335 8587
rect 9186 8558 9194 8578
rect 9214 8558 9223 8578
rect 9035 8547 9071 8548
rect 8448 8527 8489 8535
rect 8378 8521 8489 8527
rect 7704 8500 8153 8507
rect 7704 8498 7874 8500
rect 6554 8467 6664 8481
rect 6554 8464 6597 8467
rect 6554 8459 6558 8464
rect 6088 8429 6256 8431
rect 5812 8426 6256 8429
rect 5473 8402 5584 8408
rect 5473 8394 5514 8402
rect 5162 8339 5201 8383
rect 5473 8374 5481 8394
rect 5500 8374 5514 8394
rect 5473 8372 5514 8374
rect 5542 8394 5584 8402
rect 5542 8374 5558 8394
rect 5577 8374 5584 8394
rect 5542 8372 5584 8374
rect 5473 8357 5584 8372
rect 5810 8403 6256 8426
rect 5162 8315 5202 8339
rect 5502 8315 5549 8317
rect 5810 8315 5848 8403
rect 6088 8402 6256 8403
rect 6476 8437 6558 8459
rect 6587 8437 6597 8464
rect 6625 8440 6632 8467
rect 6661 8459 6664 8467
rect 6661 8440 6726 8459
rect 6625 8437 6726 8440
rect 6476 8435 6726 8437
rect 6476 8356 6513 8435
rect 6554 8422 6664 8435
rect 6628 8366 6659 8367
rect 6476 8336 6485 8356
rect 6505 8336 6513 8356
rect 6476 8326 6513 8336
rect 6572 8356 6659 8366
rect 6572 8336 6581 8356
rect 6601 8336 6659 8356
rect 6572 8327 6659 8336
rect 6572 8326 6609 8327
rect 5162 8282 5848 8315
rect 5162 8225 5201 8282
rect 5810 8280 5848 8282
rect 6628 8274 6659 8327
rect 6689 8356 6726 8435
rect 6897 8448 7290 8452
rect 6897 8431 6916 8448
rect 6936 8432 7290 8448
rect 7310 8432 7313 8452
rect 6936 8431 7313 8432
rect 6897 8427 7313 8431
rect 6897 8426 7238 8427
rect 6841 8366 6872 8367
rect 6689 8336 6698 8356
rect 6718 8336 6726 8356
rect 6689 8326 6726 8336
rect 6785 8359 6872 8366
rect 6785 8356 6846 8359
rect 6785 8336 6794 8356
rect 6814 8339 6846 8356
rect 6867 8339 6872 8359
rect 6814 8336 6872 8339
rect 6785 8329 6872 8336
rect 6897 8356 6934 8426
rect 7200 8425 7237 8426
rect 7049 8366 7085 8367
rect 6897 8336 6906 8356
rect 6926 8336 6934 8356
rect 6785 8327 6841 8329
rect 6785 8326 6822 8327
rect 6897 8326 6934 8336
rect 6993 8356 7141 8366
rect 7241 8363 7337 8365
rect 6993 8336 7002 8356
rect 7022 8336 7112 8356
rect 7132 8336 7141 8356
rect 6993 8327 7141 8336
rect 7199 8356 7337 8363
rect 7199 8336 7208 8356
rect 7228 8336 7337 8356
rect 7199 8327 7337 8336
rect 6993 8326 7030 8327
rect 7049 8275 7085 8327
rect 7104 8326 7141 8327
rect 7200 8326 7237 8327
rect 6520 8273 6561 8274
rect 6412 8266 6561 8273
rect 6412 8246 6530 8266
rect 6550 8246 6561 8266
rect 6412 8238 6561 8246
rect 6628 8270 6987 8274
rect 6628 8265 6950 8270
rect 6628 8241 6741 8265
rect 6765 8246 6950 8265
rect 6974 8246 6987 8270
rect 6765 8241 6987 8246
rect 6628 8238 6987 8241
rect 7049 8238 7084 8275
rect 7152 8272 7252 8275
rect 7152 8268 7219 8272
rect 7152 8242 7164 8268
rect 7190 8246 7219 8268
rect 7245 8246 7252 8272
rect 7190 8242 7252 8246
rect 7152 8238 7252 8242
rect 5162 8223 5210 8225
rect 5162 8205 5173 8223
rect 5191 8205 5210 8223
rect 6628 8217 6659 8238
rect 7049 8217 7085 8238
rect 6471 8216 6508 8217
rect 5162 8196 5210 8205
rect 5163 8195 5210 8196
rect 5476 8200 5586 8214
rect 5476 8197 5519 8200
rect 5476 8192 5480 8197
rect 5398 8170 5480 8192
rect 5509 8170 5519 8197
rect 5547 8173 5554 8200
rect 5583 8192 5586 8200
rect 6470 8207 6508 8216
rect 5583 8173 5648 8192
rect 6470 8187 6479 8207
rect 6499 8187 6508 8207
rect 5547 8170 5648 8173
rect 5398 8168 5648 8170
rect 5166 8132 5203 8133
rect 4784 8025 4794 8043
rect 4812 8025 4824 8043
rect 4784 8020 4824 8025
rect 5162 8129 5203 8132
rect 5162 8124 5204 8129
rect 5162 8106 5175 8124
rect 5193 8106 5204 8124
rect 5162 8092 5204 8106
rect 5242 8092 5289 8096
rect 5162 8086 5289 8092
rect 5162 8057 5250 8086
rect 5279 8057 5289 8086
rect 5398 8089 5435 8168
rect 5476 8155 5586 8168
rect 5550 8099 5581 8100
rect 5398 8069 5407 8089
rect 5427 8069 5435 8089
rect 5398 8059 5435 8069
rect 5494 8089 5581 8099
rect 5494 8069 5503 8089
rect 5523 8069 5581 8089
rect 5494 8060 5581 8069
rect 5494 8059 5531 8060
rect 5162 8053 5289 8057
rect 5162 8036 5201 8053
rect 5242 8052 5289 8053
rect 4784 8016 4821 8020
rect 5162 8018 5173 8036
rect 5191 8018 5201 8036
rect 5162 8009 5201 8018
rect 5163 8008 5200 8009
rect 5550 8007 5581 8060
rect 5611 8089 5648 8168
rect 5819 8165 6212 8185
rect 6232 8165 6235 8185
rect 6470 8179 6508 8187
rect 6574 8211 6659 8217
rect 6684 8216 6721 8217
rect 6574 8191 6582 8211
rect 6602 8191 6659 8211
rect 6574 8183 6659 8191
rect 6683 8207 6721 8216
rect 6683 8187 6692 8207
rect 6712 8187 6721 8207
rect 6574 8182 6610 8183
rect 6683 8179 6721 8187
rect 6787 8211 6872 8217
rect 6892 8216 6929 8217
rect 6787 8191 6795 8211
rect 6815 8210 6872 8211
rect 6815 8191 6844 8210
rect 6787 8190 6844 8191
rect 6865 8190 6872 8210
rect 6787 8183 6872 8190
rect 6891 8207 6929 8216
rect 6891 8187 6900 8207
rect 6920 8187 6929 8207
rect 6787 8182 6823 8183
rect 6891 8179 6929 8187
rect 6995 8211 7139 8217
rect 6995 8191 7003 8211
rect 7023 8209 7111 8211
rect 7023 8191 7052 8209
rect 6995 8188 7052 8191
rect 7079 8191 7111 8209
rect 7131 8191 7139 8211
rect 7079 8188 7139 8191
rect 6995 8183 7139 8188
rect 6995 8182 7031 8183
rect 7103 8182 7139 8183
rect 7205 8216 7242 8217
rect 7205 8215 7243 8216
rect 7205 8207 7269 8215
rect 7205 8187 7214 8207
rect 7234 8193 7269 8207
rect 7289 8193 7292 8213
rect 7234 8188 7292 8193
rect 7234 8187 7269 8188
rect 5819 8160 6235 8165
rect 5819 8159 6160 8160
rect 5763 8099 5794 8100
rect 5611 8069 5620 8089
rect 5640 8069 5648 8089
rect 5611 8059 5648 8069
rect 5707 8092 5794 8099
rect 5707 8089 5768 8092
rect 5707 8069 5716 8089
rect 5736 8072 5768 8089
rect 5789 8072 5794 8092
rect 5736 8069 5794 8072
rect 5707 8062 5794 8069
rect 5819 8089 5856 8159
rect 6122 8158 6159 8159
rect 6471 8150 6508 8179
rect 6472 8148 6508 8150
rect 6684 8148 6721 8179
rect 6472 8126 6721 8148
rect 6892 8147 6929 8179
rect 7205 8175 7269 8187
rect 7309 8149 7336 8327
rect 7704 8320 7733 8498
rect 7773 8460 7837 8472
rect 8113 8468 8150 8500
rect 8321 8499 8570 8521
rect 8321 8468 8358 8499
rect 8534 8497 8570 8499
rect 8534 8468 8571 8497
rect 8883 8488 8920 8489
rect 9186 8488 9223 8558
rect 9248 8578 9335 8585
rect 9248 8575 9306 8578
rect 9248 8555 9253 8575
rect 9274 8558 9306 8575
rect 9326 8558 9335 8578
rect 9274 8555 9335 8558
rect 9248 8548 9335 8555
rect 9394 8578 9431 8588
rect 9394 8558 9402 8578
rect 9422 8558 9431 8578
rect 9248 8547 9279 8548
rect 8882 8487 9223 8488
rect 8807 8482 9223 8487
rect 7773 8459 7808 8460
rect 7750 8454 7808 8459
rect 7750 8434 7753 8454
rect 7773 8440 7808 8454
rect 7828 8440 7837 8460
rect 7773 8432 7837 8440
rect 7799 8431 7837 8432
rect 7800 8430 7837 8431
rect 7903 8464 7939 8465
rect 8011 8464 8047 8465
rect 7903 8456 8047 8464
rect 7903 8436 7911 8456
rect 7931 8436 8019 8456
rect 8039 8436 8047 8456
rect 7903 8430 8047 8436
rect 8113 8460 8151 8468
rect 8219 8464 8255 8465
rect 8113 8440 8122 8460
rect 8142 8440 8151 8460
rect 8113 8431 8151 8440
rect 8170 8457 8255 8464
rect 8170 8437 8177 8457
rect 8198 8456 8255 8457
rect 8198 8437 8227 8456
rect 8170 8436 8227 8437
rect 8247 8436 8255 8456
rect 8113 8430 8150 8431
rect 8170 8430 8255 8436
rect 8321 8460 8359 8468
rect 8432 8464 8468 8465
rect 8321 8440 8330 8460
rect 8350 8440 8359 8460
rect 8321 8431 8359 8440
rect 8383 8456 8468 8464
rect 8383 8436 8440 8456
rect 8460 8436 8468 8456
rect 8321 8430 8358 8431
rect 8383 8430 8468 8436
rect 8534 8460 8572 8468
rect 8807 8462 8810 8482
rect 8830 8462 9223 8482
rect 9394 8479 9431 8558
rect 9461 8587 9492 8640
rect 9842 8638 9879 8639
rect 9841 8629 9880 8638
rect 9841 8611 9851 8629
rect 9869 8611 9880 8629
rect 9753 8594 9800 8595
rect 9841 8594 9880 8611
rect 9753 8590 9880 8594
rect 9511 8587 9548 8588
rect 9461 8578 9548 8587
rect 9461 8558 9519 8578
rect 9539 8558 9548 8578
rect 9461 8548 9548 8558
rect 9607 8578 9644 8588
rect 9607 8558 9615 8578
rect 9635 8558 9644 8578
rect 9461 8547 9492 8548
rect 9456 8479 9566 8492
rect 9607 8479 9644 8558
rect 9753 8561 9763 8590
rect 9792 8561 9880 8590
rect 9753 8555 9880 8561
rect 9753 8551 9800 8555
rect 9838 8541 9880 8555
rect 9838 8523 9849 8541
rect 9867 8523 9880 8541
rect 9838 8518 9880 8523
rect 9839 8515 9880 8518
rect 9839 8514 9876 8515
rect 9394 8477 9644 8479
rect 9394 8474 9495 8477
rect 8534 8440 8543 8460
rect 8563 8440 8572 8460
rect 9394 8455 9459 8474
rect 8534 8431 8572 8440
rect 9456 8447 9459 8455
rect 9488 8447 9495 8474
rect 9523 8450 9533 8477
rect 9562 8455 9644 8477
rect 9562 8450 9566 8455
rect 9523 8447 9566 8450
rect 9456 8433 9566 8447
rect 9832 8451 9879 8452
rect 9832 8442 9880 8451
rect 8534 8430 8571 8431
rect 7957 8409 7993 8430
rect 8383 8409 8414 8430
rect 9832 8424 9851 8442
rect 9869 8424 9880 8442
rect 9832 8422 9880 8424
rect 7790 8405 7890 8409
rect 7790 8401 7852 8405
rect 7790 8375 7797 8401
rect 7823 8379 7852 8401
rect 7878 8379 7890 8405
rect 7823 8375 7890 8379
rect 7790 8372 7890 8375
rect 7958 8372 7993 8409
rect 8055 8406 8414 8409
rect 8055 8401 8277 8406
rect 8055 8377 8068 8401
rect 8092 8382 8277 8401
rect 8301 8382 8414 8406
rect 8092 8377 8414 8382
rect 8055 8373 8414 8377
rect 8481 8401 8630 8409
rect 8481 8381 8492 8401
rect 8512 8381 8630 8401
rect 8481 8374 8630 8381
rect 8481 8373 8522 8374
rect 7957 8333 7993 8372
rect 7805 8320 7842 8321
rect 7901 8320 7938 8321
rect 7957 8320 7964 8333
rect 7704 8311 7843 8320
rect 7704 8291 7814 8311
rect 7834 8291 7843 8311
rect 7704 8284 7843 8291
rect 7901 8311 7964 8320
rect 7901 8291 7910 8311
rect 7930 8295 7964 8311
rect 7987 8320 7993 8333
rect 8012 8320 8049 8321
rect 7987 8311 8049 8320
rect 7987 8295 8020 8311
rect 7930 8291 8020 8295
rect 8040 8291 8049 8311
rect 7704 8282 7801 8284
rect 7704 8281 7733 8282
rect 7901 8281 8049 8291
rect 8108 8311 8145 8321
rect 8220 8320 8257 8321
rect 8201 8318 8257 8320
rect 8108 8291 8116 8311
rect 8136 8291 8145 8311
rect 7957 8280 7993 8281
rect 7805 8221 7842 8222
rect 8108 8221 8145 8291
rect 8170 8311 8257 8318
rect 8170 8308 8228 8311
rect 8170 8288 8175 8308
rect 8196 8291 8228 8308
rect 8248 8291 8257 8311
rect 8196 8288 8257 8291
rect 8170 8281 8257 8288
rect 8316 8311 8353 8321
rect 8316 8291 8324 8311
rect 8344 8291 8353 8311
rect 8170 8280 8201 8281
rect 7804 8220 8145 8221
rect 7729 8216 8145 8220
rect 7729 8215 8106 8216
rect 7729 8195 7732 8215
rect 7752 8199 8106 8215
rect 8126 8199 8145 8216
rect 7752 8195 8145 8199
rect 8316 8212 8353 8291
rect 8383 8320 8414 8373
rect 9194 8365 9232 8367
rect 9841 8365 9880 8422
rect 9194 8332 9880 8365
rect 8433 8320 8470 8321
rect 8383 8311 8470 8320
rect 8383 8291 8441 8311
rect 8461 8291 8470 8311
rect 8383 8281 8470 8291
rect 8529 8311 8566 8321
rect 8529 8291 8537 8311
rect 8557 8291 8566 8311
rect 8383 8280 8414 8281
rect 8378 8212 8488 8225
rect 8529 8212 8566 8291
rect 8316 8210 8566 8212
rect 8316 8207 8417 8210
rect 8316 8188 8381 8207
rect 8378 8180 8381 8188
rect 8410 8180 8417 8207
rect 8445 8183 8455 8210
rect 8484 8188 8566 8210
rect 8786 8244 8954 8245
rect 9194 8244 9232 8332
rect 9493 8330 9540 8332
rect 9840 8308 9880 8332
rect 8786 8221 9232 8244
rect 9458 8275 9569 8290
rect 9458 8273 9500 8275
rect 9458 8253 9465 8273
rect 9484 8253 9500 8273
rect 9458 8245 9500 8253
rect 9528 8273 9569 8275
rect 9528 8253 9542 8273
rect 9561 8253 9569 8273
rect 9841 8264 9880 8308
rect 9528 8245 9569 8253
rect 9458 8239 9569 8245
rect 8786 8218 9230 8221
rect 8786 8216 8954 8218
rect 8484 8183 8488 8188
rect 8445 8180 8488 8183
rect 8378 8166 8488 8180
rect 7168 8147 7336 8149
rect 6889 8140 7336 8147
rect 6553 8120 6664 8126
rect 6553 8112 6594 8120
rect 5971 8099 6007 8100
rect 5819 8069 5828 8089
rect 5848 8069 5856 8089
rect 5707 8060 5763 8062
rect 5707 8059 5744 8060
rect 5819 8059 5856 8069
rect 5915 8089 6063 8099
rect 6163 8096 6259 8098
rect 5915 8069 5924 8089
rect 5944 8069 6034 8089
rect 6054 8069 6063 8089
rect 5915 8060 6063 8069
rect 6121 8089 6259 8096
rect 6121 8069 6130 8089
rect 6150 8069 6259 8089
rect 6553 8092 6561 8112
rect 6580 8092 6594 8112
rect 6553 8090 6594 8092
rect 6622 8112 6664 8120
rect 6622 8092 6638 8112
rect 6657 8092 6664 8112
rect 6889 8113 6914 8140
rect 6945 8121 7336 8140
rect 6945 8113 6994 8121
rect 7168 8120 7336 8121
rect 6889 8111 6994 8113
rect 6622 8090 6664 8092
rect 6553 8075 6664 8090
rect 6121 8060 6259 8069
rect 5915 8059 5952 8060
rect 5971 8008 6007 8060
rect 6026 8059 6063 8060
rect 6122 8059 6159 8060
rect 5442 8006 5483 8007
rect 5334 7999 5483 8006
rect 4457 7997 4494 7998
rect 4407 7988 4494 7997
rect 4407 7968 4465 7988
rect 4485 7968 4494 7988
rect 4407 7958 4494 7968
rect 4553 7988 4590 7998
rect 4553 7968 4561 7988
rect 4581 7968 4590 7988
rect 5334 7979 5452 7999
rect 5472 7979 5483 7999
rect 5334 7971 5483 7979
rect 5550 8003 5909 8007
rect 5550 7998 5872 8003
rect 5550 7974 5663 7998
rect 5687 7979 5872 7998
rect 5896 7979 5909 8003
rect 5687 7974 5909 7979
rect 5550 7971 5909 7974
rect 5971 7971 6006 8008
rect 6074 8005 6174 8008
rect 6074 8001 6141 8005
rect 6074 7975 6086 8001
rect 6112 7979 6141 8001
rect 6167 7979 6174 8005
rect 6112 7975 6174 7979
rect 6074 7971 6174 7975
rect 4407 7957 4438 7958
rect 4402 7889 4512 7902
rect 4553 7889 4590 7968
rect 4787 7953 4824 7954
rect 4783 7944 4824 7953
rect 5550 7950 5581 7971
rect 5971 7950 6007 7971
rect 5393 7949 5430 7950
rect 5167 7946 5201 7947
rect 4783 7926 4796 7944
rect 4814 7926 4824 7944
rect 4783 7917 4824 7926
rect 5166 7937 5203 7946
rect 5166 7919 5175 7937
rect 5193 7919 5203 7937
rect 4783 7897 4823 7917
rect 5166 7909 5203 7919
rect 5392 7940 5430 7949
rect 5392 7920 5401 7940
rect 5421 7920 5430 7940
rect 5392 7912 5430 7920
rect 5496 7944 5581 7950
rect 5606 7949 5643 7950
rect 5496 7924 5504 7944
rect 5524 7924 5581 7944
rect 5496 7916 5581 7924
rect 5605 7940 5643 7949
rect 5605 7920 5614 7940
rect 5634 7920 5643 7940
rect 5496 7915 5532 7916
rect 5605 7912 5643 7920
rect 5709 7944 5794 7950
rect 5814 7949 5851 7950
rect 5709 7924 5717 7944
rect 5737 7943 5794 7944
rect 5737 7924 5766 7943
rect 5709 7923 5766 7924
rect 5787 7923 5794 7943
rect 5709 7916 5794 7923
rect 5813 7940 5851 7949
rect 5813 7920 5822 7940
rect 5842 7920 5851 7940
rect 5709 7915 5745 7916
rect 5813 7912 5851 7920
rect 5917 7944 6061 7950
rect 5917 7924 5925 7944
rect 5945 7943 6033 7944
rect 5945 7924 5976 7943
rect 5917 7923 5976 7924
rect 6001 7924 6033 7943
rect 6053 7924 6061 7944
rect 6001 7923 6061 7924
rect 5917 7916 6061 7923
rect 5917 7915 5953 7916
rect 6025 7915 6061 7916
rect 6127 7949 6164 7950
rect 6127 7948 6165 7949
rect 6127 7940 6191 7948
rect 6127 7920 6136 7940
rect 6156 7926 6191 7940
rect 6211 7926 6214 7946
rect 6156 7921 6214 7926
rect 6156 7920 6191 7921
rect 4340 7887 4590 7889
rect 4340 7884 4441 7887
rect 2858 7827 2922 7839
rect 3198 7835 3235 7862
rect 3406 7835 3443 7866
rect 3619 7864 3655 7866
rect 4340 7865 4405 7884
rect 3619 7835 3656 7864
rect 4402 7857 4405 7865
rect 4434 7857 4441 7884
rect 4469 7860 4479 7887
rect 4508 7865 4590 7887
rect 4698 7887 4823 7897
rect 4698 7868 4706 7887
rect 4731 7868 4823 7887
rect 4508 7860 4512 7865
rect 4698 7861 4823 7868
rect 4469 7857 4512 7860
rect 4402 7843 4512 7857
rect 2858 7826 2893 7827
rect 2835 7821 2893 7826
rect 2835 7801 2838 7821
rect 2858 7807 2893 7821
rect 2913 7807 2922 7827
rect 2858 7799 2922 7807
rect 2884 7798 2922 7799
rect 2885 7797 2922 7798
rect 2988 7831 3024 7832
rect 3096 7831 3132 7832
rect 2988 7823 3132 7831
rect 2988 7803 2996 7823
rect 3016 7820 3104 7823
rect 3016 7803 3048 7820
rect 3068 7803 3104 7820
rect 3124 7803 3132 7823
rect 2988 7797 3132 7803
rect 3198 7827 3236 7835
rect 3304 7831 3340 7832
rect 3198 7807 3207 7827
rect 3227 7807 3236 7827
rect 3198 7798 3236 7807
rect 3255 7824 3340 7831
rect 3255 7804 3262 7824
rect 3283 7823 3340 7824
rect 3283 7804 3312 7823
rect 3255 7803 3312 7804
rect 3332 7803 3340 7823
rect 3198 7797 3235 7798
rect 3255 7797 3340 7803
rect 3406 7827 3444 7835
rect 3517 7831 3553 7832
rect 3406 7807 3415 7827
rect 3435 7807 3444 7827
rect 3406 7798 3444 7807
rect 3468 7823 3553 7831
rect 3468 7803 3525 7823
rect 3545 7803 3553 7823
rect 3406 7797 3443 7798
rect 3468 7797 3553 7803
rect 3619 7827 3657 7835
rect 3619 7807 3628 7827
rect 3648 7807 3657 7827
rect 3619 7798 3657 7807
rect 4783 7813 4823 7861
rect 5167 7881 5201 7909
rect 5393 7883 5430 7912
rect 5394 7881 5430 7883
rect 5606 7881 5643 7912
rect 5167 7880 5339 7881
rect 5167 7848 5353 7880
rect 5394 7859 5643 7881
rect 5814 7880 5851 7912
rect 6127 7908 6191 7920
rect 6231 7882 6258 8060
rect 8786 8038 8813 8216
rect 8853 8178 8917 8190
rect 9193 8186 9230 8218
rect 9401 8217 9650 8239
rect 9401 8186 9438 8217
rect 9614 8215 9650 8217
rect 9614 8186 9651 8215
rect 8853 8177 8888 8178
rect 8830 8172 8888 8177
rect 8830 8152 8833 8172
rect 8853 8158 8888 8172
rect 8908 8158 8917 8178
rect 8853 8150 8917 8158
rect 8879 8149 8917 8150
rect 8880 8148 8917 8149
rect 8983 8182 9019 8183
rect 9091 8182 9127 8183
rect 8983 8177 9127 8182
rect 8983 8174 9045 8177
rect 8983 8154 8991 8174
rect 9011 8157 9045 8174
rect 9068 8174 9127 8177
rect 9068 8157 9099 8174
rect 9011 8154 9099 8157
rect 9119 8154 9127 8174
rect 8983 8148 9127 8154
rect 9193 8178 9231 8186
rect 9299 8182 9335 8183
rect 9193 8158 9202 8178
rect 9222 8158 9231 8178
rect 9193 8149 9231 8158
rect 9250 8175 9335 8182
rect 9250 8155 9257 8175
rect 9278 8174 9335 8175
rect 9278 8155 9307 8174
rect 9250 8154 9307 8155
rect 9327 8154 9335 8174
rect 9193 8148 9230 8149
rect 9250 8148 9335 8154
rect 9401 8178 9439 8186
rect 9512 8182 9548 8183
rect 9401 8158 9410 8178
rect 9430 8158 9439 8178
rect 9401 8149 9439 8158
rect 9463 8174 9548 8182
rect 9463 8154 9520 8174
rect 9540 8154 9548 8174
rect 9401 8148 9438 8149
rect 9463 8148 9548 8154
rect 9614 8178 9652 8186
rect 9614 8158 9623 8178
rect 9643 8158 9652 8178
rect 9614 8149 9652 8158
rect 9614 8148 9651 8149
rect 9037 8127 9073 8148
rect 9463 8127 9494 8148
rect 8870 8123 8970 8127
rect 8870 8119 8932 8123
rect 8870 8093 8877 8119
rect 8903 8097 8932 8119
rect 8958 8097 8970 8123
rect 8903 8093 8970 8097
rect 8870 8090 8970 8093
rect 9038 8090 9073 8127
rect 9135 8124 9494 8127
rect 9135 8119 9357 8124
rect 9135 8095 9148 8119
rect 9172 8100 9357 8119
rect 9381 8100 9494 8124
rect 9172 8095 9494 8100
rect 9135 8091 9494 8095
rect 9561 8119 9710 8127
rect 9561 8099 9572 8119
rect 9592 8099 9710 8119
rect 9561 8092 9710 8099
rect 9561 8091 9602 8092
rect 8885 8038 8922 8039
rect 8981 8038 9018 8039
rect 9037 8038 9073 8090
rect 9092 8038 9129 8039
rect 8785 8029 8923 8038
rect 8785 8009 8894 8029
rect 8914 8009 8923 8029
rect 8785 8002 8923 8009
rect 8981 8029 9129 8038
rect 8981 8009 8990 8029
rect 9010 8009 9100 8029
rect 9120 8009 9129 8029
rect 8785 8000 8881 8002
rect 8981 7999 9129 8009
rect 9188 8029 9225 8039
rect 9300 8038 9337 8039
rect 9281 8036 9337 8038
rect 9188 8009 9196 8029
rect 9216 8009 9225 8029
rect 9037 7998 9073 7999
rect 6414 7956 6524 7970
rect 6414 7953 6457 7956
rect 6414 7948 6418 7953
rect 6090 7880 6258 7882
rect 5814 7874 6258 7880
rect 5167 7816 5201 7848
rect 3619 7797 3656 7798
rect 3042 7776 3078 7797
rect 3468 7776 3499 7797
rect 4783 7795 4794 7813
rect 4812 7795 4823 7813
rect 4783 7787 4823 7795
rect 5163 7807 5201 7816
rect 5163 7789 5173 7807
rect 5191 7789 5201 7807
rect 4784 7786 4821 7787
rect 5163 7783 5201 7789
rect 5319 7785 5353 7848
rect 5475 7853 5586 7859
rect 5475 7845 5516 7853
rect 5475 7825 5483 7845
rect 5502 7825 5516 7845
rect 5475 7823 5516 7825
rect 5544 7845 5586 7853
rect 5544 7825 5560 7845
rect 5579 7825 5586 7845
rect 5544 7823 5586 7825
rect 5475 7808 5586 7823
rect 5813 7854 6258 7874
rect 5813 7785 5851 7854
rect 6090 7853 6258 7854
rect 6336 7926 6418 7948
rect 6447 7926 6457 7953
rect 6485 7929 6492 7956
rect 6521 7948 6524 7956
rect 8519 7965 8630 7980
rect 8519 7963 8561 7965
rect 6521 7929 6586 7948
rect 6485 7926 6586 7929
rect 6336 7924 6586 7926
rect 6336 7845 6373 7924
rect 6414 7911 6524 7924
rect 6488 7855 6519 7856
rect 6336 7825 6345 7845
rect 6365 7825 6373 7845
rect 6336 7815 6373 7825
rect 6432 7845 6519 7855
rect 6432 7825 6441 7845
rect 6461 7825 6519 7845
rect 6432 7816 6519 7825
rect 6432 7815 6469 7816
rect 5163 7779 5200 7783
rect 2875 7772 2975 7776
rect 2875 7768 2937 7772
rect 2875 7742 2882 7768
rect 2908 7746 2937 7768
rect 2963 7746 2975 7772
rect 2908 7742 2975 7746
rect 2875 7739 2975 7742
rect 3043 7739 3078 7776
rect 3140 7773 3499 7776
rect 3140 7768 3362 7773
rect 3140 7744 3153 7768
rect 3177 7749 3362 7768
rect 3386 7749 3499 7773
rect 3177 7744 3499 7749
rect 3140 7740 3499 7744
rect 3566 7768 3715 7776
rect 5319 7774 5851 7785
rect 3566 7748 3577 7768
rect 3597 7748 3715 7768
rect 5318 7758 5851 7774
rect 6488 7763 6519 7816
rect 6549 7845 6586 7924
rect 6757 7934 7150 7941
rect 6757 7917 6765 7934
rect 6797 7921 7150 7934
rect 7170 7921 7173 7941
rect 8252 7936 8293 7945
rect 6797 7917 7173 7921
rect 6757 7916 7173 7917
rect 7847 7934 8015 7935
rect 8252 7934 8261 7936
rect 6757 7915 7098 7916
rect 6701 7855 6732 7856
rect 6549 7825 6558 7845
rect 6578 7825 6586 7845
rect 6549 7815 6586 7825
rect 6645 7848 6732 7855
rect 6645 7845 6706 7848
rect 6645 7825 6654 7845
rect 6674 7828 6706 7845
rect 6727 7828 6732 7848
rect 6674 7825 6732 7828
rect 6645 7818 6732 7825
rect 6757 7845 6794 7915
rect 7060 7914 7097 7915
rect 7847 7914 8261 7934
rect 8287 7914 8293 7936
rect 8519 7943 8526 7963
rect 8545 7943 8561 7963
rect 8519 7935 8561 7943
rect 8589 7963 8630 7965
rect 8589 7943 8603 7963
rect 8622 7943 8630 7963
rect 8589 7935 8630 7943
rect 8885 7939 8922 7940
rect 9188 7939 9225 8009
rect 9250 8029 9337 8036
rect 9250 8026 9308 8029
rect 9250 8006 9255 8026
rect 9276 8009 9308 8026
rect 9328 8009 9337 8029
rect 9276 8006 9337 8009
rect 9250 7999 9337 8006
rect 9396 8029 9433 8039
rect 9396 8009 9404 8029
rect 9424 8009 9433 8029
rect 9250 7998 9281 7999
rect 8884 7938 9225 7939
rect 8519 7929 8630 7935
rect 8809 7933 9225 7938
rect 7847 7908 8293 7914
rect 7847 7906 8015 7908
rect 6909 7855 6945 7856
rect 6757 7825 6766 7845
rect 6786 7825 6794 7845
rect 6645 7816 6701 7818
rect 6645 7815 6682 7816
rect 6757 7815 6794 7825
rect 6853 7845 7001 7855
rect 7101 7852 7197 7854
rect 6853 7825 6862 7845
rect 6882 7840 6972 7845
rect 6882 7825 6917 7840
rect 6853 7816 6917 7825
rect 6853 7815 6890 7816
rect 6909 7799 6917 7816
rect 6938 7825 6972 7840
rect 6992 7825 7001 7845
rect 6938 7816 7001 7825
rect 7059 7845 7197 7852
rect 7059 7825 7068 7845
rect 7088 7825 7197 7845
rect 7059 7816 7197 7825
rect 6938 7799 6945 7816
rect 6964 7815 7001 7816
rect 7060 7815 7097 7816
rect 6909 7764 6945 7799
rect 6380 7762 6421 7763
rect 5318 7757 5832 7758
rect 3566 7741 3715 7748
rect 6272 7755 6421 7762
rect 4155 7745 4669 7746
rect 3566 7740 3607 7741
rect 2890 7687 2927 7688
rect 2986 7687 3023 7688
rect 3042 7687 3078 7739
rect 3097 7687 3134 7688
rect 2790 7678 2928 7687
rect 2790 7658 2899 7678
rect 2919 7658 2928 7678
rect 2790 7651 2928 7658
rect 2986 7678 3134 7687
rect 2986 7658 2995 7678
rect 3015 7658 3105 7678
rect 3125 7658 3134 7678
rect 2790 7649 2886 7651
rect 2986 7648 3134 7658
rect 3193 7678 3230 7688
rect 3305 7687 3342 7688
rect 3286 7685 3342 7687
rect 3193 7658 3201 7678
rect 3221 7658 3230 7678
rect 3042 7647 3078 7648
rect 1972 7595 2140 7597
rect 1694 7589 2140 7595
rect 762 7565 1178 7570
rect 1357 7568 1468 7574
rect 762 7564 1103 7565
rect 706 7504 737 7505
rect 554 7474 563 7494
rect 583 7474 591 7494
rect 554 7464 591 7474
rect 650 7497 737 7504
rect 650 7494 711 7497
rect 650 7474 659 7494
rect 679 7477 711 7494
rect 732 7477 737 7497
rect 679 7474 737 7477
rect 650 7467 737 7474
rect 762 7494 799 7564
rect 1065 7563 1102 7564
rect 1357 7560 1398 7568
rect 1357 7540 1365 7560
rect 1384 7540 1398 7560
rect 1357 7538 1398 7540
rect 1426 7560 1468 7568
rect 1426 7540 1442 7560
rect 1461 7540 1468 7560
rect 1694 7567 1700 7589
rect 1726 7569 2140 7589
rect 2890 7588 2927 7589
rect 3193 7588 3230 7658
rect 3255 7678 3342 7685
rect 3255 7675 3313 7678
rect 3255 7655 3260 7675
rect 3281 7658 3313 7675
rect 3333 7658 3342 7678
rect 3281 7655 3342 7658
rect 3255 7648 3342 7655
rect 3401 7678 3438 7688
rect 3401 7658 3409 7678
rect 3429 7658 3438 7678
rect 3255 7647 3286 7648
rect 2889 7587 3230 7588
rect 1726 7567 1735 7569
rect 1972 7568 2140 7569
rect 2814 7582 3230 7587
rect 1694 7558 1735 7567
rect 2814 7562 2817 7582
rect 2837 7562 3230 7582
rect 3401 7579 3438 7658
rect 3468 7687 3499 7740
rect 4136 7729 4669 7745
rect 6272 7735 6390 7755
rect 6410 7735 6421 7755
rect 4136 7718 4668 7729
rect 6272 7727 6421 7735
rect 6488 7759 6847 7763
rect 6488 7754 6810 7759
rect 6488 7730 6601 7754
rect 6625 7735 6810 7754
rect 6834 7735 6847 7759
rect 6625 7730 6847 7735
rect 6488 7727 6847 7730
rect 6909 7727 6944 7764
rect 7012 7761 7112 7764
rect 7012 7757 7079 7761
rect 7012 7731 7024 7757
rect 7050 7735 7079 7757
rect 7105 7735 7112 7761
rect 7050 7731 7112 7735
rect 7012 7727 7112 7731
rect 4787 7720 4824 7724
rect 3518 7687 3555 7688
rect 3468 7678 3555 7687
rect 3468 7658 3526 7678
rect 3546 7658 3555 7678
rect 3468 7648 3555 7658
rect 3614 7678 3651 7688
rect 3614 7658 3622 7678
rect 3642 7658 3651 7678
rect 3468 7647 3499 7648
rect 3463 7579 3573 7592
rect 3614 7579 3651 7658
rect 3401 7577 3651 7579
rect 3401 7574 3502 7577
rect 3401 7555 3466 7574
rect 1426 7538 1468 7540
rect 1357 7523 1468 7538
rect 3463 7547 3466 7555
rect 3495 7547 3502 7574
rect 3530 7550 3540 7577
rect 3569 7555 3651 7577
rect 3729 7649 3897 7650
rect 4136 7649 4174 7718
rect 3729 7629 4174 7649
rect 4401 7680 4512 7695
rect 4401 7678 4443 7680
rect 4401 7658 4408 7678
rect 4427 7658 4443 7678
rect 4401 7650 4443 7658
rect 4471 7678 4512 7680
rect 4471 7658 4485 7678
rect 4504 7658 4512 7678
rect 4471 7650 4512 7658
rect 4401 7644 4512 7650
rect 4634 7655 4668 7718
rect 4786 7714 4824 7720
rect 5166 7716 5203 7717
rect 4786 7696 4796 7714
rect 4814 7696 4824 7714
rect 4786 7687 4824 7696
rect 5164 7708 5204 7716
rect 5164 7690 5175 7708
rect 5193 7690 5204 7708
rect 6488 7706 6519 7727
rect 6909 7706 6945 7727
rect 6331 7705 6368 7706
rect 4786 7655 4820 7687
rect 3729 7623 4173 7629
rect 3729 7621 3897 7623
rect 3569 7550 3573 7555
rect 3530 7547 3573 7550
rect 3463 7533 3573 7547
rect 914 7504 950 7505
rect 762 7474 771 7494
rect 791 7474 799 7494
rect 650 7465 706 7467
rect 650 7464 687 7465
rect 762 7464 799 7474
rect 858 7494 1006 7504
rect 1106 7501 1202 7503
rect 858 7474 867 7494
rect 887 7474 977 7494
rect 997 7474 1006 7494
rect 858 7465 1006 7474
rect 1064 7494 1202 7501
rect 1064 7474 1073 7494
rect 1093 7474 1202 7494
rect 1064 7465 1202 7474
rect 858 7464 895 7465
rect 914 7413 950 7465
rect 969 7464 1006 7465
rect 1065 7464 1102 7465
rect 385 7411 426 7412
rect 277 7404 426 7411
rect 277 7384 395 7404
rect 415 7384 426 7404
rect 277 7376 426 7384
rect 493 7408 852 7412
rect 493 7403 815 7408
rect 493 7379 606 7403
rect 630 7384 815 7403
rect 839 7384 852 7408
rect 630 7379 852 7384
rect 493 7376 852 7379
rect 914 7376 949 7413
rect 1017 7410 1117 7413
rect 1017 7406 1084 7410
rect 1017 7380 1029 7406
rect 1055 7384 1084 7406
rect 1110 7384 1117 7410
rect 1055 7380 1117 7384
rect 1017 7376 1117 7380
rect 493 7355 524 7376
rect 914 7355 950 7376
rect 336 7354 373 7355
rect 335 7345 373 7354
rect 335 7325 344 7345
rect 364 7325 373 7345
rect 335 7317 373 7325
rect 439 7349 524 7355
rect 549 7354 586 7355
rect 439 7329 447 7349
rect 467 7329 524 7349
rect 439 7321 524 7329
rect 548 7345 586 7354
rect 548 7325 557 7345
rect 577 7325 586 7345
rect 439 7320 475 7321
rect 548 7317 586 7325
rect 652 7349 737 7355
rect 757 7354 794 7355
rect 652 7329 660 7349
rect 680 7348 737 7349
rect 680 7329 709 7348
rect 652 7328 709 7329
rect 730 7328 737 7348
rect 652 7321 737 7328
rect 756 7345 794 7354
rect 756 7325 765 7345
rect 785 7325 794 7345
rect 652 7320 688 7321
rect 756 7317 794 7325
rect 860 7349 1004 7355
rect 860 7329 868 7349
rect 888 7346 976 7349
rect 888 7329 919 7346
rect 860 7326 919 7329
rect 942 7329 976 7346
rect 996 7329 1004 7349
rect 942 7326 1004 7329
rect 860 7321 1004 7326
rect 860 7320 896 7321
rect 968 7320 1004 7321
rect 1070 7354 1107 7355
rect 1070 7353 1108 7354
rect 1070 7345 1134 7353
rect 1070 7325 1079 7345
rect 1099 7331 1134 7345
rect 1154 7331 1157 7351
rect 1099 7326 1157 7331
rect 1099 7325 1134 7326
rect 336 7288 373 7317
rect 337 7286 373 7288
rect 549 7286 586 7317
rect 337 7264 586 7286
rect 757 7285 794 7317
rect 1070 7313 1134 7325
rect 1174 7287 1201 7465
rect 3729 7443 3756 7621
rect 3796 7583 3860 7595
rect 4136 7591 4173 7623
rect 4344 7622 4593 7644
rect 4634 7623 4820 7655
rect 4648 7622 4820 7623
rect 4344 7591 4381 7622
rect 4557 7620 4593 7622
rect 4557 7591 4594 7620
rect 4786 7594 4820 7622
rect 5164 7642 5204 7690
rect 6330 7696 6368 7705
rect 6330 7676 6339 7696
rect 6359 7676 6368 7696
rect 6330 7668 6368 7676
rect 6434 7700 6519 7706
rect 6544 7705 6581 7706
rect 6434 7680 6442 7700
rect 6462 7680 6519 7700
rect 6434 7672 6519 7680
rect 6543 7696 6581 7705
rect 6543 7676 6552 7696
rect 6572 7676 6581 7696
rect 6434 7671 6470 7672
rect 6543 7668 6581 7676
rect 6647 7700 6732 7706
rect 6752 7705 6789 7706
rect 6647 7680 6655 7700
rect 6675 7699 6732 7700
rect 6675 7680 6704 7699
rect 6647 7679 6704 7680
rect 6725 7679 6732 7699
rect 6647 7672 6732 7679
rect 6751 7696 6789 7705
rect 6751 7676 6760 7696
rect 6780 7676 6789 7696
rect 6647 7671 6683 7672
rect 6751 7668 6789 7676
rect 6855 7700 6999 7706
rect 6855 7680 6863 7700
rect 6883 7680 6971 7700
rect 6991 7680 6999 7700
rect 6855 7672 6999 7680
rect 6855 7671 6891 7672
rect 6963 7671 6999 7672
rect 7065 7705 7102 7706
rect 7065 7704 7103 7705
rect 7065 7696 7129 7704
rect 7065 7676 7074 7696
rect 7094 7682 7129 7696
rect 7149 7682 7152 7702
rect 7094 7677 7152 7682
rect 7094 7676 7129 7677
rect 5475 7646 5585 7660
rect 5475 7643 5518 7646
rect 5164 7635 5289 7642
rect 5475 7638 5479 7643
rect 5164 7616 5256 7635
rect 5281 7616 5289 7635
rect 5164 7606 5289 7616
rect 5397 7616 5479 7638
rect 5508 7616 5518 7643
rect 5546 7619 5553 7646
rect 5582 7638 5585 7646
rect 6331 7639 6368 7668
rect 5582 7619 5647 7638
rect 6332 7637 6368 7639
rect 6544 7637 6581 7668
rect 6752 7641 6789 7668
rect 7065 7664 7129 7676
rect 5546 7616 5647 7619
rect 5397 7614 5647 7616
rect 3796 7582 3831 7583
rect 3773 7577 3831 7582
rect 3773 7557 3776 7577
rect 3796 7563 3831 7577
rect 3851 7563 3860 7583
rect 3796 7555 3860 7563
rect 3822 7554 3860 7555
rect 3823 7553 3860 7554
rect 3926 7587 3962 7588
rect 4034 7587 4070 7588
rect 3926 7580 4070 7587
rect 3926 7579 3986 7580
rect 3926 7559 3934 7579
rect 3954 7560 3986 7579
rect 4011 7579 4070 7580
rect 4011 7560 4042 7579
rect 3954 7559 4042 7560
rect 4062 7559 4070 7579
rect 3926 7553 4070 7559
rect 4136 7583 4174 7591
rect 4242 7587 4278 7588
rect 4136 7563 4145 7583
rect 4165 7563 4174 7583
rect 4136 7554 4174 7563
rect 4193 7580 4278 7587
rect 4193 7560 4200 7580
rect 4221 7579 4278 7580
rect 4221 7560 4250 7579
rect 4193 7559 4250 7560
rect 4270 7559 4278 7579
rect 4136 7553 4173 7554
rect 4193 7553 4278 7559
rect 4344 7583 4382 7591
rect 4455 7587 4491 7588
rect 4344 7563 4353 7583
rect 4373 7563 4382 7583
rect 4344 7554 4382 7563
rect 4406 7579 4491 7587
rect 4406 7559 4463 7579
rect 4483 7559 4491 7579
rect 4344 7553 4381 7554
rect 4406 7553 4491 7559
rect 4557 7583 4595 7591
rect 4557 7563 4566 7583
rect 4586 7563 4595 7583
rect 4557 7554 4595 7563
rect 4784 7584 4821 7594
rect 5164 7586 5204 7606
rect 4784 7566 4794 7584
rect 4812 7566 4821 7584
rect 4784 7557 4821 7566
rect 5163 7577 5204 7586
rect 5163 7559 5173 7577
rect 5191 7559 5204 7577
rect 4786 7556 4820 7557
rect 4557 7553 4594 7554
rect 3980 7532 4016 7553
rect 4406 7532 4437 7553
rect 5163 7550 5204 7559
rect 5163 7549 5200 7550
rect 5397 7535 5434 7614
rect 5475 7601 5585 7614
rect 5549 7545 5580 7546
rect 3813 7528 3913 7532
rect 3813 7524 3875 7528
rect 3813 7498 3820 7524
rect 3846 7502 3875 7524
rect 3901 7502 3913 7528
rect 3846 7498 3913 7502
rect 3813 7495 3913 7498
rect 3981 7495 4016 7532
rect 4078 7529 4437 7532
rect 4078 7524 4300 7529
rect 4078 7500 4091 7524
rect 4115 7505 4300 7524
rect 4324 7505 4437 7529
rect 4115 7500 4437 7505
rect 4078 7496 4437 7500
rect 4504 7524 4653 7532
rect 4504 7504 4515 7524
rect 4535 7504 4653 7524
rect 5397 7515 5406 7535
rect 5426 7515 5434 7535
rect 5397 7505 5434 7515
rect 5493 7535 5580 7545
rect 5493 7515 5502 7535
rect 5522 7515 5580 7535
rect 5493 7506 5580 7515
rect 5493 7505 5530 7506
rect 4504 7497 4653 7504
rect 4504 7496 4545 7497
rect 3828 7443 3865 7444
rect 3924 7443 3961 7444
rect 3980 7443 4016 7495
rect 4035 7443 4072 7444
rect 3728 7434 3866 7443
rect 3353 7400 3464 7415
rect 3728 7414 3837 7434
rect 3857 7414 3866 7434
rect 3728 7407 3866 7414
rect 3924 7434 4072 7443
rect 3924 7414 3933 7434
rect 3953 7414 4043 7434
rect 4063 7414 4072 7434
rect 3728 7405 3824 7407
rect 3924 7404 4072 7414
rect 4131 7434 4168 7444
rect 4243 7443 4280 7444
rect 4224 7441 4280 7443
rect 4131 7414 4139 7434
rect 4159 7414 4168 7434
rect 3980 7403 4016 7404
rect 3353 7398 3395 7400
rect 2690 7379 2760 7388
rect 2690 7370 2707 7379
rect 2681 7350 2707 7370
rect 2755 7370 2760 7379
rect 3353 7378 3360 7398
rect 3379 7378 3395 7398
rect 3353 7370 3395 7378
rect 3423 7398 3464 7400
rect 3423 7378 3437 7398
rect 3456 7378 3464 7398
rect 3423 7370 3464 7378
rect 2755 7369 2849 7370
rect 2755 7350 3125 7369
rect 3353 7364 3464 7370
rect 1468 7336 1578 7350
rect 1468 7333 1511 7336
rect 1468 7328 1472 7333
rect 1033 7285 1201 7287
rect 757 7282 1201 7285
rect 418 7258 529 7264
rect 418 7250 459 7258
rect 107 7195 146 7239
rect 418 7230 426 7250
rect 445 7230 459 7250
rect 418 7228 459 7230
rect 487 7250 529 7258
rect 487 7230 503 7250
rect 522 7230 529 7250
rect 487 7228 529 7230
rect 418 7214 529 7228
rect 755 7259 1201 7282
rect 107 7171 147 7195
rect 447 7171 494 7173
rect 755 7171 793 7259
rect 1033 7258 1201 7259
rect 1390 7306 1472 7328
rect 1501 7306 1511 7333
rect 1539 7309 1546 7336
rect 1575 7328 1578 7336
rect 2681 7343 3125 7350
rect 2681 7341 2849 7343
rect 2681 7333 2760 7341
rect 1575 7309 1640 7328
rect 1539 7306 1640 7309
rect 1390 7304 1640 7306
rect 1390 7225 1427 7304
rect 1468 7291 1578 7304
rect 1542 7235 1573 7236
rect 1390 7205 1399 7225
rect 1419 7205 1427 7225
rect 1390 7195 1427 7205
rect 1486 7225 1573 7235
rect 1486 7205 1495 7225
rect 1515 7205 1573 7225
rect 1486 7196 1573 7205
rect 1486 7195 1523 7196
rect 107 7138 793 7171
rect 1542 7143 1573 7196
rect 1603 7225 1640 7304
rect 1811 7301 2204 7321
rect 2224 7301 2227 7321
rect 1811 7296 2227 7301
rect 1811 7295 2152 7296
rect 1755 7235 1786 7236
rect 1603 7205 1612 7225
rect 1632 7205 1640 7225
rect 1603 7195 1640 7205
rect 1699 7228 1786 7235
rect 1699 7225 1760 7228
rect 1699 7205 1708 7225
rect 1728 7208 1760 7225
rect 1781 7208 1786 7228
rect 1728 7205 1786 7208
rect 1699 7198 1786 7205
rect 1811 7225 1848 7295
rect 2114 7294 2151 7295
rect 1963 7235 1999 7236
rect 1811 7205 1820 7225
rect 1840 7205 1848 7225
rect 1699 7196 1755 7198
rect 1699 7195 1736 7196
rect 1811 7195 1848 7205
rect 1907 7225 2055 7235
rect 2155 7232 2251 7234
rect 1907 7205 1916 7225
rect 1936 7205 2026 7225
rect 2046 7205 2055 7225
rect 1907 7196 2055 7205
rect 2113 7225 2251 7232
rect 2113 7205 2122 7225
rect 2142 7205 2251 7225
rect 2113 7196 2251 7205
rect 1907 7195 1944 7196
rect 1963 7144 1999 7196
rect 2018 7195 2055 7196
rect 2114 7195 2151 7196
rect 1434 7142 1475 7143
rect 106 7081 145 7138
rect 755 7136 793 7138
rect 1326 7135 1475 7142
rect 1326 7115 1444 7135
rect 1464 7115 1475 7135
rect 1326 7107 1475 7115
rect 1542 7139 1901 7143
rect 1542 7134 1864 7139
rect 1542 7110 1655 7134
rect 1679 7115 1864 7134
rect 1888 7115 1901 7139
rect 1679 7110 1901 7115
rect 1542 7107 1901 7110
rect 1963 7107 1998 7144
rect 2066 7141 2166 7144
rect 2066 7137 2133 7141
rect 2066 7111 2078 7137
rect 2104 7115 2133 7137
rect 2159 7115 2166 7141
rect 2104 7111 2166 7115
rect 2066 7107 2166 7111
rect 1542 7086 1573 7107
rect 1963 7086 1999 7107
rect 1385 7085 1422 7086
rect 106 7079 154 7081
rect 106 7061 117 7079
rect 135 7061 154 7079
rect 1384 7076 1422 7085
rect 106 7052 154 7061
rect 107 7051 154 7052
rect 420 7056 530 7070
rect 420 7053 463 7056
rect 420 7048 424 7053
rect 342 7026 424 7048
rect 453 7026 463 7053
rect 491 7029 498 7056
rect 527 7048 530 7056
rect 1384 7056 1393 7076
rect 1413 7056 1422 7076
rect 1384 7048 1422 7056
rect 1488 7080 1573 7086
rect 1598 7085 1635 7086
rect 1488 7060 1496 7080
rect 1516 7060 1573 7080
rect 1488 7052 1573 7060
rect 1597 7076 1635 7085
rect 1597 7056 1606 7076
rect 1626 7056 1635 7076
rect 1488 7051 1524 7052
rect 1597 7048 1635 7056
rect 1701 7080 1786 7086
rect 1806 7085 1843 7086
rect 1701 7060 1709 7080
rect 1729 7079 1786 7080
rect 1729 7060 1758 7079
rect 1701 7059 1758 7060
rect 1779 7059 1786 7079
rect 1701 7052 1786 7059
rect 1805 7076 1843 7085
rect 1805 7056 1814 7076
rect 1834 7056 1843 7076
rect 1701 7051 1737 7052
rect 1805 7048 1843 7056
rect 1909 7080 2053 7086
rect 1909 7060 1917 7080
rect 1937 7078 2025 7080
rect 1937 7060 1966 7078
rect 1909 7059 1966 7060
rect 1995 7060 2025 7078
rect 2045 7060 2053 7080
rect 1995 7059 2053 7060
rect 1909 7052 2053 7059
rect 1909 7051 1945 7052
rect 2017 7051 2053 7052
rect 2119 7085 2156 7086
rect 2119 7084 2157 7085
rect 2119 7076 2183 7084
rect 2119 7056 2128 7076
rect 2148 7062 2183 7076
rect 2203 7062 2206 7082
rect 2148 7057 2206 7062
rect 2148 7056 2183 7057
rect 527 7029 592 7048
rect 491 7026 592 7029
rect 342 7024 592 7026
rect 110 6988 147 6989
rect 106 6985 147 6988
rect 106 6980 148 6985
rect 106 6962 119 6980
rect 137 6962 148 6980
rect 106 6948 148 6962
rect 186 6948 233 6952
rect 106 6942 233 6948
rect 106 6913 194 6942
rect 223 6913 233 6942
rect 342 6945 379 7024
rect 420 7011 530 7024
rect 494 6955 525 6956
rect 342 6925 351 6945
rect 371 6925 379 6945
rect 342 6915 379 6925
rect 438 6945 525 6955
rect 438 6925 447 6945
rect 467 6925 525 6945
rect 438 6916 525 6925
rect 438 6915 475 6916
rect 106 6909 233 6913
rect 106 6892 145 6909
rect 186 6908 233 6909
rect 106 6874 117 6892
rect 135 6874 145 6892
rect 106 6865 145 6874
rect 107 6864 144 6865
rect 494 6863 525 6916
rect 555 6945 592 7024
rect 763 7021 1156 7041
rect 1176 7021 1179 7041
rect 763 7016 1179 7021
rect 1385 7019 1422 7048
rect 1386 7017 1422 7019
rect 1598 7017 1635 7048
rect 763 7015 1104 7016
rect 707 6955 738 6956
rect 555 6925 564 6945
rect 584 6925 592 6945
rect 555 6915 592 6925
rect 651 6948 738 6955
rect 651 6945 712 6948
rect 651 6925 660 6945
rect 680 6928 712 6945
rect 733 6928 738 6948
rect 680 6925 738 6928
rect 651 6918 738 6925
rect 763 6945 800 7015
rect 1066 7014 1103 7015
rect 1386 6995 1635 7017
rect 1806 7016 1843 7048
rect 2119 7044 2183 7056
rect 2223 7020 2250 7196
rect 2681 7163 2708 7333
rect 2748 7303 2812 7315
rect 3088 7311 3125 7343
rect 3296 7342 3545 7364
rect 3828 7344 3865 7345
rect 4131 7344 4168 7414
rect 4193 7434 4280 7441
rect 4193 7431 4251 7434
rect 4193 7411 4198 7431
rect 4219 7414 4251 7431
rect 4271 7414 4280 7434
rect 4219 7411 4280 7414
rect 4193 7404 4280 7411
rect 4339 7434 4376 7444
rect 4339 7414 4347 7434
rect 4367 7414 4376 7434
rect 4193 7403 4224 7404
rect 3827 7343 4168 7344
rect 3296 7311 3333 7342
rect 3509 7340 3545 7342
rect 3509 7311 3546 7340
rect 3752 7338 4168 7343
rect 3752 7318 3755 7338
rect 3775 7318 4168 7338
rect 4339 7335 4376 7414
rect 4406 7443 4437 7496
rect 4787 7494 4824 7495
rect 4786 7485 4825 7494
rect 4786 7467 4796 7485
rect 4814 7467 4825 7485
rect 5166 7483 5203 7487
rect 4698 7450 4745 7451
rect 4786 7450 4825 7467
rect 4698 7446 4825 7450
rect 4456 7443 4493 7444
rect 4406 7434 4493 7443
rect 4406 7414 4464 7434
rect 4484 7414 4493 7434
rect 4406 7404 4493 7414
rect 4552 7434 4589 7444
rect 4552 7414 4560 7434
rect 4580 7414 4589 7434
rect 4406 7403 4437 7404
rect 4401 7335 4511 7348
rect 4552 7335 4589 7414
rect 4698 7417 4708 7446
rect 4737 7417 4825 7446
rect 4698 7411 4825 7417
rect 4698 7407 4745 7411
rect 4783 7397 4825 7411
rect 4783 7379 4794 7397
rect 4812 7379 4825 7397
rect 4783 7374 4825 7379
rect 4784 7371 4825 7374
rect 5163 7478 5203 7483
rect 5163 7460 5175 7478
rect 5193 7460 5203 7478
rect 4784 7370 4821 7371
rect 4339 7333 4589 7335
rect 4339 7330 4440 7333
rect 4339 7311 4404 7330
rect 2748 7302 2783 7303
rect 2725 7297 2783 7302
rect 2725 7277 2728 7297
rect 2748 7283 2783 7297
rect 2803 7283 2812 7303
rect 2748 7275 2812 7283
rect 2774 7274 2812 7275
rect 2775 7273 2812 7274
rect 2878 7307 2914 7308
rect 2986 7307 3022 7308
rect 2878 7299 3022 7307
rect 2878 7279 2886 7299
rect 2906 7279 2994 7299
rect 3014 7279 3022 7299
rect 2878 7273 3022 7279
rect 3088 7303 3126 7311
rect 3194 7307 3230 7308
rect 3088 7283 3097 7303
rect 3117 7283 3126 7303
rect 3088 7274 3126 7283
rect 3145 7300 3230 7307
rect 3145 7280 3152 7300
rect 3173 7299 3230 7300
rect 3173 7280 3202 7299
rect 3145 7279 3202 7280
rect 3222 7279 3230 7299
rect 3088 7273 3125 7274
rect 3145 7273 3230 7279
rect 3296 7303 3334 7311
rect 3407 7307 3443 7308
rect 3296 7283 3305 7303
rect 3325 7283 3334 7303
rect 3296 7274 3334 7283
rect 3358 7299 3443 7307
rect 3358 7279 3415 7299
rect 3435 7279 3443 7299
rect 3296 7273 3333 7274
rect 3358 7273 3443 7279
rect 3509 7303 3547 7311
rect 3509 7283 3518 7303
rect 3538 7283 3547 7303
rect 4401 7303 4404 7311
rect 4433 7303 4440 7330
rect 4468 7306 4478 7333
rect 4507 7311 4589 7333
rect 4507 7306 4511 7311
rect 4468 7303 4511 7306
rect 4401 7289 4511 7303
rect 4777 7307 4824 7308
rect 4777 7298 4825 7307
rect 3509 7274 3547 7283
rect 4777 7280 4796 7298
rect 4814 7280 4825 7298
rect 4777 7278 4825 7280
rect 3509 7273 3546 7274
rect 2932 7252 2968 7273
rect 3358 7252 3389 7273
rect 2765 7248 2865 7252
rect 2765 7244 2827 7248
rect 2765 7218 2772 7244
rect 2798 7222 2827 7244
rect 2853 7222 2865 7248
rect 2798 7218 2865 7222
rect 2765 7215 2865 7218
rect 2933 7215 2968 7252
rect 3030 7249 3389 7252
rect 3030 7244 3252 7249
rect 3030 7220 3043 7244
rect 3067 7225 3252 7244
rect 3276 7225 3389 7249
rect 3067 7220 3389 7225
rect 3030 7216 3389 7220
rect 3456 7244 3605 7252
rect 3456 7224 3467 7244
rect 3487 7224 3605 7244
rect 3456 7217 3605 7224
rect 4138 7221 4176 7223
rect 4786 7221 4825 7278
rect 5163 7280 5203 7460
rect 5549 7453 5580 7506
rect 5610 7535 5647 7614
rect 5818 7611 6211 7631
rect 6231 7611 6234 7631
rect 6332 7615 6581 7637
rect 6750 7636 6791 7641
rect 7169 7638 7196 7816
rect 7847 7728 7874 7906
rect 8252 7903 8293 7908
rect 8462 7907 8711 7929
rect 8809 7913 8812 7933
rect 8832 7913 9225 7933
rect 9396 7930 9433 8009
rect 9463 8038 9494 8091
rect 9840 8084 9880 8264
rect 9840 8066 9850 8084
rect 9868 8066 9880 8084
rect 9840 8061 9880 8066
rect 9840 8057 9877 8061
rect 9513 8038 9550 8039
rect 9463 8029 9550 8038
rect 9463 8009 9521 8029
rect 9541 8009 9550 8029
rect 9463 7999 9550 8009
rect 9609 8029 9646 8039
rect 9609 8009 9617 8029
rect 9637 8009 9646 8029
rect 9463 7998 9494 7999
rect 9458 7930 9568 7943
rect 9609 7930 9646 8009
rect 9843 7994 9880 7995
rect 9839 7985 9880 7994
rect 9839 7967 9852 7985
rect 9870 7967 9880 7985
rect 9839 7958 9880 7967
rect 9839 7938 9879 7958
rect 9396 7928 9646 7930
rect 9396 7925 9497 7928
rect 7914 7868 7978 7880
rect 8254 7876 8291 7903
rect 8462 7876 8499 7907
rect 8675 7905 8711 7907
rect 9396 7906 9461 7925
rect 8675 7876 8712 7905
rect 9458 7898 9461 7906
rect 9490 7898 9497 7925
rect 9525 7901 9535 7928
rect 9564 7906 9646 7928
rect 9754 7928 9879 7938
rect 9754 7909 9762 7928
rect 9787 7909 9879 7928
rect 9564 7901 9568 7906
rect 9754 7902 9879 7909
rect 9525 7898 9568 7901
rect 9458 7884 9568 7898
rect 7914 7867 7949 7868
rect 7891 7862 7949 7867
rect 7891 7842 7894 7862
rect 7914 7848 7949 7862
rect 7969 7848 7978 7868
rect 7914 7840 7978 7848
rect 7940 7839 7978 7840
rect 7941 7838 7978 7839
rect 8044 7872 8080 7873
rect 8152 7872 8188 7873
rect 8044 7864 8188 7872
rect 8044 7844 8052 7864
rect 8072 7861 8160 7864
rect 8072 7844 8104 7861
rect 8124 7844 8160 7861
rect 8180 7844 8188 7864
rect 8044 7838 8188 7844
rect 8254 7868 8292 7876
rect 8360 7872 8396 7873
rect 8254 7848 8263 7868
rect 8283 7848 8292 7868
rect 8254 7839 8292 7848
rect 8311 7865 8396 7872
rect 8311 7845 8318 7865
rect 8339 7864 8396 7865
rect 8339 7845 8368 7864
rect 8311 7844 8368 7845
rect 8388 7844 8396 7864
rect 8254 7838 8291 7839
rect 8311 7838 8396 7844
rect 8462 7868 8500 7876
rect 8573 7872 8609 7873
rect 8462 7848 8471 7868
rect 8491 7848 8500 7868
rect 8462 7839 8500 7848
rect 8524 7864 8609 7872
rect 8524 7844 8581 7864
rect 8601 7844 8609 7864
rect 8462 7838 8499 7839
rect 8524 7838 8609 7844
rect 8675 7868 8713 7876
rect 8675 7848 8684 7868
rect 8704 7848 8713 7868
rect 8675 7839 8713 7848
rect 9839 7854 9879 7902
rect 8675 7838 8712 7839
rect 8098 7817 8134 7838
rect 8524 7817 8555 7838
rect 9839 7836 9850 7854
rect 9868 7836 9879 7854
rect 9839 7828 9879 7836
rect 9840 7827 9877 7828
rect 7931 7813 8031 7817
rect 7931 7809 7993 7813
rect 7931 7783 7938 7809
rect 7964 7787 7993 7809
rect 8019 7787 8031 7813
rect 7964 7783 8031 7787
rect 7931 7780 8031 7783
rect 8099 7780 8134 7817
rect 8196 7814 8555 7817
rect 8196 7809 8418 7814
rect 8196 7785 8209 7809
rect 8233 7790 8418 7809
rect 8442 7790 8555 7814
rect 8233 7785 8555 7790
rect 8196 7781 8555 7785
rect 8622 7809 8771 7817
rect 8622 7789 8633 7809
rect 8653 7789 8771 7809
rect 8622 7782 8771 7789
rect 9211 7786 9725 7787
rect 8622 7781 8663 7782
rect 7946 7728 7983 7729
rect 8042 7728 8079 7729
rect 8098 7728 8134 7780
rect 8153 7728 8190 7729
rect 7846 7719 7984 7728
rect 7846 7699 7955 7719
rect 7975 7699 7984 7719
rect 7846 7692 7984 7699
rect 8042 7719 8190 7728
rect 8042 7699 8051 7719
rect 8071 7699 8161 7719
rect 8181 7699 8190 7719
rect 7846 7690 7942 7692
rect 8042 7689 8190 7699
rect 8249 7719 8286 7729
rect 8361 7728 8398 7729
rect 8342 7726 8398 7728
rect 8249 7699 8257 7719
rect 8277 7699 8286 7719
rect 8098 7688 8134 7689
rect 7028 7636 7196 7638
rect 6750 7630 7196 7636
rect 5818 7606 6234 7611
rect 6413 7609 6524 7615
rect 5818 7605 6159 7606
rect 5762 7545 5793 7546
rect 5610 7515 5619 7535
rect 5639 7515 5647 7535
rect 5610 7505 5647 7515
rect 5706 7538 5793 7545
rect 5706 7535 5767 7538
rect 5706 7515 5715 7535
rect 5735 7518 5767 7535
rect 5788 7518 5793 7538
rect 5735 7515 5793 7518
rect 5706 7508 5793 7515
rect 5818 7535 5855 7605
rect 6121 7604 6158 7605
rect 6413 7601 6454 7609
rect 6413 7581 6421 7601
rect 6440 7581 6454 7601
rect 6413 7579 6454 7581
rect 6482 7601 6524 7609
rect 6482 7581 6498 7601
rect 6517 7581 6524 7601
rect 6750 7608 6756 7630
rect 6782 7610 7196 7630
rect 7946 7629 7983 7630
rect 8249 7629 8286 7699
rect 8311 7719 8398 7726
rect 8311 7716 8369 7719
rect 8311 7696 8316 7716
rect 8337 7699 8369 7716
rect 8389 7699 8398 7719
rect 8337 7696 8398 7699
rect 8311 7689 8398 7696
rect 8457 7719 8494 7729
rect 8457 7699 8465 7719
rect 8485 7699 8494 7719
rect 8311 7688 8342 7689
rect 7945 7628 8286 7629
rect 6782 7608 6791 7610
rect 7028 7609 7196 7610
rect 7870 7623 8286 7628
rect 6750 7599 6791 7608
rect 7870 7603 7873 7623
rect 7893 7603 8286 7623
rect 8457 7620 8494 7699
rect 8524 7728 8555 7781
rect 9192 7770 9725 7786
rect 9192 7759 9724 7770
rect 9843 7761 9880 7765
rect 8574 7728 8611 7729
rect 8524 7719 8611 7728
rect 8524 7699 8582 7719
rect 8602 7699 8611 7719
rect 8524 7689 8611 7699
rect 8670 7719 8707 7729
rect 8670 7699 8678 7719
rect 8698 7699 8707 7719
rect 8524 7688 8555 7689
rect 8519 7620 8629 7633
rect 8670 7620 8707 7699
rect 8457 7618 8707 7620
rect 8457 7615 8558 7618
rect 8457 7596 8522 7615
rect 6482 7579 6524 7581
rect 6413 7564 6524 7579
rect 8519 7588 8522 7596
rect 8551 7588 8558 7615
rect 8586 7591 8596 7618
rect 8625 7596 8707 7618
rect 8785 7690 8953 7691
rect 9192 7690 9230 7759
rect 8785 7670 9230 7690
rect 9457 7721 9568 7736
rect 9457 7719 9499 7721
rect 9457 7699 9464 7719
rect 9483 7699 9499 7719
rect 9457 7691 9499 7699
rect 9527 7719 9568 7721
rect 9527 7699 9541 7719
rect 9560 7699 9568 7719
rect 9527 7691 9568 7699
rect 9457 7685 9568 7691
rect 9690 7696 9724 7759
rect 9842 7755 9880 7761
rect 9842 7737 9852 7755
rect 9870 7737 9880 7755
rect 9842 7728 9880 7737
rect 9842 7696 9876 7728
rect 8785 7664 9229 7670
rect 8785 7662 8953 7664
rect 8625 7591 8629 7596
rect 8586 7588 8629 7591
rect 8519 7574 8629 7588
rect 5970 7545 6006 7546
rect 5818 7515 5827 7535
rect 5847 7515 5855 7535
rect 5706 7506 5762 7508
rect 5706 7505 5743 7506
rect 5818 7505 5855 7515
rect 5914 7535 6062 7545
rect 6162 7542 6258 7544
rect 5914 7515 5923 7535
rect 5943 7515 6033 7535
rect 6053 7515 6062 7535
rect 5914 7506 6062 7515
rect 6120 7535 6258 7542
rect 6120 7515 6129 7535
rect 6149 7515 6258 7535
rect 6120 7506 6258 7515
rect 5914 7505 5951 7506
rect 5970 7454 6006 7506
rect 6025 7505 6062 7506
rect 6121 7505 6158 7506
rect 5441 7452 5482 7453
rect 5333 7445 5482 7452
rect 5333 7425 5451 7445
rect 5471 7425 5482 7445
rect 5333 7417 5482 7425
rect 5549 7449 5908 7453
rect 5549 7444 5871 7449
rect 5549 7420 5662 7444
rect 5686 7425 5871 7444
rect 5895 7425 5908 7449
rect 5686 7420 5908 7425
rect 5549 7417 5908 7420
rect 5970 7417 6005 7454
rect 6073 7451 6173 7454
rect 6073 7447 6140 7451
rect 6073 7421 6085 7447
rect 6111 7425 6140 7447
rect 6166 7425 6173 7451
rect 6111 7421 6173 7425
rect 6073 7417 6173 7421
rect 5549 7396 5580 7417
rect 5970 7396 6006 7417
rect 5392 7395 5429 7396
rect 5391 7386 5429 7395
rect 5391 7366 5400 7386
rect 5420 7366 5429 7386
rect 5391 7358 5429 7366
rect 5495 7390 5580 7396
rect 5605 7395 5642 7396
rect 5495 7370 5503 7390
rect 5523 7370 5580 7390
rect 5495 7362 5580 7370
rect 5604 7386 5642 7395
rect 5604 7366 5613 7386
rect 5633 7366 5642 7386
rect 5495 7361 5531 7362
rect 5604 7358 5642 7366
rect 5708 7390 5793 7396
rect 5813 7395 5850 7396
rect 5708 7370 5716 7390
rect 5736 7389 5793 7390
rect 5736 7370 5765 7389
rect 5708 7369 5765 7370
rect 5786 7369 5793 7389
rect 5708 7362 5793 7369
rect 5812 7386 5850 7395
rect 5812 7366 5821 7386
rect 5841 7366 5850 7386
rect 5708 7361 5744 7362
rect 5812 7358 5850 7366
rect 5916 7390 6060 7396
rect 5916 7370 5924 7390
rect 5944 7387 6032 7390
rect 5944 7370 5975 7387
rect 5916 7367 5975 7370
rect 5998 7370 6032 7387
rect 6052 7370 6060 7390
rect 5998 7367 6060 7370
rect 5916 7362 6060 7367
rect 5916 7361 5952 7362
rect 6024 7361 6060 7362
rect 6126 7395 6163 7396
rect 6126 7394 6164 7395
rect 6126 7386 6190 7394
rect 6126 7366 6135 7386
rect 6155 7372 6190 7386
rect 6210 7372 6213 7392
rect 6155 7367 6213 7372
rect 6155 7366 6190 7367
rect 5392 7329 5429 7358
rect 5393 7327 5429 7329
rect 5605 7327 5642 7358
rect 5393 7305 5642 7327
rect 5813 7326 5850 7358
rect 6126 7354 6190 7366
rect 6230 7328 6257 7506
rect 8785 7484 8812 7662
rect 8852 7624 8916 7636
rect 9192 7632 9229 7664
rect 9400 7663 9649 7685
rect 9690 7664 9876 7696
rect 9704 7663 9876 7664
rect 9400 7632 9437 7663
rect 9613 7661 9649 7663
rect 9613 7632 9650 7661
rect 9842 7635 9876 7663
rect 8852 7623 8887 7624
rect 8829 7618 8887 7623
rect 8829 7598 8832 7618
rect 8852 7604 8887 7618
rect 8907 7604 8916 7624
rect 8852 7596 8916 7604
rect 8878 7595 8916 7596
rect 8879 7594 8916 7595
rect 8982 7628 9018 7629
rect 9090 7628 9126 7629
rect 8982 7621 9126 7628
rect 8982 7620 9042 7621
rect 8982 7600 8990 7620
rect 9010 7601 9042 7620
rect 9067 7620 9126 7621
rect 9067 7601 9098 7620
rect 9010 7600 9098 7601
rect 9118 7600 9126 7620
rect 8982 7594 9126 7600
rect 9192 7624 9230 7632
rect 9298 7628 9334 7629
rect 9192 7604 9201 7624
rect 9221 7604 9230 7624
rect 9192 7595 9230 7604
rect 9249 7621 9334 7628
rect 9249 7601 9256 7621
rect 9277 7620 9334 7621
rect 9277 7601 9306 7620
rect 9249 7600 9306 7601
rect 9326 7600 9334 7620
rect 9192 7594 9229 7595
rect 9249 7594 9334 7600
rect 9400 7624 9438 7632
rect 9511 7628 9547 7629
rect 9400 7604 9409 7624
rect 9429 7604 9438 7624
rect 9400 7595 9438 7604
rect 9462 7620 9547 7628
rect 9462 7600 9519 7620
rect 9539 7600 9547 7620
rect 9400 7594 9437 7595
rect 9462 7594 9547 7600
rect 9613 7624 9651 7632
rect 9613 7604 9622 7624
rect 9642 7604 9651 7624
rect 9613 7595 9651 7604
rect 9840 7625 9877 7635
rect 9840 7607 9850 7625
rect 9868 7607 9877 7625
rect 9840 7598 9877 7607
rect 9842 7597 9876 7598
rect 9613 7594 9650 7595
rect 9036 7573 9072 7594
rect 9462 7573 9493 7594
rect 8869 7569 8969 7573
rect 8869 7565 8931 7569
rect 8869 7539 8876 7565
rect 8902 7543 8931 7565
rect 8957 7543 8969 7569
rect 8902 7539 8969 7543
rect 8869 7536 8969 7539
rect 9037 7536 9072 7573
rect 9134 7570 9493 7573
rect 9134 7565 9356 7570
rect 9134 7541 9147 7565
rect 9171 7546 9356 7565
rect 9380 7546 9493 7570
rect 9171 7541 9493 7546
rect 9134 7537 9493 7541
rect 9560 7565 9709 7573
rect 9560 7545 9571 7565
rect 9591 7545 9709 7565
rect 9560 7538 9709 7545
rect 9560 7537 9601 7538
rect 8884 7484 8921 7485
rect 8980 7484 9017 7485
rect 9036 7484 9072 7536
rect 9091 7484 9128 7485
rect 8784 7475 8922 7484
rect 8409 7441 8520 7456
rect 8784 7455 8893 7475
rect 8913 7455 8922 7475
rect 8784 7448 8922 7455
rect 8980 7475 9128 7484
rect 8980 7455 8989 7475
rect 9009 7455 9099 7475
rect 9119 7455 9128 7475
rect 8784 7446 8880 7448
rect 8980 7445 9128 7455
rect 9187 7475 9224 7485
rect 9299 7484 9336 7485
rect 9280 7482 9336 7484
rect 9187 7455 9195 7475
rect 9215 7455 9224 7475
rect 9036 7444 9072 7445
rect 8409 7439 8451 7441
rect 7746 7420 7816 7429
rect 7746 7411 7763 7420
rect 7737 7391 7763 7411
rect 7811 7411 7816 7420
rect 8409 7419 8416 7439
rect 8435 7419 8451 7439
rect 8409 7411 8451 7419
rect 8479 7439 8520 7441
rect 8479 7419 8493 7439
rect 8512 7419 8520 7439
rect 8479 7411 8520 7419
rect 7811 7410 7905 7411
rect 7811 7391 8181 7410
rect 8409 7405 8520 7411
rect 6524 7377 6634 7391
rect 6524 7374 6567 7377
rect 6524 7369 6528 7374
rect 6089 7326 6257 7328
rect 5813 7323 6257 7326
rect 5474 7299 5585 7305
rect 5474 7291 5515 7299
rect 5163 7236 5202 7280
rect 5474 7271 5482 7291
rect 5501 7271 5515 7291
rect 5474 7269 5515 7271
rect 5543 7291 5585 7299
rect 5543 7271 5559 7291
rect 5578 7271 5585 7291
rect 5543 7269 5585 7271
rect 5474 7255 5585 7269
rect 5811 7300 6257 7323
rect 3456 7216 3497 7217
rect 2932 7175 2968 7215
rect 2780 7163 2817 7164
rect 2876 7163 2913 7164
rect 2932 7163 2937 7175
rect 2680 7154 2818 7163
rect 2680 7134 2789 7154
rect 2809 7134 2818 7154
rect 2680 7127 2818 7134
rect 2876 7154 2937 7163
rect 2876 7134 2885 7154
rect 2905 7143 2937 7154
rect 2964 7163 2968 7175
rect 2987 7163 3024 7164
rect 2964 7154 3024 7163
rect 2964 7143 2995 7154
rect 2905 7134 2995 7143
rect 3015 7134 3024 7154
rect 2680 7125 2776 7127
rect 2876 7124 3024 7134
rect 3083 7154 3120 7164
rect 3195 7163 3232 7164
rect 3176 7161 3232 7163
rect 3083 7134 3091 7154
rect 3111 7134 3120 7154
rect 2932 7123 2968 7124
rect 2780 7064 2817 7065
rect 3083 7064 3120 7134
rect 3145 7154 3232 7161
rect 3145 7151 3203 7154
rect 3145 7131 3150 7151
rect 3171 7134 3203 7151
rect 3223 7134 3232 7154
rect 3171 7131 3232 7134
rect 3145 7124 3232 7131
rect 3291 7154 3328 7164
rect 3291 7134 3299 7154
rect 3319 7134 3328 7154
rect 3145 7123 3176 7124
rect 2779 7063 3120 7064
rect 2704 7058 3120 7063
rect 2704 7040 2707 7058
rect 2727 7056 3120 7058
rect 2727 7040 3097 7056
rect 2745 7038 3097 7040
rect 3088 7036 3097 7038
rect 3118 7036 3120 7056
rect 3088 7024 3120 7036
rect 3291 7055 3328 7134
rect 3358 7163 3389 7216
rect 4138 7188 4824 7221
rect 3408 7163 3445 7164
rect 3358 7154 3445 7163
rect 3358 7134 3416 7154
rect 3436 7134 3445 7154
rect 3358 7124 3445 7134
rect 3504 7154 3541 7164
rect 3504 7134 3512 7154
rect 3532 7134 3541 7154
rect 3358 7123 3389 7124
rect 3353 7055 3463 7068
rect 3504 7055 3541 7134
rect 3291 7053 3541 7055
rect 3291 7050 3392 7053
rect 3291 7031 3356 7050
rect 2131 7018 2250 7020
rect 2082 7016 2250 7018
rect 1467 6989 1578 6995
rect 1806 6990 2250 7016
rect 3353 7023 3356 7031
rect 3385 7023 3392 7050
rect 3420 7026 3430 7053
rect 3459 7031 3541 7053
rect 3730 7100 3898 7101
rect 4138 7100 4176 7188
rect 4437 7186 4484 7188
rect 4784 7164 4824 7188
rect 5163 7212 5203 7236
rect 5503 7212 5550 7214
rect 5811 7212 5849 7300
rect 6089 7299 6257 7300
rect 6446 7347 6528 7369
rect 6557 7347 6567 7374
rect 6595 7350 6602 7377
rect 6631 7369 6634 7377
rect 7737 7384 8181 7391
rect 7737 7382 7905 7384
rect 7737 7374 7816 7382
rect 6631 7350 6696 7369
rect 6595 7347 6696 7350
rect 6446 7345 6696 7347
rect 6446 7266 6483 7345
rect 6524 7332 6634 7345
rect 6598 7276 6629 7277
rect 6446 7246 6455 7266
rect 6475 7246 6483 7266
rect 6446 7236 6483 7246
rect 6542 7266 6629 7276
rect 6542 7246 6551 7266
rect 6571 7246 6629 7266
rect 6542 7237 6629 7246
rect 6542 7236 6579 7237
rect 5163 7179 5849 7212
rect 6598 7184 6629 7237
rect 6659 7266 6696 7345
rect 6867 7342 7260 7362
rect 7280 7342 7283 7362
rect 6867 7337 7283 7342
rect 6867 7336 7208 7337
rect 6811 7276 6842 7277
rect 6659 7246 6668 7266
rect 6688 7246 6696 7266
rect 6659 7236 6696 7246
rect 6755 7269 6842 7276
rect 6755 7266 6816 7269
rect 6755 7246 6764 7266
rect 6784 7249 6816 7266
rect 6837 7249 6842 7269
rect 6784 7246 6842 7249
rect 6755 7239 6842 7246
rect 6867 7266 6904 7336
rect 7170 7335 7207 7336
rect 7019 7276 7055 7277
rect 6867 7246 6876 7266
rect 6896 7246 6904 7266
rect 6755 7237 6811 7239
rect 6755 7236 6792 7237
rect 6867 7236 6904 7246
rect 6963 7266 7111 7276
rect 7211 7273 7307 7275
rect 6963 7246 6972 7266
rect 6992 7246 7082 7266
rect 7102 7246 7111 7266
rect 6963 7237 7111 7246
rect 7169 7266 7307 7273
rect 7169 7246 7178 7266
rect 7198 7246 7307 7266
rect 7169 7237 7307 7246
rect 6963 7236 7000 7237
rect 7019 7185 7055 7237
rect 7074 7236 7111 7237
rect 7170 7236 7207 7237
rect 6490 7183 6531 7184
rect 3730 7077 4176 7100
rect 4402 7131 4513 7145
rect 4402 7129 4444 7131
rect 4402 7109 4409 7129
rect 4428 7109 4444 7129
rect 4402 7101 4444 7109
rect 4472 7129 4513 7131
rect 4472 7109 4486 7129
rect 4505 7109 4513 7129
rect 4785 7120 4824 7164
rect 4472 7101 4513 7109
rect 4402 7095 4513 7101
rect 3730 7074 4174 7077
rect 3730 7072 3898 7074
rect 3459 7026 3463 7031
rect 3420 7023 3463 7026
rect 3353 7009 3463 7023
rect 2082 6989 2250 6990
rect 1467 6981 1508 6989
rect 1467 6961 1475 6981
rect 1494 6961 1508 6981
rect 1467 6959 1508 6961
rect 1536 6981 1578 6989
rect 2131 6988 2239 6989
rect 1536 6961 1552 6981
rect 1571 6961 1578 6981
rect 1536 6959 1578 6961
rect 915 6955 951 6956
rect 763 6925 772 6945
rect 792 6925 800 6945
rect 651 6916 707 6918
rect 651 6915 688 6916
rect 763 6915 800 6925
rect 859 6945 1007 6955
rect 1107 6952 1203 6954
rect 859 6925 868 6945
rect 888 6925 978 6945
rect 998 6925 1007 6945
rect 859 6916 1007 6925
rect 1065 6945 1203 6952
rect 1065 6925 1074 6945
rect 1094 6925 1203 6945
rect 1467 6944 1578 6959
rect 2169 6987 2239 6988
rect 1065 6916 1203 6925
rect 859 6915 896 6916
rect 915 6864 951 6916
rect 970 6915 1007 6916
rect 1066 6915 1103 6916
rect 386 6862 427 6863
rect 278 6855 427 6862
rect 278 6835 396 6855
rect 416 6835 427 6855
rect 278 6827 427 6835
rect 494 6859 853 6863
rect 494 6854 816 6859
rect 494 6830 607 6854
rect 631 6835 816 6854
rect 840 6835 853 6859
rect 631 6830 853 6835
rect 494 6827 853 6830
rect 915 6827 950 6864
rect 1018 6861 1118 6864
rect 1018 6857 1085 6861
rect 1018 6831 1030 6857
rect 1056 6835 1085 6857
rect 1111 6835 1118 6861
rect 1056 6831 1118 6835
rect 1018 6827 1118 6831
rect 494 6806 525 6827
rect 915 6806 951 6827
rect 337 6805 374 6806
rect 111 6802 145 6803
rect 110 6793 147 6802
rect 110 6775 119 6793
rect 137 6775 147 6793
rect 110 6765 147 6775
rect 336 6796 374 6805
rect 336 6776 345 6796
rect 365 6776 374 6796
rect 336 6768 374 6776
rect 440 6800 525 6806
rect 550 6805 587 6806
rect 440 6780 448 6800
rect 468 6780 525 6800
rect 440 6772 525 6780
rect 549 6796 587 6805
rect 549 6776 558 6796
rect 578 6776 587 6796
rect 440 6771 476 6772
rect 549 6768 587 6776
rect 653 6800 738 6806
rect 758 6805 795 6806
rect 653 6780 661 6800
rect 681 6799 738 6800
rect 681 6780 710 6799
rect 653 6779 710 6780
rect 731 6779 738 6799
rect 653 6772 738 6779
rect 757 6796 795 6805
rect 757 6776 766 6796
rect 786 6776 795 6796
rect 653 6771 689 6772
rect 757 6768 795 6776
rect 861 6800 1005 6806
rect 861 6780 869 6800
rect 889 6799 977 6800
rect 889 6780 920 6799
rect 861 6779 920 6780
rect 945 6780 977 6799
rect 997 6780 1005 6800
rect 945 6779 1005 6780
rect 861 6772 1005 6779
rect 861 6771 897 6772
rect 969 6771 1005 6772
rect 1071 6805 1108 6806
rect 1071 6804 1109 6805
rect 1071 6796 1135 6804
rect 1071 6776 1080 6796
rect 1100 6782 1135 6796
rect 1155 6782 1158 6802
rect 1100 6777 1158 6782
rect 1100 6776 1135 6777
rect 111 6737 145 6765
rect 337 6739 374 6768
rect 338 6737 374 6739
rect 550 6737 587 6768
rect 111 6736 283 6737
rect 111 6704 297 6736
rect 338 6715 587 6737
rect 758 6736 795 6768
rect 1071 6764 1135 6776
rect 1175 6738 1202 6916
rect 2169 6880 2230 6987
rect 3730 6894 3757 7072
rect 3797 7034 3861 7046
rect 4137 7042 4174 7074
rect 4345 7073 4594 7095
rect 4345 7042 4382 7073
rect 4558 7071 4594 7073
rect 4558 7042 4595 7071
rect 3797 7033 3832 7034
rect 3774 7028 3832 7033
rect 3774 7008 3777 7028
rect 3797 7014 3832 7028
rect 3852 7014 3861 7034
rect 3797 7006 3861 7014
rect 3823 7005 3861 7006
rect 3824 7004 3861 7005
rect 3927 7038 3963 7039
rect 4035 7038 4071 7039
rect 3927 7033 4071 7038
rect 3927 7030 3989 7033
rect 3927 7010 3935 7030
rect 3955 7013 3989 7030
rect 4012 7030 4071 7033
rect 4012 7013 4043 7030
rect 3955 7010 4043 7013
rect 4063 7010 4071 7030
rect 3927 7004 4071 7010
rect 4137 7034 4175 7042
rect 4243 7038 4279 7039
rect 4137 7014 4146 7034
rect 4166 7014 4175 7034
rect 4137 7005 4175 7014
rect 4194 7031 4279 7038
rect 4194 7011 4201 7031
rect 4222 7030 4279 7031
rect 4222 7011 4251 7030
rect 4194 7010 4251 7011
rect 4271 7010 4279 7030
rect 4137 7004 4174 7005
rect 4194 7004 4279 7010
rect 4345 7034 4383 7042
rect 4456 7038 4492 7039
rect 4345 7014 4354 7034
rect 4374 7014 4383 7034
rect 4345 7005 4383 7014
rect 4407 7030 4492 7038
rect 4407 7010 4464 7030
rect 4484 7010 4492 7030
rect 4345 7004 4382 7005
rect 4407 7004 4492 7010
rect 4558 7034 4596 7042
rect 4558 7014 4567 7034
rect 4587 7014 4596 7034
rect 4558 7005 4596 7014
rect 4558 7004 4595 7005
rect 3981 6983 4017 7004
rect 4407 6983 4438 7004
rect 3814 6979 3914 6983
rect 3814 6975 3876 6979
rect 3814 6949 3821 6975
rect 3847 6953 3876 6975
rect 3902 6953 3914 6979
rect 3847 6949 3914 6953
rect 3814 6946 3914 6949
rect 3982 6946 4017 6983
rect 4079 6980 4438 6983
rect 4079 6975 4301 6980
rect 4079 6951 4092 6975
rect 4116 6956 4301 6975
rect 4325 6956 4438 6980
rect 4116 6951 4438 6956
rect 4079 6947 4438 6951
rect 4505 6975 4654 6983
rect 4505 6955 4516 6975
rect 4536 6955 4654 6975
rect 4505 6948 4654 6955
rect 4505 6947 4546 6948
rect 3829 6894 3866 6895
rect 3925 6894 3962 6895
rect 3981 6894 4017 6946
rect 4036 6894 4073 6895
rect 3729 6885 3867 6894
rect 2169 6869 2239 6880
rect 2169 6860 2176 6869
rect 2171 6840 2176 6860
rect 2224 6840 2239 6869
rect 3729 6865 3838 6885
rect 3858 6865 3867 6885
rect 3729 6858 3867 6865
rect 3925 6885 4073 6894
rect 3925 6865 3934 6885
rect 3954 6865 4044 6885
rect 4064 6865 4073 6885
rect 3729 6856 3825 6858
rect 3925 6855 4073 6865
rect 4132 6885 4169 6895
rect 4244 6894 4281 6895
rect 4225 6892 4281 6894
rect 4132 6865 4140 6885
rect 4160 6865 4169 6885
rect 3981 6854 4017 6855
rect 2171 6831 2239 6840
rect 1358 6812 1468 6826
rect 1358 6809 1401 6812
rect 1358 6804 1362 6809
rect 1034 6736 1202 6738
rect 758 6730 1202 6736
rect 111 6672 145 6704
rect 107 6663 145 6672
rect 107 6645 117 6663
rect 135 6645 145 6663
rect 107 6639 145 6645
rect 263 6641 297 6704
rect 419 6709 530 6715
rect 419 6701 460 6709
rect 419 6681 427 6701
rect 446 6681 460 6701
rect 419 6679 460 6681
rect 488 6701 530 6709
rect 488 6681 504 6701
rect 523 6681 530 6701
rect 488 6679 530 6681
rect 419 6664 530 6679
rect 757 6710 1202 6730
rect 757 6641 795 6710
rect 1034 6709 1202 6710
rect 1280 6782 1362 6804
rect 1391 6782 1401 6809
rect 1429 6785 1436 6812
rect 1465 6804 1468 6812
rect 3463 6821 3574 6836
rect 3463 6819 3505 6821
rect 1465 6785 1530 6804
rect 1429 6782 1530 6785
rect 1280 6780 1530 6782
rect 1280 6701 1317 6780
rect 1358 6767 1468 6780
rect 1432 6711 1463 6712
rect 1280 6681 1289 6701
rect 1309 6681 1317 6701
rect 1280 6671 1317 6681
rect 1376 6701 1463 6711
rect 1376 6681 1385 6701
rect 1405 6681 1463 6701
rect 1376 6672 1463 6681
rect 1376 6671 1413 6672
rect 107 6635 144 6639
rect 263 6630 795 6641
rect 262 6614 795 6630
rect 1432 6619 1463 6672
rect 1493 6701 1530 6780
rect 1701 6777 2094 6797
rect 2114 6777 2117 6797
rect 3196 6792 3237 6801
rect 1701 6772 2117 6777
rect 2791 6790 2959 6791
rect 3196 6790 3205 6792
rect 1701 6771 2042 6772
rect 1645 6711 1676 6712
rect 1493 6681 1502 6701
rect 1522 6681 1530 6701
rect 1493 6671 1530 6681
rect 1589 6704 1676 6711
rect 1589 6701 1650 6704
rect 1589 6681 1598 6701
rect 1618 6684 1650 6701
rect 1671 6684 1676 6704
rect 1618 6681 1676 6684
rect 1589 6674 1676 6681
rect 1701 6701 1738 6771
rect 2004 6770 2041 6771
rect 2791 6770 3205 6790
rect 3231 6770 3237 6792
rect 3463 6799 3470 6819
rect 3489 6799 3505 6819
rect 3463 6791 3505 6799
rect 3533 6819 3574 6821
rect 3533 6799 3547 6819
rect 3566 6799 3574 6819
rect 3533 6791 3574 6799
rect 3829 6795 3866 6796
rect 4132 6795 4169 6865
rect 4194 6885 4281 6892
rect 4194 6882 4252 6885
rect 4194 6862 4199 6882
rect 4220 6865 4252 6882
rect 4272 6865 4281 6885
rect 4220 6862 4281 6865
rect 4194 6855 4281 6862
rect 4340 6885 4377 6895
rect 4340 6865 4348 6885
rect 4368 6865 4377 6885
rect 4194 6854 4225 6855
rect 3828 6794 4169 6795
rect 3463 6785 3574 6791
rect 3753 6789 4169 6794
rect 2791 6764 3237 6770
rect 2791 6762 2959 6764
rect 1853 6711 1889 6712
rect 1701 6681 1710 6701
rect 1730 6681 1738 6701
rect 1589 6672 1645 6674
rect 1589 6671 1626 6672
rect 1701 6671 1738 6681
rect 1797 6701 1945 6711
rect 2045 6708 2141 6710
rect 1797 6681 1806 6701
rect 1826 6681 1916 6701
rect 1936 6681 1945 6701
rect 1797 6672 1945 6681
rect 2003 6701 2141 6708
rect 2003 6681 2012 6701
rect 2032 6681 2141 6701
rect 2003 6672 2141 6681
rect 1797 6671 1834 6672
rect 1853 6620 1889 6672
rect 1908 6671 1945 6672
rect 2004 6671 2041 6672
rect 1324 6618 1365 6619
rect 262 6613 776 6614
rect 1216 6611 1365 6618
rect 1216 6591 1334 6611
rect 1354 6591 1365 6611
rect 1216 6583 1365 6591
rect 1432 6615 1791 6619
rect 1432 6610 1754 6615
rect 1432 6586 1545 6610
rect 1569 6591 1754 6610
rect 1778 6591 1791 6615
rect 1569 6586 1791 6591
rect 1432 6583 1791 6586
rect 1853 6583 1888 6620
rect 1956 6617 2056 6620
rect 1956 6613 2023 6617
rect 1956 6587 1968 6613
rect 1994 6591 2023 6613
rect 2049 6591 2056 6617
rect 1994 6587 2056 6591
rect 1956 6583 2056 6587
rect 110 6572 147 6573
rect 108 6564 148 6572
rect 108 6546 119 6564
rect 137 6546 148 6564
rect 1432 6562 1463 6583
rect 1853 6562 1889 6583
rect 1275 6561 1312 6562
rect 108 6498 148 6546
rect 1274 6552 1312 6561
rect 1274 6532 1283 6552
rect 1303 6532 1312 6552
rect 1274 6524 1312 6532
rect 1378 6556 1463 6562
rect 1488 6561 1525 6562
rect 1378 6536 1386 6556
rect 1406 6536 1463 6556
rect 1378 6528 1463 6536
rect 1487 6552 1525 6561
rect 1487 6532 1496 6552
rect 1516 6532 1525 6552
rect 1378 6527 1414 6528
rect 1487 6524 1525 6532
rect 1591 6556 1676 6562
rect 1696 6561 1733 6562
rect 1591 6536 1599 6556
rect 1619 6555 1676 6556
rect 1619 6536 1648 6555
rect 1591 6535 1648 6536
rect 1669 6535 1676 6555
rect 1591 6528 1676 6535
rect 1695 6552 1733 6561
rect 1695 6532 1704 6552
rect 1724 6532 1733 6552
rect 1591 6527 1627 6528
rect 1695 6524 1733 6532
rect 1799 6556 1943 6562
rect 1799 6536 1807 6556
rect 1827 6539 1863 6556
rect 1883 6539 1915 6556
rect 1827 6536 1915 6539
rect 1935 6536 1943 6556
rect 1799 6528 1943 6536
rect 1799 6527 1835 6528
rect 1907 6527 1943 6528
rect 2009 6561 2046 6562
rect 2009 6560 2047 6561
rect 2009 6552 2073 6560
rect 2009 6532 2018 6552
rect 2038 6538 2073 6552
rect 2093 6538 2096 6558
rect 2038 6533 2096 6538
rect 2038 6532 2073 6533
rect 419 6502 529 6516
rect 419 6499 462 6502
rect 108 6491 233 6498
rect 419 6494 423 6499
rect 108 6472 200 6491
rect 225 6472 233 6491
rect 108 6462 233 6472
rect 341 6472 423 6494
rect 452 6472 462 6499
rect 490 6475 497 6502
rect 526 6494 529 6502
rect 1275 6495 1312 6524
rect 526 6475 591 6494
rect 1276 6493 1312 6495
rect 1488 6493 1525 6524
rect 1696 6497 1733 6524
rect 2009 6520 2073 6532
rect 490 6472 591 6475
rect 341 6470 591 6472
rect 108 6442 148 6462
rect 107 6433 148 6442
rect 107 6415 117 6433
rect 135 6415 148 6433
rect 107 6406 148 6415
rect 107 6405 144 6406
rect 341 6391 378 6470
rect 419 6457 529 6470
rect 493 6401 524 6402
rect 341 6371 350 6391
rect 370 6371 378 6391
rect 341 6361 378 6371
rect 437 6391 524 6401
rect 437 6371 446 6391
rect 466 6371 524 6391
rect 437 6362 524 6371
rect 437 6361 474 6362
rect 110 6339 147 6343
rect 107 6334 147 6339
rect 107 6316 119 6334
rect 137 6316 147 6334
rect 107 6136 147 6316
rect 493 6309 524 6362
rect 554 6391 591 6470
rect 762 6467 1155 6487
rect 1175 6467 1178 6487
rect 1276 6471 1525 6493
rect 1694 6492 1735 6497
rect 2113 6494 2140 6672
rect 2791 6584 2818 6762
rect 3196 6759 3237 6764
rect 3406 6763 3655 6785
rect 3753 6769 3756 6789
rect 3776 6769 4169 6789
rect 4340 6786 4377 6865
rect 4407 6894 4438 6947
rect 4784 6940 4824 7120
rect 5162 7122 5201 7179
rect 5811 7177 5849 7179
rect 6382 7176 6531 7183
rect 6382 7156 6500 7176
rect 6520 7156 6531 7176
rect 6382 7148 6531 7156
rect 6598 7180 6957 7184
rect 6598 7175 6920 7180
rect 6598 7151 6711 7175
rect 6735 7156 6920 7175
rect 6944 7156 6957 7180
rect 6735 7151 6957 7156
rect 6598 7148 6957 7151
rect 7019 7148 7054 7185
rect 7122 7182 7222 7185
rect 7122 7178 7189 7182
rect 7122 7152 7134 7178
rect 7160 7156 7189 7178
rect 7215 7156 7222 7182
rect 7160 7152 7222 7156
rect 7122 7148 7222 7152
rect 6598 7127 6629 7148
rect 7019 7127 7055 7148
rect 6441 7126 6478 7127
rect 5162 7120 5210 7122
rect 5162 7102 5173 7120
rect 5191 7102 5210 7120
rect 6440 7117 6478 7126
rect 5162 7093 5210 7102
rect 5163 7092 5210 7093
rect 5476 7097 5586 7111
rect 5476 7094 5519 7097
rect 5476 7089 5480 7094
rect 5398 7067 5480 7089
rect 5509 7067 5519 7094
rect 5547 7070 5554 7097
rect 5583 7089 5586 7097
rect 6440 7097 6449 7117
rect 6469 7097 6478 7117
rect 6440 7089 6478 7097
rect 6544 7121 6629 7127
rect 6654 7126 6691 7127
rect 6544 7101 6552 7121
rect 6572 7101 6629 7121
rect 6544 7093 6629 7101
rect 6653 7117 6691 7126
rect 6653 7097 6662 7117
rect 6682 7097 6691 7117
rect 6544 7092 6580 7093
rect 6653 7089 6691 7097
rect 6757 7121 6842 7127
rect 6862 7126 6899 7127
rect 6757 7101 6765 7121
rect 6785 7120 6842 7121
rect 6785 7101 6814 7120
rect 6757 7100 6814 7101
rect 6835 7100 6842 7120
rect 6757 7093 6842 7100
rect 6861 7117 6899 7126
rect 6861 7097 6870 7117
rect 6890 7097 6899 7117
rect 6757 7092 6793 7093
rect 6861 7089 6899 7097
rect 6965 7121 7109 7127
rect 6965 7101 6973 7121
rect 6993 7119 7081 7121
rect 6993 7101 7022 7119
rect 6965 7100 7022 7101
rect 7051 7101 7081 7119
rect 7101 7101 7109 7121
rect 7051 7100 7109 7101
rect 6965 7093 7109 7100
rect 6965 7092 7001 7093
rect 7073 7092 7109 7093
rect 7175 7126 7212 7127
rect 7175 7125 7213 7126
rect 7175 7117 7239 7125
rect 7175 7097 7184 7117
rect 7204 7103 7239 7117
rect 7259 7103 7262 7123
rect 7204 7098 7262 7103
rect 7204 7097 7239 7098
rect 5583 7070 5648 7089
rect 5547 7067 5648 7070
rect 5398 7065 5648 7067
rect 5166 7029 5203 7030
rect 4784 6922 4794 6940
rect 4812 6922 4824 6940
rect 4784 6917 4824 6922
rect 5162 7026 5203 7029
rect 5162 7021 5204 7026
rect 5162 7003 5175 7021
rect 5193 7003 5204 7021
rect 5162 6989 5204 7003
rect 5242 6989 5289 6993
rect 5162 6983 5289 6989
rect 5162 6954 5250 6983
rect 5279 6954 5289 6983
rect 5398 6986 5435 7065
rect 5476 7052 5586 7065
rect 5550 6996 5581 6997
rect 5398 6966 5407 6986
rect 5427 6966 5435 6986
rect 5398 6956 5435 6966
rect 5494 6986 5581 6996
rect 5494 6966 5503 6986
rect 5523 6966 5581 6986
rect 5494 6957 5581 6966
rect 5494 6956 5531 6957
rect 5162 6950 5289 6954
rect 5162 6933 5201 6950
rect 5242 6949 5289 6950
rect 4784 6913 4821 6917
rect 5162 6915 5173 6933
rect 5191 6915 5201 6933
rect 5162 6906 5201 6915
rect 5163 6905 5200 6906
rect 5550 6904 5581 6957
rect 5611 6986 5648 7065
rect 5819 7062 6212 7082
rect 6232 7062 6235 7082
rect 5819 7057 6235 7062
rect 6441 7060 6478 7089
rect 6442 7058 6478 7060
rect 6654 7058 6691 7089
rect 5819 7056 6160 7057
rect 5763 6996 5794 6997
rect 5611 6966 5620 6986
rect 5640 6966 5648 6986
rect 5611 6956 5648 6966
rect 5707 6989 5794 6996
rect 5707 6986 5768 6989
rect 5707 6966 5716 6986
rect 5736 6969 5768 6986
rect 5789 6969 5794 6989
rect 5736 6966 5794 6969
rect 5707 6959 5794 6966
rect 5819 6986 5856 7056
rect 6122 7055 6159 7056
rect 6442 7036 6691 7058
rect 6862 7057 6899 7089
rect 7175 7085 7239 7097
rect 7279 7061 7306 7237
rect 7737 7204 7764 7374
rect 7804 7344 7868 7356
rect 8144 7352 8181 7384
rect 8352 7383 8601 7405
rect 8884 7385 8921 7386
rect 9187 7385 9224 7455
rect 9249 7475 9336 7482
rect 9249 7472 9307 7475
rect 9249 7452 9254 7472
rect 9275 7455 9307 7472
rect 9327 7455 9336 7475
rect 9275 7452 9336 7455
rect 9249 7445 9336 7452
rect 9395 7475 9432 7485
rect 9395 7455 9403 7475
rect 9423 7455 9432 7475
rect 9249 7444 9280 7445
rect 8883 7384 9224 7385
rect 8352 7352 8389 7383
rect 8565 7381 8601 7383
rect 8565 7352 8602 7381
rect 8808 7379 9224 7384
rect 8808 7359 8811 7379
rect 8831 7359 9224 7379
rect 9395 7376 9432 7455
rect 9462 7484 9493 7537
rect 9843 7535 9880 7536
rect 9842 7526 9881 7535
rect 9842 7508 9852 7526
rect 9870 7508 9881 7526
rect 9754 7491 9801 7492
rect 9842 7491 9881 7508
rect 9754 7487 9881 7491
rect 9512 7484 9549 7485
rect 9462 7475 9549 7484
rect 9462 7455 9520 7475
rect 9540 7455 9549 7475
rect 9462 7445 9549 7455
rect 9608 7475 9645 7485
rect 9608 7455 9616 7475
rect 9636 7455 9645 7475
rect 9462 7444 9493 7445
rect 9457 7376 9567 7389
rect 9608 7376 9645 7455
rect 9754 7458 9764 7487
rect 9793 7458 9881 7487
rect 9754 7452 9881 7458
rect 9754 7448 9801 7452
rect 9839 7438 9881 7452
rect 9839 7420 9850 7438
rect 9868 7420 9881 7438
rect 9839 7415 9881 7420
rect 9840 7412 9881 7415
rect 9840 7411 9877 7412
rect 9395 7374 9645 7376
rect 9395 7371 9496 7374
rect 9395 7352 9460 7371
rect 7804 7343 7839 7344
rect 7781 7338 7839 7343
rect 7781 7318 7784 7338
rect 7804 7324 7839 7338
rect 7859 7324 7868 7344
rect 7804 7316 7868 7324
rect 7830 7315 7868 7316
rect 7831 7314 7868 7315
rect 7934 7348 7970 7349
rect 8042 7348 8078 7349
rect 7934 7340 8078 7348
rect 7934 7320 7942 7340
rect 7962 7320 8050 7340
rect 8070 7320 8078 7340
rect 7934 7314 8078 7320
rect 8144 7344 8182 7352
rect 8250 7348 8286 7349
rect 8144 7324 8153 7344
rect 8173 7324 8182 7344
rect 8144 7315 8182 7324
rect 8201 7341 8286 7348
rect 8201 7321 8208 7341
rect 8229 7340 8286 7341
rect 8229 7321 8258 7340
rect 8201 7320 8258 7321
rect 8278 7320 8286 7340
rect 8144 7314 8181 7315
rect 8201 7314 8286 7320
rect 8352 7344 8390 7352
rect 8463 7348 8499 7349
rect 8352 7324 8361 7344
rect 8381 7324 8390 7344
rect 8352 7315 8390 7324
rect 8414 7340 8499 7348
rect 8414 7320 8471 7340
rect 8491 7320 8499 7340
rect 8352 7314 8389 7315
rect 8414 7314 8499 7320
rect 8565 7344 8603 7352
rect 8565 7324 8574 7344
rect 8594 7324 8603 7344
rect 9457 7344 9460 7352
rect 9489 7344 9496 7371
rect 9524 7347 9534 7374
rect 9563 7352 9645 7374
rect 9563 7347 9567 7352
rect 9524 7344 9567 7347
rect 9457 7330 9567 7344
rect 9833 7348 9880 7349
rect 9833 7339 9881 7348
rect 8565 7315 8603 7324
rect 9833 7321 9852 7339
rect 9870 7321 9881 7339
rect 9833 7319 9881 7321
rect 8565 7314 8602 7315
rect 7988 7293 8024 7314
rect 8414 7293 8445 7314
rect 7821 7289 7921 7293
rect 7821 7285 7883 7289
rect 7821 7259 7828 7285
rect 7854 7263 7883 7285
rect 7909 7263 7921 7289
rect 7854 7259 7921 7263
rect 7821 7256 7921 7259
rect 7989 7256 8024 7293
rect 8086 7290 8445 7293
rect 8086 7285 8308 7290
rect 8086 7261 8099 7285
rect 8123 7266 8308 7285
rect 8332 7266 8445 7290
rect 8123 7261 8445 7266
rect 8086 7257 8445 7261
rect 8512 7285 8661 7293
rect 8512 7265 8523 7285
rect 8543 7265 8661 7285
rect 8512 7258 8661 7265
rect 9194 7262 9232 7264
rect 9842 7262 9881 7319
rect 8512 7257 8553 7258
rect 7988 7216 8024 7256
rect 7836 7204 7873 7205
rect 7932 7204 7969 7205
rect 7988 7204 7993 7216
rect 7736 7195 7874 7204
rect 7736 7175 7845 7195
rect 7865 7175 7874 7195
rect 7736 7168 7874 7175
rect 7932 7195 7993 7204
rect 7932 7175 7941 7195
rect 7961 7184 7993 7195
rect 8020 7204 8024 7216
rect 8043 7204 8080 7205
rect 8020 7195 8080 7204
rect 8020 7184 8051 7195
rect 7961 7175 8051 7184
rect 8071 7175 8080 7195
rect 7736 7166 7832 7168
rect 7932 7165 8080 7175
rect 8139 7195 8176 7205
rect 8251 7204 8288 7205
rect 8232 7202 8288 7204
rect 8139 7175 8147 7195
rect 8167 7175 8176 7195
rect 7988 7164 8024 7165
rect 7836 7105 7873 7106
rect 8139 7105 8176 7175
rect 8201 7195 8288 7202
rect 8201 7192 8259 7195
rect 8201 7172 8206 7192
rect 8227 7175 8259 7192
rect 8279 7175 8288 7195
rect 8227 7172 8288 7175
rect 8201 7165 8288 7172
rect 8347 7195 8384 7205
rect 8347 7175 8355 7195
rect 8375 7175 8384 7195
rect 8201 7164 8232 7165
rect 7835 7104 8176 7105
rect 7760 7099 8176 7104
rect 7760 7081 7763 7099
rect 7783 7097 8176 7099
rect 7783 7081 8153 7097
rect 7801 7079 8153 7081
rect 8144 7077 8153 7079
rect 8174 7077 8176 7097
rect 8144 7065 8176 7077
rect 8347 7096 8384 7175
rect 8414 7204 8445 7257
rect 9194 7229 9880 7262
rect 8464 7204 8501 7205
rect 8414 7195 8501 7204
rect 8414 7175 8472 7195
rect 8492 7175 8501 7195
rect 8414 7165 8501 7175
rect 8560 7195 8597 7205
rect 8560 7175 8568 7195
rect 8588 7175 8597 7195
rect 8414 7164 8445 7165
rect 8409 7096 8519 7109
rect 8560 7096 8597 7175
rect 8347 7094 8597 7096
rect 8347 7091 8448 7094
rect 8347 7072 8412 7091
rect 7187 7059 7306 7061
rect 7138 7057 7306 7059
rect 6523 7030 6634 7036
rect 6862 7031 7306 7057
rect 8409 7064 8412 7072
rect 8441 7064 8448 7091
rect 8476 7067 8486 7094
rect 8515 7072 8597 7094
rect 8786 7141 8954 7142
rect 9194 7141 9232 7229
rect 9493 7227 9540 7229
rect 9840 7205 9880 7229
rect 8786 7118 9232 7141
rect 9458 7172 9569 7186
rect 9458 7170 9500 7172
rect 9458 7150 9465 7170
rect 9484 7150 9500 7170
rect 9458 7142 9500 7150
rect 9528 7170 9569 7172
rect 9528 7150 9542 7170
rect 9561 7150 9569 7170
rect 9841 7161 9880 7205
rect 9528 7142 9569 7150
rect 9458 7136 9569 7142
rect 8786 7115 9230 7118
rect 8786 7113 8954 7115
rect 8515 7067 8519 7072
rect 8476 7064 8519 7067
rect 8409 7050 8519 7064
rect 7138 7030 7306 7031
rect 6523 7022 6564 7030
rect 6523 7002 6531 7022
rect 6550 7002 6564 7022
rect 6523 7000 6564 7002
rect 6592 7022 6634 7030
rect 7187 7029 7295 7030
rect 6592 7002 6608 7022
rect 6627 7002 6634 7022
rect 6592 7000 6634 7002
rect 5971 6996 6007 6997
rect 5819 6966 5828 6986
rect 5848 6966 5856 6986
rect 5707 6957 5763 6959
rect 5707 6956 5744 6957
rect 5819 6956 5856 6966
rect 5915 6986 6063 6996
rect 6163 6993 6259 6995
rect 5915 6966 5924 6986
rect 5944 6966 6034 6986
rect 6054 6966 6063 6986
rect 5915 6957 6063 6966
rect 6121 6986 6259 6993
rect 6121 6966 6130 6986
rect 6150 6966 6259 6986
rect 6523 6985 6634 7000
rect 7225 7028 7295 7029
rect 6121 6957 6259 6966
rect 5915 6956 5952 6957
rect 5971 6905 6007 6957
rect 6026 6956 6063 6957
rect 6122 6956 6159 6957
rect 5442 6903 5483 6904
rect 5334 6896 5483 6903
rect 4457 6894 4494 6895
rect 4407 6885 4494 6894
rect 4407 6865 4465 6885
rect 4485 6865 4494 6885
rect 4407 6855 4494 6865
rect 4553 6885 4590 6895
rect 4553 6865 4561 6885
rect 4581 6865 4590 6885
rect 5334 6876 5452 6896
rect 5472 6876 5483 6896
rect 5334 6868 5483 6876
rect 5550 6900 5909 6904
rect 5550 6895 5872 6900
rect 5550 6871 5663 6895
rect 5687 6876 5872 6895
rect 5896 6876 5909 6900
rect 5687 6871 5909 6876
rect 5550 6868 5909 6871
rect 5971 6868 6006 6905
rect 6074 6902 6174 6905
rect 6074 6898 6141 6902
rect 6074 6872 6086 6898
rect 6112 6876 6141 6898
rect 6167 6876 6174 6902
rect 6112 6872 6174 6876
rect 6074 6868 6174 6872
rect 4407 6854 4438 6855
rect 4402 6786 4512 6799
rect 4553 6786 4590 6865
rect 4787 6850 4824 6851
rect 4783 6841 4824 6850
rect 5550 6847 5581 6868
rect 5971 6847 6007 6868
rect 5393 6846 5430 6847
rect 5167 6843 5201 6844
rect 4783 6823 4796 6841
rect 4814 6823 4824 6841
rect 4783 6814 4824 6823
rect 5166 6834 5203 6843
rect 5166 6816 5175 6834
rect 5193 6816 5203 6834
rect 4783 6794 4823 6814
rect 5166 6806 5203 6816
rect 5392 6837 5430 6846
rect 5392 6817 5401 6837
rect 5421 6817 5430 6837
rect 5392 6809 5430 6817
rect 5496 6841 5581 6847
rect 5606 6846 5643 6847
rect 5496 6821 5504 6841
rect 5524 6821 5581 6841
rect 5496 6813 5581 6821
rect 5605 6837 5643 6846
rect 5605 6817 5614 6837
rect 5634 6817 5643 6837
rect 5496 6812 5532 6813
rect 5605 6809 5643 6817
rect 5709 6841 5794 6847
rect 5814 6846 5851 6847
rect 5709 6821 5717 6841
rect 5737 6840 5794 6841
rect 5737 6821 5766 6840
rect 5709 6820 5766 6821
rect 5787 6820 5794 6840
rect 5709 6813 5794 6820
rect 5813 6837 5851 6846
rect 5813 6817 5822 6837
rect 5842 6817 5851 6837
rect 5709 6812 5745 6813
rect 5813 6809 5851 6817
rect 5917 6841 6061 6847
rect 5917 6821 5925 6841
rect 5945 6840 6033 6841
rect 5945 6821 5976 6840
rect 5917 6820 5976 6821
rect 6001 6821 6033 6840
rect 6053 6821 6061 6841
rect 6001 6820 6061 6821
rect 5917 6813 6061 6820
rect 5917 6812 5953 6813
rect 6025 6812 6061 6813
rect 6127 6846 6164 6847
rect 6127 6845 6165 6846
rect 6127 6837 6191 6845
rect 6127 6817 6136 6837
rect 6156 6823 6191 6837
rect 6211 6823 6214 6843
rect 6156 6818 6214 6823
rect 6156 6817 6191 6818
rect 4340 6784 4590 6786
rect 4340 6781 4441 6784
rect 2858 6724 2922 6736
rect 3198 6732 3235 6759
rect 3406 6732 3443 6763
rect 3619 6761 3655 6763
rect 4340 6762 4405 6781
rect 3619 6732 3656 6761
rect 4402 6754 4405 6762
rect 4434 6754 4441 6781
rect 4469 6757 4479 6784
rect 4508 6762 4590 6784
rect 4698 6784 4823 6794
rect 4698 6765 4706 6784
rect 4731 6765 4823 6784
rect 4508 6757 4512 6762
rect 4698 6758 4823 6765
rect 4469 6754 4512 6757
rect 4402 6740 4512 6754
rect 2858 6723 2893 6724
rect 2835 6718 2893 6723
rect 2835 6698 2838 6718
rect 2858 6704 2893 6718
rect 2913 6704 2922 6724
rect 2858 6696 2922 6704
rect 2884 6695 2922 6696
rect 2885 6694 2922 6695
rect 2988 6728 3024 6729
rect 3096 6728 3132 6729
rect 2988 6720 3132 6728
rect 2988 6700 2996 6720
rect 3016 6700 3104 6720
rect 3124 6700 3132 6720
rect 2988 6694 3132 6700
rect 3198 6724 3236 6732
rect 3304 6728 3340 6729
rect 3198 6704 3207 6724
rect 3227 6704 3236 6724
rect 3198 6695 3236 6704
rect 3255 6721 3340 6728
rect 3255 6701 3262 6721
rect 3283 6720 3340 6721
rect 3283 6701 3312 6720
rect 3255 6700 3312 6701
rect 3332 6700 3340 6720
rect 3198 6694 3235 6695
rect 3255 6694 3340 6700
rect 3406 6724 3444 6732
rect 3517 6728 3553 6729
rect 3406 6704 3415 6724
rect 3435 6704 3444 6724
rect 3406 6695 3444 6704
rect 3468 6720 3553 6728
rect 3468 6700 3525 6720
rect 3545 6700 3553 6720
rect 3406 6694 3443 6695
rect 3468 6694 3553 6700
rect 3619 6724 3657 6732
rect 3619 6704 3628 6724
rect 3648 6704 3657 6724
rect 3619 6695 3657 6704
rect 4783 6710 4823 6758
rect 5167 6778 5201 6806
rect 5393 6780 5430 6809
rect 5394 6778 5430 6780
rect 5606 6778 5643 6809
rect 5167 6777 5339 6778
rect 5167 6745 5353 6777
rect 5394 6756 5643 6778
rect 5814 6777 5851 6809
rect 6127 6805 6191 6817
rect 6231 6779 6258 6957
rect 7225 6921 7286 7028
rect 8786 6935 8813 7113
rect 8853 7075 8917 7087
rect 9193 7083 9230 7115
rect 9401 7114 9650 7136
rect 9401 7083 9438 7114
rect 9614 7112 9650 7114
rect 9614 7083 9651 7112
rect 8853 7074 8888 7075
rect 8830 7069 8888 7074
rect 8830 7049 8833 7069
rect 8853 7055 8888 7069
rect 8908 7055 8917 7075
rect 8853 7047 8917 7055
rect 8879 7046 8917 7047
rect 8880 7045 8917 7046
rect 8983 7079 9019 7080
rect 9091 7079 9127 7080
rect 8983 7074 9127 7079
rect 8983 7071 9045 7074
rect 8983 7051 8991 7071
rect 9011 7054 9045 7071
rect 9068 7071 9127 7074
rect 9068 7054 9099 7071
rect 9011 7051 9099 7054
rect 9119 7051 9127 7071
rect 8983 7045 9127 7051
rect 9193 7075 9231 7083
rect 9299 7079 9335 7080
rect 9193 7055 9202 7075
rect 9222 7055 9231 7075
rect 9193 7046 9231 7055
rect 9250 7072 9335 7079
rect 9250 7052 9257 7072
rect 9278 7071 9335 7072
rect 9278 7052 9307 7071
rect 9250 7051 9307 7052
rect 9327 7051 9335 7071
rect 9193 7045 9230 7046
rect 9250 7045 9335 7051
rect 9401 7075 9439 7083
rect 9512 7079 9548 7080
rect 9401 7055 9410 7075
rect 9430 7055 9439 7075
rect 9401 7046 9439 7055
rect 9463 7071 9548 7079
rect 9463 7051 9520 7071
rect 9540 7051 9548 7071
rect 9401 7045 9438 7046
rect 9463 7045 9548 7051
rect 9614 7075 9652 7083
rect 9614 7055 9623 7075
rect 9643 7055 9652 7075
rect 9614 7046 9652 7055
rect 9614 7045 9651 7046
rect 9037 7024 9073 7045
rect 9463 7024 9494 7045
rect 8870 7020 8970 7024
rect 8870 7016 8932 7020
rect 8870 6990 8877 7016
rect 8903 6994 8932 7016
rect 8958 6994 8970 7020
rect 8903 6990 8970 6994
rect 8870 6987 8970 6990
rect 9038 6987 9073 7024
rect 9135 7021 9494 7024
rect 9135 7016 9357 7021
rect 9135 6992 9148 7016
rect 9172 6997 9357 7016
rect 9381 6997 9494 7021
rect 9172 6992 9494 6997
rect 9135 6988 9494 6992
rect 9561 7016 9710 7024
rect 9561 6996 9572 7016
rect 9592 6996 9710 7016
rect 9561 6989 9710 6996
rect 9561 6988 9602 6989
rect 8885 6935 8922 6936
rect 8981 6935 9018 6936
rect 9037 6935 9073 6987
rect 9092 6935 9129 6936
rect 8785 6926 8923 6935
rect 7225 6910 7295 6921
rect 7225 6901 7232 6910
rect 7227 6881 7232 6901
rect 7280 6881 7295 6910
rect 8785 6906 8894 6926
rect 8914 6906 8923 6926
rect 8785 6899 8923 6906
rect 8981 6926 9129 6935
rect 8981 6906 8990 6926
rect 9010 6906 9100 6926
rect 9120 6906 9129 6926
rect 8785 6897 8881 6899
rect 8981 6896 9129 6906
rect 9188 6926 9225 6936
rect 9300 6935 9337 6936
rect 9281 6933 9337 6935
rect 9188 6906 9196 6926
rect 9216 6906 9225 6926
rect 9037 6895 9073 6896
rect 7227 6872 7295 6881
rect 6414 6853 6524 6867
rect 6414 6850 6457 6853
rect 6414 6845 6418 6850
rect 6090 6777 6258 6779
rect 5814 6771 6258 6777
rect 5167 6713 5201 6745
rect 3619 6694 3656 6695
rect 3042 6673 3078 6694
rect 3468 6673 3499 6694
rect 4783 6692 4794 6710
rect 4812 6692 4823 6710
rect 4783 6684 4823 6692
rect 5163 6704 5201 6713
rect 5163 6686 5173 6704
rect 5191 6686 5201 6704
rect 4784 6683 4821 6684
rect 5163 6680 5201 6686
rect 5319 6682 5353 6745
rect 5475 6750 5586 6756
rect 5475 6742 5516 6750
rect 5475 6722 5483 6742
rect 5502 6722 5516 6742
rect 5475 6720 5516 6722
rect 5544 6742 5586 6750
rect 5544 6722 5560 6742
rect 5579 6722 5586 6742
rect 5544 6720 5586 6722
rect 5475 6705 5586 6720
rect 5813 6751 6258 6771
rect 5813 6682 5851 6751
rect 6090 6750 6258 6751
rect 6336 6823 6418 6845
rect 6447 6823 6457 6850
rect 6485 6826 6492 6853
rect 6521 6845 6524 6853
rect 8519 6862 8630 6877
rect 8519 6860 8561 6862
rect 6521 6826 6586 6845
rect 6485 6823 6586 6826
rect 6336 6821 6586 6823
rect 6336 6742 6373 6821
rect 6414 6808 6524 6821
rect 6488 6752 6519 6753
rect 6336 6722 6345 6742
rect 6365 6722 6373 6742
rect 6336 6712 6373 6722
rect 6432 6742 6519 6752
rect 6432 6722 6441 6742
rect 6461 6722 6519 6742
rect 6432 6713 6519 6722
rect 6432 6712 6469 6713
rect 5163 6676 5200 6680
rect 2875 6669 2975 6673
rect 2875 6665 2937 6669
rect 2875 6639 2882 6665
rect 2908 6643 2937 6665
rect 2963 6643 2975 6669
rect 2908 6639 2975 6643
rect 2875 6636 2975 6639
rect 3043 6636 3078 6673
rect 3140 6670 3499 6673
rect 3140 6665 3362 6670
rect 3140 6641 3153 6665
rect 3177 6646 3362 6665
rect 3386 6646 3499 6670
rect 3177 6641 3499 6646
rect 3140 6637 3499 6641
rect 3566 6665 3715 6673
rect 5319 6671 5851 6682
rect 3566 6645 3577 6665
rect 3597 6645 3715 6665
rect 5318 6655 5851 6671
rect 6488 6660 6519 6713
rect 6549 6742 6586 6821
rect 6757 6818 7150 6838
rect 7170 6818 7173 6838
rect 8252 6833 8293 6842
rect 6757 6813 7173 6818
rect 7847 6831 8015 6832
rect 8252 6831 8261 6833
rect 6757 6812 7098 6813
rect 6701 6752 6732 6753
rect 6549 6722 6558 6742
rect 6578 6722 6586 6742
rect 6549 6712 6586 6722
rect 6645 6745 6732 6752
rect 6645 6742 6706 6745
rect 6645 6722 6654 6742
rect 6674 6725 6706 6742
rect 6727 6725 6732 6745
rect 6674 6722 6732 6725
rect 6645 6715 6732 6722
rect 6757 6742 6794 6812
rect 7060 6811 7097 6812
rect 7847 6811 8261 6831
rect 8287 6811 8293 6833
rect 8519 6840 8526 6860
rect 8545 6840 8561 6860
rect 8519 6832 8561 6840
rect 8589 6860 8630 6862
rect 8589 6840 8603 6860
rect 8622 6840 8630 6860
rect 8589 6832 8630 6840
rect 8885 6836 8922 6837
rect 9188 6836 9225 6906
rect 9250 6926 9337 6933
rect 9250 6923 9308 6926
rect 9250 6903 9255 6923
rect 9276 6906 9308 6923
rect 9328 6906 9337 6926
rect 9276 6903 9337 6906
rect 9250 6896 9337 6903
rect 9396 6926 9433 6936
rect 9396 6906 9404 6926
rect 9424 6906 9433 6926
rect 9250 6895 9281 6896
rect 8884 6835 9225 6836
rect 8519 6826 8630 6832
rect 8809 6830 9225 6835
rect 7847 6805 8293 6811
rect 7847 6803 8015 6805
rect 6909 6752 6945 6753
rect 6757 6722 6766 6742
rect 6786 6722 6794 6742
rect 6645 6713 6701 6715
rect 6645 6712 6682 6713
rect 6757 6712 6794 6722
rect 6853 6742 7001 6752
rect 7101 6749 7197 6751
rect 6853 6722 6862 6742
rect 6882 6722 6972 6742
rect 6992 6722 7001 6742
rect 6853 6713 7001 6722
rect 7059 6742 7197 6749
rect 7059 6722 7068 6742
rect 7088 6722 7197 6742
rect 7059 6713 7197 6722
rect 6853 6712 6890 6713
rect 6909 6661 6945 6713
rect 6964 6712 7001 6713
rect 7060 6712 7097 6713
rect 6380 6659 6421 6660
rect 5318 6654 5832 6655
rect 3566 6638 3715 6645
rect 6272 6652 6421 6659
rect 4155 6642 4669 6643
rect 3566 6637 3607 6638
rect 3042 6601 3078 6636
rect 2890 6584 2927 6585
rect 2986 6584 3023 6585
rect 3042 6584 3049 6601
rect 2790 6575 2928 6584
rect 2790 6555 2899 6575
rect 2919 6555 2928 6575
rect 2790 6548 2928 6555
rect 2986 6575 3049 6584
rect 2986 6555 2995 6575
rect 3015 6560 3049 6575
rect 3070 6584 3078 6601
rect 3097 6584 3134 6585
rect 3070 6575 3134 6584
rect 3070 6560 3105 6575
rect 3015 6555 3105 6560
rect 3125 6555 3134 6575
rect 2790 6546 2886 6548
rect 2986 6545 3134 6555
rect 3193 6575 3230 6585
rect 3305 6584 3342 6585
rect 3286 6582 3342 6584
rect 3193 6555 3201 6575
rect 3221 6555 3230 6575
rect 3042 6544 3078 6545
rect 1972 6492 2140 6494
rect 1694 6486 2140 6492
rect 762 6462 1178 6467
rect 1357 6465 1468 6471
rect 762 6461 1103 6462
rect 706 6401 737 6402
rect 554 6371 563 6391
rect 583 6371 591 6391
rect 554 6361 591 6371
rect 650 6394 737 6401
rect 650 6391 711 6394
rect 650 6371 659 6391
rect 679 6374 711 6391
rect 732 6374 737 6394
rect 679 6371 737 6374
rect 650 6364 737 6371
rect 762 6391 799 6461
rect 1065 6460 1102 6461
rect 1357 6457 1398 6465
rect 1357 6437 1365 6457
rect 1384 6437 1398 6457
rect 1357 6435 1398 6437
rect 1426 6457 1468 6465
rect 1426 6437 1442 6457
rect 1461 6437 1468 6457
rect 1694 6464 1700 6486
rect 1726 6466 2140 6486
rect 2890 6485 2927 6486
rect 3193 6485 3230 6555
rect 3255 6575 3342 6582
rect 3255 6572 3313 6575
rect 3255 6552 3260 6572
rect 3281 6555 3313 6572
rect 3333 6555 3342 6575
rect 3281 6552 3342 6555
rect 3255 6545 3342 6552
rect 3401 6575 3438 6585
rect 3401 6555 3409 6575
rect 3429 6555 3438 6575
rect 3255 6544 3286 6545
rect 2889 6484 3230 6485
rect 1726 6464 1735 6466
rect 1972 6465 2140 6466
rect 2814 6483 3230 6484
rect 2814 6479 3190 6483
rect 1694 6455 1735 6464
rect 2814 6459 2817 6479
rect 2837 6466 3190 6479
rect 3222 6466 3230 6483
rect 2837 6459 3230 6466
rect 3401 6476 3438 6555
rect 3468 6584 3499 6637
rect 4136 6626 4669 6642
rect 6272 6632 6390 6652
rect 6410 6632 6421 6652
rect 4136 6615 4668 6626
rect 6272 6624 6421 6632
rect 6488 6656 6847 6660
rect 6488 6651 6810 6656
rect 6488 6627 6601 6651
rect 6625 6632 6810 6651
rect 6834 6632 6847 6656
rect 6625 6627 6847 6632
rect 6488 6624 6847 6627
rect 6909 6624 6944 6661
rect 7012 6658 7112 6661
rect 7012 6654 7079 6658
rect 7012 6628 7024 6654
rect 7050 6632 7079 6654
rect 7105 6632 7112 6658
rect 7050 6628 7112 6632
rect 7012 6624 7112 6628
rect 4787 6617 4824 6621
rect 3518 6584 3555 6585
rect 3468 6575 3555 6584
rect 3468 6555 3526 6575
rect 3546 6555 3555 6575
rect 3468 6545 3555 6555
rect 3614 6575 3651 6585
rect 3614 6555 3622 6575
rect 3642 6555 3651 6575
rect 3468 6544 3499 6545
rect 3463 6476 3573 6489
rect 3614 6476 3651 6555
rect 3401 6474 3651 6476
rect 3401 6471 3502 6474
rect 3401 6452 3466 6471
rect 1426 6435 1468 6437
rect 1357 6420 1468 6435
rect 3463 6444 3466 6452
rect 3495 6444 3502 6471
rect 3530 6447 3540 6474
rect 3569 6452 3651 6474
rect 3729 6546 3897 6547
rect 4136 6546 4174 6615
rect 3729 6526 4174 6546
rect 4401 6577 4512 6592
rect 4401 6575 4443 6577
rect 4401 6555 4408 6575
rect 4427 6555 4443 6575
rect 4401 6547 4443 6555
rect 4471 6575 4512 6577
rect 4471 6555 4485 6575
rect 4504 6555 4512 6575
rect 4471 6547 4512 6555
rect 4401 6541 4512 6547
rect 4634 6552 4668 6615
rect 4786 6611 4824 6617
rect 5166 6613 5203 6614
rect 4786 6593 4796 6611
rect 4814 6593 4824 6611
rect 4786 6584 4824 6593
rect 5164 6605 5204 6613
rect 5164 6587 5175 6605
rect 5193 6587 5204 6605
rect 6488 6603 6519 6624
rect 6909 6603 6945 6624
rect 6331 6602 6368 6603
rect 4786 6552 4820 6584
rect 3729 6520 4173 6526
rect 3729 6518 3897 6520
rect 3569 6447 3573 6452
rect 3530 6444 3573 6447
rect 3463 6430 3573 6444
rect 914 6401 950 6402
rect 762 6371 771 6391
rect 791 6371 799 6391
rect 650 6362 706 6364
rect 650 6361 687 6362
rect 762 6361 799 6371
rect 858 6391 1006 6401
rect 1106 6398 1202 6400
rect 858 6371 867 6391
rect 887 6371 977 6391
rect 997 6371 1006 6391
rect 858 6362 1006 6371
rect 1064 6391 1202 6398
rect 1064 6371 1073 6391
rect 1093 6371 1202 6391
rect 1064 6362 1202 6371
rect 858 6361 895 6362
rect 914 6310 950 6362
rect 969 6361 1006 6362
rect 1065 6361 1102 6362
rect 385 6308 426 6309
rect 277 6301 426 6308
rect 277 6281 395 6301
rect 415 6281 426 6301
rect 277 6273 426 6281
rect 493 6305 852 6309
rect 493 6300 815 6305
rect 493 6276 606 6300
rect 630 6281 815 6300
rect 839 6281 852 6305
rect 630 6276 852 6281
rect 493 6273 852 6276
rect 914 6273 949 6310
rect 1017 6307 1117 6310
rect 1017 6303 1084 6307
rect 1017 6277 1029 6303
rect 1055 6281 1084 6303
rect 1110 6281 1117 6307
rect 1055 6277 1117 6281
rect 1017 6273 1117 6277
rect 493 6252 524 6273
rect 914 6252 950 6273
rect 336 6251 373 6252
rect 335 6242 373 6251
rect 335 6222 344 6242
rect 364 6222 373 6242
rect 335 6214 373 6222
rect 439 6246 524 6252
rect 549 6251 586 6252
rect 439 6226 447 6246
rect 467 6226 524 6246
rect 439 6218 524 6226
rect 548 6242 586 6251
rect 548 6222 557 6242
rect 577 6222 586 6242
rect 439 6217 475 6218
rect 548 6214 586 6222
rect 652 6246 737 6252
rect 757 6251 794 6252
rect 652 6226 660 6246
rect 680 6245 737 6246
rect 680 6226 709 6245
rect 652 6225 709 6226
rect 730 6225 737 6245
rect 652 6218 737 6225
rect 756 6242 794 6251
rect 756 6222 765 6242
rect 785 6222 794 6242
rect 652 6217 688 6218
rect 756 6214 794 6222
rect 860 6246 1004 6252
rect 860 6226 868 6246
rect 888 6243 976 6246
rect 888 6226 919 6243
rect 860 6223 919 6226
rect 942 6226 976 6243
rect 996 6226 1004 6246
rect 942 6223 1004 6226
rect 860 6218 1004 6223
rect 860 6217 896 6218
rect 968 6217 1004 6218
rect 1070 6251 1107 6252
rect 1070 6250 1108 6251
rect 1070 6242 1134 6250
rect 1070 6222 1079 6242
rect 1099 6228 1134 6242
rect 1154 6228 1157 6248
rect 1099 6223 1157 6228
rect 1099 6222 1134 6223
rect 336 6185 373 6214
rect 337 6183 373 6185
rect 549 6183 586 6214
rect 337 6161 586 6183
rect 757 6182 794 6214
rect 1070 6210 1134 6222
rect 1174 6184 1201 6362
rect 3729 6340 3756 6518
rect 3796 6480 3860 6492
rect 4136 6488 4173 6520
rect 4344 6519 4593 6541
rect 4634 6520 4820 6552
rect 4648 6519 4820 6520
rect 4344 6488 4381 6519
rect 4557 6517 4593 6519
rect 4557 6488 4594 6517
rect 4786 6491 4820 6519
rect 5164 6539 5204 6587
rect 6330 6593 6368 6602
rect 6330 6573 6339 6593
rect 6359 6573 6368 6593
rect 6330 6565 6368 6573
rect 6434 6597 6519 6603
rect 6544 6602 6581 6603
rect 6434 6577 6442 6597
rect 6462 6577 6519 6597
rect 6434 6569 6519 6577
rect 6543 6593 6581 6602
rect 6543 6573 6552 6593
rect 6572 6573 6581 6593
rect 6434 6568 6470 6569
rect 6543 6565 6581 6573
rect 6647 6597 6732 6603
rect 6752 6602 6789 6603
rect 6647 6577 6655 6597
rect 6675 6596 6732 6597
rect 6675 6577 6704 6596
rect 6647 6576 6704 6577
rect 6725 6576 6732 6596
rect 6647 6569 6732 6576
rect 6751 6593 6789 6602
rect 6751 6573 6760 6593
rect 6780 6573 6789 6593
rect 6647 6568 6683 6569
rect 6751 6565 6789 6573
rect 6855 6597 6999 6603
rect 6855 6577 6863 6597
rect 6883 6580 6919 6597
rect 6939 6580 6971 6597
rect 6883 6577 6971 6580
rect 6991 6577 6999 6597
rect 6855 6569 6999 6577
rect 6855 6568 6891 6569
rect 6963 6568 6999 6569
rect 7065 6602 7102 6603
rect 7065 6601 7103 6602
rect 7065 6593 7129 6601
rect 7065 6573 7074 6593
rect 7094 6579 7129 6593
rect 7149 6579 7152 6599
rect 7094 6574 7152 6579
rect 7094 6573 7129 6574
rect 5475 6543 5585 6557
rect 5475 6540 5518 6543
rect 5164 6532 5289 6539
rect 5475 6535 5479 6540
rect 5164 6513 5256 6532
rect 5281 6513 5289 6532
rect 5164 6503 5289 6513
rect 5397 6513 5479 6535
rect 5508 6513 5518 6540
rect 5546 6516 5553 6543
rect 5582 6535 5585 6543
rect 6331 6536 6368 6565
rect 5582 6516 5647 6535
rect 6332 6534 6368 6536
rect 6544 6534 6581 6565
rect 6752 6538 6789 6565
rect 7065 6561 7129 6573
rect 5546 6513 5647 6516
rect 5397 6511 5647 6513
rect 3796 6479 3831 6480
rect 3773 6474 3831 6479
rect 3773 6454 3776 6474
rect 3796 6460 3831 6474
rect 3851 6460 3860 6480
rect 3796 6452 3860 6460
rect 3822 6451 3860 6452
rect 3823 6450 3860 6451
rect 3926 6484 3962 6485
rect 4034 6484 4070 6485
rect 3926 6477 4070 6484
rect 3926 6476 3986 6477
rect 3926 6456 3934 6476
rect 3954 6457 3986 6476
rect 4011 6476 4070 6477
rect 4011 6457 4042 6476
rect 3954 6456 4042 6457
rect 4062 6456 4070 6476
rect 3926 6450 4070 6456
rect 4136 6480 4174 6488
rect 4242 6484 4278 6485
rect 4136 6460 4145 6480
rect 4165 6460 4174 6480
rect 4136 6451 4174 6460
rect 4193 6477 4278 6484
rect 4193 6457 4200 6477
rect 4221 6476 4278 6477
rect 4221 6457 4250 6476
rect 4193 6456 4250 6457
rect 4270 6456 4278 6476
rect 4136 6450 4173 6451
rect 4193 6450 4278 6456
rect 4344 6480 4382 6488
rect 4455 6484 4491 6485
rect 4344 6460 4353 6480
rect 4373 6460 4382 6480
rect 4344 6451 4382 6460
rect 4406 6476 4491 6484
rect 4406 6456 4463 6476
rect 4483 6456 4491 6476
rect 4344 6450 4381 6451
rect 4406 6450 4491 6456
rect 4557 6480 4595 6488
rect 4557 6460 4566 6480
rect 4586 6460 4595 6480
rect 4557 6451 4595 6460
rect 4784 6481 4821 6491
rect 5164 6483 5204 6503
rect 4784 6463 4794 6481
rect 4812 6463 4821 6481
rect 4784 6454 4821 6463
rect 5163 6474 5204 6483
rect 5163 6456 5173 6474
rect 5191 6456 5204 6474
rect 4786 6453 4820 6454
rect 4557 6450 4594 6451
rect 3980 6429 4016 6450
rect 4406 6429 4437 6450
rect 5163 6447 5204 6456
rect 5163 6446 5200 6447
rect 5397 6432 5434 6511
rect 5475 6498 5585 6511
rect 5549 6442 5580 6443
rect 3813 6425 3913 6429
rect 3813 6421 3875 6425
rect 3813 6395 3820 6421
rect 3846 6399 3875 6421
rect 3901 6399 3913 6425
rect 3846 6395 3913 6399
rect 3813 6392 3913 6395
rect 3981 6392 4016 6429
rect 4078 6426 4437 6429
rect 4078 6421 4300 6426
rect 4078 6397 4091 6421
rect 4115 6402 4300 6421
rect 4324 6402 4437 6426
rect 4115 6397 4437 6402
rect 4078 6393 4437 6397
rect 4504 6421 4653 6429
rect 4504 6401 4515 6421
rect 4535 6401 4653 6421
rect 5397 6412 5406 6432
rect 5426 6412 5434 6432
rect 5397 6402 5434 6412
rect 5493 6432 5580 6442
rect 5493 6412 5502 6432
rect 5522 6412 5580 6432
rect 5493 6403 5580 6412
rect 5493 6402 5530 6403
rect 4504 6394 4653 6401
rect 4504 6393 4545 6394
rect 3828 6340 3865 6341
rect 3924 6340 3961 6341
rect 3980 6340 4016 6392
rect 4035 6340 4072 6341
rect 3728 6331 3866 6340
rect 3323 6310 3434 6325
rect 3323 6308 3365 6310
rect 2993 6287 3098 6289
rect 2651 6279 2819 6280
rect 2993 6279 3042 6287
rect 2651 6260 3042 6279
rect 3073 6260 3098 6287
rect 3323 6288 3330 6308
rect 3349 6288 3365 6308
rect 3323 6280 3365 6288
rect 3393 6308 3434 6310
rect 3393 6288 3407 6308
rect 3426 6288 3434 6308
rect 3728 6311 3837 6331
rect 3857 6311 3866 6331
rect 3728 6304 3866 6311
rect 3924 6331 4072 6340
rect 3924 6311 3933 6331
rect 3953 6311 4043 6331
rect 4063 6311 4072 6331
rect 3728 6302 3824 6304
rect 3924 6301 4072 6311
rect 4131 6331 4168 6341
rect 4243 6340 4280 6341
rect 4224 6338 4280 6340
rect 4131 6311 4139 6331
rect 4159 6311 4168 6331
rect 3980 6300 4016 6301
rect 3393 6280 3434 6288
rect 3323 6274 3434 6280
rect 2651 6253 3098 6260
rect 2651 6251 2819 6253
rect 1499 6220 1609 6234
rect 1499 6217 1542 6220
rect 1499 6212 1503 6217
rect 1033 6182 1201 6184
rect 757 6179 1201 6182
rect 418 6155 529 6161
rect 418 6147 459 6155
rect 107 6092 146 6136
rect 418 6127 426 6147
rect 445 6127 459 6147
rect 418 6125 459 6127
rect 487 6147 529 6155
rect 487 6127 503 6147
rect 522 6127 529 6147
rect 487 6125 529 6127
rect 418 6110 529 6125
rect 755 6156 1201 6179
rect 107 6068 147 6092
rect 447 6068 494 6070
rect 755 6068 793 6156
rect 1033 6155 1201 6156
rect 1421 6190 1503 6212
rect 1532 6190 1542 6217
rect 1570 6193 1577 6220
rect 1606 6212 1609 6220
rect 1606 6193 1671 6212
rect 1570 6190 1671 6193
rect 1421 6188 1671 6190
rect 1421 6109 1458 6188
rect 1499 6175 1609 6188
rect 1573 6119 1604 6120
rect 1421 6089 1430 6109
rect 1450 6089 1458 6109
rect 1421 6079 1458 6089
rect 1517 6109 1604 6119
rect 1517 6089 1526 6109
rect 1546 6089 1604 6109
rect 1517 6080 1604 6089
rect 1517 6079 1554 6080
rect 107 6035 793 6068
rect 107 5978 146 6035
rect 755 6033 793 6035
rect 1573 6027 1604 6080
rect 1634 6109 1671 6188
rect 1842 6201 2235 6205
rect 1842 6184 1861 6201
rect 1881 6185 2235 6201
rect 2255 6185 2258 6205
rect 1881 6184 2258 6185
rect 1842 6180 2258 6184
rect 1842 6179 2183 6180
rect 1786 6119 1817 6120
rect 1634 6089 1643 6109
rect 1663 6089 1671 6109
rect 1634 6079 1671 6089
rect 1730 6112 1817 6119
rect 1730 6109 1791 6112
rect 1730 6089 1739 6109
rect 1759 6092 1791 6109
rect 1812 6092 1817 6112
rect 1759 6089 1817 6092
rect 1730 6082 1817 6089
rect 1842 6109 1879 6179
rect 2145 6178 2182 6179
rect 1994 6119 2030 6120
rect 1842 6089 1851 6109
rect 1871 6089 1879 6109
rect 1730 6080 1786 6082
rect 1730 6079 1767 6080
rect 1842 6079 1879 6089
rect 1938 6109 2086 6119
rect 2254 6118 2283 6119
rect 2186 6116 2283 6118
rect 1938 6089 1947 6109
rect 1967 6105 2057 6109
rect 1967 6089 2000 6105
rect 1938 6080 2000 6089
rect 1938 6079 1975 6080
rect 1994 6067 2000 6080
rect 2023 6089 2057 6105
rect 2077 6089 2086 6109
rect 2023 6080 2086 6089
rect 2144 6109 2283 6116
rect 2144 6089 2153 6109
rect 2173 6089 2283 6109
rect 2144 6080 2283 6089
rect 2023 6067 2030 6080
rect 2049 6079 2086 6080
rect 2145 6079 2182 6080
rect 1994 6028 2030 6067
rect 1465 6026 1506 6027
rect 1357 6019 1506 6026
rect 1357 5999 1475 6019
rect 1495 5999 1506 6019
rect 1357 5991 1506 5999
rect 1573 6023 1932 6027
rect 1573 6018 1895 6023
rect 1573 5994 1686 6018
rect 1710 5999 1895 6018
rect 1919 5999 1932 6023
rect 1710 5994 1932 5999
rect 1573 5991 1932 5994
rect 1994 5991 2029 6028
rect 2097 6025 2197 6028
rect 2097 6021 2164 6025
rect 2097 5995 2109 6021
rect 2135 5999 2164 6021
rect 2190 5999 2197 6025
rect 2135 5995 2197 5999
rect 2097 5991 2197 5995
rect 107 5976 155 5978
rect 107 5958 118 5976
rect 136 5958 155 5976
rect 1573 5970 1604 5991
rect 1994 5970 2030 5991
rect 1416 5969 1453 5970
rect 107 5949 155 5958
rect 108 5948 155 5949
rect 421 5953 531 5967
rect 421 5950 464 5953
rect 421 5945 425 5950
rect 343 5923 425 5945
rect 454 5923 464 5950
rect 492 5926 499 5953
rect 528 5945 531 5953
rect 1415 5960 1453 5969
rect 528 5926 593 5945
rect 1415 5940 1424 5960
rect 1444 5940 1453 5960
rect 492 5923 593 5926
rect 343 5921 593 5923
rect 111 5885 148 5886
rect 107 5882 148 5885
rect 107 5877 149 5882
rect 107 5859 120 5877
rect 138 5859 149 5877
rect 107 5845 149 5859
rect 187 5845 234 5849
rect 107 5839 234 5845
rect 107 5810 195 5839
rect 224 5810 234 5839
rect 343 5842 380 5921
rect 421 5908 531 5921
rect 495 5852 526 5853
rect 343 5822 352 5842
rect 372 5822 380 5842
rect 343 5812 380 5822
rect 439 5842 526 5852
rect 439 5822 448 5842
rect 468 5822 526 5842
rect 439 5813 526 5822
rect 439 5812 476 5813
rect 107 5806 234 5810
rect 107 5789 146 5806
rect 187 5805 234 5806
rect 107 5771 118 5789
rect 136 5771 146 5789
rect 107 5762 146 5771
rect 108 5761 145 5762
rect 495 5760 526 5813
rect 556 5842 593 5921
rect 764 5918 1157 5938
rect 1177 5918 1180 5938
rect 1415 5932 1453 5940
rect 1519 5964 1604 5970
rect 1629 5969 1666 5970
rect 1519 5944 1527 5964
rect 1547 5944 1604 5964
rect 1519 5936 1604 5944
rect 1628 5960 1666 5969
rect 1628 5940 1637 5960
rect 1657 5940 1666 5960
rect 1519 5935 1555 5936
rect 1628 5932 1666 5940
rect 1732 5964 1817 5970
rect 1837 5969 1874 5970
rect 1732 5944 1740 5964
rect 1760 5963 1817 5964
rect 1760 5944 1789 5963
rect 1732 5943 1789 5944
rect 1810 5943 1817 5963
rect 1732 5936 1817 5943
rect 1836 5960 1874 5969
rect 1836 5940 1845 5960
rect 1865 5940 1874 5960
rect 1732 5935 1768 5936
rect 1836 5932 1874 5940
rect 1940 5964 2084 5970
rect 1940 5944 1948 5964
rect 1968 5944 2056 5964
rect 2076 5944 2084 5964
rect 1940 5936 2084 5944
rect 1940 5935 1976 5936
rect 2048 5935 2084 5936
rect 2150 5969 2187 5970
rect 2150 5968 2188 5969
rect 2150 5960 2214 5968
rect 2150 5940 2159 5960
rect 2179 5946 2214 5960
rect 2234 5946 2237 5966
rect 2179 5941 2237 5946
rect 2179 5940 2214 5941
rect 764 5913 1180 5918
rect 764 5912 1105 5913
rect 708 5852 739 5853
rect 556 5822 565 5842
rect 585 5822 593 5842
rect 556 5812 593 5822
rect 652 5845 739 5852
rect 652 5842 713 5845
rect 652 5822 661 5842
rect 681 5825 713 5842
rect 734 5825 739 5845
rect 681 5822 739 5825
rect 652 5815 739 5822
rect 764 5842 801 5912
rect 1067 5911 1104 5912
rect 1416 5903 1453 5932
rect 1417 5901 1453 5903
rect 1629 5901 1666 5932
rect 1417 5879 1666 5901
rect 1837 5900 1874 5932
rect 2150 5928 2214 5940
rect 2254 5902 2283 6080
rect 2651 6073 2678 6251
rect 2718 6213 2782 6225
rect 3058 6221 3095 6253
rect 3266 6252 3515 6274
rect 3266 6221 3303 6252
rect 3479 6250 3515 6252
rect 3479 6221 3516 6250
rect 3828 6241 3865 6242
rect 4131 6241 4168 6311
rect 4193 6331 4280 6338
rect 4193 6328 4251 6331
rect 4193 6308 4198 6328
rect 4219 6311 4251 6328
rect 4271 6311 4280 6331
rect 4219 6308 4280 6311
rect 4193 6301 4280 6308
rect 4339 6331 4376 6341
rect 4339 6311 4347 6331
rect 4367 6311 4376 6331
rect 4193 6300 4224 6301
rect 3827 6240 4168 6241
rect 3752 6235 4168 6240
rect 2718 6212 2753 6213
rect 2695 6207 2753 6212
rect 2695 6187 2698 6207
rect 2718 6193 2753 6207
rect 2773 6193 2782 6213
rect 2718 6185 2782 6193
rect 2744 6184 2782 6185
rect 2745 6183 2782 6184
rect 2848 6217 2884 6218
rect 2956 6217 2992 6218
rect 2848 6212 2992 6217
rect 2848 6209 2908 6212
rect 2848 6189 2856 6209
rect 2876 6191 2908 6209
rect 2935 6209 2992 6212
rect 2935 6191 2964 6209
rect 2876 6189 2964 6191
rect 2984 6189 2992 6209
rect 2848 6183 2992 6189
rect 3058 6213 3096 6221
rect 3164 6217 3200 6218
rect 3058 6193 3067 6213
rect 3087 6193 3096 6213
rect 3058 6184 3096 6193
rect 3115 6210 3200 6217
rect 3115 6190 3122 6210
rect 3143 6209 3200 6210
rect 3143 6190 3172 6209
rect 3115 6189 3172 6190
rect 3192 6189 3200 6209
rect 3058 6183 3095 6184
rect 3115 6183 3200 6189
rect 3266 6213 3304 6221
rect 3377 6217 3413 6218
rect 3266 6193 3275 6213
rect 3295 6193 3304 6213
rect 3266 6184 3304 6193
rect 3328 6209 3413 6217
rect 3328 6189 3385 6209
rect 3405 6189 3413 6209
rect 3266 6183 3303 6184
rect 3328 6183 3413 6189
rect 3479 6213 3517 6221
rect 3752 6215 3755 6235
rect 3775 6215 4168 6235
rect 4339 6232 4376 6311
rect 4406 6340 4437 6393
rect 4787 6391 4824 6392
rect 4786 6382 4825 6391
rect 4786 6364 4796 6382
rect 4814 6364 4825 6382
rect 5166 6380 5203 6384
rect 4698 6347 4745 6348
rect 4786 6347 4825 6364
rect 4698 6343 4825 6347
rect 4456 6340 4493 6341
rect 4406 6331 4493 6340
rect 4406 6311 4464 6331
rect 4484 6311 4493 6331
rect 4406 6301 4493 6311
rect 4552 6331 4589 6341
rect 4552 6311 4560 6331
rect 4580 6311 4589 6331
rect 4406 6300 4437 6301
rect 4401 6232 4511 6245
rect 4552 6232 4589 6311
rect 4698 6314 4708 6343
rect 4737 6314 4825 6343
rect 4698 6308 4825 6314
rect 4698 6304 4745 6308
rect 4783 6294 4825 6308
rect 4783 6276 4794 6294
rect 4812 6276 4825 6294
rect 4783 6271 4825 6276
rect 4784 6268 4825 6271
rect 5163 6375 5203 6380
rect 5163 6357 5175 6375
rect 5193 6357 5203 6375
rect 4784 6267 4821 6268
rect 4339 6230 4589 6232
rect 4339 6227 4440 6230
rect 3479 6193 3488 6213
rect 3508 6193 3517 6213
rect 4339 6208 4404 6227
rect 3479 6184 3517 6193
rect 4401 6200 4404 6208
rect 4433 6200 4440 6227
rect 4468 6203 4478 6230
rect 4507 6208 4589 6230
rect 4507 6203 4511 6208
rect 4468 6200 4511 6203
rect 4401 6186 4511 6200
rect 4777 6204 4824 6205
rect 4777 6195 4825 6204
rect 3479 6183 3516 6184
rect 2902 6162 2938 6183
rect 3328 6162 3359 6183
rect 4777 6177 4796 6195
rect 4814 6177 4825 6195
rect 4777 6175 4825 6177
rect 2735 6158 2835 6162
rect 2735 6154 2797 6158
rect 2735 6128 2742 6154
rect 2768 6132 2797 6154
rect 2823 6132 2835 6158
rect 2768 6128 2835 6132
rect 2735 6125 2835 6128
rect 2903 6125 2938 6162
rect 3000 6159 3359 6162
rect 3000 6154 3222 6159
rect 3000 6130 3013 6154
rect 3037 6135 3222 6154
rect 3246 6135 3359 6159
rect 3037 6130 3359 6135
rect 3000 6126 3359 6130
rect 3426 6154 3575 6162
rect 3426 6134 3437 6154
rect 3457 6134 3575 6154
rect 3426 6127 3575 6134
rect 3426 6126 3467 6127
rect 2750 6073 2787 6074
rect 2846 6073 2883 6074
rect 2902 6073 2938 6125
rect 2957 6073 2994 6074
rect 2650 6064 2788 6073
rect 2650 6044 2759 6064
rect 2779 6044 2788 6064
rect 2650 6037 2788 6044
rect 2846 6064 2994 6073
rect 2846 6044 2855 6064
rect 2875 6044 2965 6064
rect 2985 6044 2994 6064
rect 2650 6035 2746 6037
rect 2846 6034 2994 6044
rect 3053 6064 3090 6074
rect 3165 6073 3202 6074
rect 3146 6071 3202 6073
rect 3053 6044 3061 6064
rect 3081 6044 3090 6064
rect 2902 6033 2938 6034
rect 2750 5974 2787 5975
rect 3053 5974 3090 6044
rect 3115 6064 3202 6071
rect 3115 6061 3173 6064
rect 3115 6041 3120 6061
rect 3141 6044 3173 6061
rect 3193 6044 3202 6064
rect 3141 6041 3202 6044
rect 3115 6034 3202 6041
rect 3261 6064 3298 6074
rect 3261 6044 3269 6064
rect 3289 6044 3298 6064
rect 3115 6033 3146 6034
rect 2749 5973 3090 5974
rect 2674 5969 3090 5973
rect 2674 5968 3051 5969
rect 2674 5948 2677 5968
rect 2697 5952 3051 5968
rect 3071 5952 3090 5969
rect 2697 5948 3090 5952
rect 3261 5965 3298 6044
rect 3328 6073 3359 6126
rect 4139 6118 4177 6120
rect 4786 6118 4825 6175
rect 4139 6085 4825 6118
rect 3378 6073 3415 6074
rect 3328 6064 3415 6073
rect 3328 6044 3386 6064
rect 3406 6044 3415 6064
rect 3328 6034 3415 6044
rect 3474 6064 3511 6074
rect 3474 6044 3482 6064
rect 3502 6044 3511 6064
rect 3328 6033 3359 6034
rect 3323 5965 3433 5978
rect 3474 5965 3511 6044
rect 3261 5963 3511 5965
rect 3261 5960 3362 5963
rect 3261 5941 3326 5960
rect 3323 5933 3326 5941
rect 3355 5933 3362 5960
rect 3390 5936 3400 5963
rect 3429 5941 3511 5963
rect 3731 5997 3899 5998
rect 4139 5997 4177 6085
rect 4438 6083 4485 6085
rect 4785 6061 4825 6085
rect 3731 5974 4177 5997
rect 4403 6028 4514 6043
rect 4403 6026 4445 6028
rect 4403 6006 4410 6026
rect 4429 6006 4445 6026
rect 4403 5998 4445 6006
rect 4473 6026 4514 6028
rect 4473 6006 4487 6026
rect 4506 6006 4514 6026
rect 4786 6017 4825 6061
rect 4473 5998 4514 6006
rect 4403 5992 4514 5998
rect 3731 5971 4175 5974
rect 3731 5969 3899 5971
rect 3429 5936 3433 5941
rect 3390 5933 3433 5936
rect 3323 5919 3433 5933
rect 2113 5900 2283 5902
rect 1834 5893 2283 5900
rect 1498 5873 1609 5879
rect 1498 5865 1539 5873
rect 916 5852 952 5853
rect 764 5822 773 5842
rect 793 5822 801 5842
rect 652 5813 708 5815
rect 652 5812 689 5813
rect 764 5812 801 5822
rect 860 5842 1008 5852
rect 1108 5849 1204 5851
rect 860 5822 869 5842
rect 889 5822 979 5842
rect 999 5822 1008 5842
rect 860 5813 1008 5822
rect 1066 5842 1204 5849
rect 1066 5822 1075 5842
rect 1095 5822 1204 5842
rect 1498 5845 1506 5865
rect 1525 5845 1539 5865
rect 1498 5843 1539 5845
rect 1567 5865 1609 5873
rect 1567 5845 1583 5865
rect 1602 5845 1609 5865
rect 1834 5866 1859 5893
rect 1890 5874 2283 5893
rect 1890 5866 1939 5874
rect 2113 5873 2283 5874
rect 1834 5864 1939 5866
rect 1567 5843 1609 5845
rect 1498 5828 1609 5843
rect 1066 5813 1204 5822
rect 860 5812 897 5813
rect 916 5761 952 5813
rect 971 5812 1008 5813
rect 1067 5812 1104 5813
rect 387 5759 428 5760
rect 279 5752 428 5759
rect 279 5732 397 5752
rect 417 5732 428 5752
rect 279 5724 428 5732
rect 495 5756 854 5760
rect 495 5751 817 5756
rect 495 5727 608 5751
rect 632 5732 817 5751
rect 841 5732 854 5756
rect 632 5727 854 5732
rect 495 5724 854 5727
rect 916 5724 951 5761
rect 1019 5758 1119 5761
rect 1019 5754 1086 5758
rect 1019 5728 1031 5754
rect 1057 5732 1086 5754
rect 1112 5732 1119 5758
rect 1057 5728 1119 5732
rect 1019 5724 1119 5728
rect 495 5703 526 5724
rect 916 5703 952 5724
rect 338 5702 375 5703
rect 112 5699 146 5700
rect 111 5690 148 5699
rect 111 5672 120 5690
rect 138 5672 148 5690
rect 111 5662 148 5672
rect 337 5693 375 5702
rect 337 5673 346 5693
rect 366 5673 375 5693
rect 337 5665 375 5673
rect 441 5697 526 5703
rect 551 5702 588 5703
rect 441 5677 449 5697
rect 469 5677 526 5697
rect 441 5669 526 5677
rect 550 5693 588 5702
rect 550 5673 559 5693
rect 579 5673 588 5693
rect 441 5668 477 5669
rect 550 5665 588 5673
rect 654 5697 739 5703
rect 759 5702 796 5703
rect 654 5677 662 5697
rect 682 5696 739 5697
rect 682 5677 711 5696
rect 654 5676 711 5677
rect 732 5676 739 5696
rect 654 5669 739 5676
rect 758 5693 796 5702
rect 758 5673 767 5693
rect 787 5673 796 5693
rect 654 5668 690 5669
rect 758 5665 796 5673
rect 862 5697 1006 5703
rect 862 5677 870 5697
rect 890 5696 978 5697
rect 890 5677 921 5696
rect 862 5676 921 5677
rect 946 5677 978 5696
rect 998 5677 1006 5697
rect 946 5676 1006 5677
rect 862 5669 1006 5676
rect 862 5668 898 5669
rect 970 5668 1006 5669
rect 1072 5702 1109 5703
rect 1072 5701 1110 5702
rect 1072 5693 1136 5701
rect 1072 5673 1081 5693
rect 1101 5679 1136 5693
rect 1156 5679 1159 5699
rect 1101 5674 1159 5679
rect 1101 5673 1136 5674
rect 112 5634 146 5662
rect 338 5636 375 5665
rect 339 5634 375 5636
rect 551 5634 588 5665
rect 112 5633 284 5634
rect 112 5601 298 5633
rect 339 5612 588 5634
rect 759 5633 796 5665
rect 1072 5661 1136 5673
rect 1176 5635 1203 5813
rect 3731 5791 3758 5969
rect 3798 5931 3862 5943
rect 4138 5939 4175 5971
rect 4346 5970 4595 5992
rect 4346 5939 4383 5970
rect 4559 5968 4595 5970
rect 4559 5939 4596 5968
rect 3798 5930 3833 5931
rect 3775 5925 3833 5930
rect 3775 5905 3778 5925
rect 3798 5911 3833 5925
rect 3853 5911 3862 5931
rect 3798 5903 3862 5911
rect 3824 5902 3862 5903
rect 3825 5901 3862 5902
rect 3928 5935 3964 5936
rect 4036 5935 4072 5936
rect 3928 5930 4072 5935
rect 3928 5927 3990 5930
rect 3928 5907 3936 5927
rect 3956 5910 3990 5927
rect 4013 5927 4072 5930
rect 4013 5910 4044 5927
rect 3956 5907 4044 5910
rect 4064 5907 4072 5927
rect 3928 5901 4072 5907
rect 4138 5931 4176 5939
rect 4244 5935 4280 5936
rect 4138 5911 4147 5931
rect 4167 5911 4176 5931
rect 4138 5902 4176 5911
rect 4195 5928 4280 5935
rect 4195 5908 4202 5928
rect 4223 5927 4280 5928
rect 4223 5908 4252 5927
rect 4195 5907 4252 5908
rect 4272 5907 4280 5927
rect 4138 5901 4175 5902
rect 4195 5901 4280 5907
rect 4346 5931 4384 5939
rect 4457 5935 4493 5936
rect 4346 5911 4355 5931
rect 4375 5911 4384 5931
rect 4346 5902 4384 5911
rect 4408 5927 4493 5935
rect 4408 5907 4465 5927
rect 4485 5907 4493 5927
rect 4346 5901 4383 5902
rect 4408 5901 4493 5907
rect 4559 5931 4597 5939
rect 4559 5911 4568 5931
rect 4588 5911 4597 5931
rect 4559 5902 4597 5911
rect 4559 5901 4596 5902
rect 3982 5880 4018 5901
rect 4408 5880 4439 5901
rect 3815 5876 3915 5880
rect 3815 5872 3877 5876
rect 3815 5846 3822 5872
rect 3848 5850 3877 5872
rect 3903 5850 3915 5876
rect 3848 5846 3915 5850
rect 3815 5843 3915 5846
rect 3983 5843 4018 5880
rect 4080 5877 4439 5880
rect 4080 5872 4302 5877
rect 4080 5848 4093 5872
rect 4117 5853 4302 5872
rect 4326 5853 4439 5877
rect 4117 5848 4439 5853
rect 4080 5844 4439 5848
rect 4506 5872 4655 5880
rect 4506 5852 4517 5872
rect 4537 5852 4655 5872
rect 4506 5845 4655 5852
rect 4506 5844 4547 5845
rect 3830 5791 3867 5792
rect 3926 5791 3963 5792
rect 3982 5791 4018 5843
rect 4037 5791 4074 5792
rect 3730 5782 3868 5791
rect 3730 5762 3839 5782
rect 3859 5762 3868 5782
rect 3730 5755 3868 5762
rect 3926 5782 4074 5791
rect 3926 5762 3935 5782
rect 3955 5762 4045 5782
rect 4065 5762 4074 5782
rect 3730 5753 3826 5755
rect 3926 5752 4074 5762
rect 4133 5782 4170 5792
rect 4245 5791 4282 5792
rect 4226 5789 4282 5791
rect 4133 5762 4141 5782
rect 4161 5762 4170 5782
rect 3982 5751 4018 5752
rect 1359 5709 1469 5723
rect 1359 5706 1402 5709
rect 1359 5701 1363 5706
rect 1035 5633 1203 5635
rect 759 5627 1203 5633
rect 112 5569 146 5601
rect 108 5560 146 5569
rect 108 5542 118 5560
rect 136 5542 146 5560
rect 108 5536 146 5542
rect 264 5538 298 5601
rect 420 5606 531 5612
rect 420 5598 461 5606
rect 420 5578 428 5598
rect 447 5578 461 5598
rect 420 5576 461 5578
rect 489 5598 531 5606
rect 489 5578 505 5598
rect 524 5578 531 5598
rect 489 5576 531 5578
rect 420 5561 531 5576
rect 758 5607 1203 5627
rect 758 5538 796 5607
rect 1035 5606 1203 5607
rect 1281 5679 1363 5701
rect 1392 5679 1402 5706
rect 1430 5682 1437 5709
rect 1466 5701 1469 5709
rect 3464 5718 3575 5733
rect 3464 5716 3506 5718
rect 1466 5682 1531 5701
rect 1430 5679 1531 5682
rect 1281 5677 1531 5679
rect 1281 5598 1318 5677
rect 1359 5664 1469 5677
rect 1433 5608 1464 5609
rect 1281 5578 1290 5598
rect 1310 5578 1318 5598
rect 1281 5568 1318 5578
rect 1377 5598 1464 5608
rect 1377 5578 1386 5598
rect 1406 5578 1464 5598
rect 1377 5569 1464 5578
rect 1377 5568 1414 5569
rect 108 5532 145 5536
rect 264 5527 796 5538
rect 263 5511 796 5527
rect 1433 5516 1464 5569
rect 1494 5598 1531 5677
rect 1702 5687 2095 5694
rect 1702 5670 1710 5687
rect 1742 5674 2095 5687
rect 2115 5674 2118 5694
rect 3197 5689 3238 5698
rect 1742 5670 2118 5674
rect 1702 5669 2118 5670
rect 2792 5687 2960 5688
rect 3197 5687 3206 5689
rect 1702 5668 2043 5669
rect 1646 5608 1677 5609
rect 1494 5578 1503 5598
rect 1523 5578 1531 5598
rect 1494 5568 1531 5578
rect 1590 5601 1677 5608
rect 1590 5598 1651 5601
rect 1590 5578 1599 5598
rect 1619 5581 1651 5598
rect 1672 5581 1677 5601
rect 1619 5578 1677 5581
rect 1590 5571 1677 5578
rect 1702 5598 1739 5668
rect 2005 5667 2042 5668
rect 2792 5667 3206 5687
rect 3232 5667 3238 5689
rect 3464 5696 3471 5716
rect 3490 5696 3506 5716
rect 3464 5688 3506 5696
rect 3534 5716 3575 5718
rect 3534 5696 3548 5716
rect 3567 5696 3575 5716
rect 3534 5688 3575 5696
rect 3830 5692 3867 5693
rect 4133 5692 4170 5762
rect 4195 5782 4282 5789
rect 4195 5779 4253 5782
rect 4195 5759 4200 5779
rect 4221 5762 4253 5779
rect 4273 5762 4282 5782
rect 4221 5759 4282 5762
rect 4195 5752 4282 5759
rect 4341 5782 4378 5792
rect 4341 5762 4349 5782
rect 4369 5762 4378 5782
rect 4195 5751 4226 5752
rect 3829 5691 4170 5692
rect 3464 5682 3575 5688
rect 3754 5686 4170 5691
rect 2792 5661 3238 5667
rect 2792 5659 2960 5661
rect 1854 5608 1890 5609
rect 1702 5578 1711 5598
rect 1731 5578 1739 5598
rect 1590 5569 1646 5571
rect 1590 5568 1627 5569
rect 1702 5568 1739 5578
rect 1798 5598 1946 5608
rect 2046 5605 2142 5607
rect 1798 5578 1807 5598
rect 1827 5593 1917 5598
rect 1827 5578 1862 5593
rect 1798 5569 1862 5578
rect 1798 5568 1835 5569
rect 1854 5552 1862 5569
rect 1883 5578 1917 5593
rect 1937 5578 1946 5598
rect 1883 5569 1946 5578
rect 2004 5598 2142 5605
rect 2004 5578 2013 5598
rect 2033 5578 2142 5598
rect 2004 5569 2142 5578
rect 1883 5552 1890 5569
rect 1909 5568 1946 5569
rect 2005 5568 2042 5569
rect 1854 5517 1890 5552
rect 1325 5515 1366 5516
rect 263 5510 777 5511
rect 1217 5508 1366 5515
rect 1217 5488 1335 5508
rect 1355 5488 1366 5508
rect 1217 5480 1366 5488
rect 1433 5512 1792 5516
rect 1433 5507 1755 5512
rect 1433 5483 1546 5507
rect 1570 5488 1755 5507
rect 1779 5488 1792 5512
rect 1570 5483 1792 5488
rect 1433 5480 1792 5483
rect 1854 5480 1889 5517
rect 1957 5514 2057 5517
rect 1957 5510 2024 5514
rect 1957 5484 1969 5510
rect 1995 5488 2024 5510
rect 2050 5488 2057 5514
rect 1995 5484 2057 5488
rect 1957 5480 2057 5484
rect 111 5469 148 5470
rect 109 5461 149 5469
rect 109 5443 120 5461
rect 138 5443 149 5461
rect 1433 5459 1464 5480
rect 1854 5459 1890 5480
rect 1276 5458 1313 5459
rect 109 5395 149 5443
rect 1275 5449 1313 5458
rect 1275 5429 1284 5449
rect 1304 5429 1313 5449
rect 1275 5421 1313 5429
rect 1379 5453 1464 5459
rect 1489 5458 1526 5459
rect 1379 5433 1387 5453
rect 1407 5433 1464 5453
rect 1379 5425 1464 5433
rect 1488 5449 1526 5458
rect 1488 5429 1497 5449
rect 1517 5429 1526 5449
rect 1379 5424 1415 5425
rect 1488 5421 1526 5429
rect 1592 5453 1677 5459
rect 1697 5458 1734 5459
rect 1592 5433 1600 5453
rect 1620 5452 1677 5453
rect 1620 5433 1649 5452
rect 1592 5432 1649 5433
rect 1670 5432 1677 5452
rect 1592 5425 1677 5432
rect 1696 5449 1734 5458
rect 1696 5429 1705 5449
rect 1725 5429 1734 5449
rect 1592 5424 1628 5425
rect 1696 5421 1734 5429
rect 1800 5453 1944 5459
rect 1800 5433 1808 5453
rect 1828 5433 1916 5453
rect 1936 5433 1944 5453
rect 1800 5425 1944 5433
rect 1800 5424 1836 5425
rect 1908 5424 1944 5425
rect 2010 5458 2047 5459
rect 2010 5457 2048 5458
rect 2010 5449 2074 5457
rect 2010 5429 2019 5449
rect 2039 5435 2074 5449
rect 2094 5435 2097 5455
rect 2039 5430 2097 5435
rect 2039 5429 2074 5430
rect 420 5399 530 5413
rect 420 5396 463 5399
rect 109 5388 234 5395
rect 420 5391 424 5396
rect 109 5369 201 5388
rect 226 5369 234 5388
rect 109 5359 234 5369
rect 342 5369 424 5391
rect 453 5369 463 5396
rect 491 5372 498 5399
rect 527 5391 530 5399
rect 1276 5392 1313 5421
rect 527 5372 592 5391
rect 1277 5390 1313 5392
rect 1489 5390 1526 5421
rect 1697 5394 1734 5421
rect 2010 5417 2074 5429
rect 491 5369 592 5372
rect 342 5367 592 5369
rect 109 5339 149 5359
rect 108 5330 149 5339
rect 108 5312 118 5330
rect 136 5312 149 5330
rect 108 5303 149 5312
rect 108 5302 145 5303
rect 342 5288 379 5367
rect 420 5354 530 5367
rect 494 5298 525 5299
rect 342 5268 351 5288
rect 371 5268 379 5288
rect 342 5258 379 5268
rect 438 5288 525 5298
rect 438 5268 447 5288
rect 467 5268 525 5288
rect 438 5259 525 5268
rect 438 5258 475 5259
rect 111 5236 148 5240
rect 108 5231 148 5236
rect 108 5213 120 5231
rect 138 5213 148 5231
rect 108 5033 148 5213
rect 494 5206 525 5259
rect 555 5288 592 5367
rect 763 5364 1156 5384
rect 1176 5364 1179 5384
rect 1277 5368 1526 5390
rect 1695 5389 1736 5394
rect 2114 5391 2141 5569
rect 2792 5481 2819 5659
rect 3197 5656 3238 5661
rect 3407 5660 3656 5682
rect 3754 5666 3757 5686
rect 3777 5666 4170 5686
rect 4341 5683 4378 5762
rect 4408 5791 4439 5844
rect 4785 5837 4825 6017
rect 5163 6177 5203 6357
rect 5549 6350 5580 6403
rect 5610 6432 5647 6511
rect 5818 6508 6211 6528
rect 6231 6508 6234 6528
rect 6332 6512 6581 6534
rect 6750 6533 6791 6538
rect 7169 6535 7196 6713
rect 7847 6625 7874 6803
rect 8252 6800 8293 6805
rect 8462 6804 8711 6826
rect 8809 6810 8812 6830
rect 8832 6810 9225 6830
rect 9396 6827 9433 6906
rect 9463 6935 9494 6988
rect 9840 6981 9880 7161
rect 9840 6963 9850 6981
rect 9868 6963 9880 6981
rect 9840 6958 9880 6963
rect 9840 6954 9877 6958
rect 9513 6935 9550 6936
rect 9463 6926 9550 6935
rect 9463 6906 9521 6926
rect 9541 6906 9550 6926
rect 9463 6896 9550 6906
rect 9609 6926 9646 6936
rect 9609 6906 9617 6926
rect 9637 6906 9646 6926
rect 9463 6895 9494 6896
rect 9458 6827 9568 6840
rect 9609 6827 9646 6906
rect 9843 6891 9880 6892
rect 9839 6882 9880 6891
rect 9839 6864 9852 6882
rect 9870 6864 9880 6882
rect 9839 6855 9880 6864
rect 9839 6835 9879 6855
rect 9396 6825 9646 6827
rect 9396 6822 9497 6825
rect 7914 6765 7978 6777
rect 8254 6773 8291 6800
rect 8462 6773 8499 6804
rect 8675 6802 8711 6804
rect 9396 6803 9461 6822
rect 8675 6773 8712 6802
rect 9458 6795 9461 6803
rect 9490 6795 9497 6822
rect 9525 6798 9535 6825
rect 9564 6803 9646 6825
rect 9754 6825 9879 6835
rect 9754 6806 9762 6825
rect 9787 6806 9879 6825
rect 9564 6798 9568 6803
rect 9754 6799 9879 6806
rect 9525 6795 9568 6798
rect 9458 6781 9568 6795
rect 7914 6764 7949 6765
rect 7891 6759 7949 6764
rect 7891 6739 7894 6759
rect 7914 6745 7949 6759
rect 7969 6745 7978 6765
rect 7914 6737 7978 6745
rect 7940 6736 7978 6737
rect 7941 6735 7978 6736
rect 8044 6769 8080 6770
rect 8152 6769 8188 6770
rect 8044 6761 8188 6769
rect 8044 6741 8052 6761
rect 8072 6741 8160 6761
rect 8180 6741 8188 6761
rect 8044 6735 8188 6741
rect 8254 6765 8292 6773
rect 8360 6769 8396 6770
rect 8254 6745 8263 6765
rect 8283 6745 8292 6765
rect 8254 6736 8292 6745
rect 8311 6762 8396 6769
rect 8311 6742 8318 6762
rect 8339 6761 8396 6762
rect 8339 6742 8368 6761
rect 8311 6741 8368 6742
rect 8388 6741 8396 6761
rect 8254 6735 8291 6736
rect 8311 6735 8396 6741
rect 8462 6765 8500 6773
rect 8573 6769 8609 6770
rect 8462 6745 8471 6765
rect 8491 6745 8500 6765
rect 8462 6736 8500 6745
rect 8524 6761 8609 6769
rect 8524 6741 8581 6761
rect 8601 6741 8609 6761
rect 8462 6735 8499 6736
rect 8524 6735 8609 6741
rect 8675 6765 8713 6773
rect 8675 6745 8684 6765
rect 8704 6745 8713 6765
rect 8675 6736 8713 6745
rect 9839 6751 9879 6799
rect 8675 6735 8712 6736
rect 8098 6714 8134 6735
rect 8524 6714 8555 6735
rect 9839 6733 9850 6751
rect 9868 6733 9879 6751
rect 9839 6725 9879 6733
rect 9840 6724 9877 6725
rect 7931 6710 8031 6714
rect 7931 6706 7993 6710
rect 7931 6680 7938 6706
rect 7964 6684 7993 6706
rect 8019 6684 8031 6710
rect 7964 6680 8031 6684
rect 7931 6677 8031 6680
rect 8099 6677 8134 6714
rect 8196 6711 8555 6714
rect 8196 6706 8418 6711
rect 8196 6682 8209 6706
rect 8233 6687 8418 6706
rect 8442 6687 8555 6711
rect 8233 6682 8555 6687
rect 8196 6678 8555 6682
rect 8622 6706 8771 6714
rect 8622 6686 8633 6706
rect 8653 6686 8771 6706
rect 8622 6679 8771 6686
rect 9211 6683 9725 6684
rect 8622 6678 8663 6679
rect 8098 6642 8134 6677
rect 7946 6625 7983 6626
rect 8042 6625 8079 6626
rect 8098 6625 8105 6642
rect 7846 6616 7984 6625
rect 7846 6596 7955 6616
rect 7975 6596 7984 6616
rect 7846 6589 7984 6596
rect 8042 6616 8105 6625
rect 8042 6596 8051 6616
rect 8071 6601 8105 6616
rect 8126 6625 8134 6642
rect 8153 6625 8190 6626
rect 8126 6616 8190 6625
rect 8126 6601 8161 6616
rect 8071 6596 8161 6601
rect 8181 6596 8190 6616
rect 7846 6587 7942 6589
rect 8042 6586 8190 6596
rect 8249 6616 8286 6626
rect 8361 6625 8398 6626
rect 8342 6623 8398 6625
rect 8249 6596 8257 6616
rect 8277 6596 8286 6616
rect 8098 6585 8134 6586
rect 7028 6533 7196 6535
rect 6750 6527 7196 6533
rect 5818 6503 6234 6508
rect 6413 6506 6524 6512
rect 5818 6502 6159 6503
rect 5762 6442 5793 6443
rect 5610 6412 5619 6432
rect 5639 6412 5647 6432
rect 5610 6402 5647 6412
rect 5706 6435 5793 6442
rect 5706 6432 5767 6435
rect 5706 6412 5715 6432
rect 5735 6415 5767 6432
rect 5788 6415 5793 6435
rect 5735 6412 5793 6415
rect 5706 6405 5793 6412
rect 5818 6432 5855 6502
rect 6121 6501 6158 6502
rect 6413 6498 6454 6506
rect 6413 6478 6421 6498
rect 6440 6478 6454 6498
rect 6413 6476 6454 6478
rect 6482 6498 6524 6506
rect 6482 6478 6498 6498
rect 6517 6478 6524 6498
rect 6750 6505 6756 6527
rect 6782 6507 7196 6527
rect 7946 6526 7983 6527
rect 8249 6526 8286 6596
rect 8311 6616 8398 6623
rect 8311 6613 8369 6616
rect 8311 6593 8316 6613
rect 8337 6596 8369 6613
rect 8389 6596 8398 6616
rect 8337 6593 8398 6596
rect 8311 6586 8398 6593
rect 8457 6616 8494 6626
rect 8457 6596 8465 6616
rect 8485 6596 8494 6616
rect 8311 6585 8342 6586
rect 7945 6525 8286 6526
rect 6782 6505 6791 6507
rect 7028 6506 7196 6507
rect 7870 6524 8286 6525
rect 7870 6520 8246 6524
rect 6750 6496 6791 6505
rect 7870 6500 7873 6520
rect 7893 6507 8246 6520
rect 8278 6507 8286 6524
rect 7893 6500 8286 6507
rect 8457 6517 8494 6596
rect 8524 6625 8555 6678
rect 9192 6667 9725 6683
rect 9192 6656 9724 6667
rect 9843 6658 9880 6662
rect 8574 6625 8611 6626
rect 8524 6616 8611 6625
rect 8524 6596 8582 6616
rect 8602 6596 8611 6616
rect 8524 6586 8611 6596
rect 8670 6616 8707 6626
rect 8670 6596 8678 6616
rect 8698 6596 8707 6616
rect 8524 6585 8555 6586
rect 8519 6517 8629 6530
rect 8670 6517 8707 6596
rect 8457 6515 8707 6517
rect 8457 6512 8558 6515
rect 8457 6493 8522 6512
rect 6482 6476 6524 6478
rect 6413 6461 6524 6476
rect 8519 6485 8522 6493
rect 8551 6485 8558 6512
rect 8586 6488 8596 6515
rect 8625 6493 8707 6515
rect 8785 6587 8953 6588
rect 9192 6587 9230 6656
rect 8785 6567 9230 6587
rect 9457 6618 9568 6633
rect 9457 6616 9499 6618
rect 9457 6596 9464 6616
rect 9483 6596 9499 6616
rect 9457 6588 9499 6596
rect 9527 6616 9568 6618
rect 9527 6596 9541 6616
rect 9560 6596 9568 6616
rect 9527 6588 9568 6596
rect 9457 6582 9568 6588
rect 9690 6593 9724 6656
rect 9842 6652 9880 6658
rect 9842 6634 9852 6652
rect 9870 6634 9880 6652
rect 9842 6625 9880 6634
rect 9842 6593 9876 6625
rect 8785 6561 9229 6567
rect 8785 6559 8953 6561
rect 8625 6488 8629 6493
rect 8586 6485 8629 6488
rect 8519 6471 8629 6485
rect 5970 6442 6006 6443
rect 5818 6412 5827 6432
rect 5847 6412 5855 6432
rect 5706 6403 5762 6405
rect 5706 6402 5743 6403
rect 5818 6402 5855 6412
rect 5914 6432 6062 6442
rect 6162 6439 6258 6441
rect 5914 6412 5923 6432
rect 5943 6412 6033 6432
rect 6053 6412 6062 6432
rect 5914 6403 6062 6412
rect 6120 6432 6258 6439
rect 6120 6412 6129 6432
rect 6149 6412 6258 6432
rect 6120 6403 6258 6412
rect 5914 6402 5951 6403
rect 5970 6351 6006 6403
rect 6025 6402 6062 6403
rect 6121 6402 6158 6403
rect 5441 6349 5482 6350
rect 5333 6342 5482 6349
rect 5333 6322 5451 6342
rect 5471 6322 5482 6342
rect 5333 6314 5482 6322
rect 5549 6346 5908 6350
rect 5549 6341 5871 6346
rect 5549 6317 5662 6341
rect 5686 6322 5871 6341
rect 5895 6322 5908 6346
rect 5686 6317 5908 6322
rect 5549 6314 5908 6317
rect 5970 6314 6005 6351
rect 6073 6348 6173 6351
rect 6073 6344 6140 6348
rect 6073 6318 6085 6344
rect 6111 6322 6140 6344
rect 6166 6322 6173 6348
rect 6111 6318 6173 6322
rect 6073 6314 6173 6318
rect 5549 6293 5580 6314
rect 5970 6293 6006 6314
rect 5392 6292 5429 6293
rect 5391 6283 5429 6292
rect 5391 6263 5400 6283
rect 5420 6263 5429 6283
rect 5391 6255 5429 6263
rect 5495 6287 5580 6293
rect 5605 6292 5642 6293
rect 5495 6267 5503 6287
rect 5523 6267 5580 6287
rect 5495 6259 5580 6267
rect 5604 6283 5642 6292
rect 5604 6263 5613 6283
rect 5633 6263 5642 6283
rect 5495 6258 5531 6259
rect 5604 6255 5642 6263
rect 5708 6287 5793 6293
rect 5813 6292 5850 6293
rect 5708 6267 5716 6287
rect 5736 6286 5793 6287
rect 5736 6267 5765 6286
rect 5708 6266 5765 6267
rect 5786 6266 5793 6286
rect 5708 6259 5793 6266
rect 5812 6283 5850 6292
rect 5812 6263 5821 6283
rect 5841 6263 5850 6283
rect 5708 6258 5744 6259
rect 5812 6255 5850 6263
rect 5916 6287 6060 6293
rect 5916 6267 5924 6287
rect 5944 6284 6032 6287
rect 5944 6267 5975 6284
rect 5916 6264 5975 6267
rect 5998 6267 6032 6284
rect 6052 6267 6060 6287
rect 5998 6264 6060 6267
rect 5916 6259 6060 6264
rect 5916 6258 5952 6259
rect 6024 6258 6060 6259
rect 6126 6292 6163 6293
rect 6126 6291 6164 6292
rect 6126 6283 6190 6291
rect 6126 6263 6135 6283
rect 6155 6269 6190 6283
rect 6210 6269 6213 6289
rect 6155 6264 6213 6269
rect 6155 6263 6190 6264
rect 5392 6226 5429 6255
rect 5393 6224 5429 6226
rect 5605 6224 5642 6255
rect 5393 6202 5642 6224
rect 5813 6223 5850 6255
rect 6126 6251 6190 6263
rect 6230 6225 6257 6403
rect 8785 6381 8812 6559
rect 8852 6521 8916 6533
rect 9192 6529 9229 6561
rect 9400 6560 9649 6582
rect 9690 6561 9876 6593
rect 9704 6560 9876 6561
rect 9400 6529 9437 6560
rect 9613 6558 9649 6560
rect 9613 6529 9650 6558
rect 9842 6532 9876 6560
rect 8852 6520 8887 6521
rect 8829 6515 8887 6520
rect 8829 6495 8832 6515
rect 8852 6501 8887 6515
rect 8907 6501 8916 6521
rect 8852 6493 8916 6501
rect 8878 6492 8916 6493
rect 8879 6491 8916 6492
rect 8982 6525 9018 6526
rect 9090 6525 9126 6526
rect 8982 6518 9126 6525
rect 8982 6517 9042 6518
rect 8982 6497 8990 6517
rect 9010 6498 9042 6517
rect 9067 6517 9126 6518
rect 9067 6498 9098 6517
rect 9010 6497 9098 6498
rect 9118 6497 9126 6517
rect 8982 6491 9126 6497
rect 9192 6521 9230 6529
rect 9298 6525 9334 6526
rect 9192 6501 9201 6521
rect 9221 6501 9230 6521
rect 9192 6492 9230 6501
rect 9249 6518 9334 6525
rect 9249 6498 9256 6518
rect 9277 6517 9334 6518
rect 9277 6498 9306 6517
rect 9249 6497 9306 6498
rect 9326 6497 9334 6517
rect 9192 6491 9229 6492
rect 9249 6491 9334 6497
rect 9400 6521 9438 6529
rect 9511 6525 9547 6526
rect 9400 6501 9409 6521
rect 9429 6501 9438 6521
rect 9400 6492 9438 6501
rect 9462 6517 9547 6525
rect 9462 6497 9519 6517
rect 9539 6497 9547 6517
rect 9400 6491 9437 6492
rect 9462 6491 9547 6497
rect 9613 6521 9651 6529
rect 9613 6501 9622 6521
rect 9642 6501 9651 6521
rect 9613 6492 9651 6501
rect 9840 6522 9877 6532
rect 9840 6504 9850 6522
rect 9868 6504 9877 6522
rect 9840 6495 9877 6504
rect 9842 6494 9876 6495
rect 9613 6491 9650 6492
rect 9036 6470 9072 6491
rect 9462 6470 9493 6491
rect 8869 6466 8969 6470
rect 8869 6462 8931 6466
rect 8869 6436 8876 6462
rect 8902 6440 8931 6462
rect 8957 6440 8969 6466
rect 8902 6436 8969 6440
rect 8869 6433 8969 6436
rect 9037 6433 9072 6470
rect 9134 6467 9493 6470
rect 9134 6462 9356 6467
rect 9134 6438 9147 6462
rect 9171 6443 9356 6462
rect 9380 6443 9493 6467
rect 9171 6438 9493 6443
rect 9134 6434 9493 6438
rect 9560 6462 9709 6470
rect 9560 6442 9571 6462
rect 9591 6442 9709 6462
rect 9560 6435 9709 6442
rect 9560 6434 9601 6435
rect 8884 6381 8921 6382
rect 8980 6381 9017 6382
rect 9036 6381 9072 6433
rect 9091 6381 9128 6382
rect 8784 6372 8922 6381
rect 8379 6351 8490 6366
rect 8379 6349 8421 6351
rect 8049 6328 8154 6330
rect 7707 6320 7875 6321
rect 8049 6320 8098 6328
rect 7707 6301 8098 6320
rect 8129 6301 8154 6328
rect 8379 6329 8386 6349
rect 8405 6329 8421 6349
rect 8379 6321 8421 6329
rect 8449 6349 8490 6351
rect 8449 6329 8463 6349
rect 8482 6329 8490 6349
rect 8784 6352 8893 6372
rect 8913 6352 8922 6372
rect 8784 6345 8922 6352
rect 8980 6372 9128 6381
rect 8980 6352 8989 6372
rect 9009 6352 9099 6372
rect 9119 6352 9128 6372
rect 8784 6343 8880 6345
rect 8980 6342 9128 6352
rect 9187 6372 9224 6382
rect 9299 6381 9336 6382
rect 9280 6379 9336 6381
rect 9187 6352 9195 6372
rect 9215 6352 9224 6372
rect 9036 6341 9072 6342
rect 8449 6321 8490 6329
rect 8379 6315 8490 6321
rect 7707 6294 8154 6301
rect 7707 6292 7875 6294
rect 6555 6261 6665 6275
rect 6555 6258 6598 6261
rect 6555 6253 6559 6258
rect 6089 6223 6257 6225
rect 5813 6220 6257 6223
rect 5474 6196 5585 6202
rect 5474 6188 5515 6196
rect 5163 6133 5202 6177
rect 5474 6168 5482 6188
rect 5501 6168 5515 6188
rect 5474 6166 5515 6168
rect 5543 6188 5585 6196
rect 5543 6168 5559 6188
rect 5578 6168 5585 6188
rect 5543 6166 5585 6168
rect 5474 6151 5585 6166
rect 5811 6197 6257 6220
rect 5163 6109 5203 6133
rect 5503 6109 5550 6111
rect 5811 6109 5849 6197
rect 6089 6196 6257 6197
rect 6477 6231 6559 6253
rect 6588 6231 6598 6258
rect 6626 6234 6633 6261
rect 6662 6253 6665 6261
rect 6662 6234 6727 6253
rect 6626 6231 6727 6234
rect 6477 6229 6727 6231
rect 6477 6150 6514 6229
rect 6555 6216 6665 6229
rect 6629 6160 6660 6161
rect 6477 6130 6486 6150
rect 6506 6130 6514 6150
rect 6477 6120 6514 6130
rect 6573 6150 6660 6160
rect 6573 6130 6582 6150
rect 6602 6130 6660 6150
rect 6573 6121 6660 6130
rect 6573 6120 6610 6121
rect 5163 6076 5849 6109
rect 5163 6019 5202 6076
rect 5811 6074 5849 6076
rect 6629 6068 6660 6121
rect 6690 6150 6727 6229
rect 6898 6242 7291 6246
rect 6898 6225 6917 6242
rect 6937 6226 7291 6242
rect 7311 6226 7314 6246
rect 6937 6225 7314 6226
rect 6898 6221 7314 6225
rect 6898 6220 7239 6221
rect 6842 6160 6873 6161
rect 6690 6130 6699 6150
rect 6719 6130 6727 6150
rect 6690 6120 6727 6130
rect 6786 6153 6873 6160
rect 6786 6150 6847 6153
rect 6786 6130 6795 6150
rect 6815 6133 6847 6150
rect 6868 6133 6873 6153
rect 6815 6130 6873 6133
rect 6786 6123 6873 6130
rect 6898 6150 6935 6220
rect 7201 6219 7238 6220
rect 7050 6160 7086 6161
rect 6898 6130 6907 6150
rect 6927 6130 6935 6150
rect 6786 6121 6842 6123
rect 6786 6120 6823 6121
rect 6898 6120 6935 6130
rect 6994 6150 7142 6160
rect 7310 6159 7339 6160
rect 7242 6157 7339 6159
rect 6994 6130 7003 6150
rect 7023 6146 7113 6150
rect 7023 6130 7056 6146
rect 6994 6121 7056 6130
rect 6994 6120 7031 6121
rect 7050 6108 7056 6121
rect 7079 6130 7113 6146
rect 7133 6130 7142 6150
rect 7079 6121 7142 6130
rect 7200 6150 7339 6157
rect 7200 6130 7209 6150
rect 7229 6130 7339 6150
rect 7200 6121 7339 6130
rect 7079 6108 7086 6121
rect 7105 6120 7142 6121
rect 7201 6120 7238 6121
rect 7050 6069 7086 6108
rect 6521 6067 6562 6068
rect 6413 6060 6562 6067
rect 6413 6040 6531 6060
rect 6551 6040 6562 6060
rect 6413 6032 6562 6040
rect 6629 6064 6988 6068
rect 6629 6059 6951 6064
rect 6629 6035 6742 6059
rect 6766 6040 6951 6059
rect 6975 6040 6988 6064
rect 6766 6035 6988 6040
rect 6629 6032 6988 6035
rect 7050 6032 7085 6069
rect 7153 6066 7253 6069
rect 7153 6062 7220 6066
rect 7153 6036 7165 6062
rect 7191 6040 7220 6062
rect 7246 6040 7253 6066
rect 7191 6036 7253 6040
rect 7153 6032 7253 6036
rect 5163 6017 5211 6019
rect 5163 5999 5174 6017
rect 5192 5999 5211 6017
rect 6629 6011 6660 6032
rect 7050 6011 7086 6032
rect 6472 6010 6509 6011
rect 5163 5990 5211 5999
rect 5164 5989 5211 5990
rect 5477 5994 5587 6008
rect 5477 5991 5520 5994
rect 5477 5986 5481 5991
rect 5399 5964 5481 5986
rect 5510 5964 5520 5991
rect 5548 5967 5555 5994
rect 5584 5986 5587 5994
rect 6471 6001 6509 6010
rect 5584 5967 5649 5986
rect 6471 5981 6480 6001
rect 6500 5981 6509 6001
rect 5548 5964 5649 5967
rect 5399 5962 5649 5964
rect 5167 5926 5204 5927
rect 4785 5819 4795 5837
rect 4813 5819 4825 5837
rect 4785 5814 4825 5819
rect 5163 5923 5204 5926
rect 5163 5918 5205 5923
rect 5163 5900 5176 5918
rect 5194 5900 5205 5918
rect 5163 5886 5205 5900
rect 5243 5886 5290 5890
rect 5163 5880 5290 5886
rect 5163 5851 5251 5880
rect 5280 5851 5290 5880
rect 5399 5883 5436 5962
rect 5477 5949 5587 5962
rect 5551 5893 5582 5894
rect 5399 5863 5408 5883
rect 5428 5863 5436 5883
rect 5399 5853 5436 5863
rect 5495 5883 5582 5893
rect 5495 5863 5504 5883
rect 5524 5863 5582 5883
rect 5495 5854 5582 5863
rect 5495 5853 5532 5854
rect 5163 5847 5290 5851
rect 5163 5830 5202 5847
rect 5243 5846 5290 5847
rect 4785 5810 4822 5814
rect 5163 5812 5174 5830
rect 5192 5812 5202 5830
rect 5163 5803 5202 5812
rect 5164 5802 5201 5803
rect 5551 5801 5582 5854
rect 5612 5883 5649 5962
rect 5820 5959 6213 5979
rect 6233 5959 6236 5979
rect 6471 5973 6509 5981
rect 6575 6005 6660 6011
rect 6685 6010 6722 6011
rect 6575 5985 6583 6005
rect 6603 5985 6660 6005
rect 6575 5977 6660 5985
rect 6684 6001 6722 6010
rect 6684 5981 6693 6001
rect 6713 5981 6722 6001
rect 6575 5976 6611 5977
rect 6684 5973 6722 5981
rect 6788 6005 6873 6011
rect 6893 6010 6930 6011
rect 6788 5985 6796 6005
rect 6816 6004 6873 6005
rect 6816 5985 6845 6004
rect 6788 5984 6845 5985
rect 6866 5984 6873 6004
rect 6788 5977 6873 5984
rect 6892 6001 6930 6010
rect 6892 5981 6901 6001
rect 6921 5981 6930 6001
rect 6788 5976 6824 5977
rect 6892 5973 6930 5981
rect 6996 6005 7140 6011
rect 6996 5985 7004 6005
rect 7024 5985 7112 6005
rect 7132 5985 7140 6005
rect 6996 5977 7140 5985
rect 6996 5976 7032 5977
rect 7104 5976 7140 5977
rect 7206 6010 7243 6011
rect 7206 6009 7244 6010
rect 7206 6001 7270 6009
rect 7206 5981 7215 6001
rect 7235 5987 7270 6001
rect 7290 5987 7293 6007
rect 7235 5982 7293 5987
rect 7235 5981 7270 5982
rect 5820 5954 6236 5959
rect 5820 5953 6161 5954
rect 5764 5893 5795 5894
rect 5612 5863 5621 5883
rect 5641 5863 5649 5883
rect 5612 5853 5649 5863
rect 5708 5886 5795 5893
rect 5708 5883 5769 5886
rect 5708 5863 5717 5883
rect 5737 5866 5769 5883
rect 5790 5866 5795 5886
rect 5737 5863 5795 5866
rect 5708 5856 5795 5863
rect 5820 5883 5857 5953
rect 6123 5952 6160 5953
rect 6472 5944 6509 5973
rect 6473 5942 6509 5944
rect 6685 5942 6722 5973
rect 6473 5920 6722 5942
rect 6893 5941 6930 5973
rect 7206 5969 7270 5981
rect 7310 5943 7339 6121
rect 7707 6114 7734 6292
rect 7774 6254 7838 6266
rect 8114 6262 8151 6294
rect 8322 6293 8571 6315
rect 8322 6262 8359 6293
rect 8535 6291 8571 6293
rect 8535 6262 8572 6291
rect 8884 6282 8921 6283
rect 9187 6282 9224 6352
rect 9249 6372 9336 6379
rect 9249 6369 9307 6372
rect 9249 6349 9254 6369
rect 9275 6352 9307 6369
rect 9327 6352 9336 6372
rect 9275 6349 9336 6352
rect 9249 6342 9336 6349
rect 9395 6372 9432 6382
rect 9395 6352 9403 6372
rect 9423 6352 9432 6372
rect 9249 6341 9280 6342
rect 8883 6281 9224 6282
rect 8808 6276 9224 6281
rect 7774 6253 7809 6254
rect 7751 6248 7809 6253
rect 7751 6228 7754 6248
rect 7774 6234 7809 6248
rect 7829 6234 7838 6254
rect 7774 6226 7838 6234
rect 7800 6225 7838 6226
rect 7801 6224 7838 6225
rect 7904 6258 7940 6259
rect 8012 6258 8048 6259
rect 7904 6253 8048 6258
rect 7904 6250 7964 6253
rect 7904 6230 7912 6250
rect 7932 6232 7964 6250
rect 7991 6250 8048 6253
rect 7991 6232 8020 6250
rect 7932 6230 8020 6232
rect 8040 6230 8048 6250
rect 7904 6224 8048 6230
rect 8114 6254 8152 6262
rect 8220 6258 8256 6259
rect 8114 6234 8123 6254
rect 8143 6234 8152 6254
rect 8114 6225 8152 6234
rect 8171 6251 8256 6258
rect 8171 6231 8178 6251
rect 8199 6250 8256 6251
rect 8199 6231 8228 6250
rect 8171 6230 8228 6231
rect 8248 6230 8256 6250
rect 8114 6224 8151 6225
rect 8171 6224 8256 6230
rect 8322 6254 8360 6262
rect 8433 6258 8469 6259
rect 8322 6234 8331 6254
rect 8351 6234 8360 6254
rect 8322 6225 8360 6234
rect 8384 6250 8469 6258
rect 8384 6230 8441 6250
rect 8461 6230 8469 6250
rect 8322 6224 8359 6225
rect 8384 6224 8469 6230
rect 8535 6254 8573 6262
rect 8808 6256 8811 6276
rect 8831 6256 9224 6276
rect 9395 6273 9432 6352
rect 9462 6381 9493 6434
rect 9843 6432 9880 6433
rect 9842 6423 9881 6432
rect 9842 6405 9852 6423
rect 9870 6405 9881 6423
rect 9754 6388 9801 6389
rect 9842 6388 9881 6405
rect 9754 6384 9881 6388
rect 9512 6381 9549 6382
rect 9462 6372 9549 6381
rect 9462 6352 9520 6372
rect 9540 6352 9549 6372
rect 9462 6342 9549 6352
rect 9608 6372 9645 6382
rect 9608 6352 9616 6372
rect 9636 6352 9645 6372
rect 9462 6341 9493 6342
rect 9457 6273 9567 6286
rect 9608 6273 9645 6352
rect 9754 6355 9764 6384
rect 9793 6355 9881 6384
rect 9754 6349 9881 6355
rect 9754 6345 9801 6349
rect 9839 6335 9881 6349
rect 9839 6317 9850 6335
rect 9868 6317 9881 6335
rect 9839 6312 9881 6317
rect 9840 6309 9881 6312
rect 9840 6308 9877 6309
rect 9395 6271 9645 6273
rect 9395 6268 9496 6271
rect 8535 6234 8544 6254
rect 8564 6234 8573 6254
rect 9395 6249 9460 6268
rect 8535 6225 8573 6234
rect 9457 6241 9460 6249
rect 9489 6241 9496 6268
rect 9524 6244 9534 6271
rect 9563 6249 9645 6271
rect 9563 6244 9567 6249
rect 9524 6241 9567 6244
rect 9457 6227 9567 6241
rect 9833 6245 9880 6246
rect 9833 6236 9881 6245
rect 8535 6224 8572 6225
rect 7958 6203 7994 6224
rect 8384 6203 8415 6224
rect 9833 6218 9852 6236
rect 9870 6218 9881 6236
rect 9833 6216 9881 6218
rect 7791 6199 7891 6203
rect 7791 6195 7853 6199
rect 7791 6169 7798 6195
rect 7824 6173 7853 6195
rect 7879 6173 7891 6199
rect 7824 6169 7891 6173
rect 7791 6166 7891 6169
rect 7959 6166 7994 6203
rect 8056 6200 8415 6203
rect 8056 6195 8278 6200
rect 8056 6171 8069 6195
rect 8093 6176 8278 6195
rect 8302 6176 8415 6200
rect 8093 6171 8415 6176
rect 8056 6167 8415 6171
rect 8482 6195 8631 6203
rect 8482 6175 8493 6195
rect 8513 6175 8631 6195
rect 8482 6168 8631 6175
rect 8482 6167 8523 6168
rect 7806 6114 7843 6115
rect 7902 6114 7939 6115
rect 7958 6114 7994 6166
rect 8013 6114 8050 6115
rect 7706 6105 7844 6114
rect 7706 6085 7815 6105
rect 7835 6085 7844 6105
rect 7706 6078 7844 6085
rect 7902 6105 8050 6114
rect 7902 6085 7911 6105
rect 7931 6085 8021 6105
rect 8041 6085 8050 6105
rect 7706 6076 7802 6078
rect 7902 6075 8050 6085
rect 8109 6105 8146 6115
rect 8221 6114 8258 6115
rect 8202 6112 8258 6114
rect 8109 6085 8117 6105
rect 8137 6085 8146 6105
rect 7958 6074 7994 6075
rect 7806 6015 7843 6016
rect 8109 6015 8146 6085
rect 8171 6105 8258 6112
rect 8171 6102 8229 6105
rect 8171 6082 8176 6102
rect 8197 6085 8229 6102
rect 8249 6085 8258 6105
rect 8197 6082 8258 6085
rect 8171 6075 8258 6082
rect 8317 6105 8354 6115
rect 8317 6085 8325 6105
rect 8345 6085 8354 6105
rect 8171 6074 8202 6075
rect 7805 6014 8146 6015
rect 7730 6010 8146 6014
rect 7730 6009 8107 6010
rect 7730 5989 7733 6009
rect 7753 5993 8107 6009
rect 8127 5993 8146 6010
rect 7753 5989 8146 5993
rect 8317 6006 8354 6085
rect 8384 6114 8415 6167
rect 9195 6159 9233 6161
rect 9842 6159 9881 6216
rect 9195 6126 9881 6159
rect 8434 6114 8471 6115
rect 8384 6105 8471 6114
rect 8384 6085 8442 6105
rect 8462 6085 8471 6105
rect 8384 6075 8471 6085
rect 8530 6105 8567 6115
rect 8530 6085 8538 6105
rect 8558 6085 8567 6105
rect 8384 6074 8415 6075
rect 8379 6006 8489 6019
rect 8530 6006 8567 6085
rect 8317 6004 8567 6006
rect 8317 6001 8418 6004
rect 8317 5982 8382 6001
rect 8379 5974 8382 5982
rect 8411 5974 8418 6001
rect 8446 5977 8456 6004
rect 8485 5982 8567 6004
rect 8787 6038 8955 6039
rect 9195 6038 9233 6126
rect 9494 6124 9541 6126
rect 9841 6102 9881 6126
rect 8787 6015 9233 6038
rect 9459 6069 9570 6084
rect 9459 6067 9501 6069
rect 9459 6047 9466 6067
rect 9485 6047 9501 6067
rect 9459 6039 9501 6047
rect 9529 6067 9570 6069
rect 9529 6047 9543 6067
rect 9562 6047 9570 6067
rect 9842 6058 9881 6102
rect 9529 6039 9570 6047
rect 9459 6033 9570 6039
rect 8787 6012 9231 6015
rect 8787 6010 8955 6012
rect 8485 5977 8489 5982
rect 8446 5974 8489 5977
rect 8379 5960 8489 5974
rect 7169 5941 7339 5943
rect 6890 5934 7339 5941
rect 6554 5914 6665 5920
rect 6554 5906 6595 5914
rect 5972 5893 6008 5894
rect 5820 5863 5829 5883
rect 5849 5863 5857 5883
rect 5708 5854 5764 5856
rect 5708 5853 5745 5854
rect 5820 5853 5857 5863
rect 5916 5883 6064 5893
rect 6164 5890 6260 5892
rect 5916 5863 5925 5883
rect 5945 5863 6035 5883
rect 6055 5863 6064 5883
rect 5916 5854 6064 5863
rect 6122 5883 6260 5890
rect 6122 5863 6131 5883
rect 6151 5863 6260 5883
rect 6554 5886 6562 5906
rect 6581 5886 6595 5906
rect 6554 5884 6595 5886
rect 6623 5906 6665 5914
rect 6623 5886 6639 5906
rect 6658 5886 6665 5906
rect 6890 5907 6915 5934
rect 6946 5915 7339 5934
rect 6946 5907 6995 5915
rect 7169 5914 7339 5915
rect 6890 5905 6995 5907
rect 6623 5884 6665 5886
rect 6554 5869 6665 5884
rect 6122 5854 6260 5863
rect 5916 5853 5953 5854
rect 5972 5802 6008 5854
rect 6027 5853 6064 5854
rect 6123 5853 6160 5854
rect 5443 5800 5484 5801
rect 5335 5793 5484 5800
rect 4458 5791 4495 5792
rect 4408 5782 4495 5791
rect 4408 5762 4466 5782
rect 4486 5762 4495 5782
rect 4408 5752 4495 5762
rect 4554 5782 4591 5792
rect 4554 5762 4562 5782
rect 4582 5762 4591 5782
rect 5335 5773 5453 5793
rect 5473 5773 5484 5793
rect 5335 5765 5484 5773
rect 5551 5797 5910 5801
rect 5551 5792 5873 5797
rect 5551 5768 5664 5792
rect 5688 5773 5873 5792
rect 5897 5773 5910 5797
rect 5688 5768 5910 5773
rect 5551 5765 5910 5768
rect 5972 5765 6007 5802
rect 6075 5799 6175 5802
rect 6075 5795 6142 5799
rect 6075 5769 6087 5795
rect 6113 5773 6142 5795
rect 6168 5773 6175 5799
rect 6113 5769 6175 5773
rect 6075 5765 6175 5769
rect 4408 5751 4439 5752
rect 4403 5683 4513 5696
rect 4554 5683 4591 5762
rect 4788 5747 4825 5748
rect 4784 5738 4825 5747
rect 5551 5744 5582 5765
rect 5972 5744 6008 5765
rect 5394 5743 5431 5744
rect 5168 5740 5202 5741
rect 4784 5720 4797 5738
rect 4815 5720 4825 5738
rect 4784 5711 4825 5720
rect 5167 5731 5204 5740
rect 5167 5713 5176 5731
rect 5194 5713 5204 5731
rect 4784 5691 4824 5711
rect 5167 5703 5204 5713
rect 5393 5734 5431 5743
rect 5393 5714 5402 5734
rect 5422 5714 5431 5734
rect 5393 5706 5431 5714
rect 5497 5738 5582 5744
rect 5607 5743 5644 5744
rect 5497 5718 5505 5738
rect 5525 5718 5582 5738
rect 5497 5710 5582 5718
rect 5606 5734 5644 5743
rect 5606 5714 5615 5734
rect 5635 5714 5644 5734
rect 5497 5709 5533 5710
rect 5606 5706 5644 5714
rect 5710 5738 5795 5744
rect 5815 5743 5852 5744
rect 5710 5718 5718 5738
rect 5738 5737 5795 5738
rect 5738 5718 5767 5737
rect 5710 5717 5767 5718
rect 5788 5717 5795 5737
rect 5710 5710 5795 5717
rect 5814 5734 5852 5743
rect 5814 5714 5823 5734
rect 5843 5714 5852 5734
rect 5710 5709 5746 5710
rect 5814 5706 5852 5714
rect 5918 5738 6062 5744
rect 5918 5718 5926 5738
rect 5946 5737 6034 5738
rect 5946 5718 5977 5737
rect 5918 5717 5977 5718
rect 6002 5718 6034 5737
rect 6054 5718 6062 5738
rect 6002 5717 6062 5718
rect 5918 5710 6062 5717
rect 5918 5709 5954 5710
rect 6026 5709 6062 5710
rect 6128 5743 6165 5744
rect 6128 5742 6166 5743
rect 6128 5734 6192 5742
rect 6128 5714 6137 5734
rect 6157 5720 6192 5734
rect 6212 5720 6215 5740
rect 6157 5715 6215 5720
rect 6157 5714 6192 5715
rect 4341 5681 4591 5683
rect 4341 5678 4442 5681
rect 2859 5621 2923 5633
rect 3199 5629 3236 5656
rect 3407 5629 3444 5660
rect 3620 5658 3656 5660
rect 4341 5659 4406 5678
rect 3620 5629 3657 5658
rect 4403 5651 4406 5659
rect 4435 5651 4442 5678
rect 4470 5654 4480 5681
rect 4509 5659 4591 5681
rect 4699 5681 4824 5691
rect 4699 5662 4707 5681
rect 4732 5662 4824 5681
rect 4509 5654 4513 5659
rect 4699 5655 4824 5662
rect 4470 5651 4513 5654
rect 4403 5637 4513 5651
rect 2859 5620 2894 5621
rect 2836 5615 2894 5620
rect 2836 5595 2839 5615
rect 2859 5601 2894 5615
rect 2914 5601 2923 5621
rect 2859 5593 2923 5601
rect 2885 5592 2923 5593
rect 2886 5591 2923 5592
rect 2989 5625 3025 5626
rect 3097 5625 3133 5626
rect 2989 5617 3133 5625
rect 2989 5597 2997 5617
rect 3017 5614 3105 5617
rect 3017 5597 3049 5614
rect 3069 5597 3105 5614
rect 3125 5597 3133 5617
rect 2989 5591 3133 5597
rect 3199 5621 3237 5629
rect 3305 5625 3341 5626
rect 3199 5601 3208 5621
rect 3228 5601 3237 5621
rect 3199 5592 3237 5601
rect 3256 5618 3341 5625
rect 3256 5598 3263 5618
rect 3284 5617 3341 5618
rect 3284 5598 3313 5617
rect 3256 5597 3313 5598
rect 3333 5597 3341 5617
rect 3199 5591 3236 5592
rect 3256 5591 3341 5597
rect 3407 5621 3445 5629
rect 3518 5625 3554 5626
rect 3407 5601 3416 5621
rect 3436 5601 3445 5621
rect 3407 5592 3445 5601
rect 3469 5617 3554 5625
rect 3469 5597 3526 5617
rect 3546 5597 3554 5617
rect 3407 5591 3444 5592
rect 3469 5591 3554 5597
rect 3620 5621 3658 5629
rect 3620 5601 3629 5621
rect 3649 5601 3658 5621
rect 3620 5592 3658 5601
rect 4784 5607 4824 5655
rect 5168 5675 5202 5703
rect 5394 5677 5431 5706
rect 5395 5675 5431 5677
rect 5607 5675 5644 5706
rect 5168 5674 5340 5675
rect 5168 5642 5354 5674
rect 5395 5653 5644 5675
rect 5815 5674 5852 5706
rect 6128 5702 6192 5714
rect 6232 5676 6259 5854
rect 8787 5832 8814 6010
rect 8854 5972 8918 5984
rect 9194 5980 9231 6012
rect 9402 6011 9651 6033
rect 9402 5980 9439 6011
rect 9615 6009 9651 6011
rect 9615 5980 9652 6009
rect 8854 5971 8889 5972
rect 8831 5966 8889 5971
rect 8831 5946 8834 5966
rect 8854 5952 8889 5966
rect 8909 5952 8918 5972
rect 8854 5944 8918 5952
rect 8880 5943 8918 5944
rect 8881 5942 8918 5943
rect 8984 5976 9020 5977
rect 9092 5976 9128 5977
rect 8984 5971 9128 5976
rect 8984 5968 9046 5971
rect 8984 5948 8992 5968
rect 9012 5951 9046 5968
rect 9069 5968 9128 5971
rect 9069 5951 9100 5968
rect 9012 5948 9100 5951
rect 9120 5948 9128 5968
rect 8984 5942 9128 5948
rect 9194 5972 9232 5980
rect 9300 5976 9336 5977
rect 9194 5952 9203 5972
rect 9223 5952 9232 5972
rect 9194 5943 9232 5952
rect 9251 5969 9336 5976
rect 9251 5949 9258 5969
rect 9279 5968 9336 5969
rect 9279 5949 9308 5968
rect 9251 5948 9308 5949
rect 9328 5948 9336 5968
rect 9194 5942 9231 5943
rect 9251 5942 9336 5948
rect 9402 5972 9440 5980
rect 9513 5976 9549 5977
rect 9402 5952 9411 5972
rect 9431 5952 9440 5972
rect 9402 5943 9440 5952
rect 9464 5968 9549 5976
rect 9464 5948 9521 5968
rect 9541 5948 9549 5968
rect 9402 5942 9439 5943
rect 9464 5942 9549 5948
rect 9615 5972 9653 5980
rect 9615 5952 9624 5972
rect 9644 5952 9653 5972
rect 9615 5943 9653 5952
rect 9615 5942 9652 5943
rect 9038 5921 9074 5942
rect 9464 5921 9495 5942
rect 8871 5917 8971 5921
rect 8871 5913 8933 5917
rect 8871 5887 8878 5913
rect 8904 5891 8933 5913
rect 8959 5891 8971 5917
rect 8904 5887 8971 5891
rect 8871 5884 8971 5887
rect 9039 5884 9074 5921
rect 9136 5918 9495 5921
rect 9136 5913 9358 5918
rect 9136 5889 9149 5913
rect 9173 5894 9358 5913
rect 9382 5894 9495 5918
rect 9173 5889 9495 5894
rect 9136 5885 9495 5889
rect 9562 5913 9711 5921
rect 9562 5893 9573 5913
rect 9593 5893 9711 5913
rect 9562 5886 9711 5893
rect 9562 5885 9603 5886
rect 8886 5832 8923 5833
rect 8982 5832 9019 5833
rect 9038 5832 9074 5884
rect 9093 5832 9130 5833
rect 8786 5823 8924 5832
rect 8786 5803 8895 5823
rect 8915 5803 8924 5823
rect 8786 5796 8924 5803
rect 8982 5823 9130 5832
rect 8982 5803 8991 5823
rect 9011 5803 9101 5823
rect 9121 5803 9130 5823
rect 8786 5794 8882 5796
rect 8982 5793 9130 5803
rect 9189 5823 9226 5833
rect 9301 5832 9338 5833
rect 9282 5830 9338 5832
rect 9189 5803 9197 5823
rect 9217 5803 9226 5823
rect 9038 5792 9074 5793
rect 6415 5750 6525 5764
rect 6415 5747 6458 5750
rect 6415 5742 6419 5747
rect 6091 5674 6259 5676
rect 5815 5668 6259 5674
rect 5168 5610 5202 5642
rect 3620 5591 3657 5592
rect 3043 5570 3079 5591
rect 3469 5570 3500 5591
rect 4784 5589 4795 5607
rect 4813 5589 4824 5607
rect 4784 5581 4824 5589
rect 5164 5601 5202 5610
rect 5164 5583 5174 5601
rect 5192 5583 5202 5601
rect 4785 5580 4822 5581
rect 5164 5577 5202 5583
rect 5320 5579 5354 5642
rect 5476 5647 5587 5653
rect 5476 5639 5517 5647
rect 5476 5619 5484 5639
rect 5503 5619 5517 5639
rect 5476 5617 5517 5619
rect 5545 5639 5587 5647
rect 5545 5619 5561 5639
rect 5580 5619 5587 5639
rect 5545 5617 5587 5619
rect 5476 5602 5587 5617
rect 5814 5648 6259 5668
rect 5814 5579 5852 5648
rect 6091 5647 6259 5648
rect 6337 5720 6419 5742
rect 6448 5720 6458 5747
rect 6486 5723 6493 5750
rect 6522 5742 6525 5750
rect 8520 5759 8631 5774
rect 8520 5757 8562 5759
rect 6522 5723 6587 5742
rect 6486 5720 6587 5723
rect 6337 5718 6587 5720
rect 6337 5639 6374 5718
rect 6415 5705 6525 5718
rect 6489 5649 6520 5650
rect 6337 5619 6346 5639
rect 6366 5619 6374 5639
rect 6337 5609 6374 5619
rect 6433 5639 6520 5649
rect 6433 5619 6442 5639
rect 6462 5619 6520 5639
rect 6433 5610 6520 5619
rect 6433 5609 6470 5610
rect 5164 5573 5201 5577
rect 2876 5566 2976 5570
rect 2876 5562 2938 5566
rect 2876 5536 2883 5562
rect 2909 5540 2938 5562
rect 2964 5540 2976 5566
rect 2909 5536 2976 5540
rect 2876 5533 2976 5536
rect 3044 5533 3079 5570
rect 3141 5567 3500 5570
rect 3141 5562 3363 5567
rect 3141 5538 3154 5562
rect 3178 5543 3363 5562
rect 3387 5543 3500 5567
rect 3178 5538 3500 5543
rect 3141 5534 3500 5538
rect 3567 5562 3716 5570
rect 5320 5568 5852 5579
rect 3567 5542 3578 5562
rect 3598 5542 3716 5562
rect 5319 5552 5852 5568
rect 6489 5557 6520 5610
rect 6550 5639 6587 5718
rect 6758 5728 7151 5735
rect 6758 5711 6766 5728
rect 6798 5715 7151 5728
rect 7171 5715 7174 5735
rect 8253 5730 8294 5739
rect 6798 5711 7174 5715
rect 6758 5710 7174 5711
rect 7848 5728 8016 5729
rect 8253 5728 8262 5730
rect 6758 5709 7099 5710
rect 6702 5649 6733 5650
rect 6550 5619 6559 5639
rect 6579 5619 6587 5639
rect 6550 5609 6587 5619
rect 6646 5642 6733 5649
rect 6646 5639 6707 5642
rect 6646 5619 6655 5639
rect 6675 5622 6707 5639
rect 6728 5622 6733 5642
rect 6675 5619 6733 5622
rect 6646 5612 6733 5619
rect 6758 5639 6795 5709
rect 7061 5708 7098 5709
rect 7848 5708 8262 5728
rect 8288 5708 8294 5730
rect 8520 5737 8527 5757
rect 8546 5737 8562 5757
rect 8520 5729 8562 5737
rect 8590 5757 8631 5759
rect 8590 5737 8604 5757
rect 8623 5737 8631 5757
rect 8590 5729 8631 5737
rect 8886 5733 8923 5734
rect 9189 5733 9226 5803
rect 9251 5823 9338 5830
rect 9251 5820 9309 5823
rect 9251 5800 9256 5820
rect 9277 5803 9309 5820
rect 9329 5803 9338 5823
rect 9277 5800 9338 5803
rect 9251 5793 9338 5800
rect 9397 5823 9434 5833
rect 9397 5803 9405 5823
rect 9425 5803 9434 5823
rect 9251 5792 9282 5793
rect 8885 5732 9226 5733
rect 8520 5723 8631 5729
rect 8810 5727 9226 5732
rect 7848 5702 8294 5708
rect 7848 5700 8016 5702
rect 6910 5649 6946 5650
rect 6758 5619 6767 5639
rect 6787 5619 6795 5639
rect 6646 5610 6702 5612
rect 6646 5609 6683 5610
rect 6758 5609 6795 5619
rect 6854 5639 7002 5649
rect 7102 5646 7198 5648
rect 6854 5619 6863 5639
rect 6883 5634 6973 5639
rect 6883 5619 6918 5634
rect 6854 5610 6918 5619
rect 6854 5609 6891 5610
rect 6910 5593 6918 5610
rect 6939 5619 6973 5634
rect 6993 5619 7002 5639
rect 6939 5610 7002 5619
rect 7060 5639 7198 5646
rect 7060 5619 7069 5639
rect 7089 5619 7198 5639
rect 7060 5610 7198 5619
rect 6939 5593 6946 5610
rect 6965 5609 7002 5610
rect 7061 5609 7098 5610
rect 6910 5558 6946 5593
rect 6381 5556 6422 5557
rect 5319 5551 5833 5552
rect 3567 5535 3716 5542
rect 6273 5549 6422 5556
rect 4156 5539 4670 5540
rect 3567 5534 3608 5535
rect 2891 5481 2928 5482
rect 2987 5481 3024 5482
rect 3043 5481 3079 5533
rect 3098 5481 3135 5482
rect 2791 5472 2929 5481
rect 2791 5452 2900 5472
rect 2920 5452 2929 5472
rect 2791 5445 2929 5452
rect 2987 5472 3135 5481
rect 2987 5452 2996 5472
rect 3016 5452 3106 5472
rect 3126 5452 3135 5472
rect 2791 5443 2887 5445
rect 2987 5442 3135 5452
rect 3194 5472 3231 5482
rect 3306 5481 3343 5482
rect 3287 5479 3343 5481
rect 3194 5452 3202 5472
rect 3222 5452 3231 5472
rect 3043 5441 3079 5442
rect 1973 5389 2141 5391
rect 1695 5383 2141 5389
rect 763 5359 1179 5364
rect 1358 5362 1469 5368
rect 763 5358 1104 5359
rect 707 5298 738 5299
rect 555 5268 564 5288
rect 584 5268 592 5288
rect 555 5258 592 5268
rect 651 5291 738 5298
rect 651 5288 712 5291
rect 651 5268 660 5288
rect 680 5271 712 5288
rect 733 5271 738 5291
rect 680 5268 738 5271
rect 651 5261 738 5268
rect 763 5288 800 5358
rect 1066 5357 1103 5358
rect 1358 5354 1399 5362
rect 1358 5334 1366 5354
rect 1385 5334 1399 5354
rect 1358 5332 1399 5334
rect 1427 5354 1469 5362
rect 1427 5334 1443 5354
rect 1462 5334 1469 5354
rect 1695 5361 1701 5383
rect 1727 5363 2141 5383
rect 2891 5382 2928 5383
rect 3194 5382 3231 5452
rect 3256 5472 3343 5479
rect 3256 5469 3314 5472
rect 3256 5449 3261 5469
rect 3282 5452 3314 5469
rect 3334 5452 3343 5472
rect 3282 5449 3343 5452
rect 3256 5442 3343 5449
rect 3402 5472 3439 5482
rect 3402 5452 3410 5472
rect 3430 5452 3439 5472
rect 3256 5441 3287 5442
rect 2890 5381 3231 5382
rect 1727 5361 1736 5363
rect 1973 5362 2141 5363
rect 2815 5376 3231 5381
rect 1695 5352 1736 5361
rect 2815 5356 2818 5376
rect 2838 5356 3231 5376
rect 3402 5373 3439 5452
rect 3469 5481 3500 5534
rect 4137 5523 4670 5539
rect 6273 5529 6391 5549
rect 6411 5529 6422 5549
rect 4137 5512 4669 5523
rect 6273 5521 6422 5529
rect 6489 5553 6848 5557
rect 6489 5548 6811 5553
rect 6489 5524 6602 5548
rect 6626 5529 6811 5548
rect 6835 5529 6848 5553
rect 6626 5524 6848 5529
rect 6489 5521 6848 5524
rect 6910 5521 6945 5558
rect 7013 5555 7113 5558
rect 7013 5551 7080 5555
rect 7013 5525 7025 5551
rect 7051 5529 7080 5551
rect 7106 5529 7113 5555
rect 7051 5525 7113 5529
rect 7013 5521 7113 5525
rect 4788 5514 4825 5518
rect 3519 5481 3556 5482
rect 3469 5472 3556 5481
rect 3469 5452 3527 5472
rect 3547 5452 3556 5472
rect 3469 5442 3556 5452
rect 3615 5472 3652 5482
rect 3615 5452 3623 5472
rect 3643 5452 3652 5472
rect 3469 5441 3500 5442
rect 3464 5373 3574 5386
rect 3615 5373 3652 5452
rect 3402 5371 3652 5373
rect 3402 5368 3503 5371
rect 3402 5349 3467 5368
rect 3464 5341 3467 5349
rect 3496 5341 3503 5368
rect 3531 5344 3541 5371
rect 3570 5349 3652 5371
rect 3730 5443 3898 5444
rect 4137 5443 4175 5512
rect 3730 5423 4175 5443
rect 4402 5474 4513 5489
rect 4402 5472 4444 5474
rect 4402 5452 4409 5472
rect 4428 5452 4444 5472
rect 4402 5444 4444 5452
rect 4472 5472 4513 5474
rect 4472 5452 4486 5472
rect 4505 5452 4513 5472
rect 4472 5444 4513 5452
rect 4402 5438 4513 5444
rect 4635 5449 4669 5512
rect 4787 5508 4825 5514
rect 5167 5510 5204 5511
rect 4787 5490 4797 5508
rect 4815 5490 4825 5508
rect 4787 5481 4825 5490
rect 5165 5502 5205 5510
rect 5165 5484 5176 5502
rect 5194 5484 5205 5502
rect 6489 5500 6520 5521
rect 6910 5500 6946 5521
rect 6332 5499 6369 5500
rect 4787 5449 4821 5481
rect 3730 5417 4174 5423
rect 3730 5415 3898 5417
rect 3570 5344 3574 5349
rect 3531 5341 3574 5344
rect 1427 5332 1469 5334
rect 1358 5317 1469 5332
rect 2554 5323 2602 5337
rect 3464 5327 3574 5341
rect 915 5298 951 5299
rect 763 5268 772 5288
rect 792 5268 800 5288
rect 651 5259 707 5261
rect 651 5258 688 5259
rect 763 5258 800 5268
rect 859 5288 1007 5298
rect 1107 5295 1203 5297
rect 859 5268 868 5288
rect 888 5268 978 5288
rect 998 5268 1007 5288
rect 859 5259 1007 5268
rect 1065 5288 1203 5295
rect 1065 5268 1074 5288
rect 1094 5268 1203 5288
rect 1065 5259 1203 5268
rect 2554 5283 2567 5323
rect 2594 5283 2602 5323
rect 2554 5265 2602 5283
rect 859 5258 896 5259
rect 915 5207 951 5259
rect 970 5258 1007 5259
rect 1066 5258 1103 5259
rect 386 5205 427 5206
rect 278 5198 427 5205
rect 278 5178 396 5198
rect 416 5178 427 5198
rect 278 5170 427 5178
rect 494 5202 853 5206
rect 494 5197 816 5202
rect 494 5173 607 5197
rect 631 5178 816 5197
rect 840 5178 853 5202
rect 631 5173 853 5178
rect 494 5170 853 5173
rect 915 5170 950 5207
rect 1018 5204 1118 5207
rect 1018 5200 1085 5204
rect 1018 5174 1030 5200
rect 1056 5178 1085 5200
rect 1111 5178 1118 5204
rect 1056 5174 1118 5178
rect 1018 5170 1118 5174
rect 494 5149 525 5170
rect 915 5149 951 5170
rect 337 5148 374 5149
rect 336 5139 374 5148
rect 336 5119 345 5139
rect 365 5119 374 5139
rect 336 5111 374 5119
rect 440 5143 525 5149
rect 550 5148 587 5149
rect 440 5123 448 5143
rect 468 5123 525 5143
rect 440 5115 525 5123
rect 549 5139 587 5148
rect 549 5119 558 5139
rect 578 5119 587 5139
rect 440 5114 476 5115
rect 549 5111 587 5119
rect 653 5143 738 5149
rect 758 5148 795 5149
rect 653 5123 661 5143
rect 681 5142 738 5143
rect 681 5123 710 5142
rect 653 5122 710 5123
rect 731 5122 738 5142
rect 653 5115 738 5122
rect 757 5139 795 5148
rect 757 5119 766 5139
rect 786 5119 795 5139
rect 653 5114 689 5115
rect 757 5111 795 5119
rect 861 5143 1005 5149
rect 861 5123 869 5143
rect 889 5140 977 5143
rect 889 5123 920 5140
rect 861 5120 920 5123
rect 943 5123 977 5140
rect 997 5123 1005 5143
rect 943 5120 1005 5123
rect 861 5115 1005 5120
rect 861 5114 897 5115
rect 969 5114 1005 5115
rect 1071 5148 1108 5149
rect 1071 5147 1109 5148
rect 1071 5139 1135 5147
rect 1071 5119 1080 5139
rect 1100 5125 1135 5139
rect 1155 5125 1158 5145
rect 1100 5120 1158 5125
rect 1100 5119 1135 5120
rect 337 5082 374 5111
rect 338 5080 374 5082
rect 550 5080 587 5111
rect 338 5058 587 5080
rect 758 5079 795 5111
rect 1071 5107 1135 5119
rect 1175 5081 1202 5259
rect 2549 5158 2602 5265
rect 3730 5237 3757 5415
rect 3797 5377 3861 5389
rect 4137 5385 4174 5417
rect 4345 5416 4594 5438
rect 4635 5417 4821 5449
rect 4649 5416 4821 5417
rect 4345 5385 4382 5416
rect 4558 5414 4594 5416
rect 4558 5385 4595 5414
rect 4787 5388 4821 5416
rect 5165 5436 5205 5484
rect 6331 5490 6369 5499
rect 6331 5470 6340 5490
rect 6360 5470 6369 5490
rect 6331 5462 6369 5470
rect 6435 5494 6520 5500
rect 6545 5499 6582 5500
rect 6435 5474 6443 5494
rect 6463 5474 6520 5494
rect 6435 5466 6520 5474
rect 6544 5490 6582 5499
rect 6544 5470 6553 5490
rect 6573 5470 6582 5490
rect 6435 5465 6471 5466
rect 6544 5462 6582 5470
rect 6648 5494 6733 5500
rect 6753 5499 6790 5500
rect 6648 5474 6656 5494
rect 6676 5493 6733 5494
rect 6676 5474 6705 5493
rect 6648 5473 6705 5474
rect 6726 5473 6733 5493
rect 6648 5466 6733 5473
rect 6752 5490 6790 5499
rect 6752 5470 6761 5490
rect 6781 5470 6790 5490
rect 6648 5465 6684 5466
rect 6752 5462 6790 5470
rect 6856 5494 7000 5500
rect 6856 5474 6864 5494
rect 6884 5474 6972 5494
rect 6992 5474 7000 5494
rect 6856 5466 7000 5474
rect 6856 5465 6892 5466
rect 6964 5465 7000 5466
rect 7066 5499 7103 5500
rect 7066 5498 7104 5499
rect 7066 5490 7130 5498
rect 7066 5470 7075 5490
rect 7095 5476 7130 5490
rect 7150 5476 7153 5496
rect 7095 5471 7153 5476
rect 7095 5470 7130 5471
rect 5476 5440 5586 5454
rect 5476 5437 5519 5440
rect 5165 5429 5290 5436
rect 5476 5432 5480 5437
rect 5165 5410 5257 5429
rect 5282 5410 5290 5429
rect 5165 5400 5290 5410
rect 5398 5410 5480 5432
rect 5509 5410 5519 5437
rect 5547 5413 5554 5440
rect 5583 5432 5586 5440
rect 6332 5433 6369 5462
rect 5583 5413 5648 5432
rect 6333 5431 6369 5433
rect 6545 5431 6582 5462
rect 6753 5435 6790 5462
rect 7066 5458 7130 5470
rect 5547 5410 5648 5413
rect 5398 5408 5648 5410
rect 3797 5376 3832 5377
rect 3774 5371 3832 5376
rect 3774 5351 3777 5371
rect 3797 5357 3832 5371
rect 3852 5357 3861 5377
rect 3797 5349 3861 5357
rect 3823 5348 3861 5349
rect 3824 5347 3861 5348
rect 3927 5381 3963 5382
rect 4035 5381 4071 5382
rect 3927 5374 4071 5381
rect 3927 5373 3987 5374
rect 3927 5353 3935 5373
rect 3955 5354 3987 5373
rect 4012 5373 4071 5374
rect 4012 5354 4043 5373
rect 3955 5353 4043 5354
rect 4063 5353 4071 5373
rect 3927 5347 4071 5353
rect 4137 5377 4175 5385
rect 4243 5381 4279 5382
rect 4137 5357 4146 5377
rect 4166 5357 4175 5377
rect 4137 5348 4175 5357
rect 4194 5374 4279 5381
rect 4194 5354 4201 5374
rect 4222 5373 4279 5374
rect 4222 5354 4251 5373
rect 4194 5353 4251 5354
rect 4271 5353 4279 5373
rect 4137 5347 4174 5348
rect 4194 5347 4279 5353
rect 4345 5377 4383 5385
rect 4456 5381 4492 5382
rect 4345 5357 4354 5377
rect 4374 5357 4383 5377
rect 4345 5348 4383 5357
rect 4407 5373 4492 5381
rect 4407 5353 4464 5373
rect 4484 5353 4492 5373
rect 4345 5347 4382 5348
rect 4407 5347 4492 5353
rect 4558 5377 4596 5385
rect 4558 5357 4567 5377
rect 4587 5357 4596 5377
rect 4558 5348 4596 5357
rect 4785 5378 4822 5388
rect 5165 5380 5205 5400
rect 4785 5360 4795 5378
rect 4813 5360 4822 5378
rect 4785 5351 4822 5360
rect 5164 5371 5205 5380
rect 5164 5353 5174 5371
rect 5192 5353 5205 5371
rect 4787 5350 4821 5351
rect 4558 5347 4595 5348
rect 3981 5326 4017 5347
rect 4407 5326 4438 5347
rect 5164 5344 5205 5353
rect 5164 5343 5201 5344
rect 5398 5329 5435 5408
rect 5476 5395 5586 5408
rect 5550 5339 5581 5340
rect 3814 5322 3914 5326
rect 3814 5318 3876 5322
rect 3814 5292 3821 5318
rect 3847 5296 3876 5318
rect 3902 5296 3914 5322
rect 3847 5292 3914 5296
rect 3814 5289 3914 5292
rect 3982 5289 4017 5326
rect 4079 5323 4438 5326
rect 4079 5318 4301 5323
rect 4079 5294 4092 5318
rect 4116 5299 4301 5318
rect 4325 5299 4438 5323
rect 4116 5294 4438 5299
rect 4079 5290 4438 5294
rect 4505 5318 4654 5326
rect 4505 5298 4516 5318
rect 4536 5298 4654 5318
rect 5398 5309 5407 5329
rect 5427 5309 5435 5329
rect 5398 5299 5435 5309
rect 5494 5329 5581 5339
rect 5494 5309 5503 5329
rect 5523 5309 5581 5329
rect 5494 5300 5581 5309
rect 5494 5299 5531 5300
rect 4505 5291 4654 5298
rect 4505 5290 4546 5291
rect 3829 5237 3866 5238
rect 3925 5237 3962 5238
rect 3981 5237 4017 5289
rect 4036 5237 4073 5238
rect 3729 5228 3867 5237
rect 3729 5208 3838 5228
rect 3858 5208 3867 5228
rect 3355 5188 3466 5203
rect 3729 5201 3867 5208
rect 3925 5228 4073 5237
rect 3925 5208 3934 5228
rect 3954 5208 4044 5228
rect 4064 5208 4073 5228
rect 3729 5199 3825 5201
rect 3925 5198 4073 5208
rect 4132 5228 4169 5238
rect 4244 5237 4281 5238
rect 4225 5235 4281 5237
rect 4132 5208 4140 5228
rect 4160 5208 4169 5228
rect 3981 5197 4017 5198
rect 3355 5186 3397 5188
rect 3355 5166 3362 5186
rect 3381 5166 3397 5186
rect 3355 5158 3397 5166
rect 3425 5186 3466 5188
rect 3425 5166 3439 5186
rect 3458 5166 3466 5186
rect 3425 5158 3466 5166
rect 2549 5157 2851 5158
rect 1468 5136 1578 5150
rect 1468 5133 1511 5136
rect 1468 5128 1472 5133
rect 1034 5079 1202 5081
rect 758 5076 1202 5079
rect 419 5052 530 5058
rect 419 5044 460 5052
rect 108 4989 147 5033
rect 419 5024 427 5044
rect 446 5024 460 5044
rect 419 5022 460 5024
rect 488 5044 530 5052
rect 488 5024 504 5044
rect 523 5024 530 5044
rect 488 5023 530 5024
rect 756 5053 1202 5076
rect 488 5022 531 5023
rect 419 5003 531 5022
rect 108 4965 148 4989
rect 448 4965 495 4966
rect 756 4965 794 5053
rect 1034 5052 1202 5053
rect 1390 5106 1472 5128
rect 1501 5106 1511 5133
rect 1539 5109 1546 5136
rect 1575 5128 1578 5136
rect 2549 5131 3127 5157
rect 3355 5152 3466 5158
rect 2549 5129 2851 5131
rect 2549 5128 2735 5129
rect 1575 5109 1640 5128
rect 1539 5106 1640 5109
rect 1390 5104 1640 5106
rect 1390 5025 1427 5104
rect 1468 5091 1578 5104
rect 1542 5035 1573 5036
rect 1390 5005 1399 5025
rect 1419 5005 1427 5025
rect 1390 4995 1427 5005
rect 1486 5025 1573 5035
rect 1486 5005 1495 5025
rect 1515 5005 1573 5025
rect 1486 4996 1573 5005
rect 1486 4995 1523 4996
rect 108 4955 794 4965
rect 104 4932 794 4955
rect 1542 4943 1573 4996
rect 1603 5025 1640 5104
rect 1811 5101 2204 5121
rect 2224 5101 2227 5121
rect 2549 5120 2602 5128
rect 1811 5096 2227 5101
rect 1811 5095 2152 5096
rect 1755 5035 1786 5036
rect 1603 5005 1612 5025
rect 1632 5005 1640 5025
rect 1603 4995 1640 5005
rect 1699 5028 1786 5035
rect 1699 5025 1760 5028
rect 1699 5005 1708 5025
rect 1728 5008 1760 5025
rect 1781 5008 1786 5028
rect 1728 5005 1786 5008
rect 1699 4998 1786 5005
rect 1811 5025 1848 5095
rect 2114 5094 2151 5095
rect 1963 5035 1999 5036
rect 1811 5005 1820 5025
rect 1840 5005 1848 5025
rect 1699 4996 1755 4998
rect 1699 4995 1736 4996
rect 1811 4995 1848 5005
rect 1907 5025 2055 5035
rect 2155 5032 2251 5034
rect 1907 5005 1916 5025
rect 1936 5005 2026 5025
rect 2046 5005 2055 5025
rect 1907 4996 2055 5005
rect 2113 5025 2251 5032
rect 2113 5005 2122 5025
rect 2142 5005 2251 5025
rect 2113 4996 2251 5005
rect 1907 4995 1944 4996
rect 1963 4944 1999 4996
rect 2018 4995 2055 4996
rect 2114 4995 2151 4996
rect 1434 4942 1475 4943
rect 104 4913 146 4932
rect 756 4930 794 4932
rect 1326 4935 1475 4942
rect 107 4875 146 4913
rect 1326 4915 1444 4935
rect 1464 4915 1475 4935
rect 1326 4907 1475 4915
rect 1542 4939 1901 4943
rect 1542 4934 1864 4939
rect 1542 4910 1655 4934
rect 1679 4915 1864 4934
rect 1888 4915 1901 4939
rect 1679 4910 1901 4915
rect 1542 4907 1901 4910
rect 1963 4907 1998 4944
rect 2066 4941 2166 4944
rect 2066 4937 2133 4941
rect 2066 4911 2078 4937
rect 2104 4915 2133 4937
rect 2159 4915 2166 4941
rect 2104 4911 2166 4915
rect 2066 4907 2166 4911
rect 1542 4886 1573 4907
rect 1963 4886 1999 4907
rect 1385 4885 1422 4886
rect 1384 4876 1422 4885
rect 107 4873 155 4875
rect 107 4855 118 4873
rect 136 4855 155 4873
rect 107 4846 155 4855
rect 108 4845 155 4846
rect 421 4850 531 4864
rect 421 4847 464 4850
rect 421 4842 425 4847
rect 343 4820 425 4842
rect 454 4820 464 4847
rect 492 4823 499 4850
rect 528 4842 531 4850
rect 1384 4856 1393 4876
rect 1413 4856 1422 4876
rect 1384 4848 1422 4856
rect 1488 4880 1573 4886
rect 1598 4885 1635 4886
rect 1488 4860 1496 4880
rect 1516 4860 1573 4880
rect 1488 4852 1573 4860
rect 1597 4876 1635 4885
rect 1597 4856 1606 4876
rect 1626 4856 1635 4876
rect 1488 4851 1524 4852
rect 1597 4848 1635 4856
rect 1701 4880 1786 4886
rect 1806 4885 1843 4886
rect 1701 4860 1709 4880
rect 1729 4879 1786 4880
rect 1729 4860 1758 4879
rect 1701 4859 1758 4860
rect 1779 4859 1786 4879
rect 1701 4852 1786 4859
rect 1805 4876 1843 4885
rect 1805 4856 1814 4876
rect 1834 4856 1843 4876
rect 1701 4851 1737 4852
rect 1805 4848 1843 4856
rect 1909 4882 2053 4886
rect 1909 4880 1966 4882
rect 1909 4860 1917 4880
rect 1937 4860 1966 4880
rect 1909 4858 1966 4860
rect 1992 4880 2053 4882
rect 1992 4860 2025 4880
rect 2045 4860 2053 4880
rect 1992 4858 2053 4860
rect 1909 4852 2053 4858
rect 1909 4851 1945 4852
rect 2017 4851 2053 4852
rect 2119 4885 2156 4886
rect 2119 4884 2157 4885
rect 2119 4876 2183 4884
rect 2119 4856 2128 4876
rect 2148 4862 2183 4876
rect 2203 4862 2206 4882
rect 2148 4857 2206 4862
rect 2148 4856 2183 4857
rect 528 4823 593 4842
rect 492 4820 593 4823
rect 343 4818 593 4820
rect 111 4782 148 4783
rect 107 4779 148 4782
rect 107 4774 149 4779
rect 107 4756 120 4774
rect 138 4756 149 4774
rect 107 4742 149 4756
rect 187 4742 234 4746
rect 107 4736 234 4742
rect 107 4707 195 4736
rect 224 4707 234 4736
rect 343 4739 380 4818
rect 421 4805 531 4818
rect 495 4749 526 4750
rect 343 4719 352 4739
rect 372 4719 380 4739
rect 343 4709 380 4719
rect 439 4739 526 4749
rect 439 4719 448 4739
rect 468 4719 526 4739
rect 439 4710 526 4719
rect 439 4709 476 4710
rect 107 4703 234 4707
rect 107 4686 146 4703
rect 187 4702 234 4703
rect 107 4668 118 4686
rect 136 4668 146 4686
rect 107 4659 146 4668
rect 108 4658 145 4659
rect 495 4657 526 4710
rect 556 4739 593 4818
rect 764 4815 1157 4835
rect 1177 4815 1180 4835
rect 1385 4819 1422 4848
rect 764 4810 1180 4815
rect 1386 4817 1422 4819
rect 1598 4817 1635 4848
rect 764 4809 1105 4810
rect 708 4749 739 4750
rect 556 4719 565 4739
rect 585 4719 593 4739
rect 556 4709 593 4719
rect 652 4742 739 4749
rect 652 4739 713 4742
rect 652 4719 661 4739
rect 681 4722 713 4739
rect 734 4722 739 4742
rect 681 4719 739 4722
rect 652 4712 739 4719
rect 764 4739 801 4809
rect 1067 4808 1104 4809
rect 1386 4795 1635 4817
rect 1806 4816 1843 4848
rect 2119 4844 2183 4856
rect 2223 4819 2250 4996
rect 2683 4951 2710 5128
rect 2750 5091 2814 5103
rect 3090 5099 3127 5131
rect 3298 5130 3547 5152
rect 3829 5138 3866 5139
rect 4132 5138 4169 5208
rect 4194 5228 4281 5235
rect 4194 5225 4252 5228
rect 4194 5205 4199 5225
rect 4220 5208 4252 5225
rect 4272 5208 4281 5228
rect 4220 5205 4281 5208
rect 4194 5198 4281 5205
rect 4340 5228 4377 5238
rect 4340 5208 4348 5228
rect 4368 5208 4377 5228
rect 4194 5197 4225 5198
rect 3828 5137 4169 5138
rect 3298 5099 3335 5130
rect 3511 5128 3547 5130
rect 3753 5132 4169 5137
rect 3511 5099 3548 5128
rect 3753 5112 3756 5132
rect 3776 5112 4169 5132
rect 4340 5129 4377 5208
rect 4407 5237 4438 5290
rect 4788 5288 4825 5289
rect 4787 5279 4826 5288
rect 4787 5261 4797 5279
rect 4815 5261 4826 5279
rect 5167 5277 5204 5281
rect 4699 5244 4746 5245
rect 4787 5244 4826 5261
rect 4699 5240 4826 5244
rect 4457 5237 4494 5238
rect 4407 5228 4494 5237
rect 4407 5208 4465 5228
rect 4485 5208 4494 5228
rect 4407 5198 4494 5208
rect 4553 5228 4590 5238
rect 4553 5208 4561 5228
rect 4581 5208 4590 5228
rect 4407 5197 4438 5198
rect 4402 5129 4512 5142
rect 4553 5129 4590 5208
rect 4699 5211 4709 5240
rect 4738 5211 4826 5240
rect 4699 5205 4826 5211
rect 4699 5201 4746 5205
rect 4784 5191 4826 5205
rect 4784 5173 4795 5191
rect 4813 5173 4826 5191
rect 4784 5168 4826 5173
rect 4785 5165 4826 5168
rect 5164 5272 5204 5277
rect 5164 5254 5176 5272
rect 5194 5254 5204 5272
rect 4785 5164 4822 5165
rect 4340 5127 4590 5129
rect 4340 5124 4441 5127
rect 4340 5105 4405 5124
rect 2750 5090 2785 5091
rect 2727 5085 2785 5090
rect 2727 5065 2730 5085
rect 2750 5071 2785 5085
rect 2805 5071 2814 5091
rect 2750 5063 2814 5071
rect 2776 5062 2814 5063
rect 2777 5061 2814 5062
rect 2880 5095 2916 5096
rect 2988 5095 3024 5096
rect 2880 5088 3024 5095
rect 2880 5087 2937 5088
rect 2880 5067 2888 5087
rect 2908 5068 2937 5087
rect 2962 5087 3024 5088
rect 2962 5068 2996 5087
rect 2908 5067 2996 5068
rect 3016 5067 3024 5087
rect 2880 5061 3024 5067
rect 3090 5091 3128 5099
rect 3196 5095 3232 5096
rect 3090 5071 3099 5091
rect 3119 5071 3128 5091
rect 3090 5062 3128 5071
rect 3147 5088 3232 5095
rect 3147 5068 3154 5088
rect 3175 5087 3232 5088
rect 3175 5068 3204 5087
rect 3147 5067 3204 5068
rect 3224 5067 3232 5087
rect 3090 5061 3127 5062
rect 3147 5061 3232 5067
rect 3298 5091 3336 5099
rect 3409 5095 3445 5096
rect 3298 5071 3307 5091
rect 3327 5071 3336 5091
rect 3298 5062 3336 5071
rect 3360 5087 3445 5095
rect 3360 5067 3417 5087
rect 3437 5067 3445 5087
rect 3298 5061 3335 5062
rect 3360 5061 3445 5067
rect 3511 5091 3549 5099
rect 3511 5071 3520 5091
rect 3540 5071 3549 5091
rect 4402 5097 4405 5105
rect 4434 5097 4441 5124
rect 4469 5100 4479 5127
rect 4508 5105 4590 5127
rect 4508 5100 4512 5105
rect 4469 5097 4512 5100
rect 4402 5083 4512 5097
rect 4778 5101 4825 5102
rect 4778 5092 4826 5101
rect 4778 5074 4797 5092
rect 4815 5074 4826 5092
rect 4778 5072 4826 5074
rect 3511 5062 3549 5071
rect 3511 5061 3548 5062
rect 2934 5040 2970 5061
rect 3360 5040 3391 5061
rect 2767 5036 2867 5040
rect 2767 5032 2829 5036
rect 2767 5006 2774 5032
rect 2800 5010 2829 5032
rect 2855 5010 2867 5036
rect 2800 5006 2867 5010
rect 2767 5003 2867 5006
rect 2935 5003 2970 5040
rect 3032 5037 3391 5040
rect 3032 5032 3254 5037
rect 3032 5008 3045 5032
rect 3069 5013 3254 5032
rect 3278 5013 3391 5037
rect 3069 5008 3391 5013
rect 3032 5004 3391 5008
rect 3458 5032 3607 5040
rect 3458 5012 3469 5032
rect 3489 5012 3607 5032
rect 4787 5034 4826 5072
rect 5164 5074 5204 5254
rect 5550 5247 5581 5300
rect 5611 5329 5648 5408
rect 5819 5405 6212 5425
rect 6232 5405 6235 5425
rect 6333 5409 6582 5431
rect 6751 5430 6792 5435
rect 7170 5432 7197 5610
rect 7848 5522 7875 5700
rect 8253 5697 8294 5702
rect 8463 5701 8712 5723
rect 8810 5707 8813 5727
rect 8833 5707 9226 5727
rect 9397 5724 9434 5803
rect 9464 5832 9495 5885
rect 9841 5878 9881 6058
rect 9841 5860 9851 5878
rect 9869 5860 9881 5878
rect 9841 5855 9881 5860
rect 9841 5851 9878 5855
rect 9514 5832 9551 5833
rect 9464 5823 9551 5832
rect 9464 5803 9522 5823
rect 9542 5803 9551 5823
rect 9464 5793 9551 5803
rect 9610 5823 9647 5833
rect 9610 5803 9618 5823
rect 9638 5803 9647 5823
rect 9464 5792 9495 5793
rect 9459 5724 9569 5737
rect 9610 5724 9647 5803
rect 9844 5788 9881 5789
rect 9840 5779 9881 5788
rect 9840 5761 9853 5779
rect 9871 5761 9881 5779
rect 9840 5752 9881 5761
rect 9840 5732 9880 5752
rect 9397 5722 9647 5724
rect 9397 5719 9498 5722
rect 7915 5662 7979 5674
rect 8255 5670 8292 5697
rect 8463 5670 8500 5701
rect 8676 5699 8712 5701
rect 9397 5700 9462 5719
rect 8676 5670 8713 5699
rect 9459 5692 9462 5700
rect 9491 5692 9498 5719
rect 9526 5695 9536 5722
rect 9565 5700 9647 5722
rect 9755 5722 9880 5732
rect 9755 5703 9763 5722
rect 9788 5703 9880 5722
rect 9565 5695 9569 5700
rect 9755 5696 9880 5703
rect 9526 5692 9569 5695
rect 9459 5678 9569 5692
rect 7915 5661 7950 5662
rect 7892 5656 7950 5661
rect 7892 5636 7895 5656
rect 7915 5642 7950 5656
rect 7970 5642 7979 5662
rect 7915 5634 7979 5642
rect 7941 5633 7979 5634
rect 7942 5632 7979 5633
rect 8045 5666 8081 5667
rect 8153 5666 8189 5667
rect 8045 5658 8189 5666
rect 8045 5638 8053 5658
rect 8073 5655 8161 5658
rect 8073 5638 8105 5655
rect 8125 5638 8161 5655
rect 8181 5638 8189 5658
rect 8045 5632 8189 5638
rect 8255 5662 8293 5670
rect 8361 5666 8397 5667
rect 8255 5642 8264 5662
rect 8284 5642 8293 5662
rect 8255 5633 8293 5642
rect 8312 5659 8397 5666
rect 8312 5639 8319 5659
rect 8340 5658 8397 5659
rect 8340 5639 8369 5658
rect 8312 5638 8369 5639
rect 8389 5638 8397 5658
rect 8255 5632 8292 5633
rect 8312 5632 8397 5638
rect 8463 5662 8501 5670
rect 8574 5666 8610 5667
rect 8463 5642 8472 5662
rect 8492 5642 8501 5662
rect 8463 5633 8501 5642
rect 8525 5658 8610 5666
rect 8525 5638 8582 5658
rect 8602 5638 8610 5658
rect 8463 5632 8500 5633
rect 8525 5632 8610 5638
rect 8676 5662 8714 5670
rect 8676 5642 8685 5662
rect 8705 5642 8714 5662
rect 8676 5633 8714 5642
rect 9840 5648 9880 5696
rect 8676 5632 8713 5633
rect 8099 5611 8135 5632
rect 8525 5611 8556 5632
rect 9840 5630 9851 5648
rect 9869 5630 9880 5648
rect 9840 5622 9880 5630
rect 9841 5621 9878 5622
rect 7932 5607 8032 5611
rect 7932 5603 7994 5607
rect 7932 5577 7939 5603
rect 7965 5581 7994 5603
rect 8020 5581 8032 5607
rect 7965 5577 8032 5581
rect 7932 5574 8032 5577
rect 8100 5574 8135 5611
rect 8197 5608 8556 5611
rect 8197 5603 8419 5608
rect 8197 5579 8210 5603
rect 8234 5584 8419 5603
rect 8443 5584 8556 5608
rect 8234 5579 8556 5584
rect 8197 5575 8556 5579
rect 8623 5603 8772 5611
rect 8623 5583 8634 5603
rect 8654 5583 8772 5603
rect 8623 5576 8772 5583
rect 9212 5580 9726 5581
rect 8623 5575 8664 5576
rect 7947 5522 7984 5523
rect 8043 5522 8080 5523
rect 8099 5522 8135 5574
rect 8154 5522 8191 5523
rect 7847 5513 7985 5522
rect 7847 5493 7956 5513
rect 7976 5493 7985 5513
rect 7847 5486 7985 5493
rect 8043 5513 8191 5522
rect 8043 5493 8052 5513
rect 8072 5493 8162 5513
rect 8182 5493 8191 5513
rect 7847 5484 7943 5486
rect 8043 5483 8191 5493
rect 8250 5513 8287 5523
rect 8362 5522 8399 5523
rect 8343 5520 8399 5522
rect 8250 5493 8258 5513
rect 8278 5493 8287 5513
rect 8099 5482 8135 5483
rect 7029 5430 7197 5432
rect 6751 5424 7197 5430
rect 5819 5400 6235 5405
rect 6414 5403 6525 5409
rect 5819 5399 6160 5400
rect 5763 5339 5794 5340
rect 5611 5309 5620 5329
rect 5640 5309 5648 5329
rect 5611 5299 5648 5309
rect 5707 5332 5794 5339
rect 5707 5329 5768 5332
rect 5707 5309 5716 5329
rect 5736 5312 5768 5329
rect 5789 5312 5794 5332
rect 5736 5309 5794 5312
rect 5707 5302 5794 5309
rect 5819 5329 5856 5399
rect 6122 5398 6159 5399
rect 6414 5395 6455 5403
rect 6414 5375 6422 5395
rect 6441 5375 6455 5395
rect 6414 5373 6455 5375
rect 6483 5395 6525 5403
rect 6483 5375 6499 5395
rect 6518 5375 6525 5395
rect 6751 5402 6757 5424
rect 6783 5404 7197 5424
rect 7947 5423 7984 5424
rect 8250 5423 8287 5493
rect 8312 5513 8399 5520
rect 8312 5510 8370 5513
rect 8312 5490 8317 5510
rect 8338 5493 8370 5510
rect 8390 5493 8399 5513
rect 8338 5490 8399 5493
rect 8312 5483 8399 5490
rect 8458 5513 8495 5523
rect 8458 5493 8466 5513
rect 8486 5493 8495 5513
rect 8312 5482 8343 5483
rect 7946 5422 8287 5423
rect 6783 5402 6792 5404
rect 7029 5403 7197 5404
rect 7871 5417 8287 5422
rect 6751 5393 6792 5402
rect 7871 5397 7874 5417
rect 7894 5397 8287 5417
rect 8458 5414 8495 5493
rect 8525 5522 8556 5575
rect 9193 5564 9726 5580
rect 9193 5553 9725 5564
rect 9844 5555 9881 5559
rect 8575 5522 8612 5523
rect 8525 5513 8612 5522
rect 8525 5493 8583 5513
rect 8603 5493 8612 5513
rect 8525 5483 8612 5493
rect 8671 5513 8708 5523
rect 8671 5493 8679 5513
rect 8699 5493 8708 5513
rect 8525 5482 8556 5483
rect 8520 5414 8630 5427
rect 8671 5414 8708 5493
rect 8458 5412 8708 5414
rect 8458 5409 8559 5412
rect 8458 5390 8523 5409
rect 8520 5382 8523 5390
rect 8552 5382 8559 5409
rect 8587 5385 8597 5412
rect 8626 5390 8708 5412
rect 8786 5484 8954 5485
rect 9193 5484 9231 5553
rect 8786 5464 9231 5484
rect 9458 5515 9569 5530
rect 9458 5513 9500 5515
rect 9458 5493 9465 5513
rect 9484 5493 9500 5513
rect 9458 5485 9500 5493
rect 9528 5513 9569 5515
rect 9528 5493 9542 5513
rect 9561 5493 9569 5513
rect 9528 5485 9569 5493
rect 9458 5479 9569 5485
rect 9691 5490 9725 5553
rect 9843 5549 9881 5555
rect 9843 5531 9853 5549
rect 9871 5531 9881 5549
rect 9843 5522 9881 5531
rect 9843 5490 9877 5522
rect 8786 5458 9230 5464
rect 8786 5456 8954 5458
rect 8626 5385 8630 5390
rect 8587 5382 8630 5385
rect 6483 5373 6525 5375
rect 6414 5358 6525 5373
rect 7610 5364 7658 5378
rect 8520 5368 8630 5382
rect 5971 5339 6007 5340
rect 5819 5309 5828 5329
rect 5848 5309 5856 5329
rect 5707 5300 5763 5302
rect 5707 5299 5744 5300
rect 5819 5299 5856 5309
rect 5915 5329 6063 5339
rect 6163 5336 6259 5338
rect 5915 5309 5924 5329
rect 5944 5309 6034 5329
rect 6054 5309 6063 5329
rect 5915 5300 6063 5309
rect 6121 5329 6259 5336
rect 6121 5309 6130 5329
rect 6150 5309 6259 5329
rect 6121 5300 6259 5309
rect 7610 5324 7623 5364
rect 7650 5324 7658 5364
rect 7610 5306 7658 5324
rect 5915 5299 5952 5300
rect 5971 5248 6007 5300
rect 6026 5299 6063 5300
rect 6122 5299 6159 5300
rect 5442 5246 5483 5247
rect 5334 5239 5483 5246
rect 5334 5219 5452 5239
rect 5472 5219 5483 5239
rect 5334 5211 5483 5219
rect 5550 5243 5909 5247
rect 5550 5238 5872 5243
rect 5550 5214 5663 5238
rect 5687 5219 5872 5238
rect 5896 5219 5909 5243
rect 5687 5214 5909 5219
rect 5550 5211 5909 5214
rect 5971 5211 6006 5248
rect 6074 5245 6174 5248
rect 6074 5241 6141 5245
rect 6074 5215 6086 5241
rect 6112 5219 6141 5241
rect 6167 5219 6174 5245
rect 6112 5215 6174 5219
rect 6074 5211 6174 5215
rect 5550 5190 5581 5211
rect 5971 5190 6007 5211
rect 5393 5189 5430 5190
rect 5392 5180 5430 5189
rect 5392 5160 5401 5180
rect 5421 5160 5430 5180
rect 5392 5152 5430 5160
rect 5496 5184 5581 5190
rect 5606 5189 5643 5190
rect 5496 5164 5504 5184
rect 5524 5164 5581 5184
rect 5496 5156 5581 5164
rect 5605 5180 5643 5189
rect 5605 5160 5614 5180
rect 5634 5160 5643 5180
rect 5496 5155 5532 5156
rect 5605 5152 5643 5160
rect 5709 5184 5794 5190
rect 5814 5189 5851 5190
rect 5709 5164 5717 5184
rect 5737 5183 5794 5184
rect 5737 5164 5766 5183
rect 5709 5163 5766 5164
rect 5787 5163 5794 5183
rect 5709 5156 5794 5163
rect 5813 5180 5851 5189
rect 5813 5160 5822 5180
rect 5842 5160 5851 5180
rect 5709 5155 5745 5156
rect 5813 5152 5851 5160
rect 5917 5184 6061 5190
rect 5917 5164 5925 5184
rect 5945 5181 6033 5184
rect 5945 5164 5976 5181
rect 5917 5161 5976 5164
rect 5999 5164 6033 5181
rect 6053 5164 6061 5184
rect 5999 5161 6061 5164
rect 5917 5156 6061 5161
rect 5917 5155 5953 5156
rect 6025 5155 6061 5156
rect 6127 5189 6164 5190
rect 6127 5188 6165 5189
rect 6127 5180 6191 5188
rect 6127 5160 6136 5180
rect 6156 5166 6191 5180
rect 6211 5166 6214 5186
rect 6156 5161 6214 5166
rect 6156 5160 6191 5161
rect 5393 5123 5430 5152
rect 5394 5121 5430 5123
rect 5606 5121 5643 5152
rect 5394 5099 5643 5121
rect 5814 5120 5851 5152
rect 6127 5148 6191 5160
rect 6231 5122 6258 5300
rect 7605 5199 7658 5306
rect 8786 5278 8813 5456
rect 8853 5418 8917 5430
rect 9193 5426 9230 5458
rect 9401 5457 9650 5479
rect 9691 5458 9877 5490
rect 9705 5457 9877 5458
rect 9401 5426 9438 5457
rect 9614 5455 9650 5457
rect 9614 5426 9651 5455
rect 9843 5429 9877 5457
rect 8853 5417 8888 5418
rect 8830 5412 8888 5417
rect 8830 5392 8833 5412
rect 8853 5398 8888 5412
rect 8908 5398 8917 5418
rect 8853 5390 8917 5398
rect 8879 5389 8917 5390
rect 8880 5388 8917 5389
rect 8983 5422 9019 5423
rect 9091 5422 9127 5423
rect 8983 5415 9127 5422
rect 8983 5414 9043 5415
rect 8983 5394 8991 5414
rect 9011 5395 9043 5414
rect 9068 5414 9127 5415
rect 9068 5395 9099 5414
rect 9011 5394 9099 5395
rect 9119 5394 9127 5414
rect 8983 5388 9127 5394
rect 9193 5418 9231 5426
rect 9299 5422 9335 5423
rect 9193 5398 9202 5418
rect 9222 5398 9231 5418
rect 9193 5389 9231 5398
rect 9250 5415 9335 5422
rect 9250 5395 9257 5415
rect 9278 5414 9335 5415
rect 9278 5395 9307 5414
rect 9250 5394 9307 5395
rect 9327 5394 9335 5414
rect 9193 5388 9230 5389
rect 9250 5388 9335 5394
rect 9401 5418 9439 5426
rect 9512 5422 9548 5423
rect 9401 5398 9410 5418
rect 9430 5398 9439 5418
rect 9401 5389 9439 5398
rect 9463 5414 9548 5422
rect 9463 5394 9520 5414
rect 9540 5394 9548 5414
rect 9401 5388 9438 5389
rect 9463 5388 9548 5394
rect 9614 5418 9652 5426
rect 9614 5398 9623 5418
rect 9643 5398 9652 5418
rect 9614 5389 9652 5398
rect 9841 5419 9878 5429
rect 9841 5401 9851 5419
rect 9869 5401 9878 5419
rect 9841 5392 9878 5401
rect 9843 5391 9877 5392
rect 9614 5388 9651 5389
rect 9037 5367 9073 5388
rect 9463 5367 9494 5388
rect 8870 5363 8970 5367
rect 8870 5359 8932 5363
rect 8870 5333 8877 5359
rect 8903 5337 8932 5359
rect 8958 5337 8970 5363
rect 8903 5333 8970 5337
rect 8870 5330 8970 5333
rect 9038 5330 9073 5367
rect 9135 5364 9494 5367
rect 9135 5359 9357 5364
rect 9135 5335 9148 5359
rect 9172 5340 9357 5359
rect 9381 5340 9494 5364
rect 9172 5335 9494 5340
rect 9135 5331 9494 5335
rect 9561 5359 9710 5367
rect 9561 5339 9572 5359
rect 9592 5339 9710 5359
rect 9561 5332 9710 5339
rect 9561 5331 9602 5332
rect 8885 5278 8922 5279
rect 8981 5278 9018 5279
rect 9037 5278 9073 5330
rect 9092 5278 9129 5279
rect 8785 5269 8923 5278
rect 8785 5249 8894 5269
rect 8914 5249 8923 5269
rect 8411 5229 8522 5244
rect 8785 5242 8923 5249
rect 8981 5269 9129 5278
rect 8981 5249 8990 5269
rect 9010 5249 9100 5269
rect 9120 5249 9129 5269
rect 8785 5240 8881 5242
rect 8981 5239 9129 5249
rect 9188 5269 9225 5279
rect 9300 5278 9337 5279
rect 9281 5276 9337 5278
rect 9188 5249 9196 5269
rect 9216 5249 9225 5269
rect 9037 5238 9073 5239
rect 8411 5227 8453 5229
rect 8411 5207 8418 5227
rect 8437 5207 8453 5227
rect 8411 5199 8453 5207
rect 8481 5227 8522 5229
rect 8481 5207 8495 5227
rect 8514 5207 8522 5227
rect 8481 5199 8522 5207
rect 7605 5198 7907 5199
rect 6524 5177 6634 5191
rect 6524 5174 6567 5177
rect 6524 5169 6528 5174
rect 6090 5120 6258 5122
rect 5814 5117 6258 5120
rect 5475 5093 5586 5099
rect 5475 5085 5516 5093
rect 3458 5005 3607 5012
rect 4139 5015 4177 5017
rect 4787 5015 4829 5034
rect 3458 5004 3499 5005
rect 2934 4999 2970 5003
rect 2934 4970 2971 4999
rect 2782 4951 2819 4952
rect 2878 4951 2915 4952
rect 2934 4951 2970 4970
rect 2989 4951 3026 4952
rect 2682 4942 2820 4951
rect 2682 4922 2791 4942
rect 2811 4922 2820 4942
rect 2682 4915 2820 4922
rect 2878 4942 3026 4951
rect 2878 4922 2887 4942
rect 2907 4922 2997 4942
rect 3017 4922 3026 4942
rect 2682 4913 2778 4915
rect 2878 4912 3026 4922
rect 3085 4942 3122 4952
rect 3197 4951 3234 4952
rect 3178 4949 3234 4951
rect 3085 4922 3093 4942
rect 3113 4922 3122 4942
rect 2934 4911 2970 4912
rect 2782 4852 2819 4853
rect 3085 4852 3122 4922
rect 3147 4942 3234 4949
rect 3147 4939 3205 4942
rect 3147 4919 3152 4939
rect 3173 4922 3205 4939
rect 3225 4922 3234 4942
rect 3173 4919 3234 4922
rect 3147 4912 3234 4919
rect 3293 4942 3330 4952
rect 3293 4922 3301 4942
rect 3321 4922 3330 4942
rect 3147 4911 3178 4912
rect 2781 4851 3122 4852
rect 2706 4846 3122 4851
rect 2331 4819 2384 4827
rect 2706 4826 2709 4846
rect 2729 4826 3122 4846
rect 3293 4843 3330 4922
rect 3360 4951 3391 5004
rect 4139 4992 4829 5015
rect 5164 5030 5203 5074
rect 5475 5065 5483 5085
rect 5502 5065 5516 5085
rect 5475 5063 5516 5065
rect 5544 5085 5586 5093
rect 5544 5065 5560 5085
rect 5579 5065 5586 5085
rect 5544 5064 5586 5065
rect 5812 5094 6258 5117
rect 5544 5063 5587 5064
rect 5475 5044 5587 5063
rect 5164 5006 5204 5030
rect 5504 5006 5551 5007
rect 5812 5006 5850 5094
rect 6090 5093 6258 5094
rect 6446 5147 6528 5169
rect 6557 5147 6567 5174
rect 6595 5150 6602 5177
rect 6631 5169 6634 5177
rect 7605 5172 8183 5198
rect 8411 5193 8522 5199
rect 7605 5170 7907 5172
rect 7605 5169 7791 5170
rect 6631 5150 6696 5169
rect 6595 5147 6696 5150
rect 6446 5145 6696 5147
rect 6446 5066 6483 5145
rect 6524 5132 6634 5145
rect 6598 5076 6629 5077
rect 6446 5046 6455 5066
rect 6475 5046 6483 5066
rect 6446 5036 6483 5046
rect 6542 5066 6629 5076
rect 6542 5046 6551 5066
rect 6571 5046 6629 5066
rect 6542 5037 6629 5046
rect 6542 5036 6579 5037
rect 5164 4996 5850 5006
rect 4139 4982 4825 4992
rect 3410 4951 3447 4952
rect 3360 4942 3447 4951
rect 3360 4922 3418 4942
rect 3438 4922 3447 4942
rect 3360 4912 3447 4922
rect 3506 4942 3543 4952
rect 3506 4922 3514 4942
rect 3534 4922 3543 4942
rect 3360 4911 3391 4912
rect 3355 4843 3465 4856
rect 3506 4843 3543 4922
rect 3293 4841 3543 4843
rect 3293 4838 3394 4841
rect 3293 4819 3358 4838
rect 2198 4818 2384 4819
rect 2082 4816 2384 4818
rect 1467 4789 1578 4795
rect 1806 4790 2384 4816
rect 3355 4811 3358 4819
rect 3387 4811 3394 4838
rect 3422 4814 3432 4841
rect 3461 4819 3543 4841
rect 3731 4894 3899 4895
rect 4139 4894 4177 4982
rect 4438 4981 4485 4982
rect 4785 4958 4825 4982
rect 4402 4925 4514 4944
rect 4402 4924 4445 4925
rect 3731 4871 4177 4894
rect 4403 4923 4445 4924
rect 4403 4903 4410 4923
rect 4429 4903 4445 4923
rect 4403 4895 4445 4903
rect 4473 4923 4514 4925
rect 4473 4903 4487 4923
rect 4506 4903 4514 4923
rect 4786 4914 4825 4958
rect 5160 4973 5850 4996
rect 6598 4984 6629 5037
rect 6659 5066 6696 5145
rect 6867 5142 7260 5162
rect 7280 5142 7283 5162
rect 7605 5161 7658 5169
rect 6867 5137 7283 5142
rect 6867 5136 7208 5137
rect 6811 5076 6842 5077
rect 6659 5046 6668 5066
rect 6688 5046 6696 5066
rect 6659 5036 6696 5046
rect 6755 5069 6842 5076
rect 6755 5066 6816 5069
rect 6755 5046 6764 5066
rect 6784 5049 6816 5066
rect 6837 5049 6842 5069
rect 6784 5046 6842 5049
rect 6755 5039 6842 5046
rect 6867 5066 6904 5136
rect 7170 5135 7207 5136
rect 7019 5076 7055 5077
rect 6867 5046 6876 5066
rect 6896 5046 6904 5066
rect 6755 5037 6811 5039
rect 6755 5036 6792 5037
rect 6867 5036 6904 5046
rect 6963 5066 7111 5076
rect 7211 5073 7307 5075
rect 6963 5046 6972 5066
rect 6992 5046 7082 5066
rect 7102 5046 7111 5066
rect 6963 5037 7111 5046
rect 7169 5066 7307 5073
rect 7169 5046 7178 5066
rect 7198 5046 7307 5066
rect 7169 5037 7307 5046
rect 6963 5036 7000 5037
rect 7019 4985 7055 5037
rect 7074 5036 7111 5037
rect 7170 5036 7207 5037
rect 6490 4983 6531 4984
rect 5160 4954 5202 4973
rect 5812 4971 5850 4973
rect 6382 4976 6531 4983
rect 4473 4895 4514 4903
rect 4403 4889 4514 4895
rect 3731 4868 4175 4871
rect 3731 4866 3899 4868
rect 3461 4814 3465 4819
rect 3422 4811 3465 4814
rect 3355 4797 3465 4811
rect 2082 4789 2384 4790
rect 1467 4781 1508 4789
rect 1467 4761 1475 4781
rect 1494 4761 1508 4781
rect 1467 4759 1508 4761
rect 1536 4781 1578 4789
rect 1536 4761 1552 4781
rect 1571 4761 1578 4781
rect 1536 4759 1578 4761
rect 916 4749 952 4750
rect 764 4719 773 4739
rect 793 4719 801 4739
rect 652 4710 708 4712
rect 652 4709 689 4710
rect 764 4709 801 4719
rect 860 4739 1008 4749
rect 1108 4746 1204 4748
rect 860 4719 869 4739
rect 889 4719 979 4739
rect 999 4719 1008 4739
rect 860 4710 1008 4719
rect 1066 4739 1204 4746
rect 1467 4744 1578 4759
rect 1066 4719 1075 4739
rect 1095 4719 1204 4739
rect 1066 4710 1204 4719
rect 860 4709 897 4710
rect 916 4658 952 4710
rect 971 4709 1008 4710
rect 1067 4709 1104 4710
rect 387 4656 428 4657
rect 279 4649 428 4656
rect 279 4629 397 4649
rect 417 4629 428 4649
rect 279 4621 428 4629
rect 495 4653 854 4657
rect 495 4648 817 4653
rect 495 4624 608 4648
rect 632 4629 817 4648
rect 841 4629 854 4653
rect 632 4624 854 4629
rect 495 4621 854 4624
rect 916 4621 951 4658
rect 1019 4655 1119 4658
rect 1019 4651 1086 4655
rect 1019 4625 1031 4651
rect 1057 4629 1086 4651
rect 1112 4629 1119 4655
rect 1057 4625 1119 4629
rect 1019 4621 1119 4625
rect 495 4600 526 4621
rect 916 4600 952 4621
rect 338 4599 375 4600
rect 112 4596 146 4597
rect 111 4587 148 4596
rect 111 4569 120 4587
rect 138 4569 148 4587
rect 111 4559 148 4569
rect 337 4590 375 4599
rect 337 4570 346 4590
rect 366 4570 375 4590
rect 337 4562 375 4570
rect 441 4594 526 4600
rect 551 4599 588 4600
rect 441 4574 449 4594
rect 469 4574 526 4594
rect 441 4566 526 4574
rect 550 4590 588 4599
rect 550 4570 559 4590
rect 579 4570 588 4590
rect 441 4565 477 4566
rect 550 4562 588 4570
rect 654 4594 739 4600
rect 759 4599 796 4600
rect 654 4574 662 4594
rect 682 4593 739 4594
rect 682 4574 711 4593
rect 654 4573 711 4574
rect 732 4573 739 4593
rect 654 4566 739 4573
rect 758 4590 796 4599
rect 758 4570 767 4590
rect 787 4570 796 4590
rect 654 4565 690 4566
rect 758 4562 796 4570
rect 862 4594 1006 4600
rect 862 4574 870 4594
rect 890 4593 978 4594
rect 890 4574 921 4593
rect 862 4573 921 4574
rect 946 4574 978 4593
rect 998 4574 1006 4594
rect 946 4573 1006 4574
rect 862 4566 1006 4573
rect 862 4565 898 4566
rect 970 4565 1006 4566
rect 1072 4599 1109 4600
rect 1072 4598 1110 4599
rect 1072 4590 1136 4598
rect 1072 4570 1081 4590
rect 1101 4576 1136 4590
rect 1156 4576 1159 4596
rect 1101 4571 1159 4576
rect 1101 4570 1136 4571
rect 112 4531 146 4559
rect 338 4533 375 4562
rect 339 4531 375 4533
rect 551 4531 588 4562
rect 112 4530 284 4531
rect 112 4498 298 4530
rect 339 4509 588 4531
rect 759 4530 796 4562
rect 1072 4558 1136 4570
rect 1176 4532 1203 4710
rect 2331 4682 2384 4789
rect 3731 4688 3758 4866
rect 3798 4828 3862 4840
rect 4138 4836 4175 4868
rect 4346 4867 4595 4889
rect 4346 4836 4383 4867
rect 4559 4865 4595 4867
rect 4559 4836 4596 4865
rect 3798 4827 3833 4828
rect 3775 4822 3833 4827
rect 3775 4802 3778 4822
rect 3798 4808 3833 4822
rect 3853 4808 3862 4828
rect 3798 4800 3862 4808
rect 3824 4799 3862 4800
rect 3825 4798 3862 4799
rect 3928 4832 3964 4833
rect 4036 4832 4072 4833
rect 3928 4827 4072 4832
rect 3928 4824 3990 4827
rect 3928 4804 3936 4824
rect 3956 4807 3990 4824
rect 4013 4824 4072 4827
rect 4013 4807 4044 4824
rect 3956 4804 4044 4807
rect 4064 4804 4072 4824
rect 3928 4798 4072 4804
rect 4138 4828 4176 4836
rect 4244 4832 4280 4833
rect 4138 4808 4147 4828
rect 4167 4808 4176 4828
rect 4138 4799 4176 4808
rect 4195 4825 4280 4832
rect 4195 4805 4202 4825
rect 4223 4824 4280 4825
rect 4223 4805 4252 4824
rect 4195 4804 4252 4805
rect 4272 4804 4280 4824
rect 4138 4798 4175 4799
rect 4195 4798 4280 4804
rect 4346 4828 4384 4836
rect 4457 4832 4493 4833
rect 4346 4808 4355 4828
rect 4375 4808 4384 4828
rect 4346 4799 4384 4808
rect 4408 4824 4493 4832
rect 4408 4804 4465 4824
rect 4485 4804 4493 4824
rect 4346 4798 4383 4799
rect 4408 4798 4493 4804
rect 4559 4828 4597 4836
rect 4559 4808 4568 4828
rect 4588 4808 4597 4828
rect 4559 4799 4597 4808
rect 4559 4798 4596 4799
rect 3982 4777 4018 4798
rect 4408 4777 4439 4798
rect 3815 4773 3915 4777
rect 3815 4769 3877 4773
rect 3815 4743 3822 4769
rect 3848 4747 3877 4769
rect 3903 4747 3915 4773
rect 3848 4743 3915 4747
rect 3815 4740 3915 4743
rect 3983 4740 4018 4777
rect 4080 4774 4439 4777
rect 4080 4769 4302 4774
rect 4080 4745 4093 4769
rect 4117 4750 4302 4769
rect 4326 4750 4439 4774
rect 4117 4745 4439 4750
rect 4080 4741 4439 4745
rect 4506 4769 4655 4777
rect 4506 4749 4517 4769
rect 4537 4749 4655 4769
rect 4506 4742 4655 4749
rect 4506 4741 4547 4742
rect 3830 4688 3867 4689
rect 3926 4688 3963 4689
rect 3982 4688 4018 4740
rect 4037 4688 4074 4689
rect 2331 4664 2379 4682
rect 2331 4624 2339 4664
rect 2366 4624 2379 4664
rect 3730 4679 3868 4688
rect 3730 4659 3839 4679
rect 3859 4659 3868 4679
rect 3730 4652 3868 4659
rect 3926 4679 4074 4688
rect 3926 4659 3935 4679
rect 3955 4659 4045 4679
rect 4065 4659 4074 4679
rect 3730 4650 3826 4652
rect 3926 4649 4074 4659
rect 4133 4679 4170 4689
rect 4245 4688 4282 4689
rect 4226 4686 4282 4688
rect 4133 4659 4141 4679
rect 4161 4659 4170 4679
rect 3982 4648 4018 4649
rect 1359 4606 1469 4620
rect 2331 4610 2379 4624
rect 3464 4615 3575 4630
rect 3464 4613 3506 4615
rect 1359 4603 1402 4606
rect 1359 4598 1363 4603
rect 1035 4530 1203 4532
rect 759 4524 1203 4530
rect 112 4466 146 4498
rect 108 4457 146 4466
rect 108 4439 118 4457
rect 136 4439 146 4457
rect 108 4433 146 4439
rect 264 4435 298 4498
rect 420 4503 531 4509
rect 420 4495 461 4503
rect 420 4475 428 4495
rect 447 4475 461 4495
rect 420 4473 461 4475
rect 489 4495 531 4503
rect 489 4475 505 4495
rect 524 4475 531 4495
rect 489 4473 531 4475
rect 420 4458 531 4473
rect 758 4504 1203 4524
rect 758 4435 796 4504
rect 1035 4503 1203 4504
rect 1281 4576 1363 4598
rect 1392 4576 1402 4603
rect 1430 4579 1437 4606
rect 1466 4598 1469 4606
rect 1466 4579 1531 4598
rect 1430 4576 1531 4579
rect 1281 4574 1531 4576
rect 1281 4495 1318 4574
rect 1359 4561 1469 4574
rect 1433 4505 1464 4506
rect 1281 4475 1290 4495
rect 1310 4475 1318 4495
rect 1281 4465 1318 4475
rect 1377 4495 1464 4505
rect 1377 4475 1386 4495
rect 1406 4475 1464 4495
rect 1377 4466 1464 4475
rect 1377 4465 1414 4466
rect 108 4429 145 4433
rect 264 4424 796 4435
rect 263 4408 796 4424
rect 1433 4413 1464 4466
rect 1494 4495 1531 4574
rect 1702 4571 2095 4591
rect 2115 4571 2118 4591
rect 3197 4586 3238 4595
rect 1702 4566 2118 4571
rect 2792 4584 2960 4585
rect 3197 4584 3206 4586
rect 1702 4565 2043 4566
rect 1646 4505 1677 4506
rect 1494 4475 1503 4495
rect 1523 4475 1531 4495
rect 1494 4465 1531 4475
rect 1590 4498 1677 4505
rect 1590 4495 1651 4498
rect 1590 4475 1599 4495
rect 1619 4478 1651 4495
rect 1672 4478 1677 4498
rect 1619 4475 1677 4478
rect 1590 4468 1677 4475
rect 1702 4495 1739 4565
rect 2005 4564 2042 4565
rect 2792 4564 3206 4584
rect 3232 4564 3238 4586
rect 3464 4593 3471 4613
rect 3490 4593 3506 4613
rect 3464 4585 3506 4593
rect 3534 4613 3575 4615
rect 3534 4593 3548 4613
rect 3567 4593 3575 4613
rect 3534 4585 3575 4593
rect 3830 4589 3867 4590
rect 4133 4589 4170 4659
rect 4195 4679 4282 4686
rect 4195 4676 4253 4679
rect 4195 4656 4200 4676
rect 4221 4659 4253 4676
rect 4273 4659 4282 4679
rect 4221 4656 4282 4659
rect 4195 4649 4282 4656
rect 4341 4679 4378 4689
rect 4341 4659 4349 4679
rect 4369 4659 4378 4679
rect 4195 4648 4226 4649
rect 3829 4588 4170 4589
rect 3464 4579 3575 4585
rect 3754 4583 4170 4588
rect 2792 4558 3238 4564
rect 2792 4556 2960 4558
rect 1854 4505 1890 4506
rect 1702 4475 1711 4495
rect 1731 4475 1739 4495
rect 1590 4466 1646 4468
rect 1590 4465 1627 4466
rect 1702 4465 1739 4475
rect 1798 4495 1946 4505
rect 2046 4502 2142 4504
rect 1798 4475 1807 4495
rect 1827 4475 1917 4495
rect 1937 4475 1946 4495
rect 1798 4466 1946 4475
rect 2004 4495 2142 4502
rect 2004 4475 2013 4495
rect 2033 4475 2142 4495
rect 2004 4466 2142 4475
rect 1798 4465 1835 4466
rect 1854 4414 1890 4466
rect 1909 4465 1946 4466
rect 2005 4465 2042 4466
rect 1325 4412 1366 4413
rect 263 4407 777 4408
rect 1217 4405 1366 4412
rect 1217 4385 1335 4405
rect 1355 4385 1366 4405
rect 1217 4377 1366 4385
rect 1433 4409 1792 4413
rect 1433 4404 1755 4409
rect 1433 4380 1546 4404
rect 1570 4385 1755 4404
rect 1779 4385 1792 4409
rect 1570 4380 1792 4385
rect 1433 4377 1792 4380
rect 1854 4377 1889 4414
rect 1957 4411 2057 4414
rect 1957 4407 2024 4411
rect 1957 4381 1969 4407
rect 1995 4385 2024 4407
rect 2050 4385 2057 4411
rect 1995 4381 2057 4385
rect 1957 4377 2057 4381
rect 111 4366 148 4367
rect 109 4358 149 4366
rect 109 4340 120 4358
rect 138 4340 149 4358
rect 1433 4356 1464 4377
rect 1854 4356 1890 4377
rect 1276 4355 1313 4356
rect 109 4292 149 4340
rect 1275 4346 1313 4355
rect 1275 4326 1284 4346
rect 1304 4326 1313 4346
rect 1275 4318 1313 4326
rect 1379 4350 1464 4356
rect 1489 4355 1526 4356
rect 1379 4330 1387 4350
rect 1407 4330 1464 4350
rect 1379 4322 1464 4330
rect 1488 4346 1526 4355
rect 1488 4326 1497 4346
rect 1517 4326 1526 4346
rect 1379 4321 1415 4322
rect 1488 4318 1526 4326
rect 1592 4350 1677 4356
rect 1697 4355 1734 4356
rect 1592 4330 1600 4350
rect 1620 4349 1677 4350
rect 1620 4330 1649 4349
rect 1592 4329 1649 4330
rect 1670 4329 1677 4349
rect 1592 4322 1677 4329
rect 1696 4346 1734 4355
rect 1696 4326 1705 4346
rect 1725 4326 1734 4346
rect 1592 4321 1628 4322
rect 1696 4318 1734 4326
rect 1800 4350 1944 4356
rect 1800 4330 1808 4350
rect 1828 4333 1864 4350
rect 1884 4333 1916 4350
rect 1828 4330 1916 4333
rect 1936 4330 1944 4350
rect 1800 4322 1944 4330
rect 1800 4321 1836 4322
rect 1908 4321 1944 4322
rect 2010 4355 2047 4356
rect 2010 4354 2048 4355
rect 2010 4346 2074 4354
rect 2010 4326 2019 4346
rect 2039 4332 2074 4346
rect 2094 4332 2097 4352
rect 2039 4327 2097 4332
rect 2039 4326 2074 4327
rect 420 4296 530 4310
rect 420 4293 463 4296
rect 109 4285 234 4292
rect 420 4288 424 4293
rect 109 4266 201 4285
rect 226 4266 234 4285
rect 109 4256 234 4266
rect 342 4266 424 4288
rect 453 4266 463 4293
rect 491 4269 498 4296
rect 527 4288 530 4296
rect 1276 4289 1313 4318
rect 527 4269 592 4288
rect 1277 4287 1313 4289
rect 1489 4287 1526 4318
rect 1697 4291 1734 4318
rect 2010 4314 2074 4326
rect 491 4266 592 4269
rect 342 4264 592 4266
rect 109 4236 149 4256
rect 108 4227 149 4236
rect 108 4209 118 4227
rect 136 4209 149 4227
rect 108 4200 149 4209
rect 108 4199 145 4200
rect 342 4185 379 4264
rect 420 4251 530 4264
rect 494 4195 525 4196
rect 342 4165 351 4185
rect 371 4165 379 4185
rect 342 4155 379 4165
rect 438 4185 525 4195
rect 438 4165 447 4185
rect 467 4165 525 4185
rect 438 4156 525 4165
rect 438 4155 475 4156
rect 111 4133 148 4137
rect 108 4128 148 4133
rect 108 4110 120 4128
rect 138 4110 148 4128
rect 108 3930 148 4110
rect 494 4103 525 4156
rect 555 4185 592 4264
rect 763 4261 1156 4281
rect 1176 4261 1179 4281
rect 1277 4265 1526 4287
rect 1695 4286 1736 4291
rect 2114 4288 2141 4466
rect 2792 4378 2819 4556
rect 3197 4553 3238 4558
rect 3407 4557 3656 4579
rect 3754 4563 3757 4583
rect 3777 4563 4170 4583
rect 4341 4580 4378 4659
rect 4408 4688 4439 4741
rect 4785 4734 4825 4914
rect 5163 4916 5202 4954
rect 6382 4956 6500 4976
rect 6520 4956 6531 4976
rect 6382 4948 6531 4956
rect 6598 4980 6957 4984
rect 6598 4975 6920 4980
rect 6598 4951 6711 4975
rect 6735 4956 6920 4975
rect 6944 4956 6957 4980
rect 6735 4951 6957 4956
rect 6598 4948 6957 4951
rect 7019 4948 7054 4985
rect 7122 4982 7222 4985
rect 7122 4978 7189 4982
rect 7122 4952 7134 4978
rect 7160 4956 7189 4978
rect 7215 4956 7222 4982
rect 7160 4952 7222 4956
rect 7122 4948 7222 4952
rect 6598 4927 6629 4948
rect 7019 4927 7055 4948
rect 6441 4926 6478 4927
rect 6440 4917 6478 4926
rect 5163 4914 5211 4916
rect 5163 4896 5174 4914
rect 5192 4896 5211 4914
rect 5163 4887 5211 4896
rect 5164 4886 5211 4887
rect 5477 4891 5587 4905
rect 5477 4888 5520 4891
rect 5477 4883 5481 4888
rect 5399 4861 5481 4883
rect 5510 4861 5520 4888
rect 5548 4864 5555 4891
rect 5584 4883 5587 4891
rect 6440 4897 6449 4917
rect 6469 4897 6478 4917
rect 6440 4889 6478 4897
rect 6544 4921 6629 4927
rect 6654 4926 6691 4927
rect 6544 4901 6552 4921
rect 6572 4901 6629 4921
rect 6544 4893 6629 4901
rect 6653 4917 6691 4926
rect 6653 4897 6662 4917
rect 6682 4897 6691 4917
rect 6544 4892 6580 4893
rect 6653 4889 6691 4897
rect 6757 4921 6842 4927
rect 6862 4926 6899 4927
rect 6757 4901 6765 4921
rect 6785 4920 6842 4921
rect 6785 4901 6814 4920
rect 6757 4900 6814 4901
rect 6835 4900 6842 4920
rect 6757 4893 6842 4900
rect 6861 4917 6899 4926
rect 6861 4897 6870 4917
rect 6890 4897 6899 4917
rect 6757 4892 6793 4893
rect 6861 4889 6899 4897
rect 6965 4923 7109 4927
rect 6965 4921 7022 4923
rect 6965 4901 6973 4921
rect 6993 4901 7022 4921
rect 6965 4899 7022 4901
rect 7048 4921 7109 4923
rect 7048 4901 7081 4921
rect 7101 4901 7109 4921
rect 7048 4899 7109 4901
rect 6965 4893 7109 4899
rect 6965 4892 7001 4893
rect 7073 4892 7109 4893
rect 7175 4926 7212 4927
rect 7175 4925 7213 4926
rect 7175 4917 7239 4925
rect 7175 4897 7184 4917
rect 7204 4903 7239 4917
rect 7259 4903 7262 4923
rect 7204 4898 7262 4903
rect 7204 4897 7239 4898
rect 5584 4864 5649 4883
rect 5548 4861 5649 4864
rect 5399 4859 5649 4861
rect 5167 4823 5204 4824
rect 4785 4716 4795 4734
rect 4813 4716 4825 4734
rect 4785 4711 4825 4716
rect 5163 4820 5204 4823
rect 5163 4815 5205 4820
rect 5163 4797 5176 4815
rect 5194 4797 5205 4815
rect 5163 4783 5205 4797
rect 5243 4783 5290 4787
rect 5163 4777 5290 4783
rect 5163 4748 5251 4777
rect 5280 4748 5290 4777
rect 5399 4780 5436 4859
rect 5477 4846 5587 4859
rect 5551 4790 5582 4791
rect 5399 4760 5408 4780
rect 5428 4760 5436 4780
rect 5399 4750 5436 4760
rect 5495 4780 5582 4790
rect 5495 4760 5504 4780
rect 5524 4760 5582 4780
rect 5495 4751 5582 4760
rect 5495 4750 5532 4751
rect 5163 4744 5290 4748
rect 5163 4727 5202 4744
rect 5243 4743 5290 4744
rect 4785 4707 4822 4711
rect 5163 4709 5174 4727
rect 5192 4709 5202 4727
rect 5163 4700 5202 4709
rect 5164 4699 5201 4700
rect 5551 4698 5582 4751
rect 5612 4780 5649 4859
rect 5820 4856 6213 4876
rect 6233 4856 6236 4876
rect 6441 4860 6478 4889
rect 5820 4851 6236 4856
rect 6442 4858 6478 4860
rect 6654 4858 6691 4889
rect 5820 4850 6161 4851
rect 5764 4790 5795 4791
rect 5612 4760 5621 4780
rect 5641 4760 5649 4780
rect 5612 4750 5649 4760
rect 5708 4783 5795 4790
rect 5708 4780 5769 4783
rect 5708 4760 5717 4780
rect 5737 4763 5769 4780
rect 5790 4763 5795 4783
rect 5737 4760 5795 4763
rect 5708 4753 5795 4760
rect 5820 4780 5857 4850
rect 6123 4849 6160 4850
rect 6442 4836 6691 4858
rect 6862 4857 6899 4889
rect 7175 4885 7239 4897
rect 7279 4860 7306 5037
rect 7739 4992 7766 5169
rect 7806 5132 7870 5144
rect 8146 5140 8183 5172
rect 8354 5171 8603 5193
rect 8885 5179 8922 5180
rect 9188 5179 9225 5249
rect 9250 5269 9337 5276
rect 9250 5266 9308 5269
rect 9250 5246 9255 5266
rect 9276 5249 9308 5266
rect 9328 5249 9337 5269
rect 9276 5246 9337 5249
rect 9250 5239 9337 5246
rect 9396 5269 9433 5279
rect 9396 5249 9404 5269
rect 9424 5249 9433 5269
rect 9250 5238 9281 5239
rect 8884 5178 9225 5179
rect 8354 5140 8391 5171
rect 8567 5169 8603 5171
rect 8809 5173 9225 5178
rect 8567 5140 8604 5169
rect 8809 5153 8812 5173
rect 8832 5153 9225 5173
rect 9396 5170 9433 5249
rect 9463 5278 9494 5331
rect 9844 5329 9881 5330
rect 9843 5320 9882 5329
rect 9843 5302 9853 5320
rect 9871 5302 9882 5320
rect 9755 5285 9802 5286
rect 9843 5285 9882 5302
rect 9755 5281 9882 5285
rect 9513 5278 9550 5279
rect 9463 5269 9550 5278
rect 9463 5249 9521 5269
rect 9541 5249 9550 5269
rect 9463 5239 9550 5249
rect 9609 5269 9646 5279
rect 9609 5249 9617 5269
rect 9637 5249 9646 5269
rect 9463 5238 9494 5239
rect 9458 5170 9568 5183
rect 9609 5170 9646 5249
rect 9755 5252 9765 5281
rect 9794 5252 9882 5281
rect 9755 5246 9882 5252
rect 9755 5242 9802 5246
rect 9840 5232 9882 5246
rect 9840 5214 9851 5232
rect 9869 5214 9882 5232
rect 9840 5209 9882 5214
rect 9841 5206 9882 5209
rect 9841 5205 9878 5206
rect 9396 5168 9646 5170
rect 9396 5165 9497 5168
rect 9396 5146 9461 5165
rect 7806 5131 7841 5132
rect 7783 5126 7841 5131
rect 7783 5106 7786 5126
rect 7806 5112 7841 5126
rect 7861 5112 7870 5132
rect 7806 5104 7870 5112
rect 7832 5103 7870 5104
rect 7833 5102 7870 5103
rect 7936 5136 7972 5137
rect 8044 5136 8080 5137
rect 7936 5129 8080 5136
rect 7936 5128 7993 5129
rect 7936 5108 7944 5128
rect 7964 5109 7993 5128
rect 8018 5128 8080 5129
rect 8018 5109 8052 5128
rect 7964 5108 8052 5109
rect 8072 5108 8080 5128
rect 7936 5102 8080 5108
rect 8146 5132 8184 5140
rect 8252 5136 8288 5137
rect 8146 5112 8155 5132
rect 8175 5112 8184 5132
rect 8146 5103 8184 5112
rect 8203 5129 8288 5136
rect 8203 5109 8210 5129
rect 8231 5128 8288 5129
rect 8231 5109 8260 5128
rect 8203 5108 8260 5109
rect 8280 5108 8288 5128
rect 8146 5102 8183 5103
rect 8203 5102 8288 5108
rect 8354 5132 8392 5140
rect 8465 5136 8501 5137
rect 8354 5112 8363 5132
rect 8383 5112 8392 5132
rect 8354 5103 8392 5112
rect 8416 5128 8501 5136
rect 8416 5108 8473 5128
rect 8493 5108 8501 5128
rect 8354 5102 8391 5103
rect 8416 5102 8501 5108
rect 8567 5132 8605 5140
rect 8567 5112 8576 5132
rect 8596 5112 8605 5132
rect 9458 5138 9461 5146
rect 9490 5138 9497 5165
rect 9525 5141 9535 5168
rect 9564 5146 9646 5168
rect 9564 5141 9568 5146
rect 9525 5138 9568 5141
rect 9458 5124 9568 5138
rect 9834 5142 9881 5143
rect 9834 5133 9882 5142
rect 9834 5115 9853 5133
rect 9871 5115 9882 5133
rect 9834 5113 9882 5115
rect 8567 5103 8605 5112
rect 8567 5102 8604 5103
rect 7990 5081 8026 5102
rect 8416 5081 8447 5102
rect 7823 5077 7923 5081
rect 7823 5073 7885 5077
rect 7823 5047 7830 5073
rect 7856 5051 7885 5073
rect 7911 5051 7923 5077
rect 7856 5047 7923 5051
rect 7823 5044 7923 5047
rect 7991 5044 8026 5081
rect 8088 5078 8447 5081
rect 8088 5073 8310 5078
rect 8088 5049 8101 5073
rect 8125 5054 8310 5073
rect 8334 5054 8447 5078
rect 8125 5049 8447 5054
rect 8088 5045 8447 5049
rect 8514 5073 8663 5081
rect 8514 5053 8525 5073
rect 8545 5053 8663 5073
rect 9843 5075 9882 5113
rect 8514 5046 8663 5053
rect 9195 5056 9233 5058
rect 9843 5056 9885 5075
rect 8514 5045 8555 5046
rect 7990 5040 8026 5044
rect 7990 5011 8027 5040
rect 7838 4992 7875 4993
rect 7934 4992 7971 4993
rect 7990 4992 8026 5011
rect 8045 4992 8082 4993
rect 7738 4983 7876 4992
rect 7738 4963 7847 4983
rect 7867 4963 7876 4983
rect 7738 4956 7876 4963
rect 7934 4983 8082 4992
rect 7934 4963 7943 4983
rect 7963 4963 8053 4983
rect 8073 4963 8082 4983
rect 7738 4954 7834 4956
rect 7934 4953 8082 4963
rect 8141 4983 8178 4993
rect 8253 4992 8290 4993
rect 8234 4990 8290 4992
rect 8141 4963 8149 4983
rect 8169 4963 8178 4983
rect 7990 4952 8026 4953
rect 7838 4893 7875 4894
rect 8141 4893 8178 4963
rect 8203 4983 8290 4990
rect 8203 4980 8261 4983
rect 8203 4960 8208 4980
rect 8229 4963 8261 4980
rect 8281 4963 8290 4983
rect 8229 4960 8290 4963
rect 8203 4953 8290 4960
rect 8349 4983 8386 4993
rect 8349 4963 8357 4983
rect 8377 4963 8386 4983
rect 8203 4952 8234 4953
rect 7837 4892 8178 4893
rect 7762 4887 8178 4892
rect 7387 4860 7440 4868
rect 7762 4867 7765 4887
rect 7785 4867 8178 4887
rect 8349 4884 8386 4963
rect 8416 4992 8447 5045
rect 9195 5033 9885 5056
rect 9195 5023 9881 5033
rect 8466 4992 8503 4993
rect 8416 4983 8503 4992
rect 8416 4963 8474 4983
rect 8494 4963 8503 4983
rect 8416 4953 8503 4963
rect 8562 4983 8599 4993
rect 8562 4963 8570 4983
rect 8590 4963 8599 4983
rect 8416 4952 8447 4953
rect 8411 4884 8521 4897
rect 8562 4884 8599 4963
rect 8349 4882 8599 4884
rect 8349 4879 8450 4882
rect 8349 4860 8414 4879
rect 7254 4859 7440 4860
rect 7138 4857 7440 4859
rect 6523 4830 6634 4836
rect 6862 4831 7440 4857
rect 8411 4852 8414 4860
rect 8443 4852 8450 4879
rect 8478 4855 8488 4882
rect 8517 4860 8599 4882
rect 8787 4935 8955 4936
rect 9195 4935 9233 5023
rect 9494 5022 9541 5023
rect 9841 4999 9881 5023
rect 9458 4966 9570 4985
rect 9458 4965 9501 4966
rect 8787 4912 9233 4935
rect 9459 4964 9501 4965
rect 9459 4944 9466 4964
rect 9485 4944 9501 4964
rect 9459 4936 9501 4944
rect 9529 4964 9570 4966
rect 9529 4944 9543 4964
rect 9562 4944 9570 4964
rect 9842 4955 9881 4999
rect 9529 4936 9570 4944
rect 9459 4930 9570 4936
rect 8787 4909 9231 4912
rect 8787 4907 8955 4909
rect 8517 4855 8521 4860
rect 8478 4852 8521 4855
rect 8411 4838 8521 4852
rect 7138 4830 7440 4831
rect 6523 4822 6564 4830
rect 6523 4802 6531 4822
rect 6550 4802 6564 4822
rect 6523 4800 6564 4802
rect 6592 4822 6634 4830
rect 6592 4802 6608 4822
rect 6627 4802 6634 4822
rect 6592 4800 6634 4802
rect 5972 4790 6008 4791
rect 5820 4760 5829 4780
rect 5849 4760 5857 4780
rect 5708 4751 5764 4753
rect 5708 4750 5745 4751
rect 5820 4750 5857 4760
rect 5916 4780 6064 4790
rect 6164 4787 6260 4789
rect 5916 4760 5925 4780
rect 5945 4760 6035 4780
rect 6055 4760 6064 4780
rect 5916 4751 6064 4760
rect 6122 4780 6260 4787
rect 6523 4785 6634 4800
rect 6122 4760 6131 4780
rect 6151 4760 6260 4780
rect 6122 4751 6260 4760
rect 5916 4750 5953 4751
rect 5972 4699 6008 4751
rect 6027 4750 6064 4751
rect 6123 4750 6160 4751
rect 5443 4697 5484 4698
rect 5335 4690 5484 4697
rect 4458 4688 4495 4689
rect 4408 4679 4495 4688
rect 4408 4659 4466 4679
rect 4486 4659 4495 4679
rect 4408 4649 4495 4659
rect 4554 4679 4591 4689
rect 4554 4659 4562 4679
rect 4582 4659 4591 4679
rect 5335 4670 5453 4690
rect 5473 4670 5484 4690
rect 5335 4662 5484 4670
rect 5551 4694 5910 4698
rect 5551 4689 5873 4694
rect 5551 4665 5664 4689
rect 5688 4670 5873 4689
rect 5897 4670 5910 4694
rect 5688 4665 5910 4670
rect 5551 4662 5910 4665
rect 5972 4662 6007 4699
rect 6075 4696 6175 4699
rect 6075 4692 6142 4696
rect 6075 4666 6087 4692
rect 6113 4670 6142 4692
rect 6168 4670 6175 4696
rect 6113 4666 6175 4670
rect 6075 4662 6175 4666
rect 4408 4648 4439 4649
rect 4403 4580 4513 4593
rect 4554 4580 4591 4659
rect 4788 4644 4825 4645
rect 4784 4635 4825 4644
rect 5551 4641 5582 4662
rect 5972 4641 6008 4662
rect 5394 4640 5431 4641
rect 5168 4637 5202 4638
rect 4784 4617 4797 4635
rect 4815 4617 4825 4635
rect 4784 4608 4825 4617
rect 5167 4628 5204 4637
rect 5167 4610 5176 4628
rect 5194 4610 5204 4628
rect 4784 4588 4824 4608
rect 5167 4600 5204 4610
rect 5393 4631 5431 4640
rect 5393 4611 5402 4631
rect 5422 4611 5431 4631
rect 5393 4603 5431 4611
rect 5497 4635 5582 4641
rect 5607 4640 5644 4641
rect 5497 4615 5505 4635
rect 5525 4615 5582 4635
rect 5497 4607 5582 4615
rect 5606 4631 5644 4640
rect 5606 4611 5615 4631
rect 5635 4611 5644 4631
rect 5497 4606 5533 4607
rect 5606 4603 5644 4611
rect 5710 4635 5795 4641
rect 5815 4640 5852 4641
rect 5710 4615 5718 4635
rect 5738 4634 5795 4635
rect 5738 4615 5767 4634
rect 5710 4614 5767 4615
rect 5788 4614 5795 4634
rect 5710 4607 5795 4614
rect 5814 4631 5852 4640
rect 5814 4611 5823 4631
rect 5843 4611 5852 4631
rect 5710 4606 5746 4607
rect 5814 4603 5852 4611
rect 5918 4635 6062 4641
rect 5918 4615 5926 4635
rect 5946 4634 6034 4635
rect 5946 4615 5977 4634
rect 5918 4614 5977 4615
rect 6002 4615 6034 4634
rect 6054 4615 6062 4635
rect 6002 4614 6062 4615
rect 5918 4607 6062 4614
rect 5918 4606 5954 4607
rect 6026 4606 6062 4607
rect 6128 4640 6165 4641
rect 6128 4639 6166 4640
rect 6128 4631 6192 4639
rect 6128 4611 6137 4631
rect 6157 4617 6192 4631
rect 6212 4617 6215 4637
rect 6157 4612 6215 4617
rect 6157 4611 6192 4612
rect 4341 4578 4591 4580
rect 4341 4575 4442 4578
rect 2859 4518 2923 4530
rect 3199 4526 3236 4553
rect 3407 4526 3444 4557
rect 3620 4555 3656 4557
rect 4341 4556 4406 4575
rect 3620 4526 3657 4555
rect 4403 4548 4406 4556
rect 4435 4548 4442 4575
rect 4470 4551 4480 4578
rect 4509 4556 4591 4578
rect 4699 4578 4824 4588
rect 4699 4559 4707 4578
rect 4732 4559 4824 4578
rect 4509 4551 4513 4556
rect 4699 4552 4824 4559
rect 4470 4548 4513 4551
rect 4403 4534 4513 4548
rect 2859 4517 2894 4518
rect 2836 4512 2894 4517
rect 2836 4492 2839 4512
rect 2859 4498 2894 4512
rect 2914 4498 2923 4518
rect 2859 4490 2923 4498
rect 2885 4489 2923 4490
rect 2886 4488 2923 4489
rect 2989 4522 3025 4523
rect 3097 4522 3133 4523
rect 2989 4514 3133 4522
rect 2989 4494 2997 4514
rect 3017 4494 3105 4514
rect 3125 4494 3133 4514
rect 2989 4488 3133 4494
rect 3199 4518 3237 4526
rect 3305 4522 3341 4523
rect 3199 4498 3208 4518
rect 3228 4498 3237 4518
rect 3199 4489 3237 4498
rect 3256 4515 3341 4522
rect 3256 4495 3263 4515
rect 3284 4514 3341 4515
rect 3284 4495 3313 4514
rect 3256 4494 3313 4495
rect 3333 4494 3341 4514
rect 3199 4488 3236 4489
rect 3256 4488 3341 4494
rect 3407 4518 3445 4526
rect 3518 4522 3554 4523
rect 3407 4498 3416 4518
rect 3436 4498 3445 4518
rect 3407 4489 3445 4498
rect 3469 4514 3554 4522
rect 3469 4494 3526 4514
rect 3546 4494 3554 4514
rect 3407 4488 3444 4489
rect 3469 4488 3554 4494
rect 3620 4518 3658 4526
rect 3620 4498 3629 4518
rect 3649 4498 3658 4518
rect 3620 4489 3658 4498
rect 4784 4504 4824 4552
rect 5168 4572 5202 4600
rect 5394 4574 5431 4603
rect 5395 4572 5431 4574
rect 5607 4572 5644 4603
rect 5168 4571 5340 4572
rect 5168 4539 5354 4571
rect 5395 4550 5644 4572
rect 5815 4571 5852 4603
rect 6128 4599 6192 4611
rect 6232 4573 6259 4751
rect 7387 4723 7440 4830
rect 8787 4729 8814 4907
rect 8854 4869 8918 4881
rect 9194 4877 9231 4909
rect 9402 4908 9651 4930
rect 9402 4877 9439 4908
rect 9615 4906 9651 4908
rect 9615 4877 9652 4906
rect 8854 4868 8889 4869
rect 8831 4863 8889 4868
rect 8831 4843 8834 4863
rect 8854 4849 8889 4863
rect 8909 4849 8918 4869
rect 8854 4841 8918 4849
rect 8880 4840 8918 4841
rect 8881 4839 8918 4840
rect 8984 4873 9020 4874
rect 9092 4873 9128 4874
rect 8984 4868 9128 4873
rect 8984 4865 9046 4868
rect 8984 4845 8992 4865
rect 9012 4848 9046 4865
rect 9069 4865 9128 4868
rect 9069 4848 9100 4865
rect 9012 4845 9100 4848
rect 9120 4845 9128 4865
rect 8984 4839 9128 4845
rect 9194 4869 9232 4877
rect 9300 4873 9336 4874
rect 9194 4849 9203 4869
rect 9223 4849 9232 4869
rect 9194 4840 9232 4849
rect 9251 4866 9336 4873
rect 9251 4846 9258 4866
rect 9279 4865 9336 4866
rect 9279 4846 9308 4865
rect 9251 4845 9308 4846
rect 9328 4845 9336 4865
rect 9194 4839 9231 4840
rect 9251 4839 9336 4845
rect 9402 4869 9440 4877
rect 9513 4873 9549 4874
rect 9402 4849 9411 4869
rect 9431 4849 9440 4869
rect 9402 4840 9440 4849
rect 9464 4865 9549 4873
rect 9464 4845 9521 4865
rect 9541 4845 9549 4865
rect 9402 4839 9439 4840
rect 9464 4839 9549 4845
rect 9615 4869 9653 4877
rect 9615 4849 9624 4869
rect 9644 4849 9653 4869
rect 9615 4840 9653 4849
rect 9615 4839 9652 4840
rect 9038 4818 9074 4839
rect 9464 4818 9495 4839
rect 8871 4814 8971 4818
rect 8871 4810 8933 4814
rect 8871 4784 8878 4810
rect 8904 4788 8933 4810
rect 8959 4788 8971 4814
rect 8904 4784 8971 4788
rect 8871 4781 8971 4784
rect 9039 4781 9074 4818
rect 9136 4815 9495 4818
rect 9136 4810 9358 4815
rect 9136 4786 9149 4810
rect 9173 4791 9358 4810
rect 9382 4791 9495 4815
rect 9173 4786 9495 4791
rect 9136 4782 9495 4786
rect 9562 4810 9711 4818
rect 9562 4790 9573 4810
rect 9593 4790 9711 4810
rect 9562 4783 9711 4790
rect 9562 4782 9603 4783
rect 8886 4729 8923 4730
rect 8982 4729 9019 4730
rect 9038 4729 9074 4781
rect 9093 4729 9130 4730
rect 7387 4705 7435 4723
rect 7387 4665 7395 4705
rect 7422 4665 7435 4705
rect 8786 4720 8924 4729
rect 8786 4700 8895 4720
rect 8915 4700 8924 4720
rect 8786 4693 8924 4700
rect 8982 4720 9130 4729
rect 8982 4700 8991 4720
rect 9011 4700 9101 4720
rect 9121 4700 9130 4720
rect 8786 4691 8882 4693
rect 8982 4690 9130 4700
rect 9189 4720 9226 4730
rect 9301 4729 9338 4730
rect 9282 4727 9338 4729
rect 9189 4700 9197 4720
rect 9217 4700 9226 4720
rect 9038 4689 9074 4690
rect 6415 4647 6525 4661
rect 7387 4651 7435 4665
rect 8520 4656 8631 4671
rect 8520 4654 8562 4656
rect 6415 4644 6458 4647
rect 6415 4639 6419 4644
rect 6091 4571 6259 4573
rect 5815 4565 6259 4571
rect 5168 4507 5202 4539
rect 3620 4488 3657 4489
rect 3043 4467 3079 4488
rect 3469 4467 3500 4488
rect 4784 4486 4795 4504
rect 4813 4486 4824 4504
rect 4784 4478 4824 4486
rect 5164 4498 5202 4507
rect 5164 4480 5174 4498
rect 5192 4480 5202 4498
rect 4785 4477 4822 4478
rect 5164 4474 5202 4480
rect 5320 4476 5354 4539
rect 5476 4544 5587 4550
rect 5476 4536 5517 4544
rect 5476 4516 5484 4536
rect 5503 4516 5517 4536
rect 5476 4514 5517 4516
rect 5545 4536 5587 4544
rect 5545 4516 5561 4536
rect 5580 4516 5587 4536
rect 5545 4514 5587 4516
rect 5476 4499 5587 4514
rect 5814 4545 6259 4565
rect 5814 4476 5852 4545
rect 6091 4544 6259 4545
rect 6337 4617 6419 4639
rect 6448 4617 6458 4644
rect 6486 4620 6493 4647
rect 6522 4639 6525 4647
rect 6522 4620 6587 4639
rect 6486 4617 6587 4620
rect 6337 4615 6587 4617
rect 6337 4536 6374 4615
rect 6415 4602 6525 4615
rect 6489 4546 6520 4547
rect 6337 4516 6346 4536
rect 6366 4516 6374 4536
rect 6337 4506 6374 4516
rect 6433 4536 6520 4546
rect 6433 4516 6442 4536
rect 6462 4516 6520 4536
rect 6433 4507 6520 4516
rect 6433 4506 6470 4507
rect 5164 4470 5201 4474
rect 2876 4463 2976 4467
rect 2876 4459 2938 4463
rect 2876 4433 2883 4459
rect 2909 4437 2938 4459
rect 2964 4437 2976 4463
rect 2909 4433 2976 4437
rect 2876 4430 2976 4433
rect 3044 4430 3079 4467
rect 3141 4464 3500 4467
rect 3141 4459 3363 4464
rect 3141 4435 3154 4459
rect 3178 4440 3363 4459
rect 3387 4440 3500 4464
rect 3178 4435 3500 4440
rect 3141 4431 3500 4435
rect 3567 4459 3716 4467
rect 5320 4465 5852 4476
rect 3567 4439 3578 4459
rect 3598 4439 3716 4459
rect 5319 4449 5852 4465
rect 6489 4454 6520 4507
rect 6550 4536 6587 4615
rect 6758 4612 7151 4632
rect 7171 4612 7174 4632
rect 8253 4627 8294 4636
rect 6758 4607 7174 4612
rect 7848 4625 8016 4626
rect 8253 4625 8262 4627
rect 6758 4606 7099 4607
rect 6702 4546 6733 4547
rect 6550 4516 6559 4536
rect 6579 4516 6587 4536
rect 6550 4506 6587 4516
rect 6646 4539 6733 4546
rect 6646 4536 6707 4539
rect 6646 4516 6655 4536
rect 6675 4519 6707 4536
rect 6728 4519 6733 4539
rect 6675 4516 6733 4519
rect 6646 4509 6733 4516
rect 6758 4536 6795 4606
rect 7061 4605 7098 4606
rect 7848 4605 8262 4625
rect 8288 4605 8294 4627
rect 8520 4634 8527 4654
rect 8546 4634 8562 4654
rect 8520 4626 8562 4634
rect 8590 4654 8631 4656
rect 8590 4634 8604 4654
rect 8623 4634 8631 4654
rect 8590 4626 8631 4634
rect 8886 4630 8923 4631
rect 9189 4630 9226 4700
rect 9251 4720 9338 4727
rect 9251 4717 9309 4720
rect 9251 4697 9256 4717
rect 9277 4700 9309 4717
rect 9329 4700 9338 4720
rect 9277 4697 9338 4700
rect 9251 4690 9338 4697
rect 9397 4720 9434 4730
rect 9397 4700 9405 4720
rect 9425 4700 9434 4720
rect 9251 4689 9282 4690
rect 8885 4629 9226 4630
rect 8520 4620 8631 4626
rect 8810 4624 9226 4629
rect 7848 4599 8294 4605
rect 7848 4597 8016 4599
rect 6910 4546 6946 4547
rect 6758 4516 6767 4536
rect 6787 4516 6795 4536
rect 6646 4507 6702 4509
rect 6646 4506 6683 4507
rect 6758 4506 6795 4516
rect 6854 4536 7002 4546
rect 7102 4543 7198 4545
rect 6854 4516 6863 4536
rect 6883 4516 6973 4536
rect 6993 4516 7002 4536
rect 6854 4507 7002 4516
rect 7060 4536 7198 4543
rect 7060 4516 7069 4536
rect 7089 4516 7198 4536
rect 7060 4507 7198 4516
rect 6854 4506 6891 4507
rect 6910 4455 6946 4507
rect 6965 4506 7002 4507
rect 7061 4506 7098 4507
rect 6381 4453 6422 4454
rect 5319 4448 5833 4449
rect 3567 4432 3716 4439
rect 6273 4446 6422 4453
rect 4156 4436 4670 4437
rect 3567 4431 3608 4432
rect 3043 4395 3079 4430
rect 2891 4378 2928 4379
rect 2987 4378 3024 4379
rect 3043 4378 3050 4395
rect 2791 4369 2929 4378
rect 2791 4349 2900 4369
rect 2920 4349 2929 4369
rect 2791 4342 2929 4349
rect 2987 4369 3050 4378
rect 2987 4349 2996 4369
rect 3016 4354 3050 4369
rect 3071 4378 3079 4395
rect 3098 4378 3135 4379
rect 3071 4369 3135 4378
rect 3071 4354 3106 4369
rect 3016 4349 3106 4354
rect 3126 4349 3135 4369
rect 2791 4340 2887 4342
rect 2987 4339 3135 4349
rect 3194 4369 3231 4379
rect 3306 4378 3343 4379
rect 3287 4376 3343 4378
rect 3194 4349 3202 4369
rect 3222 4349 3231 4369
rect 3043 4338 3079 4339
rect 1973 4286 2141 4288
rect 1695 4280 2141 4286
rect 763 4256 1179 4261
rect 1358 4259 1469 4265
rect 763 4255 1104 4256
rect 707 4195 738 4196
rect 555 4165 564 4185
rect 584 4165 592 4185
rect 555 4155 592 4165
rect 651 4188 738 4195
rect 651 4185 712 4188
rect 651 4165 660 4185
rect 680 4168 712 4185
rect 733 4168 738 4188
rect 680 4165 738 4168
rect 651 4158 738 4165
rect 763 4185 800 4255
rect 1066 4254 1103 4255
rect 1358 4251 1399 4259
rect 1358 4231 1366 4251
rect 1385 4231 1399 4251
rect 1358 4229 1399 4231
rect 1427 4251 1469 4259
rect 1427 4231 1443 4251
rect 1462 4231 1469 4251
rect 1695 4258 1701 4280
rect 1727 4260 2141 4280
rect 2891 4279 2928 4280
rect 3194 4279 3231 4349
rect 3256 4369 3343 4376
rect 3256 4366 3314 4369
rect 3256 4346 3261 4366
rect 3282 4349 3314 4366
rect 3334 4349 3343 4369
rect 3282 4346 3343 4349
rect 3256 4339 3343 4346
rect 3402 4369 3439 4379
rect 3402 4349 3410 4369
rect 3430 4349 3439 4369
rect 3256 4338 3287 4339
rect 2890 4278 3231 4279
rect 1727 4258 1736 4260
rect 1973 4259 2141 4260
rect 2815 4277 3231 4278
rect 2815 4273 3191 4277
rect 1695 4249 1736 4258
rect 2815 4253 2818 4273
rect 2838 4260 3191 4273
rect 3223 4260 3231 4277
rect 2838 4253 3231 4260
rect 3402 4270 3439 4349
rect 3469 4378 3500 4431
rect 4137 4420 4670 4436
rect 6273 4426 6391 4446
rect 6411 4426 6422 4446
rect 4137 4409 4669 4420
rect 6273 4418 6422 4426
rect 6489 4450 6848 4454
rect 6489 4445 6811 4450
rect 6489 4421 6602 4445
rect 6626 4426 6811 4445
rect 6835 4426 6848 4450
rect 6626 4421 6848 4426
rect 6489 4418 6848 4421
rect 6910 4418 6945 4455
rect 7013 4452 7113 4455
rect 7013 4448 7080 4452
rect 7013 4422 7025 4448
rect 7051 4426 7080 4448
rect 7106 4426 7113 4452
rect 7051 4422 7113 4426
rect 7013 4418 7113 4422
rect 4788 4411 4825 4415
rect 3519 4378 3556 4379
rect 3469 4369 3556 4378
rect 3469 4349 3527 4369
rect 3547 4349 3556 4369
rect 3469 4339 3556 4349
rect 3615 4369 3652 4379
rect 3615 4349 3623 4369
rect 3643 4349 3652 4369
rect 3469 4338 3500 4339
rect 3464 4270 3574 4283
rect 3615 4270 3652 4349
rect 3402 4268 3652 4270
rect 3402 4265 3503 4268
rect 3402 4246 3467 4265
rect 1427 4229 1469 4231
rect 1358 4214 1469 4229
rect 3464 4238 3467 4246
rect 3496 4238 3503 4265
rect 3531 4241 3541 4268
rect 3570 4246 3652 4268
rect 3730 4340 3898 4341
rect 4137 4340 4175 4409
rect 3730 4320 4175 4340
rect 4402 4371 4513 4386
rect 4402 4369 4444 4371
rect 4402 4349 4409 4369
rect 4428 4349 4444 4369
rect 4402 4341 4444 4349
rect 4472 4369 4513 4371
rect 4472 4349 4486 4369
rect 4505 4349 4513 4369
rect 4472 4341 4513 4349
rect 4402 4335 4513 4341
rect 4635 4346 4669 4409
rect 4787 4405 4825 4411
rect 5167 4407 5204 4408
rect 4787 4387 4797 4405
rect 4815 4387 4825 4405
rect 4787 4378 4825 4387
rect 5165 4399 5205 4407
rect 5165 4381 5176 4399
rect 5194 4381 5205 4399
rect 6489 4397 6520 4418
rect 6910 4397 6946 4418
rect 6332 4396 6369 4397
rect 4787 4346 4821 4378
rect 3730 4314 4174 4320
rect 3730 4312 3898 4314
rect 3570 4241 3574 4246
rect 3531 4238 3574 4241
rect 3464 4224 3574 4238
rect 915 4195 951 4196
rect 763 4165 772 4185
rect 792 4165 800 4185
rect 651 4156 707 4158
rect 651 4155 688 4156
rect 763 4155 800 4165
rect 859 4185 1007 4195
rect 1107 4192 1203 4194
rect 859 4165 868 4185
rect 888 4165 978 4185
rect 998 4165 1007 4185
rect 859 4156 1007 4165
rect 1065 4185 1203 4192
rect 1065 4165 1074 4185
rect 1094 4165 1203 4185
rect 1065 4156 1203 4165
rect 859 4155 896 4156
rect 915 4104 951 4156
rect 970 4155 1007 4156
rect 1066 4155 1103 4156
rect 386 4102 427 4103
rect 278 4095 427 4102
rect 278 4075 396 4095
rect 416 4075 427 4095
rect 278 4067 427 4075
rect 494 4099 853 4103
rect 494 4094 816 4099
rect 494 4070 607 4094
rect 631 4075 816 4094
rect 840 4075 853 4099
rect 631 4070 853 4075
rect 494 4067 853 4070
rect 915 4067 950 4104
rect 1018 4101 1118 4104
rect 1018 4097 1085 4101
rect 1018 4071 1030 4097
rect 1056 4075 1085 4097
rect 1111 4075 1118 4101
rect 1056 4071 1118 4075
rect 1018 4067 1118 4071
rect 494 4046 525 4067
rect 915 4046 951 4067
rect 337 4045 374 4046
rect 336 4036 374 4045
rect 336 4016 345 4036
rect 365 4016 374 4036
rect 336 4008 374 4016
rect 440 4040 525 4046
rect 550 4045 587 4046
rect 440 4020 448 4040
rect 468 4020 525 4040
rect 440 4012 525 4020
rect 549 4036 587 4045
rect 549 4016 558 4036
rect 578 4016 587 4036
rect 440 4011 476 4012
rect 549 4008 587 4016
rect 653 4040 738 4046
rect 758 4045 795 4046
rect 653 4020 661 4040
rect 681 4039 738 4040
rect 681 4020 710 4039
rect 653 4019 710 4020
rect 731 4019 738 4039
rect 653 4012 738 4019
rect 757 4036 795 4045
rect 757 4016 766 4036
rect 786 4016 795 4036
rect 653 4011 689 4012
rect 757 4008 795 4016
rect 861 4040 1005 4046
rect 861 4020 869 4040
rect 889 4037 977 4040
rect 889 4020 920 4037
rect 861 4017 920 4020
rect 943 4020 977 4037
rect 997 4020 1005 4040
rect 943 4017 1005 4020
rect 861 4012 1005 4017
rect 861 4011 897 4012
rect 969 4011 1005 4012
rect 1071 4045 1108 4046
rect 1071 4044 1109 4045
rect 1071 4036 1135 4044
rect 1071 4016 1080 4036
rect 1100 4022 1135 4036
rect 1155 4022 1158 4042
rect 1100 4017 1158 4022
rect 1100 4016 1135 4017
rect 337 3979 374 4008
rect 338 3977 374 3979
rect 550 3977 587 4008
rect 338 3955 587 3977
rect 758 3976 795 4008
rect 1071 4004 1135 4016
rect 1175 3978 1202 4156
rect 3730 4134 3757 4312
rect 3797 4274 3861 4286
rect 4137 4282 4174 4314
rect 4345 4313 4594 4335
rect 4635 4314 4821 4346
rect 4649 4313 4821 4314
rect 4345 4282 4382 4313
rect 4558 4311 4594 4313
rect 4558 4282 4595 4311
rect 4787 4285 4821 4313
rect 5165 4333 5205 4381
rect 6331 4387 6369 4396
rect 6331 4367 6340 4387
rect 6360 4367 6369 4387
rect 6331 4359 6369 4367
rect 6435 4391 6520 4397
rect 6545 4396 6582 4397
rect 6435 4371 6443 4391
rect 6463 4371 6520 4391
rect 6435 4363 6520 4371
rect 6544 4387 6582 4396
rect 6544 4367 6553 4387
rect 6573 4367 6582 4387
rect 6435 4362 6471 4363
rect 6544 4359 6582 4367
rect 6648 4391 6733 4397
rect 6753 4396 6790 4397
rect 6648 4371 6656 4391
rect 6676 4390 6733 4391
rect 6676 4371 6705 4390
rect 6648 4370 6705 4371
rect 6726 4370 6733 4390
rect 6648 4363 6733 4370
rect 6752 4387 6790 4396
rect 6752 4367 6761 4387
rect 6781 4367 6790 4387
rect 6648 4362 6684 4363
rect 6752 4359 6790 4367
rect 6856 4391 7000 4397
rect 6856 4371 6864 4391
rect 6884 4374 6920 4391
rect 6940 4374 6972 4391
rect 6884 4371 6972 4374
rect 6992 4371 7000 4391
rect 6856 4363 7000 4371
rect 6856 4362 6892 4363
rect 6964 4362 7000 4363
rect 7066 4396 7103 4397
rect 7066 4395 7104 4396
rect 7066 4387 7130 4395
rect 7066 4367 7075 4387
rect 7095 4373 7130 4387
rect 7150 4373 7153 4393
rect 7095 4368 7153 4373
rect 7095 4367 7130 4368
rect 5476 4337 5586 4351
rect 5476 4334 5519 4337
rect 5165 4326 5290 4333
rect 5476 4329 5480 4334
rect 5165 4307 5257 4326
rect 5282 4307 5290 4326
rect 5165 4297 5290 4307
rect 5398 4307 5480 4329
rect 5509 4307 5519 4334
rect 5547 4310 5554 4337
rect 5583 4329 5586 4337
rect 6332 4330 6369 4359
rect 5583 4310 5648 4329
rect 6333 4328 6369 4330
rect 6545 4328 6582 4359
rect 6753 4332 6790 4359
rect 7066 4355 7130 4367
rect 5547 4307 5648 4310
rect 5398 4305 5648 4307
rect 3797 4273 3832 4274
rect 3774 4268 3832 4273
rect 3774 4248 3777 4268
rect 3797 4254 3832 4268
rect 3852 4254 3861 4274
rect 3797 4246 3861 4254
rect 3823 4245 3861 4246
rect 3824 4244 3861 4245
rect 3927 4278 3963 4279
rect 4035 4278 4071 4279
rect 3927 4271 4071 4278
rect 3927 4270 3987 4271
rect 3927 4250 3935 4270
rect 3955 4251 3987 4270
rect 4012 4270 4071 4271
rect 4012 4251 4043 4270
rect 3955 4250 4043 4251
rect 4063 4250 4071 4270
rect 3927 4244 4071 4250
rect 4137 4274 4175 4282
rect 4243 4278 4279 4279
rect 4137 4254 4146 4274
rect 4166 4254 4175 4274
rect 4137 4245 4175 4254
rect 4194 4271 4279 4278
rect 4194 4251 4201 4271
rect 4222 4270 4279 4271
rect 4222 4251 4251 4270
rect 4194 4250 4251 4251
rect 4271 4250 4279 4270
rect 4137 4244 4174 4245
rect 4194 4244 4279 4250
rect 4345 4274 4383 4282
rect 4456 4278 4492 4279
rect 4345 4254 4354 4274
rect 4374 4254 4383 4274
rect 4345 4245 4383 4254
rect 4407 4270 4492 4278
rect 4407 4250 4464 4270
rect 4484 4250 4492 4270
rect 4345 4244 4382 4245
rect 4407 4244 4492 4250
rect 4558 4274 4596 4282
rect 4558 4254 4567 4274
rect 4587 4254 4596 4274
rect 4558 4245 4596 4254
rect 4785 4275 4822 4285
rect 5165 4277 5205 4297
rect 4785 4257 4795 4275
rect 4813 4257 4822 4275
rect 4785 4248 4822 4257
rect 5164 4268 5205 4277
rect 5164 4250 5174 4268
rect 5192 4250 5205 4268
rect 4787 4247 4821 4248
rect 4558 4244 4595 4245
rect 3981 4223 4017 4244
rect 4407 4223 4438 4244
rect 5164 4241 5205 4250
rect 5164 4240 5201 4241
rect 5398 4226 5435 4305
rect 5476 4292 5586 4305
rect 5550 4236 5581 4237
rect 3814 4219 3914 4223
rect 3814 4215 3876 4219
rect 3814 4189 3821 4215
rect 3847 4193 3876 4215
rect 3902 4193 3914 4219
rect 3847 4189 3914 4193
rect 3814 4186 3914 4189
rect 3982 4186 4017 4223
rect 4079 4220 4438 4223
rect 4079 4215 4301 4220
rect 4079 4191 4092 4215
rect 4116 4196 4301 4215
rect 4325 4196 4438 4220
rect 4116 4191 4438 4196
rect 4079 4187 4438 4191
rect 4505 4215 4654 4223
rect 4505 4195 4516 4215
rect 4536 4195 4654 4215
rect 5398 4206 5407 4226
rect 5427 4206 5435 4226
rect 5398 4196 5435 4206
rect 5494 4226 5581 4236
rect 5494 4206 5503 4226
rect 5523 4206 5581 4226
rect 5494 4197 5581 4206
rect 5494 4196 5531 4197
rect 4505 4188 4654 4195
rect 4505 4187 4546 4188
rect 3829 4134 3866 4135
rect 3925 4134 3962 4135
rect 3981 4134 4017 4186
rect 4036 4134 4073 4135
rect 3729 4125 3867 4134
rect 3324 4104 3435 4119
rect 3324 4102 3366 4104
rect 2994 4081 3099 4083
rect 2650 4073 2820 4074
rect 2994 4073 3043 4081
rect 2650 4054 3043 4073
rect 3074 4054 3099 4081
rect 3324 4082 3331 4102
rect 3350 4082 3366 4102
rect 3324 4074 3366 4082
rect 3394 4102 3435 4104
rect 3394 4082 3408 4102
rect 3427 4082 3435 4102
rect 3729 4105 3838 4125
rect 3858 4105 3867 4125
rect 3729 4098 3867 4105
rect 3925 4125 4073 4134
rect 3925 4105 3934 4125
rect 3954 4105 4044 4125
rect 4064 4105 4073 4125
rect 3729 4096 3825 4098
rect 3925 4095 4073 4105
rect 4132 4125 4169 4135
rect 4244 4134 4281 4135
rect 4225 4132 4281 4134
rect 4132 4105 4140 4125
rect 4160 4105 4169 4125
rect 3981 4094 4017 4095
rect 3394 4074 3435 4082
rect 3324 4068 3435 4074
rect 2650 4047 3099 4054
rect 2650 4045 2820 4047
rect 1500 4014 1610 4028
rect 1500 4011 1543 4014
rect 1500 4006 1504 4011
rect 1034 3976 1202 3978
rect 758 3973 1202 3976
rect 419 3949 530 3955
rect 419 3941 460 3949
rect 108 3886 147 3930
rect 419 3921 427 3941
rect 446 3921 460 3941
rect 419 3919 460 3921
rect 488 3941 530 3949
rect 488 3921 504 3941
rect 523 3921 530 3941
rect 488 3919 530 3921
rect 419 3904 530 3919
rect 756 3950 1202 3973
rect 108 3862 148 3886
rect 448 3862 495 3864
rect 756 3862 794 3950
rect 1034 3949 1202 3950
rect 1422 3984 1504 4006
rect 1533 3984 1543 4011
rect 1571 3987 1578 4014
rect 1607 4006 1610 4014
rect 1607 3987 1672 4006
rect 1571 3984 1672 3987
rect 1422 3982 1672 3984
rect 1422 3903 1459 3982
rect 1500 3969 1610 3982
rect 1574 3913 1605 3914
rect 1422 3883 1431 3903
rect 1451 3883 1459 3903
rect 1422 3873 1459 3883
rect 1518 3903 1605 3913
rect 1518 3883 1527 3903
rect 1547 3883 1605 3903
rect 1518 3874 1605 3883
rect 1518 3873 1555 3874
rect 108 3829 794 3862
rect 108 3772 147 3829
rect 756 3827 794 3829
rect 1574 3821 1605 3874
rect 1635 3903 1672 3982
rect 1843 3995 2236 3999
rect 1843 3978 1862 3995
rect 1882 3979 2236 3995
rect 2256 3979 2259 3999
rect 1882 3978 2259 3979
rect 1843 3974 2259 3978
rect 1843 3973 2184 3974
rect 1787 3913 1818 3914
rect 1635 3883 1644 3903
rect 1664 3883 1672 3903
rect 1635 3873 1672 3883
rect 1731 3906 1818 3913
rect 1731 3903 1792 3906
rect 1731 3883 1740 3903
rect 1760 3886 1792 3903
rect 1813 3886 1818 3906
rect 1760 3883 1818 3886
rect 1731 3876 1818 3883
rect 1843 3903 1880 3973
rect 2146 3972 2183 3973
rect 1995 3913 2031 3914
rect 1843 3883 1852 3903
rect 1872 3883 1880 3903
rect 1731 3874 1787 3876
rect 1731 3873 1768 3874
rect 1843 3873 1880 3883
rect 1939 3903 2087 3913
rect 2187 3910 2283 3912
rect 1939 3883 1948 3903
rect 1968 3883 2058 3903
rect 2078 3883 2087 3903
rect 1939 3874 2087 3883
rect 2145 3903 2283 3910
rect 2145 3883 2154 3903
rect 2174 3883 2283 3903
rect 2145 3874 2283 3883
rect 1939 3873 1976 3874
rect 1995 3822 2031 3874
rect 2050 3873 2087 3874
rect 2146 3873 2183 3874
rect 1466 3820 1507 3821
rect 1358 3813 1507 3820
rect 1358 3793 1476 3813
rect 1496 3793 1507 3813
rect 1358 3785 1507 3793
rect 1574 3817 1933 3821
rect 1574 3812 1896 3817
rect 1574 3788 1687 3812
rect 1711 3793 1896 3812
rect 1920 3793 1933 3817
rect 1711 3788 1933 3793
rect 1574 3785 1933 3788
rect 1995 3785 2030 3822
rect 2098 3819 2198 3822
rect 2098 3815 2165 3819
rect 2098 3789 2110 3815
rect 2136 3793 2165 3815
rect 2191 3793 2198 3819
rect 2136 3789 2198 3793
rect 2098 3785 2198 3789
rect 108 3770 156 3772
rect 108 3752 119 3770
rect 137 3752 156 3770
rect 1574 3764 1605 3785
rect 1995 3764 2031 3785
rect 1417 3763 1454 3764
rect 108 3743 156 3752
rect 109 3742 156 3743
rect 422 3747 532 3761
rect 422 3744 465 3747
rect 422 3739 426 3744
rect 344 3717 426 3739
rect 455 3717 465 3744
rect 493 3720 500 3747
rect 529 3739 532 3747
rect 1416 3754 1454 3763
rect 529 3720 594 3739
rect 1416 3734 1425 3754
rect 1445 3734 1454 3754
rect 493 3717 594 3720
rect 344 3715 594 3717
rect 112 3679 149 3680
rect 108 3676 149 3679
rect 108 3671 150 3676
rect 108 3653 121 3671
rect 139 3653 150 3671
rect 108 3639 150 3653
rect 188 3639 235 3643
rect 108 3633 235 3639
rect 108 3604 196 3633
rect 225 3604 235 3633
rect 344 3636 381 3715
rect 422 3702 532 3715
rect 496 3646 527 3647
rect 344 3616 353 3636
rect 373 3616 381 3636
rect 344 3606 381 3616
rect 440 3636 527 3646
rect 440 3616 449 3636
rect 469 3616 527 3636
rect 440 3607 527 3616
rect 440 3606 477 3607
rect 108 3600 235 3604
rect 108 3583 147 3600
rect 188 3599 235 3600
rect 108 3565 119 3583
rect 137 3565 147 3583
rect 108 3556 147 3565
rect 109 3555 146 3556
rect 496 3554 527 3607
rect 557 3636 594 3715
rect 765 3712 1158 3732
rect 1178 3712 1181 3732
rect 1416 3726 1454 3734
rect 1520 3758 1605 3764
rect 1630 3763 1667 3764
rect 1520 3738 1528 3758
rect 1548 3738 1605 3758
rect 1520 3730 1605 3738
rect 1629 3754 1667 3763
rect 1629 3734 1638 3754
rect 1658 3734 1667 3754
rect 1520 3729 1556 3730
rect 1629 3726 1667 3734
rect 1733 3758 1818 3764
rect 1838 3763 1875 3764
rect 1733 3738 1741 3758
rect 1761 3757 1818 3758
rect 1761 3738 1790 3757
rect 1733 3737 1790 3738
rect 1811 3737 1818 3757
rect 1733 3730 1818 3737
rect 1837 3754 1875 3763
rect 1837 3734 1846 3754
rect 1866 3734 1875 3754
rect 1733 3729 1769 3730
rect 1837 3726 1875 3734
rect 1941 3758 2085 3764
rect 1941 3738 1949 3758
rect 1969 3756 2057 3758
rect 1969 3738 1998 3756
rect 1941 3735 1998 3738
rect 2025 3738 2057 3756
rect 2077 3738 2085 3758
rect 2025 3735 2085 3738
rect 1941 3730 2085 3735
rect 1941 3729 1977 3730
rect 2049 3729 2085 3730
rect 2151 3763 2188 3764
rect 2151 3762 2189 3763
rect 2151 3754 2215 3762
rect 2151 3734 2160 3754
rect 2180 3740 2215 3754
rect 2235 3740 2238 3760
rect 2180 3735 2238 3740
rect 2180 3734 2215 3735
rect 765 3707 1181 3712
rect 765 3706 1106 3707
rect 709 3646 740 3647
rect 557 3616 566 3636
rect 586 3616 594 3636
rect 557 3606 594 3616
rect 653 3639 740 3646
rect 653 3636 714 3639
rect 653 3616 662 3636
rect 682 3619 714 3636
rect 735 3619 740 3639
rect 682 3616 740 3619
rect 653 3609 740 3616
rect 765 3636 802 3706
rect 1068 3705 1105 3706
rect 1417 3697 1454 3726
rect 1418 3695 1454 3697
rect 1630 3695 1667 3726
rect 1418 3673 1667 3695
rect 1838 3694 1875 3726
rect 2151 3722 2215 3734
rect 2255 3696 2282 3874
rect 2650 3867 2679 4045
rect 2719 4007 2783 4019
rect 3059 4015 3096 4047
rect 3267 4046 3516 4068
rect 3267 4015 3304 4046
rect 3480 4044 3516 4046
rect 3480 4015 3517 4044
rect 3829 4035 3866 4036
rect 4132 4035 4169 4105
rect 4194 4125 4281 4132
rect 4194 4122 4252 4125
rect 4194 4102 4199 4122
rect 4220 4105 4252 4122
rect 4272 4105 4281 4125
rect 4220 4102 4281 4105
rect 4194 4095 4281 4102
rect 4340 4125 4377 4135
rect 4340 4105 4348 4125
rect 4368 4105 4377 4125
rect 4194 4094 4225 4095
rect 3828 4034 4169 4035
rect 3753 4029 4169 4034
rect 2719 4006 2754 4007
rect 2696 4001 2754 4006
rect 2696 3981 2699 4001
rect 2719 3987 2754 4001
rect 2774 3987 2783 4007
rect 2719 3979 2783 3987
rect 2745 3978 2783 3979
rect 2746 3977 2783 3978
rect 2849 4011 2885 4012
rect 2957 4011 2993 4012
rect 2849 4003 2993 4011
rect 2849 3983 2857 4003
rect 2877 3983 2965 4003
rect 2985 3983 2993 4003
rect 2849 3977 2993 3983
rect 3059 4007 3097 4015
rect 3165 4011 3201 4012
rect 3059 3987 3068 4007
rect 3088 3987 3097 4007
rect 3059 3978 3097 3987
rect 3116 4004 3201 4011
rect 3116 3984 3123 4004
rect 3144 4003 3201 4004
rect 3144 3984 3173 4003
rect 3116 3983 3173 3984
rect 3193 3983 3201 4003
rect 3059 3977 3096 3978
rect 3116 3977 3201 3983
rect 3267 4007 3305 4015
rect 3378 4011 3414 4012
rect 3267 3987 3276 4007
rect 3296 3987 3305 4007
rect 3267 3978 3305 3987
rect 3329 4003 3414 4011
rect 3329 3983 3386 4003
rect 3406 3983 3414 4003
rect 3267 3977 3304 3978
rect 3329 3977 3414 3983
rect 3480 4007 3518 4015
rect 3753 4009 3756 4029
rect 3776 4009 4169 4029
rect 4340 4026 4377 4105
rect 4407 4134 4438 4187
rect 4788 4185 4825 4186
rect 4787 4176 4826 4185
rect 4787 4158 4797 4176
rect 4815 4158 4826 4176
rect 5167 4174 5204 4178
rect 4699 4141 4746 4142
rect 4787 4141 4826 4158
rect 4699 4137 4826 4141
rect 4457 4134 4494 4135
rect 4407 4125 4494 4134
rect 4407 4105 4465 4125
rect 4485 4105 4494 4125
rect 4407 4095 4494 4105
rect 4553 4125 4590 4135
rect 4553 4105 4561 4125
rect 4581 4105 4590 4125
rect 4407 4094 4438 4095
rect 4402 4026 4512 4039
rect 4553 4026 4590 4105
rect 4699 4108 4709 4137
rect 4738 4108 4826 4137
rect 4699 4102 4826 4108
rect 4699 4098 4746 4102
rect 4784 4088 4826 4102
rect 4784 4070 4795 4088
rect 4813 4070 4826 4088
rect 4784 4065 4826 4070
rect 4785 4062 4826 4065
rect 5164 4169 5204 4174
rect 5164 4151 5176 4169
rect 5194 4151 5204 4169
rect 4785 4061 4822 4062
rect 4340 4024 4590 4026
rect 4340 4021 4441 4024
rect 3480 3987 3489 4007
rect 3509 3987 3518 4007
rect 4340 4002 4405 4021
rect 3480 3978 3518 3987
rect 4402 3994 4405 4002
rect 4434 3994 4441 4021
rect 4469 3997 4479 4024
rect 4508 4002 4590 4024
rect 4508 3997 4512 4002
rect 4469 3994 4512 3997
rect 4402 3980 4512 3994
rect 4778 3998 4825 3999
rect 4778 3989 4826 3998
rect 3480 3977 3517 3978
rect 2903 3956 2939 3977
rect 3329 3956 3360 3977
rect 4778 3971 4797 3989
rect 4815 3971 4826 3989
rect 4778 3969 4826 3971
rect 2736 3952 2836 3956
rect 2736 3948 2798 3952
rect 2736 3922 2743 3948
rect 2769 3926 2798 3948
rect 2824 3926 2836 3952
rect 2769 3922 2836 3926
rect 2736 3919 2836 3922
rect 2904 3919 2939 3956
rect 3001 3953 3360 3956
rect 3001 3948 3223 3953
rect 3001 3924 3014 3948
rect 3038 3929 3223 3948
rect 3247 3929 3360 3953
rect 3038 3924 3360 3929
rect 3001 3920 3360 3924
rect 3427 3948 3576 3956
rect 3427 3928 3438 3948
rect 3458 3928 3576 3948
rect 3427 3921 3576 3928
rect 3427 3920 3468 3921
rect 2903 3880 2939 3919
rect 2751 3867 2788 3868
rect 2847 3867 2884 3868
rect 2903 3867 2910 3880
rect 2650 3858 2789 3867
rect 2650 3838 2760 3858
rect 2780 3838 2789 3858
rect 2650 3831 2789 3838
rect 2847 3858 2910 3867
rect 2847 3838 2856 3858
rect 2876 3842 2910 3858
rect 2933 3867 2939 3880
rect 2958 3867 2995 3868
rect 2933 3858 2995 3867
rect 2933 3842 2966 3858
rect 2876 3838 2966 3842
rect 2986 3838 2995 3858
rect 2650 3829 2747 3831
rect 2650 3828 2679 3829
rect 2847 3828 2995 3838
rect 3054 3858 3091 3868
rect 3166 3867 3203 3868
rect 3147 3865 3203 3867
rect 3054 3838 3062 3858
rect 3082 3838 3091 3858
rect 2903 3827 2939 3828
rect 2751 3768 2788 3769
rect 3054 3768 3091 3838
rect 3116 3858 3203 3865
rect 3116 3855 3174 3858
rect 3116 3835 3121 3855
rect 3142 3838 3174 3855
rect 3194 3838 3203 3858
rect 3142 3835 3203 3838
rect 3116 3828 3203 3835
rect 3262 3858 3299 3868
rect 3262 3838 3270 3858
rect 3290 3838 3299 3858
rect 3116 3827 3147 3828
rect 2750 3767 3091 3768
rect 2675 3763 3091 3767
rect 2675 3762 3052 3763
rect 2675 3742 2678 3762
rect 2698 3746 3052 3762
rect 3072 3746 3091 3763
rect 2698 3742 3091 3746
rect 3262 3759 3299 3838
rect 3329 3867 3360 3920
rect 4140 3912 4178 3914
rect 4787 3912 4826 3969
rect 4140 3879 4826 3912
rect 3379 3867 3416 3868
rect 3329 3858 3416 3867
rect 3329 3838 3387 3858
rect 3407 3838 3416 3858
rect 3329 3828 3416 3838
rect 3475 3858 3512 3868
rect 3475 3838 3483 3858
rect 3503 3838 3512 3858
rect 3329 3827 3360 3828
rect 3324 3759 3434 3772
rect 3475 3759 3512 3838
rect 3262 3757 3512 3759
rect 3262 3754 3363 3757
rect 3262 3735 3327 3754
rect 3324 3727 3327 3735
rect 3356 3727 3363 3754
rect 3391 3730 3401 3757
rect 3430 3735 3512 3757
rect 3732 3791 3900 3792
rect 4140 3791 4178 3879
rect 4439 3877 4486 3879
rect 4786 3855 4826 3879
rect 3732 3768 4178 3791
rect 4404 3822 4515 3837
rect 4404 3820 4446 3822
rect 4404 3800 4411 3820
rect 4430 3800 4446 3820
rect 4404 3792 4446 3800
rect 4474 3820 4515 3822
rect 4474 3800 4488 3820
rect 4507 3800 4515 3820
rect 4787 3811 4826 3855
rect 4474 3792 4515 3800
rect 4404 3786 4515 3792
rect 3732 3765 4176 3768
rect 3732 3763 3900 3765
rect 3430 3730 3434 3735
rect 3391 3727 3434 3730
rect 3324 3713 3434 3727
rect 2114 3694 2282 3696
rect 1835 3687 2282 3694
rect 1499 3667 1610 3673
rect 1499 3659 1540 3667
rect 917 3646 953 3647
rect 765 3616 774 3636
rect 794 3616 802 3636
rect 653 3607 709 3609
rect 653 3606 690 3607
rect 765 3606 802 3616
rect 861 3636 1009 3646
rect 1109 3643 1205 3645
rect 861 3616 870 3636
rect 890 3616 980 3636
rect 1000 3616 1009 3636
rect 861 3607 1009 3616
rect 1067 3636 1205 3643
rect 1067 3616 1076 3636
rect 1096 3616 1205 3636
rect 1499 3639 1507 3659
rect 1526 3639 1540 3659
rect 1499 3637 1540 3639
rect 1568 3659 1610 3667
rect 1568 3639 1584 3659
rect 1603 3639 1610 3659
rect 1835 3660 1860 3687
rect 1891 3668 2282 3687
rect 1891 3660 1940 3668
rect 2114 3667 2282 3668
rect 1835 3658 1940 3660
rect 1568 3637 1610 3639
rect 1499 3622 1610 3637
rect 1067 3607 1205 3616
rect 861 3606 898 3607
rect 917 3555 953 3607
rect 972 3606 1009 3607
rect 1068 3606 1105 3607
rect 388 3553 429 3554
rect 280 3546 429 3553
rect 280 3526 398 3546
rect 418 3526 429 3546
rect 280 3518 429 3526
rect 496 3550 855 3554
rect 496 3545 818 3550
rect 496 3521 609 3545
rect 633 3526 818 3545
rect 842 3526 855 3550
rect 633 3521 855 3526
rect 496 3518 855 3521
rect 917 3518 952 3555
rect 1020 3552 1120 3555
rect 1020 3548 1087 3552
rect 1020 3522 1032 3548
rect 1058 3526 1087 3548
rect 1113 3526 1120 3552
rect 1058 3522 1120 3526
rect 1020 3518 1120 3522
rect 496 3497 527 3518
rect 917 3497 953 3518
rect 339 3496 376 3497
rect 113 3493 147 3494
rect 112 3484 149 3493
rect 112 3466 121 3484
rect 139 3466 149 3484
rect 112 3456 149 3466
rect 338 3487 376 3496
rect 338 3467 347 3487
rect 367 3467 376 3487
rect 338 3459 376 3467
rect 442 3491 527 3497
rect 552 3496 589 3497
rect 442 3471 450 3491
rect 470 3471 527 3491
rect 442 3463 527 3471
rect 551 3487 589 3496
rect 551 3467 560 3487
rect 580 3467 589 3487
rect 442 3462 478 3463
rect 551 3459 589 3467
rect 655 3491 740 3497
rect 760 3496 797 3497
rect 655 3471 663 3491
rect 683 3490 740 3491
rect 683 3471 712 3490
rect 655 3470 712 3471
rect 733 3470 740 3490
rect 655 3463 740 3470
rect 759 3487 797 3496
rect 759 3467 768 3487
rect 788 3467 797 3487
rect 655 3462 691 3463
rect 759 3459 797 3467
rect 863 3491 1007 3497
rect 863 3471 871 3491
rect 891 3490 979 3491
rect 891 3471 922 3490
rect 863 3470 922 3471
rect 947 3471 979 3490
rect 999 3471 1007 3491
rect 947 3470 1007 3471
rect 863 3463 1007 3470
rect 863 3462 899 3463
rect 971 3462 1007 3463
rect 1073 3496 1110 3497
rect 1073 3495 1111 3496
rect 1073 3487 1137 3495
rect 1073 3467 1082 3487
rect 1102 3473 1137 3487
rect 1157 3473 1160 3493
rect 1102 3468 1160 3473
rect 1102 3467 1137 3468
rect 113 3428 147 3456
rect 339 3430 376 3459
rect 340 3428 376 3430
rect 552 3428 589 3459
rect 113 3427 285 3428
rect 113 3395 299 3427
rect 340 3406 589 3428
rect 760 3427 797 3459
rect 1073 3455 1137 3467
rect 1177 3429 1204 3607
rect 3732 3585 3759 3763
rect 3799 3725 3863 3737
rect 4139 3733 4176 3765
rect 4347 3764 4596 3786
rect 4347 3733 4384 3764
rect 4560 3762 4596 3764
rect 4560 3733 4597 3762
rect 3799 3724 3834 3725
rect 3776 3719 3834 3724
rect 3776 3699 3779 3719
rect 3799 3705 3834 3719
rect 3854 3705 3863 3725
rect 3799 3697 3863 3705
rect 3825 3696 3863 3697
rect 3826 3695 3863 3696
rect 3929 3729 3965 3730
rect 4037 3729 4073 3730
rect 3929 3724 4073 3729
rect 3929 3721 3991 3724
rect 3929 3701 3937 3721
rect 3957 3704 3991 3721
rect 4014 3721 4073 3724
rect 4014 3704 4045 3721
rect 3957 3701 4045 3704
rect 4065 3701 4073 3721
rect 3929 3695 4073 3701
rect 4139 3725 4177 3733
rect 4245 3729 4281 3730
rect 4139 3705 4148 3725
rect 4168 3705 4177 3725
rect 4139 3696 4177 3705
rect 4196 3722 4281 3729
rect 4196 3702 4203 3722
rect 4224 3721 4281 3722
rect 4224 3702 4253 3721
rect 4196 3701 4253 3702
rect 4273 3701 4281 3721
rect 4139 3695 4176 3696
rect 4196 3695 4281 3701
rect 4347 3725 4385 3733
rect 4458 3729 4494 3730
rect 4347 3705 4356 3725
rect 4376 3705 4385 3725
rect 4347 3696 4385 3705
rect 4409 3721 4494 3729
rect 4409 3701 4466 3721
rect 4486 3701 4494 3721
rect 4347 3695 4384 3696
rect 4409 3695 4494 3701
rect 4560 3725 4598 3733
rect 4560 3705 4569 3725
rect 4589 3705 4598 3725
rect 4560 3696 4598 3705
rect 4560 3695 4597 3696
rect 3983 3674 4019 3695
rect 4409 3674 4440 3695
rect 3816 3670 3916 3674
rect 3816 3666 3878 3670
rect 3816 3640 3823 3666
rect 3849 3644 3878 3666
rect 3904 3644 3916 3670
rect 3849 3640 3916 3644
rect 3816 3637 3916 3640
rect 3984 3637 4019 3674
rect 4081 3671 4440 3674
rect 4081 3666 4303 3671
rect 4081 3642 4094 3666
rect 4118 3647 4303 3666
rect 4327 3647 4440 3671
rect 4118 3642 4440 3647
rect 4081 3638 4440 3642
rect 4507 3666 4656 3674
rect 4507 3646 4518 3666
rect 4538 3646 4656 3666
rect 4507 3639 4656 3646
rect 4507 3638 4548 3639
rect 3831 3585 3868 3586
rect 3927 3585 3964 3586
rect 3983 3585 4019 3637
rect 4038 3585 4075 3586
rect 3731 3576 3869 3585
rect 3731 3556 3840 3576
rect 3860 3556 3869 3576
rect 3731 3549 3869 3556
rect 3927 3576 4075 3585
rect 3927 3556 3936 3576
rect 3956 3556 4046 3576
rect 4066 3556 4075 3576
rect 3731 3547 3827 3549
rect 3927 3546 4075 3556
rect 4134 3576 4171 3586
rect 4246 3585 4283 3586
rect 4227 3583 4283 3585
rect 4134 3556 4142 3576
rect 4162 3556 4171 3576
rect 3983 3545 4019 3546
rect 1360 3503 1470 3517
rect 1360 3500 1403 3503
rect 1360 3495 1364 3500
rect 1036 3427 1204 3429
rect 760 3421 1204 3427
rect 113 3363 147 3395
rect 109 3354 147 3363
rect 109 3336 119 3354
rect 137 3336 147 3354
rect 109 3330 147 3336
rect 265 3332 299 3395
rect 421 3400 532 3406
rect 421 3392 462 3400
rect 421 3372 429 3392
rect 448 3372 462 3392
rect 421 3370 462 3372
rect 490 3392 532 3400
rect 490 3372 506 3392
rect 525 3372 532 3392
rect 490 3370 532 3372
rect 421 3355 532 3370
rect 759 3401 1204 3421
rect 759 3332 797 3401
rect 1036 3400 1204 3401
rect 1282 3473 1364 3495
rect 1393 3473 1403 3500
rect 1431 3476 1438 3503
rect 1467 3495 1470 3503
rect 3465 3512 3576 3527
rect 3465 3510 3507 3512
rect 1467 3476 1532 3495
rect 1431 3473 1532 3476
rect 1282 3471 1532 3473
rect 1282 3392 1319 3471
rect 1360 3458 1470 3471
rect 1434 3402 1465 3403
rect 1282 3372 1291 3392
rect 1311 3372 1319 3392
rect 1282 3362 1319 3372
rect 1378 3392 1465 3402
rect 1378 3372 1387 3392
rect 1407 3372 1465 3392
rect 1378 3363 1465 3372
rect 1378 3362 1415 3363
rect 109 3326 146 3330
rect 265 3321 797 3332
rect 264 3305 797 3321
rect 1434 3310 1465 3363
rect 1495 3392 1532 3471
rect 1703 3481 2096 3488
rect 1703 3464 1711 3481
rect 1743 3468 2096 3481
rect 2116 3468 2119 3488
rect 3198 3483 3239 3492
rect 1743 3464 2119 3468
rect 1703 3463 2119 3464
rect 2793 3481 2961 3482
rect 3198 3481 3207 3483
rect 1703 3462 2044 3463
rect 1647 3402 1678 3403
rect 1495 3372 1504 3392
rect 1524 3372 1532 3392
rect 1495 3362 1532 3372
rect 1591 3395 1678 3402
rect 1591 3392 1652 3395
rect 1591 3372 1600 3392
rect 1620 3375 1652 3392
rect 1673 3375 1678 3395
rect 1620 3372 1678 3375
rect 1591 3365 1678 3372
rect 1703 3392 1740 3462
rect 2006 3461 2043 3462
rect 2793 3461 3207 3481
rect 3233 3461 3239 3483
rect 3465 3490 3472 3510
rect 3491 3490 3507 3510
rect 3465 3482 3507 3490
rect 3535 3510 3576 3512
rect 3535 3490 3549 3510
rect 3568 3490 3576 3510
rect 3535 3482 3576 3490
rect 3831 3486 3868 3487
rect 4134 3486 4171 3556
rect 4196 3576 4283 3583
rect 4196 3573 4254 3576
rect 4196 3553 4201 3573
rect 4222 3556 4254 3573
rect 4274 3556 4283 3576
rect 4222 3553 4283 3556
rect 4196 3546 4283 3553
rect 4342 3576 4379 3586
rect 4342 3556 4350 3576
rect 4370 3556 4379 3576
rect 4196 3545 4227 3546
rect 3830 3485 4171 3486
rect 3465 3476 3576 3482
rect 3755 3480 4171 3485
rect 2793 3455 3239 3461
rect 2793 3453 2961 3455
rect 1855 3402 1891 3403
rect 1703 3372 1712 3392
rect 1732 3372 1740 3392
rect 1591 3363 1647 3365
rect 1591 3362 1628 3363
rect 1703 3362 1740 3372
rect 1799 3392 1947 3402
rect 2047 3399 2143 3401
rect 1799 3372 1808 3392
rect 1828 3387 1918 3392
rect 1828 3372 1863 3387
rect 1799 3363 1863 3372
rect 1799 3362 1836 3363
rect 1855 3346 1863 3363
rect 1884 3372 1918 3387
rect 1938 3372 1947 3392
rect 1884 3363 1947 3372
rect 2005 3392 2143 3399
rect 2005 3372 2014 3392
rect 2034 3372 2143 3392
rect 2005 3363 2143 3372
rect 1884 3346 1891 3363
rect 1910 3362 1947 3363
rect 2006 3362 2043 3363
rect 1855 3311 1891 3346
rect 1326 3309 1367 3310
rect 264 3304 778 3305
rect 1218 3302 1367 3309
rect 1218 3282 1336 3302
rect 1356 3282 1367 3302
rect 1218 3274 1367 3282
rect 1434 3306 1793 3310
rect 1434 3301 1756 3306
rect 1434 3277 1547 3301
rect 1571 3282 1756 3301
rect 1780 3282 1793 3306
rect 1571 3277 1793 3282
rect 1434 3274 1793 3277
rect 1855 3274 1890 3311
rect 1958 3308 2058 3311
rect 1958 3304 2025 3308
rect 1958 3278 1970 3304
rect 1996 3282 2025 3304
rect 2051 3282 2058 3308
rect 1996 3278 2058 3282
rect 1958 3274 2058 3278
rect 112 3263 149 3264
rect 110 3255 150 3263
rect 110 3237 121 3255
rect 139 3237 150 3255
rect 1434 3253 1465 3274
rect 1855 3253 1891 3274
rect 1277 3252 1314 3253
rect 110 3189 150 3237
rect 1276 3243 1314 3252
rect 1276 3223 1285 3243
rect 1305 3223 1314 3243
rect 1276 3215 1314 3223
rect 1380 3247 1465 3253
rect 1490 3252 1527 3253
rect 1380 3227 1388 3247
rect 1408 3227 1465 3247
rect 1380 3219 1465 3227
rect 1489 3243 1527 3252
rect 1489 3223 1498 3243
rect 1518 3223 1527 3243
rect 1380 3218 1416 3219
rect 1489 3215 1527 3223
rect 1593 3247 1678 3253
rect 1698 3252 1735 3253
rect 1593 3227 1601 3247
rect 1621 3246 1678 3247
rect 1621 3227 1650 3246
rect 1593 3226 1650 3227
rect 1671 3226 1678 3246
rect 1593 3219 1678 3226
rect 1697 3243 1735 3252
rect 1697 3223 1706 3243
rect 1726 3223 1735 3243
rect 1593 3218 1629 3219
rect 1697 3215 1735 3223
rect 1801 3247 1945 3253
rect 1801 3227 1809 3247
rect 1829 3227 1917 3247
rect 1937 3227 1945 3247
rect 1801 3219 1945 3227
rect 1801 3218 1837 3219
rect 1909 3218 1945 3219
rect 2011 3252 2048 3253
rect 2011 3251 2049 3252
rect 2011 3243 2075 3251
rect 2011 3223 2020 3243
rect 2040 3229 2075 3243
rect 2095 3229 2098 3249
rect 2040 3224 2098 3229
rect 2040 3223 2075 3224
rect 421 3193 531 3207
rect 421 3190 464 3193
rect 110 3182 235 3189
rect 421 3185 425 3190
rect 110 3163 202 3182
rect 227 3163 235 3182
rect 110 3153 235 3163
rect 343 3163 425 3185
rect 454 3163 464 3190
rect 492 3166 499 3193
rect 528 3185 531 3193
rect 1277 3186 1314 3215
rect 528 3166 593 3185
rect 1278 3184 1314 3186
rect 1490 3184 1527 3215
rect 1698 3188 1735 3215
rect 2011 3211 2075 3223
rect 492 3163 593 3166
rect 343 3161 593 3163
rect 110 3133 150 3153
rect 109 3124 150 3133
rect 109 3106 119 3124
rect 137 3106 150 3124
rect 109 3097 150 3106
rect 109 3096 146 3097
rect 343 3082 380 3161
rect 421 3148 531 3161
rect 495 3092 526 3093
rect 343 3062 352 3082
rect 372 3062 380 3082
rect 343 3052 380 3062
rect 439 3082 526 3092
rect 439 3062 448 3082
rect 468 3062 526 3082
rect 439 3053 526 3062
rect 439 3052 476 3053
rect 112 3030 149 3034
rect 109 3025 149 3030
rect 109 3007 121 3025
rect 139 3007 149 3025
rect 109 2827 149 3007
rect 495 3000 526 3053
rect 556 3082 593 3161
rect 764 3158 1157 3178
rect 1177 3158 1180 3178
rect 1278 3162 1527 3184
rect 1696 3183 1737 3188
rect 2115 3185 2142 3363
rect 2793 3275 2820 3453
rect 3198 3450 3239 3455
rect 3408 3454 3657 3476
rect 3755 3460 3758 3480
rect 3778 3460 4171 3480
rect 4342 3477 4379 3556
rect 4409 3585 4440 3638
rect 4786 3631 4826 3811
rect 5164 3971 5204 4151
rect 5550 4144 5581 4197
rect 5611 4226 5648 4305
rect 5819 4302 6212 4322
rect 6232 4302 6235 4322
rect 6333 4306 6582 4328
rect 6751 4327 6792 4332
rect 7170 4329 7197 4507
rect 7848 4419 7875 4597
rect 8253 4594 8294 4599
rect 8463 4598 8712 4620
rect 8810 4604 8813 4624
rect 8833 4604 9226 4624
rect 9397 4621 9434 4700
rect 9464 4729 9495 4782
rect 9841 4775 9881 4955
rect 9841 4757 9851 4775
rect 9869 4757 9881 4775
rect 9841 4752 9881 4757
rect 9841 4748 9878 4752
rect 9514 4729 9551 4730
rect 9464 4720 9551 4729
rect 9464 4700 9522 4720
rect 9542 4700 9551 4720
rect 9464 4690 9551 4700
rect 9610 4720 9647 4730
rect 9610 4700 9618 4720
rect 9638 4700 9647 4720
rect 9464 4689 9495 4690
rect 9459 4621 9569 4634
rect 9610 4621 9647 4700
rect 9844 4685 9881 4686
rect 9840 4676 9881 4685
rect 9840 4658 9853 4676
rect 9871 4658 9881 4676
rect 9840 4649 9881 4658
rect 9840 4629 9880 4649
rect 9397 4619 9647 4621
rect 9397 4616 9498 4619
rect 7915 4559 7979 4571
rect 8255 4567 8292 4594
rect 8463 4567 8500 4598
rect 8676 4596 8712 4598
rect 9397 4597 9462 4616
rect 8676 4567 8713 4596
rect 9459 4589 9462 4597
rect 9491 4589 9498 4616
rect 9526 4592 9536 4619
rect 9565 4597 9647 4619
rect 9755 4619 9880 4629
rect 9755 4600 9763 4619
rect 9788 4600 9880 4619
rect 9565 4592 9569 4597
rect 9755 4593 9880 4600
rect 9526 4589 9569 4592
rect 9459 4575 9569 4589
rect 7915 4558 7950 4559
rect 7892 4553 7950 4558
rect 7892 4533 7895 4553
rect 7915 4539 7950 4553
rect 7970 4539 7979 4559
rect 7915 4531 7979 4539
rect 7941 4530 7979 4531
rect 7942 4529 7979 4530
rect 8045 4563 8081 4564
rect 8153 4563 8189 4564
rect 8045 4555 8189 4563
rect 8045 4535 8053 4555
rect 8073 4535 8161 4555
rect 8181 4535 8189 4555
rect 8045 4529 8189 4535
rect 8255 4559 8293 4567
rect 8361 4563 8397 4564
rect 8255 4539 8264 4559
rect 8284 4539 8293 4559
rect 8255 4530 8293 4539
rect 8312 4556 8397 4563
rect 8312 4536 8319 4556
rect 8340 4555 8397 4556
rect 8340 4536 8369 4555
rect 8312 4535 8369 4536
rect 8389 4535 8397 4555
rect 8255 4529 8292 4530
rect 8312 4529 8397 4535
rect 8463 4559 8501 4567
rect 8574 4563 8610 4564
rect 8463 4539 8472 4559
rect 8492 4539 8501 4559
rect 8463 4530 8501 4539
rect 8525 4555 8610 4563
rect 8525 4535 8582 4555
rect 8602 4535 8610 4555
rect 8463 4529 8500 4530
rect 8525 4529 8610 4535
rect 8676 4559 8714 4567
rect 8676 4539 8685 4559
rect 8705 4539 8714 4559
rect 8676 4530 8714 4539
rect 9840 4545 9880 4593
rect 8676 4529 8713 4530
rect 8099 4508 8135 4529
rect 8525 4508 8556 4529
rect 9840 4527 9851 4545
rect 9869 4527 9880 4545
rect 9840 4519 9880 4527
rect 9841 4518 9878 4519
rect 7932 4504 8032 4508
rect 7932 4500 7994 4504
rect 7932 4474 7939 4500
rect 7965 4478 7994 4500
rect 8020 4478 8032 4504
rect 7965 4474 8032 4478
rect 7932 4471 8032 4474
rect 8100 4471 8135 4508
rect 8197 4505 8556 4508
rect 8197 4500 8419 4505
rect 8197 4476 8210 4500
rect 8234 4481 8419 4500
rect 8443 4481 8556 4505
rect 8234 4476 8556 4481
rect 8197 4472 8556 4476
rect 8623 4500 8772 4508
rect 8623 4480 8634 4500
rect 8654 4480 8772 4500
rect 8623 4473 8772 4480
rect 9212 4477 9726 4478
rect 8623 4472 8664 4473
rect 8099 4436 8135 4471
rect 7947 4419 7984 4420
rect 8043 4419 8080 4420
rect 8099 4419 8106 4436
rect 7847 4410 7985 4419
rect 7847 4390 7956 4410
rect 7976 4390 7985 4410
rect 7847 4383 7985 4390
rect 8043 4410 8106 4419
rect 8043 4390 8052 4410
rect 8072 4395 8106 4410
rect 8127 4419 8135 4436
rect 8154 4419 8191 4420
rect 8127 4410 8191 4419
rect 8127 4395 8162 4410
rect 8072 4390 8162 4395
rect 8182 4390 8191 4410
rect 7847 4381 7943 4383
rect 8043 4380 8191 4390
rect 8250 4410 8287 4420
rect 8362 4419 8399 4420
rect 8343 4417 8399 4419
rect 8250 4390 8258 4410
rect 8278 4390 8287 4410
rect 8099 4379 8135 4380
rect 7029 4327 7197 4329
rect 6751 4321 7197 4327
rect 5819 4297 6235 4302
rect 6414 4300 6525 4306
rect 5819 4296 6160 4297
rect 5763 4236 5794 4237
rect 5611 4206 5620 4226
rect 5640 4206 5648 4226
rect 5611 4196 5648 4206
rect 5707 4229 5794 4236
rect 5707 4226 5768 4229
rect 5707 4206 5716 4226
rect 5736 4209 5768 4226
rect 5789 4209 5794 4229
rect 5736 4206 5794 4209
rect 5707 4199 5794 4206
rect 5819 4226 5856 4296
rect 6122 4295 6159 4296
rect 6414 4292 6455 4300
rect 6414 4272 6422 4292
rect 6441 4272 6455 4292
rect 6414 4270 6455 4272
rect 6483 4292 6525 4300
rect 6483 4272 6499 4292
rect 6518 4272 6525 4292
rect 6751 4299 6757 4321
rect 6783 4301 7197 4321
rect 7947 4320 7984 4321
rect 8250 4320 8287 4390
rect 8312 4410 8399 4417
rect 8312 4407 8370 4410
rect 8312 4387 8317 4407
rect 8338 4390 8370 4407
rect 8390 4390 8399 4410
rect 8338 4387 8399 4390
rect 8312 4380 8399 4387
rect 8458 4410 8495 4420
rect 8458 4390 8466 4410
rect 8486 4390 8495 4410
rect 8312 4379 8343 4380
rect 7946 4319 8287 4320
rect 6783 4299 6792 4301
rect 7029 4300 7197 4301
rect 7871 4318 8287 4319
rect 7871 4314 8247 4318
rect 6751 4290 6792 4299
rect 7871 4294 7874 4314
rect 7894 4301 8247 4314
rect 8279 4301 8287 4318
rect 7894 4294 8287 4301
rect 8458 4311 8495 4390
rect 8525 4419 8556 4472
rect 9193 4461 9726 4477
rect 9193 4450 9725 4461
rect 9844 4452 9881 4456
rect 8575 4419 8612 4420
rect 8525 4410 8612 4419
rect 8525 4390 8583 4410
rect 8603 4390 8612 4410
rect 8525 4380 8612 4390
rect 8671 4410 8708 4420
rect 8671 4390 8679 4410
rect 8699 4390 8708 4410
rect 8525 4379 8556 4380
rect 8520 4311 8630 4324
rect 8671 4311 8708 4390
rect 8458 4309 8708 4311
rect 8458 4306 8559 4309
rect 8458 4287 8523 4306
rect 6483 4270 6525 4272
rect 6414 4255 6525 4270
rect 8520 4279 8523 4287
rect 8552 4279 8559 4306
rect 8587 4282 8597 4309
rect 8626 4287 8708 4309
rect 8786 4381 8954 4382
rect 9193 4381 9231 4450
rect 8786 4361 9231 4381
rect 9458 4412 9569 4427
rect 9458 4410 9500 4412
rect 9458 4390 9465 4410
rect 9484 4390 9500 4410
rect 9458 4382 9500 4390
rect 9528 4410 9569 4412
rect 9528 4390 9542 4410
rect 9561 4390 9569 4410
rect 9528 4382 9569 4390
rect 9458 4376 9569 4382
rect 9691 4387 9725 4450
rect 9843 4446 9881 4452
rect 9843 4428 9853 4446
rect 9871 4428 9881 4446
rect 9843 4419 9881 4428
rect 9843 4387 9877 4419
rect 8786 4355 9230 4361
rect 8786 4353 8954 4355
rect 8626 4282 8630 4287
rect 8587 4279 8630 4282
rect 8520 4265 8630 4279
rect 5971 4236 6007 4237
rect 5819 4206 5828 4226
rect 5848 4206 5856 4226
rect 5707 4197 5763 4199
rect 5707 4196 5744 4197
rect 5819 4196 5856 4206
rect 5915 4226 6063 4236
rect 6163 4233 6259 4235
rect 5915 4206 5924 4226
rect 5944 4206 6034 4226
rect 6054 4206 6063 4226
rect 5915 4197 6063 4206
rect 6121 4226 6259 4233
rect 6121 4206 6130 4226
rect 6150 4206 6259 4226
rect 6121 4197 6259 4206
rect 5915 4196 5952 4197
rect 5971 4145 6007 4197
rect 6026 4196 6063 4197
rect 6122 4196 6159 4197
rect 5442 4143 5483 4144
rect 5334 4136 5483 4143
rect 5334 4116 5452 4136
rect 5472 4116 5483 4136
rect 5334 4108 5483 4116
rect 5550 4140 5909 4144
rect 5550 4135 5872 4140
rect 5550 4111 5663 4135
rect 5687 4116 5872 4135
rect 5896 4116 5909 4140
rect 5687 4111 5909 4116
rect 5550 4108 5909 4111
rect 5971 4108 6006 4145
rect 6074 4142 6174 4145
rect 6074 4138 6141 4142
rect 6074 4112 6086 4138
rect 6112 4116 6141 4138
rect 6167 4116 6174 4142
rect 6112 4112 6174 4116
rect 6074 4108 6174 4112
rect 5550 4087 5581 4108
rect 5971 4087 6007 4108
rect 5393 4086 5430 4087
rect 5392 4077 5430 4086
rect 5392 4057 5401 4077
rect 5421 4057 5430 4077
rect 5392 4049 5430 4057
rect 5496 4081 5581 4087
rect 5606 4086 5643 4087
rect 5496 4061 5504 4081
rect 5524 4061 5581 4081
rect 5496 4053 5581 4061
rect 5605 4077 5643 4086
rect 5605 4057 5614 4077
rect 5634 4057 5643 4077
rect 5496 4052 5532 4053
rect 5605 4049 5643 4057
rect 5709 4081 5794 4087
rect 5814 4086 5851 4087
rect 5709 4061 5717 4081
rect 5737 4080 5794 4081
rect 5737 4061 5766 4080
rect 5709 4060 5766 4061
rect 5787 4060 5794 4080
rect 5709 4053 5794 4060
rect 5813 4077 5851 4086
rect 5813 4057 5822 4077
rect 5842 4057 5851 4077
rect 5709 4052 5745 4053
rect 5813 4049 5851 4057
rect 5917 4081 6061 4087
rect 5917 4061 5925 4081
rect 5945 4078 6033 4081
rect 5945 4061 5976 4078
rect 5917 4058 5976 4061
rect 5999 4061 6033 4078
rect 6053 4061 6061 4081
rect 5999 4058 6061 4061
rect 5917 4053 6061 4058
rect 5917 4052 5953 4053
rect 6025 4052 6061 4053
rect 6127 4086 6164 4087
rect 6127 4085 6165 4086
rect 6127 4077 6191 4085
rect 6127 4057 6136 4077
rect 6156 4063 6191 4077
rect 6211 4063 6214 4083
rect 6156 4058 6214 4063
rect 6156 4057 6191 4058
rect 5393 4020 5430 4049
rect 5394 4018 5430 4020
rect 5606 4018 5643 4049
rect 5394 3996 5643 4018
rect 5814 4017 5851 4049
rect 6127 4045 6191 4057
rect 6231 4019 6258 4197
rect 8786 4175 8813 4353
rect 8853 4315 8917 4327
rect 9193 4323 9230 4355
rect 9401 4354 9650 4376
rect 9691 4355 9877 4387
rect 9705 4354 9877 4355
rect 9401 4323 9438 4354
rect 9614 4352 9650 4354
rect 9614 4323 9651 4352
rect 9843 4326 9877 4354
rect 8853 4314 8888 4315
rect 8830 4309 8888 4314
rect 8830 4289 8833 4309
rect 8853 4295 8888 4309
rect 8908 4295 8917 4315
rect 8853 4287 8917 4295
rect 8879 4286 8917 4287
rect 8880 4285 8917 4286
rect 8983 4319 9019 4320
rect 9091 4319 9127 4320
rect 8983 4312 9127 4319
rect 8983 4311 9043 4312
rect 8983 4291 8991 4311
rect 9011 4292 9043 4311
rect 9068 4311 9127 4312
rect 9068 4292 9099 4311
rect 9011 4291 9099 4292
rect 9119 4291 9127 4311
rect 8983 4285 9127 4291
rect 9193 4315 9231 4323
rect 9299 4319 9335 4320
rect 9193 4295 9202 4315
rect 9222 4295 9231 4315
rect 9193 4286 9231 4295
rect 9250 4312 9335 4319
rect 9250 4292 9257 4312
rect 9278 4311 9335 4312
rect 9278 4292 9307 4311
rect 9250 4291 9307 4292
rect 9327 4291 9335 4311
rect 9193 4285 9230 4286
rect 9250 4285 9335 4291
rect 9401 4315 9439 4323
rect 9512 4319 9548 4320
rect 9401 4295 9410 4315
rect 9430 4295 9439 4315
rect 9401 4286 9439 4295
rect 9463 4311 9548 4319
rect 9463 4291 9520 4311
rect 9540 4291 9548 4311
rect 9401 4285 9438 4286
rect 9463 4285 9548 4291
rect 9614 4315 9652 4323
rect 9614 4295 9623 4315
rect 9643 4295 9652 4315
rect 9614 4286 9652 4295
rect 9841 4316 9878 4326
rect 9841 4298 9851 4316
rect 9869 4298 9878 4316
rect 9841 4289 9878 4298
rect 9843 4288 9877 4289
rect 9614 4285 9651 4286
rect 9037 4264 9073 4285
rect 9463 4264 9494 4285
rect 8870 4260 8970 4264
rect 8870 4256 8932 4260
rect 8870 4230 8877 4256
rect 8903 4234 8932 4256
rect 8958 4234 8970 4260
rect 8903 4230 8970 4234
rect 8870 4227 8970 4230
rect 9038 4227 9073 4264
rect 9135 4261 9494 4264
rect 9135 4256 9357 4261
rect 9135 4232 9148 4256
rect 9172 4237 9357 4256
rect 9381 4237 9494 4261
rect 9172 4232 9494 4237
rect 9135 4228 9494 4232
rect 9561 4256 9710 4264
rect 9561 4236 9572 4256
rect 9592 4236 9710 4256
rect 9561 4229 9710 4236
rect 9561 4228 9602 4229
rect 8885 4175 8922 4176
rect 8981 4175 9018 4176
rect 9037 4175 9073 4227
rect 9092 4175 9129 4176
rect 8785 4166 8923 4175
rect 8380 4145 8491 4160
rect 8380 4143 8422 4145
rect 8050 4122 8155 4124
rect 7706 4114 7876 4115
rect 8050 4114 8099 4122
rect 7706 4095 8099 4114
rect 8130 4095 8155 4122
rect 8380 4123 8387 4143
rect 8406 4123 8422 4143
rect 8380 4115 8422 4123
rect 8450 4143 8491 4145
rect 8450 4123 8464 4143
rect 8483 4123 8491 4143
rect 8785 4146 8894 4166
rect 8914 4146 8923 4166
rect 8785 4139 8923 4146
rect 8981 4166 9129 4175
rect 8981 4146 8990 4166
rect 9010 4146 9100 4166
rect 9120 4146 9129 4166
rect 8785 4137 8881 4139
rect 8981 4136 9129 4146
rect 9188 4166 9225 4176
rect 9300 4175 9337 4176
rect 9281 4173 9337 4175
rect 9188 4146 9196 4166
rect 9216 4146 9225 4166
rect 9037 4135 9073 4136
rect 8450 4115 8491 4123
rect 8380 4109 8491 4115
rect 7706 4088 8155 4095
rect 7706 4086 7876 4088
rect 6556 4055 6666 4069
rect 6556 4052 6599 4055
rect 6556 4047 6560 4052
rect 6090 4017 6258 4019
rect 5814 4014 6258 4017
rect 5475 3990 5586 3996
rect 5475 3982 5516 3990
rect 5164 3927 5203 3971
rect 5475 3962 5483 3982
rect 5502 3962 5516 3982
rect 5475 3960 5516 3962
rect 5544 3982 5586 3990
rect 5544 3962 5560 3982
rect 5579 3962 5586 3982
rect 5544 3960 5586 3962
rect 5475 3945 5586 3960
rect 5812 3991 6258 4014
rect 5164 3903 5204 3927
rect 5504 3903 5551 3905
rect 5812 3903 5850 3991
rect 6090 3990 6258 3991
rect 6478 4025 6560 4047
rect 6589 4025 6599 4052
rect 6627 4028 6634 4055
rect 6663 4047 6666 4055
rect 6663 4028 6728 4047
rect 6627 4025 6728 4028
rect 6478 4023 6728 4025
rect 6478 3944 6515 4023
rect 6556 4010 6666 4023
rect 6630 3954 6661 3955
rect 6478 3924 6487 3944
rect 6507 3924 6515 3944
rect 6478 3914 6515 3924
rect 6574 3944 6661 3954
rect 6574 3924 6583 3944
rect 6603 3924 6661 3944
rect 6574 3915 6661 3924
rect 6574 3914 6611 3915
rect 5164 3870 5850 3903
rect 5164 3813 5203 3870
rect 5812 3868 5850 3870
rect 6630 3862 6661 3915
rect 6691 3944 6728 4023
rect 6899 4036 7292 4040
rect 6899 4019 6918 4036
rect 6938 4020 7292 4036
rect 7312 4020 7315 4040
rect 6938 4019 7315 4020
rect 6899 4015 7315 4019
rect 6899 4014 7240 4015
rect 6843 3954 6874 3955
rect 6691 3924 6700 3944
rect 6720 3924 6728 3944
rect 6691 3914 6728 3924
rect 6787 3947 6874 3954
rect 6787 3944 6848 3947
rect 6787 3924 6796 3944
rect 6816 3927 6848 3944
rect 6869 3927 6874 3947
rect 6816 3924 6874 3927
rect 6787 3917 6874 3924
rect 6899 3944 6936 4014
rect 7202 4013 7239 4014
rect 7051 3954 7087 3955
rect 6899 3924 6908 3944
rect 6928 3924 6936 3944
rect 6787 3915 6843 3917
rect 6787 3914 6824 3915
rect 6899 3914 6936 3924
rect 6995 3944 7143 3954
rect 7243 3951 7339 3953
rect 6995 3924 7004 3944
rect 7024 3924 7114 3944
rect 7134 3924 7143 3944
rect 6995 3915 7143 3924
rect 7201 3944 7339 3951
rect 7201 3924 7210 3944
rect 7230 3924 7339 3944
rect 7201 3915 7339 3924
rect 6995 3914 7032 3915
rect 7051 3863 7087 3915
rect 7106 3914 7143 3915
rect 7202 3914 7239 3915
rect 6522 3861 6563 3862
rect 6414 3854 6563 3861
rect 6414 3834 6532 3854
rect 6552 3834 6563 3854
rect 6414 3826 6563 3834
rect 6630 3858 6989 3862
rect 6630 3853 6952 3858
rect 6630 3829 6743 3853
rect 6767 3834 6952 3853
rect 6976 3834 6989 3858
rect 6767 3829 6989 3834
rect 6630 3826 6989 3829
rect 7051 3826 7086 3863
rect 7154 3860 7254 3863
rect 7154 3856 7221 3860
rect 7154 3830 7166 3856
rect 7192 3834 7221 3856
rect 7247 3834 7254 3860
rect 7192 3830 7254 3834
rect 7154 3826 7254 3830
rect 5164 3811 5212 3813
rect 5164 3793 5175 3811
rect 5193 3793 5212 3811
rect 6630 3805 6661 3826
rect 7051 3805 7087 3826
rect 6473 3804 6510 3805
rect 5164 3784 5212 3793
rect 5165 3783 5212 3784
rect 5478 3788 5588 3802
rect 5478 3785 5521 3788
rect 5478 3780 5482 3785
rect 5400 3758 5482 3780
rect 5511 3758 5521 3785
rect 5549 3761 5556 3788
rect 5585 3780 5588 3788
rect 6472 3795 6510 3804
rect 5585 3761 5650 3780
rect 6472 3775 6481 3795
rect 6501 3775 6510 3795
rect 5549 3758 5650 3761
rect 5400 3756 5650 3758
rect 5168 3720 5205 3721
rect 4786 3613 4796 3631
rect 4814 3613 4826 3631
rect 4786 3608 4826 3613
rect 5164 3717 5205 3720
rect 5164 3712 5206 3717
rect 5164 3694 5177 3712
rect 5195 3694 5206 3712
rect 5164 3680 5206 3694
rect 5244 3680 5291 3684
rect 5164 3674 5291 3680
rect 5164 3645 5252 3674
rect 5281 3645 5291 3674
rect 5400 3677 5437 3756
rect 5478 3743 5588 3756
rect 5552 3687 5583 3688
rect 5400 3657 5409 3677
rect 5429 3657 5437 3677
rect 5400 3647 5437 3657
rect 5496 3677 5583 3687
rect 5496 3657 5505 3677
rect 5525 3657 5583 3677
rect 5496 3648 5583 3657
rect 5496 3647 5533 3648
rect 5164 3641 5291 3645
rect 5164 3624 5203 3641
rect 5244 3640 5291 3641
rect 4786 3604 4823 3608
rect 5164 3606 5175 3624
rect 5193 3606 5203 3624
rect 5164 3597 5203 3606
rect 5165 3596 5202 3597
rect 5552 3595 5583 3648
rect 5613 3677 5650 3756
rect 5821 3753 6214 3773
rect 6234 3753 6237 3773
rect 6472 3767 6510 3775
rect 6576 3799 6661 3805
rect 6686 3804 6723 3805
rect 6576 3779 6584 3799
rect 6604 3779 6661 3799
rect 6576 3771 6661 3779
rect 6685 3795 6723 3804
rect 6685 3775 6694 3795
rect 6714 3775 6723 3795
rect 6576 3770 6612 3771
rect 6685 3767 6723 3775
rect 6789 3799 6874 3805
rect 6894 3804 6931 3805
rect 6789 3779 6797 3799
rect 6817 3798 6874 3799
rect 6817 3779 6846 3798
rect 6789 3778 6846 3779
rect 6867 3778 6874 3798
rect 6789 3771 6874 3778
rect 6893 3795 6931 3804
rect 6893 3775 6902 3795
rect 6922 3775 6931 3795
rect 6789 3770 6825 3771
rect 6893 3767 6931 3775
rect 6997 3799 7141 3805
rect 6997 3779 7005 3799
rect 7025 3797 7113 3799
rect 7025 3779 7054 3797
rect 6997 3776 7054 3779
rect 7081 3779 7113 3797
rect 7133 3779 7141 3799
rect 7081 3776 7141 3779
rect 6997 3771 7141 3776
rect 6997 3770 7033 3771
rect 7105 3770 7141 3771
rect 7207 3804 7244 3805
rect 7207 3803 7245 3804
rect 7207 3795 7271 3803
rect 7207 3775 7216 3795
rect 7236 3781 7271 3795
rect 7291 3781 7294 3801
rect 7236 3776 7294 3781
rect 7236 3775 7271 3776
rect 5821 3748 6237 3753
rect 5821 3747 6162 3748
rect 5765 3687 5796 3688
rect 5613 3657 5622 3677
rect 5642 3657 5650 3677
rect 5613 3647 5650 3657
rect 5709 3680 5796 3687
rect 5709 3677 5770 3680
rect 5709 3657 5718 3677
rect 5738 3660 5770 3677
rect 5791 3660 5796 3680
rect 5738 3657 5796 3660
rect 5709 3650 5796 3657
rect 5821 3677 5858 3747
rect 6124 3746 6161 3747
rect 6473 3738 6510 3767
rect 6474 3736 6510 3738
rect 6686 3736 6723 3767
rect 6474 3714 6723 3736
rect 6894 3735 6931 3767
rect 7207 3763 7271 3775
rect 7311 3737 7338 3915
rect 7706 3908 7735 4086
rect 7775 4048 7839 4060
rect 8115 4056 8152 4088
rect 8323 4087 8572 4109
rect 8323 4056 8360 4087
rect 8536 4085 8572 4087
rect 8536 4056 8573 4085
rect 8885 4076 8922 4077
rect 9188 4076 9225 4146
rect 9250 4166 9337 4173
rect 9250 4163 9308 4166
rect 9250 4143 9255 4163
rect 9276 4146 9308 4163
rect 9328 4146 9337 4166
rect 9276 4143 9337 4146
rect 9250 4136 9337 4143
rect 9396 4166 9433 4176
rect 9396 4146 9404 4166
rect 9424 4146 9433 4166
rect 9250 4135 9281 4136
rect 8884 4075 9225 4076
rect 8809 4070 9225 4075
rect 7775 4047 7810 4048
rect 7752 4042 7810 4047
rect 7752 4022 7755 4042
rect 7775 4028 7810 4042
rect 7830 4028 7839 4048
rect 7775 4020 7839 4028
rect 7801 4019 7839 4020
rect 7802 4018 7839 4019
rect 7905 4052 7941 4053
rect 8013 4052 8049 4053
rect 7905 4044 8049 4052
rect 7905 4024 7913 4044
rect 7933 4024 8021 4044
rect 8041 4024 8049 4044
rect 7905 4018 8049 4024
rect 8115 4048 8153 4056
rect 8221 4052 8257 4053
rect 8115 4028 8124 4048
rect 8144 4028 8153 4048
rect 8115 4019 8153 4028
rect 8172 4045 8257 4052
rect 8172 4025 8179 4045
rect 8200 4044 8257 4045
rect 8200 4025 8229 4044
rect 8172 4024 8229 4025
rect 8249 4024 8257 4044
rect 8115 4018 8152 4019
rect 8172 4018 8257 4024
rect 8323 4048 8361 4056
rect 8434 4052 8470 4053
rect 8323 4028 8332 4048
rect 8352 4028 8361 4048
rect 8323 4019 8361 4028
rect 8385 4044 8470 4052
rect 8385 4024 8442 4044
rect 8462 4024 8470 4044
rect 8323 4018 8360 4019
rect 8385 4018 8470 4024
rect 8536 4048 8574 4056
rect 8809 4050 8812 4070
rect 8832 4050 9225 4070
rect 9396 4067 9433 4146
rect 9463 4175 9494 4228
rect 9844 4226 9881 4227
rect 9843 4217 9882 4226
rect 9843 4199 9853 4217
rect 9871 4199 9882 4217
rect 9755 4182 9802 4183
rect 9843 4182 9882 4199
rect 9755 4178 9882 4182
rect 9513 4175 9550 4176
rect 9463 4166 9550 4175
rect 9463 4146 9521 4166
rect 9541 4146 9550 4166
rect 9463 4136 9550 4146
rect 9609 4166 9646 4176
rect 9609 4146 9617 4166
rect 9637 4146 9646 4166
rect 9463 4135 9494 4136
rect 9458 4067 9568 4080
rect 9609 4067 9646 4146
rect 9755 4149 9765 4178
rect 9794 4149 9882 4178
rect 9755 4143 9882 4149
rect 9755 4139 9802 4143
rect 9840 4129 9882 4143
rect 9840 4111 9851 4129
rect 9869 4111 9882 4129
rect 9840 4106 9882 4111
rect 9841 4103 9882 4106
rect 9841 4102 9878 4103
rect 9396 4065 9646 4067
rect 9396 4062 9497 4065
rect 8536 4028 8545 4048
rect 8565 4028 8574 4048
rect 9396 4043 9461 4062
rect 8536 4019 8574 4028
rect 9458 4035 9461 4043
rect 9490 4035 9497 4062
rect 9525 4038 9535 4065
rect 9564 4043 9646 4065
rect 9564 4038 9568 4043
rect 9525 4035 9568 4038
rect 9458 4021 9568 4035
rect 9834 4039 9881 4040
rect 9834 4030 9882 4039
rect 8536 4018 8573 4019
rect 7959 3997 7995 4018
rect 8385 3997 8416 4018
rect 9834 4012 9853 4030
rect 9871 4012 9882 4030
rect 9834 4010 9882 4012
rect 7792 3993 7892 3997
rect 7792 3989 7854 3993
rect 7792 3963 7799 3989
rect 7825 3967 7854 3989
rect 7880 3967 7892 3993
rect 7825 3963 7892 3967
rect 7792 3960 7892 3963
rect 7960 3960 7995 3997
rect 8057 3994 8416 3997
rect 8057 3989 8279 3994
rect 8057 3965 8070 3989
rect 8094 3970 8279 3989
rect 8303 3970 8416 3994
rect 8094 3965 8416 3970
rect 8057 3961 8416 3965
rect 8483 3989 8632 3997
rect 8483 3969 8494 3989
rect 8514 3969 8632 3989
rect 8483 3962 8632 3969
rect 8483 3961 8524 3962
rect 7959 3921 7995 3960
rect 7807 3908 7844 3909
rect 7903 3908 7940 3909
rect 7959 3908 7966 3921
rect 7706 3899 7845 3908
rect 7706 3879 7816 3899
rect 7836 3879 7845 3899
rect 7706 3872 7845 3879
rect 7903 3899 7966 3908
rect 7903 3879 7912 3899
rect 7932 3883 7966 3899
rect 7989 3908 7995 3921
rect 8014 3908 8051 3909
rect 7989 3899 8051 3908
rect 7989 3883 8022 3899
rect 7932 3879 8022 3883
rect 8042 3879 8051 3899
rect 7706 3870 7803 3872
rect 7706 3869 7735 3870
rect 7903 3869 8051 3879
rect 8110 3899 8147 3909
rect 8222 3908 8259 3909
rect 8203 3906 8259 3908
rect 8110 3879 8118 3899
rect 8138 3879 8147 3899
rect 7959 3868 7995 3869
rect 7807 3809 7844 3810
rect 8110 3809 8147 3879
rect 8172 3899 8259 3906
rect 8172 3896 8230 3899
rect 8172 3876 8177 3896
rect 8198 3879 8230 3896
rect 8250 3879 8259 3899
rect 8198 3876 8259 3879
rect 8172 3869 8259 3876
rect 8318 3899 8355 3909
rect 8318 3879 8326 3899
rect 8346 3879 8355 3899
rect 8172 3868 8203 3869
rect 7806 3808 8147 3809
rect 7731 3804 8147 3808
rect 7731 3803 8108 3804
rect 7731 3783 7734 3803
rect 7754 3787 8108 3803
rect 8128 3787 8147 3804
rect 7754 3783 8147 3787
rect 8318 3800 8355 3879
rect 8385 3908 8416 3961
rect 9196 3953 9234 3955
rect 9843 3953 9882 4010
rect 9196 3920 9882 3953
rect 8435 3908 8472 3909
rect 8385 3899 8472 3908
rect 8385 3879 8443 3899
rect 8463 3879 8472 3899
rect 8385 3869 8472 3879
rect 8531 3899 8568 3909
rect 8531 3879 8539 3899
rect 8559 3879 8568 3899
rect 8385 3868 8416 3869
rect 8380 3800 8490 3813
rect 8531 3800 8568 3879
rect 8318 3798 8568 3800
rect 8318 3795 8419 3798
rect 8318 3776 8383 3795
rect 8380 3768 8383 3776
rect 8412 3768 8419 3795
rect 8447 3771 8457 3798
rect 8486 3776 8568 3798
rect 8788 3832 8956 3833
rect 9196 3832 9234 3920
rect 9495 3918 9542 3920
rect 9842 3896 9882 3920
rect 8788 3809 9234 3832
rect 9460 3863 9571 3878
rect 9460 3861 9502 3863
rect 9460 3841 9467 3861
rect 9486 3841 9502 3861
rect 9460 3833 9502 3841
rect 9530 3861 9571 3863
rect 9530 3841 9544 3861
rect 9563 3841 9571 3861
rect 9843 3852 9882 3896
rect 9530 3833 9571 3841
rect 9460 3827 9571 3833
rect 8788 3806 9232 3809
rect 8788 3804 8956 3806
rect 8486 3771 8490 3776
rect 8447 3768 8490 3771
rect 8380 3754 8490 3768
rect 7170 3735 7338 3737
rect 6891 3728 7338 3735
rect 6555 3708 6666 3714
rect 6555 3700 6596 3708
rect 5973 3687 6009 3688
rect 5821 3657 5830 3677
rect 5850 3657 5858 3677
rect 5709 3648 5765 3650
rect 5709 3647 5746 3648
rect 5821 3647 5858 3657
rect 5917 3677 6065 3687
rect 6165 3684 6261 3686
rect 5917 3657 5926 3677
rect 5946 3657 6036 3677
rect 6056 3657 6065 3677
rect 5917 3648 6065 3657
rect 6123 3677 6261 3684
rect 6123 3657 6132 3677
rect 6152 3657 6261 3677
rect 6555 3680 6563 3700
rect 6582 3680 6596 3700
rect 6555 3678 6596 3680
rect 6624 3700 6666 3708
rect 6624 3680 6640 3700
rect 6659 3680 6666 3700
rect 6891 3701 6916 3728
rect 6947 3709 7338 3728
rect 6947 3701 6996 3709
rect 7170 3708 7338 3709
rect 6891 3699 6996 3701
rect 6624 3678 6666 3680
rect 6555 3663 6666 3678
rect 6123 3648 6261 3657
rect 5917 3647 5954 3648
rect 5973 3596 6009 3648
rect 6028 3647 6065 3648
rect 6124 3647 6161 3648
rect 5444 3594 5485 3595
rect 5336 3587 5485 3594
rect 4459 3585 4496 3586
rect 4409 3576 4496 3585
rect 4409 3556 4467 3576
rect 4487 3556 4496 3576
rect 4409 3546 4496 3556
rect 4555 3576 4592 3586
rect 4555 3556 4563 3576
rect 4583 3556 4592 3576
rect 5336 3567 5454 3587
rect 5474 3567 5485 3587
rect 5336 3559 5485 3567
rect 5552 3591 5911 3595
rect 5552 3586 5874 3591
rect 5552 3562 5665 3586
rect 5689 3567 5874 3586
rect 5898 3567 5911 3591
rect 5689 3562 5911 3567
rect 5552 3559 5911 3562
rect 5973 3559 6008 3596
rect 6076 3593 6176 3596
rect 6076 3589 6143 3593
rect 6076 3563 6088 3589
rect 6114 3567 6143 3589
rect 6169 3567 6176 3593
rect 6114 3563 6176 3567
rect 6076 3559 6176 3563
rect 4409 3545 4440 3546
rect 4404 3477 4514 3490
rect 4555 3477 4592 3556
rect 4789 3541 4826 3542
rect 4785 3532 4826 3541
rect 5552 3538 5583 3559
rect 5973 3538 6009 3559
rect 5395 3537 5432 3538
rect 5169 3534 5203 3535
rect 4785 3514 4798 3532
rect 4816 3514 4826 3532
rect 4785 3505 4826 3514
rect 5168 3525 5205 3534
rect 5168 3507 5177 3525
rect 5195 3507 5205 3525
rect 4785 3485 4825 3505
rect 5168 3497 5205 3507
rect 5394 3528 5432 3537
rect 5394 3508 5403 3528
rect 5423 3508 5432 3528
rect 5394 3500 5432 3508
rect 5498 3532 5583 3538
rect 5608 3537 5645 3538
rect 5498 3512 5506 3532
rect 5526 3512 5583 3532
rect 5498 3504 5583 3512
rect 5607 3528 5645 3537
rect 5607 3508 5616 3528
rect 5636 3508 5645 3528
rect 5498 3503 5534 3504
rect 5607 3500 5645 3508
rect 5711 3532 5796 3538
rect 5816 3537 5853 3538
rect 5711 3512 5719 3532
rect 5739 3531 5796 3532
rect 5739 3512 5768 3531
rect 5711 3511 5768 3512
rect 5789 3511 5796 3531
rect 5711 3504 5796 3511
rect 5815 3528 5853 3537
rect 5815 3508 5824 3528
rect 5844 3508 5853 3528
rect 5711 3503 5747 3504
rect 5815 3500 5853 3508
rect 5919 3532 6063 3538
rect 5919 3512 5927 3532
rect 5947 3531 6035 3532
rect 5947 3512 5978 3531
rect 5919 3511 5978 3512
rect 6003 3512 6035 3531
rect 6055 3512 6063 3532
rect 6003 3511 6063 3512
rect 5919 3504 6063 3511
rect 5919 3503 5955 3504
rect 6027 3503 6063 3504
rect 6129 3537 6166 3538
rect 6129 3536 6167 3537
rect 6129 3528 6193 3536
rect 6129 3508 6138 3528
rect 6158 3514 6193 3528
rect 6213 3514 6216 3534
rect 6158 3509 6216 3514
rect 6158 3508 6193 3509
rect 4342 3475 4592 3477
rect 4342 3472 4443 3475
rect 2860 3415 2924 3427
rect 3200 3423 3237 3450
rect 3408 3423 3445 3454
rect 3621 3452 3657 3454
rect 4342 3453 4407 3472
rect 3621 3423 3658 3452
rect 4404 3445 4407 3453
rect 4436 3445 4443 3472
rect 4471 3448 4481 3475
rect 4510 3453 4592 3475
rect 4700 3475 4825 3485
rect 4700 3456 4708 3475
rect 4733 3456 4825 3475
rect 4510 3448 4514 3453
rect 4700 3449 4825 3456
rect 4471 3445 4514 3448
rect 4404 3431 4514 3445
rect 2860 3414 2895 3415
rect 2837 3409 2895 3414
rect 2837 3389 2840 3409
rect 2860 3395 2895 3409
rect 2915 3395 2924 3415
rect 2860 3387 2924 3395
rect 2886 3386 2924 3387
rect 2887 3385 2924 3386
rect 2990 3419 3026 3420
rect 3098 3419 3134 3420
rect 2990 3411 3134 3419
rect 2990 3391 2998 3411
rect 3018 3408 3106 3411
rect 3018 3391 3050 3408
rect 3070 3391 3106 3408
rect 3126 3391 3134 3411
rect 2990 3385 3134 3391
rect 3200 3415 3238 3423
rect 3306 3419 3342 3420
rect 3200 3395 3209 3415
rect 3229 3395 3238 3415
rect 3200 3386 3238 3395
rect 3257 3412 3342 3419
rect 3257 3392 3264 3412
rect 3285 3411 3342 3412
rect 3285 3392 3314 3411
rect 3257 3391 3314 3392
rect 3334 3391 3342 3411
rect 3200 3385 3237 3386
rect 3257 3385 3342 3391
rect 3408 3415 3446 3423
rect 3519 3419 3555 3420
rect 3408 3395 3417 3415
rect 3437 3395 3446 3415
rect 3408 3386 3446 3395
rect 3470 3411 3555 3419
rect 3470 3391 3527 3411
rect 3547 3391 3555 3411
rect 3408 3385 3445 3386
rect 3470 3385 3555 3391
rect 3621 3415 3659 3423
rect 3621 3395 3630 3415
rect 3650 3395 3659 3415
rect 3621 3386 3659 3395
rect 4785 3401 4825 3449
rect 5169 3469 5203 3497
rect 5395 3471 5432 3500
rect 5396 3469 5432 3471
rect 5608 3469 5645 3500
rect 5169 3468 5341 3469
rect 5169 3436 5355 3468
rect 5396 3447 5645 3469
rect 5816 3468 5853 3500
rect 6129 3496 6193 3508
rect 6233 3470 6260 3648
rect 8788 3626 8815 3804
rect 8855 3766 8919 3778
rect 9195 3774 9232 3806
rect 9403 3805 9652 3827
rect 9403 3774 9440 3805
rect 9616 3803 9652 3805
rect 9616 3774 9653 3803
rect 8855 3765 8890 3766
rect 8832 3760 8890 3765
rect 8832 3740 8835 3760
rect 8855 3746 8890 3760
rect 8910 3746 8919 3766
rect 8855 3738 8919 3746
rect 8881 3737 8919 3738
rect 8882 3736 8919 3737
rect 8985 3770 9021 3771
rect 9093 3770 9129 3771
rect 8985 3765 9129 3770
rect 8985 3762 9047 3765
rect 8985 3742 8993 3762
rect 9013 3745 9047 3762
rect 9070 3762 9129 3765
rect 9070 3745 9101 3762
rect 9013 3742 9101 3745
rect 9121 3742 9129 3762
rect 8985 3736 9129 3742
rect 9195 3766 9233 3774
rect 9301 3770 9337 3771
rect 9195 3746 9204 3766
rect 9224 3746 9233 3766
rect 9195 3737 9233 3746
rect 9252 3763 9337 3770
rect 9252 3743 9259 3763
rect 9280 3762 9337 3763
rect 9280 3743 9309 3762
rect 9252 3742 9309 3743
rect 9329 3742 9337 3762
rect 9195 3736 9232 3737
rect 9252 3736 9337 3742
rect 9403 3766 9441 3774
rect 9514 3770 9550 3771
rect 9403 3746 9412 3766
rect 9432 3746 9441 3766
rect 9403 3737 9441 3746
rect 9465 3762 9550 3770
rect 9465 3742 9522 3762
rect 9542 3742 9550 3762
rect 9403 3736 9440 3737
rect 9465 3736 9550 3742
rect 9616 3766 9654 3774
rect 9616 3746 9625 3766
rect 9645 3746 9654 3766
rect 9616 3737 9654 3746
rect 9616 3736 9653 3737
rect 9039 3715 9075 3736
rect 9465 3715 9496 3736
rect 8872 3711 8972 3715
rect 8872 3707 8934 3711
rect 8872 3681 8879 3707
rect 8905 3685 8934 3707
rect 8960 3685 8972 3711
rect 8905 3681 8972 3685
rect 8872 3678 8972 3681
rect 9040 3678 9075 3715
rect 9137 3712 9496 3715
rect 9137 3707 9359 3712
rect 9137 3683 9150 3707
rect 9174 3688 9359 3707
rect 9383 3688 9496 3712
rect 9174 3683 9496 3688
rect 9137 3679 9496 3683
rect 9563 3707 9712 3715
rect 9563 3687 9574 3707
rect 9594 3687 9712 3707
rect 9563 3680 9712 3687
rect 9563 3679 9604 3680
rect 8887 3626 8924 3627
rect 8983 3626 9020 3627
rect 9039 3626 9075 3678
rect 9094 3626 9131 3627
rect 8787 3617 8925 3626
rect 8787 3597 8896 3617
rect 8916 3597 8925 3617
rect 8787 3590 8925 3597
rect 8983 3617 9131 3626
rect 8983 3597 8992 3617
rect 9012 3597 9102 3617
rect 9122 3597 9131 3617
rect 8787 3588 8883 3590
rect 8983 3587 9131 3597
rect 9190 3617 9227 3627
rect 9302 3626 9339 3627
rect 9283 3624 9339 3626
rect 9190 3597 9198 3617
rect 9218 3597 9227 3617
rect 9039 3586 9075 3587
rect 6416 3544 6526 3558
rect 6416 3541 6459 3544
rect 6416 3536 6420 3541
rect 6092 3468 6260 3470
rect 5816 3462 6260 3468
rect 5169 3404 5203 3436
rect 3621 3385 3658 3386
rect 3044 3364 3080 3385
rect 3470 3364 3501 3385
rect 4785 3383 4796 3401
rect 4814 3383 4825 3401
rect 4785 3375 4825 3383
rect 5165 3395 5203 3404
rect 5165 3377 5175 3395
rect 5193 3377 5203 3395
rect 4786 3374 4823 3375
rect 5165 3371 5203 3377
rect 5321 3373 5355 3436
rect 5477 3441 5588 3447
rect 5477 3433 5518 3441
rect 5477 3413 5485 3433
rect 5504 3413 5518 3433
rect 5477 3411 5518 3413
rect 5546 3433 5588 3441
rect 5546 3413 5562 3433
rect 5581 3413 5588 3433
rect 5546 3411 5588 3413
rect 5477 3396 5588 3411
rect 5815 3442 6260 3462
rect 5815 3373 5853 3442
rect 6092 3441 6260 3442
rect 6338 3514 6420 3536
rect 6449 3514 6459 3541
rect 6487 3517 6494 3544
rect 6523 3536 6526 3544
rect 8521 3553 8632 3568
rect 8521 3551 8563 3553
rect 6523 3517 6588 3536
rect 6487 3514 6588 3517
rect 6338 3512 6588 3514
rect 6338 3433 6375 3512
rect 6416 3499 6526 3512
rect 6490 3443 6521 3444
rect 6338 3413 6347 3433
rect 6367 3413 6375 3433
rect 6338 3403 6375 3413
rect 6434 3433 6521 3443
rect 6434 3413 6443 3433
rect 6463 3413 6521 3433
rect 6434 3404 6521 3413
rect 6434 3403 6471 3404
rect 5165 3367 5202 3371
rect 2877 3360 2977 3364
rect 2877 3356 2939 3360
rect 2877 3330 2884 3356
rect 2910 3334 2939 3356
rect 2965 3334 2977 3360
rect 2910 3330 2977 3334
rect 2877 3327 2977 3330
rect 3045 3327 3080 3364
rect 3142 3361 3501 3364
rect 3142 3356 3364 3361
rect 3142 3332 3155 3356
rect 3179 3337 3364 3356
rect 3388 3337 3501 3361
rect 3179 3332 3501 3337
rect 3142 3328 3501 3332
rect 3568 3356 3717 3364
rect 5321 3362 5853 3373
rect 3568 3336 3579 3356
rect 3599 3336 3717 3356
rect 5320 3346 5853 3362
rect 6490 3351 6521 3404
rect 6551 3433 6588 3512
rect 6759 3522 7152 3529
rect 6759 3505 6767 3522
rect 6799 3509 7152 3522
rect 7172 3509 7175 3529
rect 8254 3524 8295 3533
rect 6799 3505 7175 3509
rect 6759 3504 7175 3505
rect 7849 3522 8017 3523
rect 8254 3522 8263 3524
rect 6759 3503 7100 3504
rect 6703 3443 6734 3444
rect 6551 3413 6560 3433
rect 6580 3413 6588 3433
rect 6551 3403 6588 3413
rect 6647 3436 6734 3443
rect 6647 3433 6708 3436
rect 6647 3413 6656 3433
rect 6676 3416 6708 3433
rect 6729 3416 6734 3436
rect 6676 3413 6734 3416
rect 6647 3406 6734 3413
rect 6759 3433 6796 3503
rect 7062 3502 7099 3503
rect 7849 3502 8263 3522
rect 8289 3502 8295 3524
rect 8521 3531 8528 3551
rect 8547 3531 8563 3551
rect 8521 3523 8563 3531
rect 8591 3551 8632 3553
rect 8591 3531 8605 3551
rect 8624 3531 8632 3551
rect 8591 3523 8632 3531
rect 8887 3527 8924 3528
rect 9190 3527 9227 3597
rect 9252 3617 9339 3624
rect 9252 3614 9310 3617
rect 9252 3594 9257 3614
rect 9278 3597 9310 3614
rect 9330 3597 9339 3617
rect 9278 3594 9339 3597
rect 9252 3587 9339 3594
rect 9398 3617 9435 3627
rect 9398 3597 9406 3617
rect 9426 3597 9435 3617
rect 9252 3586 9283 3587
rect 8886 3526 9227 3527
rect 8521 3517 8632 3523
rect 8811 3521 9227 3526
rect 7849 3496 8295 3502
rect 7849 3494 8017 3496
rect 6911 3443 6947 3444
rect 6759 3413 6768 3433
rect 6788 3413 6796 3433
rect 6647 3404 6703 3406
rect 6647 3403 6684 3404
rect 6759 3403 6796 3413
rect 6855 3433 7003 3443
rect 7103 3440 7199 3442
rect 6855 3413 6864 3433
rect 6884 3428 6974 3433
rect 6884 3413 6919 3428
rect 6855 3404 6919 3413
rect 6855 3403 6892 3404
rect 6911 3387 6919 3404
rect 6940 3413 6974 3428
rect 6994 3413 7003 3433
rect 6940 3404 7003 3413
rect 7061 3433 7199 3440
rect 7061 3413 7070 3433
rect 7090 3413 7199 3433
rect 7061 3404 7199 3413
rect 6940 3387 6947 3404
rect 6966 3403 7003 3404
rect 7062 3403 7099 3404
rect 6911 3352 6947 3387
rect 6382 3350 6423 3351
rect 5320 3345 5834 3346
rect 3568 3329 3717 3336
rect 6274 3343 6423 3350
rect 4157 3333 4671 3334
rect 3568 3328 3609 3329
rect 2892 3275 2929 3276
rect 2988 3275 3025 3276
rect 3044 3275 3080 3327
rect 3099 3275 3136 3276
rect 2792 3266 2930 3275
rect 2792 3246 2901 3266
rect 2921 3246 2930 3266
rect 2792 3239 2930 3246
rect 2988 3266 3136 3275
rect 2988 3246 2997 3266
rect 3017 3246 3107 3266
rect 3127 3246 3136 3266
rect 2792 3237 2888 3239
rect 2988 3236 3136 3246
rect 3195 3266 3232 3276
rect 3307 3275 3344 3276
rect 3288 3273 3344 3275
rect 3195 3246 3203 3266
rect 3223 3246 3232 3266
rect 3044 3235 3080 3236
rect 1974 3183 2142 3185
rect 1696 3177 2142 3183
rect 764 3153 1180 3158
rect 1359 3156 1470 3162
rect 764 3152 1105 3153
rect 708 3092 739 3093
rect 556 3062 565 3082
rect 585 3062 593 3082
rect 556 3052 593 3062
rect 652 3085 739 3092
rect 652 3082 713 3085
rect 652 3062 661 3082
rect 681 3065 713 3082
rect 734 3065 739 3085
rect 681 3062 739 3065
rect 652 3055 739 3062
rect 764 3082 801 3152
rect 1067 3151 1104 3152
rect 1359 3148 1400 3156
rect 1359 3128 1367 3148
rect 1386 3128 1400 3148
rect 1359 3126 1400 3128
rect 1428 3148 1470 3156
rect 1428 3128 1444 3148
rect 1463 3128 1470 3148
rect 1696 3155 1702 3177
rect 1728 3157 2142 3177
rect 2892 3176 2929 3177
rect 3195 3176 3232 3246
rect 3257 3266 3344 3273
rect 3257 3263 3315 3266
rect 3257 3243 3262 3263
rect 3283 3246 3315 3263
rect 3335 3246 3344 3266
rect 3283 3243 3344 3246
rect 3257 3236 3344 3243
rect 3403 3266 3440 3276
rect 3403 3246 3411 3266
rect 3431 3246 3440 3266
rect 3257 3235 3288 3236
rect 2891 3175 3232 3176
rect 1728 3155 1737 3157
rect 1974 3156 2142 3157
rect 2816 3170 3232 3175
rect 1696 3146 1737 3155
rect 2816 3150 2819 3170
rect 2839 3150 3232 3170
rect 3403 3167 3440 3246
rect 3470 3275 3501 3328
rect 4138 3317 4671 3333
rect 6274 3323 6392 3343
rect 6412 3323 6423 3343
rect 4138 3306 4670 3317
rect 6274 3315 6423 3323
rect 6490 3347 6849 3351
rect 6490 3342 6812 3347
rect 6490 3318 6603 3342
rect 6627 3323 6812 3342
rect 6836 3323 6849 3347
rect 6627 3318 6849 3323
rect 6490 3315 6849 3318
rect 6911 3315 6946 3352
rect 7014 3349 7114 3352
rect 7014 3345 7081 3349
rect 7014 3319 7026 3345
rect 7052 3323 7081 3345
rect 7107 3323 7114 3349
rect 7052 3319 7114 3323
rect 7014 3315 7114 3319
rect 4789 3308 4826 3312
rect 3520 3275 3557 3276
rect 3470 3266 3557 3275
rect 3470 3246 3528 3266
rect 3548 3246 3557 3266
rect 3470 3236 3557 3246
rect 3616 3266 3653 3276
rect 3616 3246 3624 3266
rect 3644 3246 3653 3266
rect 3470 3235 3501 3236
rect 3465 3167 3575 3180
rect 3616 3167 3653 3246
rect 3403 3165 3653 3167
rect 3403 3162 3504 3165
rect 3403 3143 3468 3162
rect 1428 3126 1470 3128
rect 1359 3111 1470 3126
rect 3465 3135 3468 3143
rect 3497 3135 3504 3162
rect 3532 3138 3542 3165
rect 3571 3143 3653 3165
rect 3731 3237 3899 3238
rect 4138 3237 4176 3306
rect 3731 3217 4176 3237
rect 4403 3268 4514 3283
rect 4403 3266 4445 3268
rect 4403 3246 4410 3266
rect 4429 3246 4445 3266
rect 4403 3238 4445 3246
rect 4473 3266 4514 3268
rect 4473 3246 4487 3266
rect 4506 3246 4514 3266
rect 4473 3238 4514 3246
rect 4403 3232 4514 3238
rect 4636 3243 4670 3306
rect 4788 3302 4826 3308
rect 5168 3304 5205 3305
rect 4788 3284 4798 3302
rect 4816 3284 4826 3302
rect 4788 3275 4826 3284
rect 5166 3296 5206 3304
rect 5166 3278 5177 3296
rect 5195 3278 5206 3296
rect 6490 3294 6521 3315
rect 6911 3294 6947 3315
rect 6333 3293 6370 3294
rect 4788 3243 4822 3275
rect 3731 3211 4175 3217
rect 3731 3209 3899 3211
rect 3571 3138 3575 3143
rect 3532 3135 3575 3138
rect 3465 3121 3575 3135
rect 2694 3107 2762 3116
rect 916 3092 952 3093
rect 764 3062 773 3082
rect 793 3062 801 3082
rect 652 3053 708 3055
rect 652 3052 689 3053
rect 764 3052 801 3062
rect 860 3082 1008 3092
rect 1108 3089 1204 3091
rect 860 3062 869 3082
rect 889 3062 979 3082
rect 999 3062 1008 3082
rect 860 3053 1008 3062
rect 1066 3082 1204 3089
rect 1066 3062 1075 3082
rect 1095 3062 1204 3082
rect 2694 3078 2709 3107
rect 2757 3087 2762 3107
rect 2757 3078 2764 3087
rect 2694 3067 2764 3078
rect 1066 3053 1204 3062
rect 860 3052 897 3053
rect 916 3001 952 3053
rect 971 3052 1008 3053
rect 1067 3052 1104 3053
rect 387 2999 428 3000
rect 279 2992 428 2999
rect 279 2972 397 2992
rect 417 2972 428 2992
rect 279 2964 428 2972
rect 495 2996 854 3000
rect 495 2991 817 2996
rect 495 2967 608 2991
rect 632 2972 817 2991
rect 841 2972 854 2996
rect 632 2967 854 2972
rect 495 2964 854 2967
rect 916 2964 951 3001
rect 1019 2998 1119 3001
rect 1019 2994 1086 2998
rect 1019 2968 1031 2994
rect 1057 2972 1086 2994
rect 1112 2972 1119 2998
rect 1057 2968 1119 2972
rect 1019 2964 1119 2968
rect 495 2943 526 2964
rect 916 2943 952 2964
rect 338 2942 375 2943
rect 337 2933 375 2942
rect 337 2913 346 2933
rect 366 2913 375 2933
rect 337 2905 375 2913
rect 441 2937 526 2943
rect 551 2942 588 2943
rect 441 2917 449 2937
rect 469 2917 526 2937
rect 441 2909 526 2917
rect 550 2933 588 2942
rect 550 2913 559 2933
rect 579 2913 588 2933
rect 441 2908 477 2909
rect 550 2905 588 2913
rect 654 2937 739 2943
rect 759 2942 796 2943
rect 654 2917 662 2937
rect 682 2936 739 2937
rect 682 2917 711 2936
rect 654 2916 711 2917
rect 732 2916 739 2936
rect 654 2909 739 2916
rect 758 2933 796 2942
rect 758 2913 767 2933
rect 787 2913 796 2933
rect 654 2908 690 2909
rect 758 2905 796 2913
rect 862 2937 1006 2943
rect 862 2917 870 2937
rect 890 2934 978 2937
rect 890 2917 921 2934
rect 862 2914 921 2917
rect 944 2917 978 2934
rect 998 2917 1006 2937
rect 944 2914 1006 2917
rect 862 2909 1006 2914
rect 862 2908 898 2909
rect 970 2908 1006 2909
rect 1072 2942 1109 2943
rect 1072 2941 1110 2942
rect 1072 2933 1136 2941
rect 1072 2913 1081 2933
rect 1101 2919 1136 2933
rect 1156 2919 1159 2939
rect 1101 2914 1159 2919
rect 1101 2913 1136 2914
rect 338 2876 375 2905
rect 339 2874 375 2876
rect 551 2874 588 2905
rect 339 2852 588 2874
rect 759 2873 796 2905
rect 1072 2901 1136 2913
rect 1176 2875 1203 3053
rect 2703 2960 2764 3067
rect 3731 3031 3758 3209
rect 3798 3171 3862 3183
rect 4138 3179 4175 3211
rect 4346 3210 4595 3232
rect 4636 3211 4822 3243
rect 4650 3210 4822 3211
rect 4346 3179 4383 3210
rect 4559 3208 4595 3210
rect 4559 3179 4596 3208
rect 4788 3182 4822 3210
rect 5166 3230 5206 3278
rect 6332 3284 6370 3293
rect 6332 3264 6341 3284
rect 6361 3264 6370 3284
rect 6332 3256 6370 3264
rect 6436 3288 6521 3294
rect 6546 3293 6583 3294
rect 6436 3268 6444 3288
rect 6464 3268 6521 3288
rect 6436 3260 6521 3268
rect 6545 3284 6583 3293
rect 6545 3264 6554 3284
rect 6574 3264 6583 3284
rect 6436 3259 6472 3260
rect 6545 3256 6583 3264
rect 6649 3288 6734 3294
rect 6754 3293 6791 3294
rect 6649 3268 6657 3288
rect 6677 3287 6734 3288
rect 6677 3268 6706 3287
rect 6649 3267 6706 3268
rect 6727 3267 6734 3287
rect 6649 3260 6734 3267
rect 6753 3284 6791 3293
rect 6753 3264 6762 3284
rect 6782 3264 6791 3284
rect 6649 3259 6685 3260
rect 6753 3256 6791 3264
rect 6857 3288 7001 3294
rect 6857 3268 6865 3288
rect 6885 3268 6973 3288
rect 6993 3268 7001 3288
rect 6857 3260 7001 3268
rect 6857 3259 6893 3260
rect 6965 3259 7001 3260
rect 7067 3293 7104 3294
rect 7067 3292 7105 3293
rect 7067 3284 7131 3292
rect 7067 3264 7076 3284
rect 7096 3270 7131 3284
rect 7151 3270 7154 3290
rect 7096 3265 7154 3270
rect 7096 3264 7131 3265
rect 5477 3234 5587 3248
rect 5477 3231 5520 3234
rect 5166 3223 5291 3230
rect 5477 3226 5481 3231
rect 5166 3204 5258 3223
rect 5283 3204 5291 3223
rect 5166 3194 5291 3204
rect 5399 3204 5481 3226
rect 5510 3204 5520 3231
rect 5548 3207 5555 3234
rect 5584 3226 5587 3234
rect 6333 3227 6370 3256
rect 5584 3207 5649 3226
rect 6334 3225 6370 3227
rect 6546 3225 6583 3256
rect 6754 3229 6791 3256
rect 7067 3252 7131 3264
rect 5548 3204 5649 3207
rect 5399 3202 5649 3204
rect 3798 3170 3833 3171
rect 3775 3165 3833 3170
rect 3775 3145 3778 3165
rect 3798 3151 3833 3165
rect 3853 3151 3862 3171
rect 3798 3143 3862 3151
rect 3824 3142 3862 3143
rect 3825 3141 3862 3142
rect 3928 3175 3964 3176
rect 4036 3175 4072 3176
rect 3928 3168 4072 3175
rect 3928 3167 3988 3168
rect 3928 3147 3936 3167
rect 3956 3148 3988 3167
rect 4013 3167 4072 3168
rect 4013 3148 4044 3167
rect 3956 3147 4044 3148
rect 4064 3147 4072 3167
rect 3928 3141 4072 3147
rect 4138 3171 4176 3179
rect 4244 3175 4280 3176
rect 4138 3151 4147 3171
rect 4167 3151 4176 3171
rect 4138 3142 4176 3151
rect 4195 3168 4280 3175
rect 4195 3148 4202 3168
rect 4223 3167 4280 3168
rect 4223 3148 4252 3167
rect 4195 3147 4252 3148
rect 4272 3147 4280 3167
rect 4138 3141 4175 3142
rect 4195 3141 4280 3147
rect 4346 3171 4384 3179
rect 4457 3175 4493 3176
rect 4346 3151 4355 3171
rect 4375 3151 4384 3171
rect 4346 3142 4384 3151
rect 4408 3167 4493 3175
rect 4408 3147 4465 3167
rect 4485 3147 4493 3167
rect 4346 3141 4383 3142
rect 4408 3141 4493 3147
rect 4559 3171 4597 3179
rect 4559 3151 4568 3171
rect 4588 3151 4597 3171
rect 4559 3142 4597 3151
rect 4786 3172 4823 3182
rect 5166 3174 5206 3194
rect 4786 3154 4796 3172
rect 4814 3154 4823 3172
rect 4786 3145 4823 3154
rect 5165 3165 5206 3174
rect 5165 3147 5175 3165
rect 5193 3147 5206 3165
rect 4788 3144 4822 3145
rect 4559 3141 4596 3142
rect 3982 3120 4018 3141
rect 4408 3120 4439 3141
rect 5165 3138 5206 3147
rect 5165 3137 5202 3138
rect 5399 3123 5436 3202
rect 5477 3189 5587 3202
rect 5551 3133 5582 3134
rect 3815 3116 3915 3120
rect 3815 3112 3877 3116
rect 3815 3086 3822 3112
rect 3848 3090 3877 3112
rect 3903 3090 3915 3116
rect 3848 3086 3915 3090
rect 3815 3083 3915 3086
rect 3983 3083 4018 3120
rect 4080 3117 4439 3120
rect 4080 3112 4302 3117
rect 4080 3088 4093 3112
rect 4117 3093 4302 3112
rect 4326 3093 4439 3117
rect 4117 3088 4439 3093
rect 4080 3084 4439 3088
rect 4506 3112 4655 3120
rect 4506 3092 4517 3112
rect 4537 3092 4655 3112
rect 5399 3103 5408 3123
rect 5428 3103 5436 3123
rect 5399 3093 5436 3103
rect 5495 3123 5582 3133
rect 5495 3103 5504 3123
rect 5524 3103 5582 3123
rect 5495 3094 5582 3103
rect 5495 3093 5532 3094
rect 4506 3085 4655 3092
rect 4506 3084 4547 3085
rect 3830 3031 3867 3032
rect 3926 3031 3963 3032
rect 3982 3031 4018 3083
rect 4037 3031 4074 3032
rect 3730 3022 3868 3031
rect 2694 2959 2764 2960
rect 3355 2988 3466 3003
rect 3730 3002 3839 3022
rect 3859 3002 3868 3022
rect 3730 2995 3868 3002
rect 3926 3022 4074 3031
rect 3926 3002 3935 3022
rect 3955 3002 4045 3022
rect 4065 3002 4074 3022
rect 3730 2993 3826 2995
rect 3926 2992 4074 3002
rect 4133 3022 4170 3032
rect 4245 3031 4282 3032
rect 4226 3029 4282 3031
rect 4133 3002 4141 3022
rect 4161 3002 4170 3022
rect 3982 2991 4018 2992
rect 3355 2986 3397 2988
rect 3355 2966 3362 2986
rect 3381 2966 3397 2986
rect 2694 2958 2802 2959
rect 3355 2958 3397 2966
rect 3425 2986 3466 2988
rect 3425 2966 3439 2986
rect 3458 2966 3466 2986
rect 3425 2958 3466 2966
rect 2683 2957 2851 2958
rect 1470 2924 1580 2938
rect 1470 2921 1513 2924
rect 1470 2916 1474 2921
rect 1035 2873 1203 2875
rect 759 2870 1203 2873
rect 420 2846 531 2852
rect 420 2838 461 2846
rect 109 2783 148 2827
rect 420 2818 428 2838
rect 447 2818 461 2838
rect 420 2816 461 2818
rect 489 2838 531 2846
rect 489 2818 505 2838
rect 524 2818 531 2838
rect 489 2816 531 2818
rect 420 2802 531 2816
rect 757 2847 1203 2870
rect 109 2759 149 2783
rect 449 2759 496 2761
rect 757 2759 795 2847
rect 1035 2846 1203 2847
rect 1392 2894 1474 2916
rect 1503 2894 1513 2921
rect 1541 2897 1548 2924
rect 1577 2916 1580 2924
rect 2683 2931 3127 2957
rect 3355 2952 3466 2958
rect 2683 2929 2851 2931
rect 2683 2927 2802 2929
rect 1577 2897 1642 2916
rect 1541 2894 1642 2897
rect 1392 2892 1642 2894
rect 1392 2813 1429 2892
rect 1470 2879 1580 2892
rect 1544 2823 1575 2824
rect 1392 2793 1401 2813
rect 1421 2793 1429 2813
rect 1392 2783 1429 2793
rect 1488 2813 1575 2823
rect 1488 2793 1497 2813
rect 1517 2793 1575 2813
rect 1488 2784 1575 2793
rect 1488 2783 1525 2784
rect 109 2726 795 2759
rect 1544 2731 1575 2784
rect 1605 2813 1642 2892
rect 1813 2911 1845 2923
rect 1813 2891 1815 2911
rect 1836 2909 1845 2911
rect 1836 2907 2188 2909
rect 1836 2891 2206 2907
rect 1813 2889 2206 2891
rect 2226 2889 2229 2907
rect 1813 2884 2229 2889
rect 1813 2883 2154 2884
rect 1757 2823 1788 2824
rect 1605 2793 1614 2813
rect 1634 2793 1642 2813
rect 1605 2783 1642 2793
rect 1701 2816 1788 2823
rect 1701 2813 1762 2816
rect 1701 2793 1710 2813
rect 1730 2796 1762 2813
rect 1783 2796 1788 2816
rect 1730 2793 1788 2796
rect 1701 2786 1788 2793
rect 1813 2813 1850 2883
rect 2116 2882 2153 2883
rect 1965 2823 2001 2824
rect 1813 2793 1822 2813
rect 1842 2793 1850 2813
rect 1701 2784 1757 2786
rect 1701 2783 1738 2784
rect 1813 2783 1850 2793
rect 1909 2813 2057 2823
rect 2157 2820 2253 2822
rect 1909 2793 1918 2813
rect 1938 2804 2028 2813
rect 1938 2793 1969 2804
rect 1909 2784 1969 2793
rect 1909 2783 1946 2784
rect 1965 2772 1969 2784
rect 1996 2793 2028 2804
rect 2048 2793 2057 2813
rect 1996 2784 2057 2793
rect 2115 2813 2253 2820
rect 2115 2793 2124 2813
rect 2144 2793 2253 2813
rect 2115 2784 2253 2793
rect 1996 2772 2001 2784
rect 2020 2783 2057 2784
rect 2116 2783 2153 2784
rect 1965 2732 2001 2772
rect 1436 2730 1477 2731
rect 108 2669 147 2726
rect 757 2724 795 2726
rect 1328 2723 1477 2730
rect 1328 2703 1446 2723
rect 1466 2703 1477 2723
rect 1328 2695 1477 2703
rect 1544 2727 1903 2731
rect 1544 2722 1866 2727
rect 1544 2698 1657 2722
rect 1681 2703 1866 2722
rect 1890 2703 1903 2727
rect 1681 2698 1903 2703
rect 1544 2695 1903 2698
rect 1965 2695 2000 2732
rect 2068 2729 2168 2732
rect 2068 2725 2135 2729
rect 2068 2699 2080 2725
rect 2106 2703 2135 2725
rect 2161 2703 2168 2729
rect 2106 2699 2168 2703
rect 2068 2695 2168 2699
rect 1544 2674 1575 2695
rect 1965 2674 2001 2695
rect 1387 2673 1424 2674
rect 108 2667 156 2669
rect 108 2649 119 2667
rect 137 2649 156 2667
rect 1386 2664 1424 2673
rect 108 2640 156 2649
rect 109 2639 156 2640
rect 422 2644 532 2658
rect 422 2641 465 2644
rect 422 2636 426 2641
rect 344 2614 426 2636
rect 455 2614 465 2641
rect 493 2617 500 2644
rect 529 2636 532 2644
rect 1386 2644 1395 2664
rect 1415 2644 1424 2664
rect 1386 2636 1424 2644
rect 1490 2668 1575 2674
rect 1600 2673 1637 2674
rect 1490 2648 1498 2668
rect 1518 2648 1575 2668
rect 1490 2640 1575 2648
rect 1599 2664 1637 2673
rect 1599 2644 1608 2664
rect 1628 2644 1637 2664
rect 1490 2639 1526 2640
rect 1599 2636 1637 2644
rect 1703 2668 1788 2674
rect 1808 2673 1845 2674
rect 1703 2648 1711 2668
rect 1731 2667 1788 2668
rect 1731 2648 1760 2667
rect 1703 2647 1760 2648
rect 1781 2647 1788 2667
rect 1703 2640 1788 2647
rect 1807 2664 1845 2673
rect 1807 2644 1816 2664
rect 1836 2644 1845 2664
rect 1703 2639 1739 2640
rect 1807 2636 1845 2644
rect 1911 2668 2055 2674
rect 1911 2648 1919 2668
rect 1939 2648 2027 2668
rect 2047 2648 2055 2668
rect 1911 2640 2055 2648
rect 1911 2639 1947 2640
rect 2019 2639 2055 2640
rect 2121 2673 2158 2674
rect 2121 2672 2159 2673
rect 2121 2664 2185 2672
rect 2121 2644 2130 2664
rect 2150 2650 2185 2664
rect 2205 2650 2208 2670
rect 2150 2645 2208 2650
rect 2150 2644 2185 2645
rect 529 2617 594 2636
rect 493 2614 594 2617
rect 344 2612 594 2614
rect 112 2576 149 2577
rect 108 2573 149 2576
rect 108 2568 150 2573
rect 108 2550 121 2568
rect 139 2550 150 2568
rect 108 2536 150 2550
rect 188 2536 235 2540
rect 108 2530 235 2536
rect 108 2501 196 2530
rect 225 2501 235 2530
rect 344 2533 381 2612
rect 422 2599 532 2612
rect 496 2543 527 2544
rect 344 2513 353 2533
rect 373 2513 381 2533
rect 344 2503 381 2513
rect 440 2533 527 2543
rect 440 2513 449 2533
rect 469 2513 527 2533
rect 440 2504 527 2513
rect 440 2503 477 2504
rect 108 2497 235 2501
rect 108 2480 147 2497
rect 188 2496 235 2497
rect 108 2462 119 2480
rect 137 2462 147 2480
rect 108 2453 147 2462
rect 109 2452 146 2453
rect 496 2451 527 2504
rect 557 2533 594 2612
rect 765 2609 1158 2629
rect 1178 2609 1181 2629
rect 765 2604 1181 2609
rect 1387 2607 1424 2636
rect 1388 2605 1424 2607
rect 1600 2605 1637 2636
rect 765 2603 1106 2604
rect 709 2543 740 2544
rect 557 2513 566 2533
rect 586 2513 594 2533
rect 557 2503 594 2513
rect 653 2536 740 2543
rect 653 2533 714 2536
rect 653 2513 662 2533
rect 682 2516 714 2533
rect 735 2516 740 2536
rect 682 2513 740 2516
rect 653 2506 740 2513
rect 765 2533 802 2603
rect 1068 2602 1105 2603
rect 1388 2583 1637 2605
rect 1808 2604 1845 2636
rect 2121 2632 2185 2644
rect 2225 2614 2252 2784
rect 2683 2751 2710 2927
rect 2750 2891 2814 2903
rect 3090 2899 3127 2931
rect 3298 2930 3547 2952
rect 3830 2932 3867 2933
rect 4133 2932 4170 3002
rect 4195 3022 4282 3029
rect 4195 3019 4253 3022
rect 4195 2999 4200 3019
rect 4221 3002 4253 3019
rect 4273 3002 4282 3022
rect 4221 2999 4282 3002
rect 4195 2992 4282 2999
rect 4341 3022 4378 3032
rect 4341 3002 4349 3022
rect 4369 3002 4378 3022
rect 4195 2991 4226 2992
rect 3829 2931 4170 2932
rect 3298 2899 3335 2930
rect 3511 2928 3547 2930
rect 3511 2899 3548 2928
rect 3754 2926 4170 2931
rect 3754 2906 3757 2926
rect 3777 2906 4170 2926
rect 4341 2923 4378 3002
rect 4408 3031 4439 3084
rect 4789 3082 4826 3083
rect 4788 3073 4827 3082
rect 4788 3055 4798 3073
rect 4816 3055 4827 3073
rect 5168 3071 5205 3075
rect 4700 3038 4747 3039
rect 4788 3038 4827 3055
rect 4700 3034 4827 3038
rect 4458 3031 4495 3032
rect 4408 3022 4495 3031
rect 4408 3002 4466 3022
rect 4486 3002 4495 3022
rect 4408 2992 4495 3002
rect 4554 3022 4591 3032
rect 4554 3002 4562 3022
rect 4582 3002 4591 3022
rect 4408 2991 4439 2992
rect 4403 2923 4513 2936
rect 4554 2923 4591 3002
rect 4700 3005 4710 3034
rect 4739 3005 4827 3034
rect 4700 2999 4827 3005
rect 4700 2995 4747 2999
rect 4785 2985 4827 2999
rect 4785 2967 4796 2985
rect 4814 2967 4827 2985
rect 4785 2962 4827 2967
rect 4786 2959 4827 2962
rect 5165 3066 5205 3071
rect 5165 3048 5177 3066
rect 5195 3048 5205 3066
rect 4786 2958 4823 2959
rect 4341 2921 4591 2923
rect 4341 2918 4442 2921
rect 4341 2899 4406 2918
rect 2750 2890 2785 2891
rect 2727 2885 2785 2890
rect 2727 2865 2730 2885
rect 2750 2871 2785 2885
rect 2805 2871 2814 2891
rect 2750 2863 2814 2871
rect 2776 2862 2814 2863
rect 2777 2861 2814 2862
rect 2880 2895 2916 2896
rect 2988 2895 3024 2896
rect 2880 2888 3024 2895
rect 2880 2887 2938 2888
rect 2880 2867 2888 2887
rect 2908 2869 2938 2887
rect 2967 2887 3024 2888
rect 2967 2869 2996 2887
rect 2908 2867 2996 2869
rect 3016 2867 3024 2887
rect 2880 2861 3024 2867
rect 3090 2891 3128 2899
rect 3196 2895 3232 2896
rect 3090 2871 3099 2891
rect 3119 2871 3128 2891
rect 3090 2862 3128 2871
rect 3147 2888 3232 2895
rect 3147 2868 3154 2888
rect 3175 2887 3232 2888
rect 3175 2868 3204 2887
rect 3147 2867 3204 2868
rect 3224 2867 3232 2887
rect 3090 2861 3127 2862
rect 3147 2861 3232 2867
rect 3298 2891 3336 2899
rect 3409 2895 3445 2896
rect 3298 2871 3307 2891
rect 3327 2871 3336 2891
rect 3298 2862 3336 2871
rect 3360 2887 3445 2895
rect 3360 2867 3417 2887
rect 3437 2867 3445 2887
rect 3298 2861 3335 2862
rect 3360 2861 3445 2867
rect 3511 2891 3549 2899
rect 3511 2871 3520 2891
rect 3540 2871 3549 2891
rect 4403 2891 4406 2899
rect 4435 2891 4442 2918
rect 4470 2894 4480 2921
rect 4509 2899 4591 2921
rect 4509 2894 4513 2899
rect 4470 2891 4513 2894
rect 4403 2877 4513 2891
rect 4779 2895 4826 2896
rect 4779 2886 4827 2895
rect 3511 2862 3549 2871
rect 4779 2868 4798 2886
rect 4816 2868 4827 2886
rect 4779 2866 4827 2868
rect 3511 2861 3548 2862
rect 2934 2840 2970 2861
rect 3360 2840 3391 2861
rect 2767 2836 2867 2840
rect 2767 2832 2829 2836
rect 2767 2806 2774 2832
rect 2800 2810 2829 2832
rect 2855 2810 2867 2836
rect 2800 2806 2867 2810
rect 2767 2803 2867 2806
rect 2935 2803 2970 2840
rect 3032 2837 3391 2840
rect 3032 2832 3254 2837
rect 3032 2808 3045 2832
rect 3069 2813 3254 2832
rect 3278 2813 3391 2837
rect 3069 2808 3391 2813
rect 3032 2804 3391 2808
rect 3458 2832 3607 2840
rect 3458 2812 3469 2832
rect 3489 2812 3607 2832
rect 3458 2805 3607 2812
rect 4140 2809 4178 2811
rect 4788 2809 4827 2866
rect 5165 2868 5205 3048
rect 5551 3041 5582 3094
rect 5612 3123 5649 3202
rect 5820 3199 6213 3219
rect 6233 3199 6236 3219
rect 6334 3203 6583 3225
rect 6752 3224 6793 3229
rect 7171 3226 7198 3404
rect 7849 3316 7876 3494
rect 8254 3491 8295 3496
rect 8464 3495 8713 3517
rect 8811 3501 8814 3521
rect 8834 3501 9227 3521
rect 9398 3518 9435 3597
rect 9465 3626 9496 3679
rect 9842 3672 9882 3852
rect 9842 3654 9852 3672
rect 9870 3654 9882 3672
rect 9842 3649 9882 3654
rect 9842 3645 9879 3649
rect 9515 3626 9552 3627
rect 9465 3617 9552 3626
rect 9465 3597 9523 3617
rect 9543 3597 9552 3617
rect 9465 3587 9552 3597
rect 9611 3617 9648 3627
rect 9611 3597 9619 3617
rect 9639 3597 9648 3617
rect 9465 3586 9496 3587
rect 9460 3518 9570 3531
rect 9611 3518 9648 3597
rect 9845 3582 9882 3583
rect 9841 3573 9882 3582
rect 9841 3555 9854 3573
rect 9872 3555 9882 3573
rect 9841 3546 9882 3555
rect 9841 3526 9881 3546
rect 9398 3516 9648 3518
rect 9398 3513 9499 3516
rect 7916 3456 7980 3468
rect 8256 3464 8293 3491
rect 8464 3464 8501 3495
rect 8677 3493 8713 3495
rect 9398 3494 9463 3513
rect 8677 3464 8714 3493
rect 9460 3486 9463 3494
rect 9492 3486 9499 3513
rect 9527 3489 9537 3516
rect 9566 3494 9648 3516
rect 9756 3516 9881 3526
rect 9756 3497 9764 3516
rect 9789 3497 9881 3516
rect 9566 3489 9570 3494
rect 9756 3490 9881 3497
rect 9527 3486 9570 3489
rect 9460 3472 9570 3486
rect 7916 3455 7951 3456
rect 7893 3450 7951 3455
rect 7893 3430 7896 3450
rect 7916 3436 7951 3450
rect 7971 3436 7980 3456
rect 7916 3428 7980 3436
rect 7942 3427 7980 3428
rect 7943 3426 7980 3427
rect 8046 3460 8082 3461
rect 8154 3460 8190 3461
rect 8046 3452 8190 3460
rect 8046 3432 8054 3452
rect 8074 3449 8162 3452
rect 8074 3432 8106 3449
rect 8126 3432 8162 3449
rect 8182 3432 8190 3452
rect 8046 3426 8190 3432
rect 8256 3456 8294 3464
rect 8362 3460 8398 3461
rect 8256 3436 8265 3456
rect 8285 3436 8294 3456
rect 8256 3427 8294 3436
rect 8313 3453 8398 3460
rect 8313 3433 8320 3453
rect 8341 3452 8398 3453
rect 8341 3433 8370 3452
rect 8313 3432 8370 3433
rect 8390 3432 8398 3452
rect 8256 3426 8293 3427
rect 8313 3426 8398 3432
rect 8464 3456 8502 3464
rect 8575 3460 8611 3461
rect 8464 3436 8473 3456
rect 8493 3436 8502 3456
rect 8464 3427 8502 3436
rect 8526 3452 8611 3460
rect 8526 3432 8583 3452
rect 8603 3432 8611 3452
rect 8464 3426 8501 3427
rect 8526 3426 8611 3432
rect 8677 3456 8715 3464
rect 8677 3436 8686 3456
rect 8706 3436 8715 3456
rect 8677 3427 8715 3436
rect 9841 3442 9881 3490
rect 8677 3426 8714 3427
rect 8100 3405 8136 3426
rect 8526 3405 8557 3426
rect 9841 3424 9852 3442
rect 9870 3424 9881 3442
rect 9841 3416 9881 3424
rect 9842 3415 9879 3416
rect 7933 3401 8033 3405
rect 7933 3397 7995 3401
rect 7933 3371 7940 3397
rect 7966 3375 7995 3397
rect 8021 3375 8033 3401
rect 7966 3371 8033 3375
rect 7933 3368 8033 3371
rect 8101 3368 8136 3405
rect 8198 3402 8557 3405
rect 8198 3397 8420 3402
rect 8198 3373 8211 3397
rect 8235 3378 8420 3397
rect 8444 3378 8557 3402
rect 8235 3373 8557 3378
rect 8198 3369 8557 3373
rect 8624 3397 8773 3405
rect 8624 3377 8635 3397
rect 8655 3377 8773 3397
rect 8624 3370 8773 3377
rect 9213 3374 9727 3375
rect 8624 3369 8665 3370
rect 7948 3316 7985 3317
rect 8044 3316 8081 3317
rect 8100 3316 8136 3368
rect 8155 3316 8192 3317
rect 7848 3307 7986 3316
rect 7848 3287 7957 3307
rect 7977 3287 7986 3307
rect 7848 3280 7986 3287
rect 8044 3307 8192 3316
rect 8044 3287 8053 3307
rect 8073 3287 8163 3307
rect 8183 3287 8192 3307
rect 7848 3278 7944 3280
rect 8044 3277 8192 3287
rect 8251 3307 8288 3317
rect 8363 3316 8400 3317
rect 8344 3314 8400 3316
rect 8251 3287 8259 3307
rect 8279 3287 8288 3307
rect 8100 3276 8136 3277
rect 7030 3224 7198 3226
rect 6752 3218 7198 3224
rect 5820 3194 6236 3199
rect 6415 3197 6526 3203
rect 5820 3193 6161 3194
rect 5764 3133 5795 3134
rect 5612 3103 5621 3123
rect 5641 3103 5649 3123
rect 5612 3093 5649 3103
rect 5708 3126 5795 3133
rect 5708 3123 5769 3126
rect 5708 3103 5717 3123
rect 5737 3106 5769 3123
rect 5790 3106 5795 3126
rect 5737 3103 5795 3106
rect 5708 3096 5795 3103
rect 5820 3123 5857 3193
rect 6123 3192 6160 3193
rect 6415 3189 6456 3197
rect 6415 3169 6423 3189
rect 6442 3169 6456 3189
rect 6415 3167 6456 3169
rect 6484 3189 6526 3197
rect 6484 3169 6500 3189
rect 6519 3169 6526 3189
rect 6752 3196 6758 3218
rect 6784 3198 7198 3218
rect 7948 3217 7985 3218
rect 8251 3217 8288 3287
rect 8313 3307 8400 3314
rect 8313 3304 8371 3307
rect 8313 3284 8318 3304
rect 8339 3287 8371 3304
rect 8391 3287 8400 3307
rect 8339 3284 8400 3287
rect 8313 3277 8400 3284
rect 8459 3307 8496 3317
rect 8459 3287 8467 3307
rect 8487 3287 8496 3307
rect 8313 3276 8344 3277
rect 7947 3216 8288 3217
rect 6784 3196 6793 3198
rect 7030 3197 7198 3198
rect 7872 3211 8288 3216
rect 6752 3187 6793 3196
rect 7872 3191 7875 3211
rect 7895 3191 8288 3211
rect 8459 3208 8496 3287
rect 8526 3316 8557 3369
rect 9194 3358 9727 3374
rect 9194 3347 9726 3358
rect 9845 3349 9882 3353
rect 8576 3316 8613 3317
rect 8526 3307 8613 3316
rect 8526 3287 8584 3307
rect 8604 3287 8613 3307
rect 8526 3277 8613 3287
rect 8672 3307 8709 3317
rect 8672 3287 8680 3307
rect 8700 3287 8709 3307
rect 8526 3276 8557 3277
rect 8521 3208 8631 3221
rect 8672 3208 8709 3287
rect 8459 3206 8709 3208
rect 8459 3203 8560 3206
rect 8459 3184 8524 3203
rect 6484 3167 6526 3169
rect 6415 3152 6526 3167
rect 8521 3176 8524 3184
rect 8553 3176 8560 3203
rect 8588 3179 8598 3206
rect 8627 3184 8709 3206
rect 8787 3278 8955 3279
rect 9194 3278 9232 3347
rect 8787 3258 9232 3278
rect 9459 3309 9570 3324
rect 9459 3307 9501 3309
rect 9459 3287 9466 3307
rect 9485 3287 9501 3307
rect 9459 3279 9501 3287
rect 9529 3307 9570 3309
rect 9529 3287 9543 3307
rect 9562 3287 9570 3307
rect 9529 3279 9570 3287
rect 9459 3273 9570 3279
rect 9692 3284 9726 3347
rect 9844 3343 9882 3349
rect 9844 3325 9854 3343
rect 9872 3325 9882 3343
rect 9844 3316 9882 3325
rect 9844 3284 9878 3316
rect 8787 3252 9231 3258
rect 8787 3250 8955 3252
rect 8627 3179 8631 3184
rect 8588 3176 8631 3179
rect 8521 3162 8631 3176
rect 7750 3148 7818 3157
rect 5972 3133 6008 3134
rect 5820 3103 5829 3123
rect 5849 3103 5857 3123
rect 5708 3094 5764 3096
rect 5708 3093 5745 3094
rect 5820 3093 5857 3103
rect 5916 3123 6064 3133
rect 6164 3130 6260 3132
rect 5916 3103 5925 3123
rect 5945 3103 6035 3123
rect 6055 3103 6064 3123
rect 5916 3094 6064 3103
rect 6122 3123 6260 3130
rect 6122 3103 6131 3123
rect 6151 3103 6260 3123
rect 7750 3119 7765 3148
rect 7813 3128 7818 3148
rect 7813 3119 7820 3128
rect 7750 3108 7820 3119
rect 6122 3094 6260 3103
rect 5916 3093 5953 3094
rect 5972 3042 6008 3094
rect 6027 3093 6064 3094
rect 6123 3093 6160 3094
rect 5443 3040 5484 3041
rect 5335 3033 5484 3040
rect 5335 3013 5453 3033
rect 5473 3013 5484 3033
rect 5335 3005 5484 3013
rect 5551 3037 5910 3041
rect 5551 3032 5873 3037
rect 5551 3008 5664 3032
rect 5688 3013 5873 3032
rect 5897 3013 5910 3037
rect 5688 3008 5910 3013
rect 5551 3005 5910 3008
rect 5972 3005 6007 3042
rect 6075 3039 6175 3042
rect 6075 3035 6142 3039
rect 6075 3009 6087 3035
rect 6113 3013 6142 3035
rect 6168 3013 6175 3039
rect 6113 3009 6175 3013
rect 6075 3005 6175 3009
rect 5551 2984 5582 3005
rect 5972 2984 6008 3005
rect 5394 2983 5431 2984
rect 5393 2974 5431 2983
rect 5393 2954 5402 2974
rect 5422 2954 5431 2974
rect 5393 2946 5431 2954
rect 5497 2978 5582 2984
rect 5607 2983 5644 2984
rect 5497 2958 5505 2978
rect 5525 2958 5582 2978
rect 5497 2950 5582 2958
rect 5606 2974 5644 2983
rect 5606 2954 5615 2974
rect 5635 2954 5644 2974
rect 5497 2949 5533 2950
rect 5606 2946 5644 2954
rect 5710 2978 5795 2984
rect 5815 2983 5852 2984
rect 5710 2958 5718 2978
rect 5738 2977 5795 2978
rect 5738 2958 5767 2977
rect 5710 2957 5767 2958
rect 5788 2957 5795 2977
rect 5710 2950 5795 2957
rect 5814 2974 5852 2983
rect 5814 2954 5823 2974
rect 5843 2954 5852 2974
rect 5710 2949 5746 2950
rect 5814 2946 5852 2954
rect 5918 2978 6062 2984
rect 5918 2958 5926 2978
rect 5946 2975 6034 2978
rect 5946 2958 5977 2975
rect 5918 2955 5977 2958
rect 6000 2958 6034 2975
rect 6054 2958 6062 2978
rect 6000 2955 6062 2958
rect 5918 2950 6062 2955
rect 5918 2949 5954 2950
rect 6026 2949 6062 2950
rect 6128 2983 6165 2984
rect 6128 2982 6166 2983
rect 6128 2974 6192 2982
rect 6128 2954 6137 2974
rect 6157 2960 6192 2974
rect 6212 2960 6215 2980
rect 6157 2955 6215 2960
rect 6157 2954 6192 2955
rect 5394 2917 5431 2946
rect 5395 2915 5431 2917
rect 5607 2915 5644 2946
rect 5395 2893 5644 2915
rect 5815 2914 5852 2946
rect 6128 2942 6192 2954
rect 6232 2916 6259 3094
rect 7759 3001 7820 3108
rect 8787 3072 8814 3250
rect 8854 3212 8918 3224
rect 9194 3220 9231 3252
rect 9402 3251 9651 3273
rect 9692 3252 9878 3284
rect 9706 3251 9878 3252
rect 9402 3220 9439 3251
rect 9615 3249 9651 3251
rect 9615 3220 9652 3249
rect 9844 3223 9878 3251
rect 8854 3211 8889 3212
rect 8831 3206 8889 3211
rect 8831 3186 8834 3206
rect 8854 3192 8889 3206
rect 8909 3192 8918 3212
rect 8854 3184 8918 3192
rect 8880 3183 8918 3184
rect 8881 3182 8918 3183
rect 8984 3216 9020 3217
rect 9092 3216 9128 3217
rect 8984 3209 9128 3216
rect 8984 3208 9044 3209
rect 8984 3188 8992 3208
rect 9012 3189 9044 3208
rect 9069 3208 9128 3209
rect 9069 3189 9100 3208
rect 9012 3188 9100 3189
rect 9120 3188 9128 3208
rect 8984 3182 9128 3188
rect 9194 3212 9232 3220
rect 9300 3216 9336 3217
rect 9194 3192 9203 3212
rect 9223 3192 9232 3212
rect 9194 3183 9232 3192
rect 9251 3209 9336 3216
rect 9251 3189 9258 3209
rect 9279 3208 9336 3209
rect 9279 3189 9308 3208
rect 9251 3188 9308 3189
rect 9328 3188 9336 3208
rect 9194 3182 9231 3183
rect 9251 3182 9336 3188
rect 9402 3212 9440 3220
rect 9513 3216 9549 3217
rect 9402 3192 9411 3212
rect 9431 3192 9440 3212
rect 9402 3183 9440 3192
rect 9464 3208 9549 3216
rect 9464 3188 9521 3208
rect 9541 3188 9549 3208
rect 9402 3182 9439 3183
rect 9464 3182 9549 3188
rect 9615 3212 9653 3220
rect 9615 3192 9624 3212
rect 9644 3192 9653 3212
rect 9615 3183 9653 3192
rect 9842 3213 9879 3223
rect 9842 3195 9852 3213
rect 9870 3195 9879 3213
rect 9842 3186 9879 3195
rect 9844 3185 9878 3186
rect 9615 3182 9652 3183
rect 9038 3161 9074 3182
rect 9464 3161 9495 3182
rect 8871 3157 8971 3161
rect 8871 3153 8933 3157
rect 8871 3127 8878 3153
rect 8904 3131 8933 3153
rect 8959 3131 8971 3157
rect 8904 3127 8971 3131
rect 8871 3124 8971 3127
rect 9039 3124 9074 3161
rect 9136 3158 9495 3161
rect 9136 3153 9358 3158
rect 9136 3129 9149 3153
rect 9173 3134 9358 3153
rect 9382 3134 9495 3158
rect 9173 3129 9495 3134
rect 9136 3125 9495 3129
rect 9562 3153 9711 3161
rect 9562 3133 9573 3153
rect 9593 3133 9711 3153
rect 9562 3126 9711 3133
rect 9562 3125 9603 3126
rect 8886 3072 8923 3073
rect 8982 3072 9019 3073
rect 9038 3072 9074 3124
rect 9093 3072 9130 3073
rect 8786 3063 8924 3072
rect 7750 3000 7820 3001
rect 8411 3029 8522 3044
rect 8786 3043 8895 3063
rect 8915 3043 8924 3063
rect 8786 3036 8924 3043
rect 8982 3063 9130 3072
rect 8982 3043 8991 3063
rect 9011 3043 9101 3063
rect 9121 3043 9130 3063
rect 8786 3034 8882 3036
rect 8982 3033 9130 3043
rect 9189 3063 9226 3073
rect 9301 3072 9338 3073
rect 9282 3070 9338 3072
rect 9189 3043 9197 3063
rect 9217 3043 9226 3063
rect 9038 3032 9074 3033
rect 8411 3027 8453 3029
rect 8411 3007 8418 3027
rect 8437 3007 8453 3027
rect 7750 2999 7858 3000
rect 8411 2999 8453 3007
rect 8481 3027 8522 3029
rect 8481 3007 8495 3027
rect 8514 3007 8522 3027
rect 8481 2999 8522 3007
rect 7739 2998 7907 2999
rect 6526 2965 6636 2979
rect 6526 2962 6569 2965
rect 6526 2957 6530 2962
rect 6091 2914 6259 2916
rect 5815 2911 6259 2914
rect 5476 2887 5587 2893
rect 5476 2879 5517 2887
rect 5165 2824 5204 2868
rect 5476 2859 5484 2879
rect 5503 2859 5517 2879
rect 5476 2857 5517 2859
rect 5545 2879 5587 2887
rect 5545 2859 5561 2879
rect 5580 2859 5587 2879
rect 5545 2857 5587 2859
rect 5476 2843 5587 2857
rect 5813 2888 6259 2911
rect 3458 2804 3499 2805
rect 2782 2751 2819 2752
rect 2878 2751 2915 2752
rect 2934 2751 2970 2803
rect 2989 2751 3026 2752
rect 2682 2742 2820 2751
rect 2682 2722 2791 2742
rect 2811 2722 2820 2742
rect 2682 2715 2820 2722
rect 2878 2742 3026 2751
rect 2878 2722 2887 2742
rect 2907 2722 2997 2742
rect 3017 2722 3026 2742
rect 2682 2713 2778 2715
rect 2878 2712 3026 2722
rect 3085 2742 3122 2752
rect 3197 2751 3234 2752
rect 3178 2749 3234 2751
rect 3085 2722 3093 2742
rect 3113 2722 3122 2742
rect 2934 2711 2970 2712
rect 2782 2652 2819 2653
rect 3085 2652 3122 2722
rect 3147 2742 3234 2749
rect 3147 2739 3205 2742
rect 3147 2719 3152 2739
rect 3173 2722 3205 2739
rect 3225 2722 3234 2742
rect 3173 2719 3234 2722
rect 3147 2712 3234 2719
rect 3293 2742 3330 2752
rect 3293 2722 3301 2742
rect 3321 2722 3330 2742
rect 3147 2711 3178 2712
rect 2781 2651 3122 2652
rect 2706 2646 3122 2651
rect 2706 2626 2709 2646
rect 2729 2626 3122 2646
rect 3293 2643 3330 2722
rect 3360 2751 3391 2804
rect 4140 2776 4826 2809
rect 3410 2751 3447 2752
rect 3360 2742 3447 2751
rect 3360 2722 3418 2742
rect 3438 2722 3447 2742
rect 3360 2712 3447 2722
rect 3506 2742 3543 2752
rect 3506 2722 3514 2742
rect 3534 2722 3543 2742
rect 3360 2711 3391 2712
rect 3355 2643 3465 2656
rect 3506 2643 3543 2722
rect 3293 2641 3543 2643
rect 3293 2638 3394 2641
rect 3293 2619 3358 2638
rect 2173 2606 2252 2614
rect 2084 2604 2252 2606
rect 1808 2597 2252 2604
rect 3355 2611 3358 2619
rect 3387 2611 3394 2638
rect 3422 2614 3432 2641
rect 3461 2619 3543 2641
rect 3732 2688 3900 2689
rect 4140 2688 4178 2776
rect 4439 2774 4486 2776
rect 4786 2752 4826 2776
rect 5165 2800 5205 2824
rect 5505 2800 5552 2802
rect 5813 2800 5851 2888
rect 6091 2887 6259 2888
rect 6448 2935 6530 2957
rect 6559 2935 6569 2962
rect 6597 2938 6604 2965
rect 6633 2957 6636 2965
rect 7739 2972 8183 2998
rect 8411 2993 8522 2999
rect 7739 2970 7907 2972
rect 7739 2968 7858 2970
rect 6633 2938 6698 2957
rect 6597 2935 6698 2938
rect 6448 2933 6698 2935
rect 6448 2854 6485 2933
rect 6526 2920 6636 2933
rect 6600 2864 6631 2865
rect 6448 2834 6457 2854
rect 6477 2834 6485 2854
rect 6448 2824 6485 2834
rect 6544 2854 6631 2864
rect 6544 2834 6553 2854
rect 6573 2834 6631 2854
rect 6544 2825 6631 2834
rect 6544 2824 6581 2825
rect 5165 2767 5851 2800
rect 6600 2772 6631 2825
rect 6661 2854 6698 2933
rect 6869 2952 6901 2964
rect 6869 2932 6871 2952
rect 6892 2950 6901 2952
rect 6892 2948 7244 2950
rect 6892 2932 7262 2948
rect 6869 2930 7262 2932
rect 7282 2930 7285 2948
rect 6869 2925 7285 2930
rect 6869 2924 7210 2925
rect 6813 2864 6844 2865
rect 6661 2834 6670 2854
rect 6690 2834 6698 2854
rect 6661 2824 6698 2834
rect 6757 2857 6844 2864
rect 6757 2854 6818 2857
rect 6757 2834 6766 2854
rect 6786 2837 6818 2854
rect 6839 2837 6844 2857
rect 6786 2834 6844 2837
rect 6757 2827 6844 2834
rect 6869 2854 6906 2924
rect 7172 2923 7209 2924
rect 7021 2864 7057 2865
rect 6869 2834 6878 2854
rect 6898 2834 6906 2854
rect 6757 2825 6813 2827
rect 6757 2824 6794 2825
rect 6869 2824 6906 2834
rect 6965 2854 7113 2864
rect 7213 2861 7309 2863
rect 6965 2834 6974 2854
rect 6994 2845 7084 2854
rect 6994 2834 7025 2845
rect 6965 2825 7025 2834
rect 6965 2824 7002 2825
rect 7021 2813 7025 2825
rect 7052 2834 7084 2845
rect 7104 2834 7113 2854
rect 7052 2825 7113 2834
rect 7171 2854 7309 2861
rect 7171 2834 7180 2854
rect 7200 2834 7309 2854
rect 7171 2825 7309 2834
rect 7052 2813 7057 2825
rect 7076 2824 7113 2825
rect 7172 2824 7209 2825
rect 7021 2773 7057 2813
rect 6492 2771 6533 2772
rect 3732 2665 4178 2688
rect 4404 2719 4515 2733
rect 4404 2717 4446 2719
rect 4404 2697 4411 2717
rect 4430 2697 4446 2717
rect 4404 2689 4446 2697
rect 4474 2717 4515 2719
rect 4474 2697 4488 2717
rect 4507 2697 4515 2717
rect 4787 2708 4826 2752
rect 4474 2689 4515 2697
rect 4404 2683 4515 2689
rect 3732 2662 4176 2665
rect 3732 2660 3900 2662
rect 3461 2614 3465 2619
rect 3422 2611 3465 2614
rect 3355 2597 3465 2611
rect 1469 2577 1580 2583
rect 1808 2578 2178 2597
rect 2084 2577 2178 2578
rect 1469 2569 1510 2577
rect 1469 2549 1477 2569
rect 1496 2549 1510 2569
rect 1469 2547 1510 2549
rect 1538 2569 1580 2577
rect 1538 2549 1554 2569
rect 1573 2549 1580 2569
rect 2173 2568 2178 2577
rect 2226 2577 2252 2597
rect 2226 2568 2243 2577
rect 2173 2559 2243 2568
rect 1538 2547 1580 2549
rect 917 2543 953 2544
rect 765 2513 774 2533
rect 794 2513 802 2533
rect 653 2504 709 2506
rect 653 2503 690 2504
rect 765 2503 802 2513
rect 861 2533 1009 2543
rect 1109 2540 1205 2542
rect 861 2513 870 2533
rect 890 2513 980 2533
rect 1000 2513 1009 2533
rect 861 2504 1009 2513
rect 1067 2533 1205 2540
rect 1067 2513 1076 2533
rect 1096 2513 1205 2533
rect 1469 2532 1580 2547
rect 1067 2504 1205 2513
rect 861 2503 898 2504
rect 917 2452 953 2504
rect 972 2503 1009 2504
rect 1068 2503 1105 2504
rect 388 2450 429 2451
rect 280 2443 429 2450
rect 280 2423 398 2443
rect 418 2423 429 2443
rect 280 2415 429 2423
rect 496 2447 855 2451
rect 496 2442 818 2447
rect 496 2418 609 2442
rect 633 2423 818 2442
rect 842 2423 855 2447
rect 633 2418 855 2423
rect 496 2415 855 2418
rect 917 2415 952 2452
rect 1020 2449 1120 2452
rect 1020 2445 1087 2449
rect 1020 2419 1032 2445
rect 1058 2423 1087 2445
rect 1113 2423 1120 2449
rect 1058 2419 1120 2423
rect 1020 2415 1120 2419
rect 496 2394 527 2415
rect 917 2394 953 2415
rect 339 2393 376 2394
rect 113 2390 147 2391
rect 112 2381 149 2390
rect 112 2363 121 2381
rect 139 2363 149 2381
rect 112 2353 149 2363
rect 338 2384 376 2393
rect 338 2364 347 2384
rect 367 2364 376 2384
rect 338 2356 376 2364
rect 442 2388 527 2394
rect 552 2393 589 2394
rect 442 2368 450 2388
rect 470 2368 527 2388
rect 442 2360 527 2368
rect 551 2384 589 2393
rect 551 2364 560 2384
rect 580 2364 589 2384
rect 442 2359 478 2360
rect 551 2356 589 2364
rect 655 2388 740 2394
rect 760 2393 797 2394
rect 655 2368 663 2388
rect 683 2387 740 2388
rect 683 2368 712 2387
rect 655 2367 712 2368
rect 733 2367 740 2387
rect 655 2360 740 2367
rect 759 2384 797 2393
rect 759 2364 768 2384
rect 788 2364 797 2384
rect 655 2359 691 2360
rect 759 2356 797 2364
rect 863 2388 1007 2394
rect 863 2368 871 2388
rect 891 2387 979 2388
rect 891 2368 922 2387
rect 863 2367 922 2368
rect 947 2368 979 2387
rect 999 2368 1007 2388
rect 947 2367 1007 2368
rect 863 2360 1007 2367
rect 863 2359 899 2360
rect 971 2359 1007 2360
rect 1073 2393 1110 2394
rect 1073 2392 1111 2393
rect 1073 2384 1137 2392
rect 1073 2364 1082 2384
rect 1102 2370 1137 2384
rect 1157 2370 1160 2390
rect 1102 2365 1160 2370
rect 1102 2364 1137 2365
rect 113 2325 147 2353
rect 339 2327 376 2356
rect 340 2325 376 2327
rect 552 2325 589 2356
rect 113 2324 285 2325
rect 113 2292 299 2324
rect 340 2303 589 2325
rect 760 2324 797 2356
rect 1073 2352 1137 2364
rect 1177 2326 1204 2504
rect 3732 2482 3759 2660
rect 3799 2622 3863 2634
rect 4139 2630 4176 2662
rect 4347 2661 4596 2683
rect 4347 2630 4384 2661
rect 4560 2659 4596 2661
rect 4560 2630 4597 2659
rect 3799 2621 3834 2622
rect 3776 2616 3834 2621
rect 3776 2596 3779 2616
rect 3799 2602 3834 2616
rect 3854 2602 3863 2622
rect 3799 2594 3863 2602
rect 3825 2593 3863 2594
rect 3826 2592 3863 2593
rect 3929 2626 3965 2627
rect 4037 2626 4073 2627
rect 3929 2621 4073 2626
rect 3929 2618 3991 2621
rect 3929 2598 3937 2618
rect 3957 2601 3991 2618
rect 4014 2618 4073 2621
rect 4014 2601 4045 2618
rect 3957 2598 4045 2601
rect 4065 2598 4073 2618
rect 3929 2592 4073 2598
rect 4139 2622 4177 2630
rect 4245 2626 4281 2627
rect 4139 2602 4148 2622
rect 4168 2602 4177 2622
rect 4139 2593 4177 2602
rect 4196 2619 4281 2626
rect 4196 2599 4203 2619
rect 4224 2618 4281 2619
rect 4224 2599 4253 2618
rect 4196 2598 4253 2599
rect 4273 2598 4281 2618
rect 4139 2592 4176 2593
rect 4196 2592 4281 2598
rect 4347 2622 4385 2630
rect 4458 2626 4494 2627
rect 4347 2602 4356 2622
rect 4376 2602 4385 2622
rect 4347 2593 4385 2602
rect 4409 2618 4494 2626
rect 4409 2598 4466 2618
rect 4486 2598 4494 2618
rect 4347 2592 4384 2593
rect 4409 2592 4494 2598
rect 4560 2622 4598 2630
rect 4560 2602 4569 2622
rect 4589 2602 4598 2622
rect 4560 2593 4598 2602
rect 4560 2592 4597 2593
rect 3983 2571 4019 2592
rect 4409 2571 4440 2592
rect 3816 2567 3916 2571
rect 3816 2563 3878 2567
rect 3816 2537 3823 2563
rect 3849 2541 3878 2563
rect 3904 2541 3916 2567
rect 3849 2537 3916 2541
rect 3816 2534 3916 2537
rect 3984 2534 4019 2571
rect 4081 2568 4440 2571
rect 4081 2563 4303 2568
rect 4081 2539 4094 2563
rect 4118 2544 4303 2563
rect 4327 2544 4440 2568
rect 4118 2539 4440 2544
rect 4081 2535 4440 2539
rect 4507 2563 4656 2571
rect 4507 2543 4518 2563
rect 4538 2543 4656 2563
rect 4507 2536 4656 2543
rect 4507 2535 4548 2536
rect 3831 2482 3868 2483
rect 3927 2482 3964 2483
rect 3983 2482 4019 2534
rect 4038 2482 4075 2483
rect 3731 2473 3869 2482
rect 3731 2453 3840 2473
rect 3860 2453 3869 2473
rect 3731 2446 3869 2453
rect 3927 2473 4075 2482
rect 3927 2453 3936 2473
rect 3956 2453 4046 2473
rect 4066 2453 4075 2473
rect 3731 2444 3827 2446
rect 3927 2443 4075 2453
rect 4134 2473 4171 2483
rect 4246 2482 4283 2483
rect 4227 2480 4283 2482
rect 4134 2453 4142 2473
rect 4162 2453 4171 2473
rect 3983 2442 4019 2443
rect 1360 2400 1470 2414
rect 1360 2397 1403 2400
rect 1360 2392 1364 2397
rect 1036 2324 1204 2326
rect 760 2318 1204 2324
rect 113 2260 147 2292
rect 109 2251 147 2260
rect 109 2233 119 2251
rect 137 2233 147 2251
rect 109 2227 147 2233
rect 265 2229 299 2292
rect 421 2297 532 2303
rect 421 2289 462 2297
rect 421 2269 429 2289
rect 448 2269 462 2289
rect 421 2267 462 2269
rect 490 2289 532 2297
rect 490 2269 506 2289
rect 525 2269 532 2289
rect 490 2267 532 2269
rect 421 2252 532 2267
rect 759 2298 1204 2318
rect 759 2229 797 2298
rect 1036 2297 1204 2298
rect 1282 2370 1364 2392
rect 1393 2370 1403 2397
rect 1431 2373 1438 2400
rect 1467 2392 1470 2400
rect 3465 2409 3576 2424
rect 3465 2407 3507 2409
rect 1467 2373 1532 2392
rect 1431 2370 1532 2373
rect 1282 2368 1532 2370
rect 1282 2289 1319 2368
rect 1360 2355 1470 2368
rect 1434 2299 1465 2300
rect 1282 2269 1291 2289
rect 1311 2269 1319 2289
rect 1282 2259 1319 2269
rect 1378 2289 1465 2299
rect 1378 2269 1387 2289
rect 1407 2269 1465 2289
rect 1378 2260 1465 2269
rect 1378 2259 1415 2260
rect 109 2223 146 2227
rect 265 2218 797 2229
rect 264 2202 797 2218
rect 1434 2207 1465 2260
rect 1495 2289 1532 2368
rect 1703 2365 2096 2385
rect 2116 2365 2119 2385
rect 3198 2380 3239 2389
rect 1703 2360 2119 2365
rect 2793 2378 2961 2379
rect 3198 2378 3207 2380
rect 1703 2359 2044 2360
rect 1647 2299 1678 2300
rect 1495 2269 1504 2289
rect 1524 2269 1532 2289
rect 1495 2259 1532 2269
rect 1591 2292 1678 2299
rect 1591 2289 1652 2292
rect 1591 2269 1600 2289
rect 1620 2272 1652 2289
rect 1673 2272 1678 2292
rect 1620 2269 1678 2272
rect 1591 2262 1678 2269
rect 1703 2289 1740 2359
rect 2006 2358 2043 2359
rect 2793 2358 3207 2378
rect 3233 2358 3239 2380
rect 3465 2387 3472 2407
rect 3491 2387 3507 2407
rect 3465 2379 3507 2387
rect 3535 2407 3576 2409
rect 3535 2387 3549 2407
rect 3568 2387 3576 2407
rect 3535 2379 3576 2387
rect 3831 2383 3868 2384
rect 4134 2383 4171 2453
rect 4196 2473 4283 2480
rect 4196 2470 4254 2473
rect 4196 2450 4201 2470
rect 4222 2453 4254 2470
rect 4274 2453 4283 2473
rect 4222 2450 4283 2453
rect 4196 2443 4283 2450
rect 4342 2473 4379 2483
rect 4342 2453 4350 2473
rect 4370 2453 4379 2473
rect 4196 2442 4227 2443
rect 3830 2382 4171 2383
rect 3465 2373 3576 2379
rect 3755 2377 4171 2382
rect 2793 2352 3239 2358
rect 2793 2350 2961 2352
rect 1855 2299 1891 2300
rect 1703 2269 1712 2289
rect 1732 2269 1740 2289
rect 1591 2260 1647 2262
rect 1591 2259 1628 2260
rect 1703 2259 1740 2269
rect 1799 2289 1947 2299
rect 2047 2296 2143 2298
rect 1799 2269 1808 2289
rect 1828 2269 1918 2289
rect 1938 2269 1947 2289
rect 1799 2260 1947 2269
rect 2005 2289 2143 2296
rect 2005 2269 2014 2289
rect 2034 2269 2143 2289
rect 2005 2260 2143 2269
rect 1799 2259 1836 2260
rect 1855 2208 1891 2260
rect 1910 2259 1947 2260
rect 2006 2259 2043 2260
rect 1326 2206 1367 2207
rect 264 2201 778 2202
rect 1218 2199 1367 2206
rect 1218 2179 1336 2199
rect 1356 2179 1367 2199
rect 1218 2171 1367 2179
rect 1434 2203 1793 2207
rect 1434 2198 1756 2203
rect 1434 2174 1547 2198
rect 1571 2179 1756 2198
rect 1780 2179 1793 2203
rect 1571 2174 1793 2179
rect 1434 2171 1793 2174
rect 1855 2171 1890 2208
rect 1958 2205 2058 2208
rect 1958 2201 2025 2205
rect 1958 2175 1970 2201
rect 1996 2179 2025 2201
rect 2051 2179 2058 2205
rect 1996 2175 2058 2179
rect 1958 2171 2058 2175
rect 112 2160 149 2161
rect 110 2152 150 2160
rect 110 2134 121 2152
rect 139 2134 150 2152
rect 1434 2150 1465 2171
rect 1855 2150 1891 2171
rect 1277 2149 1314 2150
rect 110 2086 150 2134
rect 1276 2140 1314 2149
rect 1276 2120 1285 2140
rect 1305 2120 1314 2140
rect 1276 2112 1314 2120
rect 1380 2144 1465 2150
rect 1490 2149 1527 2150
rect 1380 2124 1388 2144
rect 1408 2124 1465 2144
rect 1380 2116 1465 2124
rect 1489 2140 1527 2149
rect 1489 2120 1498 2140
rect 1518 2120 1527 2140
rect 1380 2115 1416 2116
rect 1489 2112 1527 2120
rect 1593 2144 1678 2150
rect 1698 2149 1735 2150
rect 1593 2124 1601 2144
rect 1621 2143 1678 2144
rect 1621 2124 1650 2143
rect 1593 2123 1650 2124
rect 1671 2123 1678 2143
rect 1593 2116 1678 2123
rect 1697 2140 1735 2149
rect 1697 2120 1706 2140
rect 1726 2120 1735 2140
rect 1593 2115 1629 2116
rect 1697 2112 1735 2120
rect 1801 2144 1945 2150
rect 1801 2124 1809 2144
rect 1829 2127 1865 2144
rect 1885 2127 1917 2144
rect 1829 2124 1917 2127
rect 1937 2124 1945 2144
rect 1801 2116 1945 2124
rect 1801 2115 1837 2116
rect 1909 2115 1945 2116
rect 2011 2149 2048 2150
rect 2011 2148 2049 2149
rect 2011 2140 2075 2148
rect 2011 2120 2020 2140
rect 2040 2126 2075 2140
rect 2095 2126 2098 2146
rect 2040 2121 2098 2126
rect 2040 2120 2075 2121
rect 421 2090 531 2104
rect 421 2087 464 2090
rect 110 2079 235 2086
rect 421 2082 425 2087
rect 110 2060 202 2079
rect 227 2060 235 2079
rect 110 2050 235 2060
rect 343 2060 425 2082
rect 454 2060 464 2087
rect 492 2063 499 2090
rect 528 2082 531 2090
rect 1277 2083 1314 2112
rect 528 2063 593 2082
rect 1278 2081 1314 2083
rect 1490 2081 1527 2112
rect 1698 2085 1735 2112
rect 2011 2108 2075 2120
rect 492 2060 593 2063
rect 343 2058 593 2060
rect 110 2030 150 2050
rect 109 2021 150 2030
rect 109 2003 119 2021
rect 137 2003 150 2021
rect 109 1994 150 2003
rect 109 1993 146 1994
rect 343 1979 380 2058
rect 421 2045 531 2058
rect 495 1989 526 1990
rect 343 1959 352 1979
rect 372 1959 380 1979
rect 343 1949 380 1959
rect 439 1979 526 1989
rect 439 1959 448 1979
rect 468 1959 526 1979
rect 439 1950 526 1959
rect 439 1949 476 1950
rect 112 1927 149 1931
rect 109 1922 149 1927
rect 109 1904 121 1922
rect 139 1904 149 1922
rect 109 1724 149 1904
rect 495 1897 526 1950
rect 556 1979 593 2058
rect 764 2055 1157 2075
rect 1177 2055 1180 2075
rect 1278 2059 1527 2081
rect 1696 2080 1737 2085
rect 2115 2082 2142 2260
rect 2793 2172 2820 2350
rect 3198 2347 3239 2352
rect 3408 2351 3657 2373
rect 3755 2357 3758 2377
rect 3778 2357 4171 2377
rect 4342 2374 4379 2453
rect 4409 2482 4440 2535
rect 4786 2528 4826 2708
rect 5164 2710 5203 2767
rect 5813 2765 5851 2767
rect 6384 2764 6533 2771
rect 6384 2744 6502 2764
rect 6522 2744 6533 2764
rect 6384 2736 6533 2744
rect 6600 2768 6959 2772
rect 6600 2763 6922 2768
rect 6600 2739 6713 2763
rect 6737 2744 6922 2763
rect 6946 2744 6959 2768
rect 6737 2739 6959 2744
rect 6600 2736 6959 2739
rect 7021 2736 7056 2773
rect 7124 2770 7224 2773
rect 7124 2766 7191 2770
rect 7124 2740 7136 2766
rect 7162 2744 7191 2766
rect 7217 2744 7224 2770
rect 7162 2740 7224 2744
rect 7124 2736 7224 2740
rect 6600 2715 6631 2736
rect 7021 2715 7057 2736
rect 6443 2714 6480 2715
rect 5164 2708 5212 2710
rect 5164 2690 5175 2708
rect 5193 2690 5212 2708
rect 6442 2705 6480 2714
rect 5164 2681 5212 2690
rect 5165 2680 5212 2681
rect 5478 2685 5588 2699
rect 5478 2682 5521 2685
rect 5478 2677 5482 2682
rect 5400 2655 5482 2677
rect 5511 2655 5521 2682
rect 5549 2658 5556 2685
rect 5585 2677 5588 2685
rect 6442 2685 6451 2705
rect 6471 2685 6480 2705
rect 6442 2677 6480 2685
rect 6546 2709 6631 2715
rect 6656 2714 6693 2715
rect 6546 2689 6554 2709
rect 6574 2689 6631 2709
rect 6546 2681 6631 2689
rect 6655 2705 6693 2714
rect 6655 2685 6664 2705
rect 6684 2685 6693 2705
rect 6546 2680 6582 2681
rect 6655 2677 6693 2685
rect 6759 2709 6844 2715
rect 6864 2714 6901 2715
rect 6759 2689 6767 2709
rect 6787 2708 6844 2709
rect 6787 2689 6816 2708
rect 6759 2688 6816 2689
rect 6837 2688 6844 2708
rect 6759 2681 6844 2688
rect 6863 2705 6901 2714
rect 6863 2685 6872 2705
rect 6892 2685 6901 2705
rect 6759 2680 6795 2681
rect 6863 2677 6901 2685
rect 6967 2709 7111 2715
rect 6967 2689 6975 2709
rect 6995 2689 7083 2709
rect 7103 2689 7111 2709
rect 6967 2681 7111 2689
rect 6967 2680 7003 2681
rect 7075 2680 7111 2681
rect 7177 2714 7214 2715
rect 7177 2713 7215 2714
rect 7177 2705 7241 2713
rect 7177 2685 7186 2705
rect 7206 2691 7241 2705
rect 7261 2691 7264 2711
rect 7206 2686 7264 2691
rect 7206 2685 7241 2686
rect 5585 2658 5650 2677
rect 5549 2655 5650 2658
rect 5400 2653 5650 2655
rect 5168 2617 5205 2618
rect 4786 2510 4796 2528
rect 4814 2510 4826 2528
rect 4786 2505 4826 2510
rect 5164 2614 5205 2617
rect 5164 2609 5206 2614
rect 5164 2591 5177 2609
rect 5195 2591 5206 2609
rect 5164 2577 5206 2591
rect 5244 2577 5291 2581
rect 5164 2571 5291 2577
rect 5164 2542 5252 2571
rect 5281 2542 5291 2571
rect 5400 2574 5437 2653
rect 5478 2640 5588 2653
rect 5552 2584 5583 2585
rect 5400 2554 5409 2574
rect 5429 2554 5437 2574
rect 5400 2544 5437 2554
rect 5496 2574 5583 2584
rect 5496 2554 5505 2574
rect 5525 2554 5583 2574
rect 5496 2545 5583 2554
rect 5496 2544 5533 2545
rect 5164 2538 5291 2542
rect 5164 2521 5203 2538
rect 5244 2537 5291 2538
rect 4786 2501 4823 2505
rect 5164 2503 5175 2521
rect 5193 2503 5203 2521
rect 5164 2494 5203 2503
rect 5165 2493 5202 2494
rect 5552 2492 5583 2545
rect 5613 2574 5650 2653
rect 5821 2650 6214 2670
rect 6234 2650 6237 2670
rect 5821 2645 6237 2650
rect 6443 2648 6480 2677
rect 6444 2646 6480 2648
rect 6656 2646 6693 2677
rect 5821 2644 6162 2645
rect 5765 2584 5796 2585
rect 5613 2554 5622 2574
rect 5642 2554 5650 2574
rect 5613 2544 5650 2554
rect 5709 2577 5796 2584
rect 5709 2574 5770 2577
rect 5709 2554 5718 2574
rect 5738 2557 5770 2574
rect 5791 2557 5796 2577
rect 5738 2554 5796 2557
rect 5709 2547 5796 2554
rect 5821 2574 5858 2644
rect 6124 2643 6161 2644
rect 6444 2624 6693 2646
rect 6864 2645 6901 2677
rect 7177 2673 7241 2685
rect 7281 2655 7308 2825
rect 7739 2792 7766 2968
rect 7806 2932 7870 2944
rect 8146 2940 8183 2972
rect 8354 2971 8603 2993
rect 8886 2973 8923 2974
rect 9189 2973 9226 3043
rect 9251 3063 9338 3070
rect 9251 3060 9309 3063
rect 9251 3040 9256 3060
rect 9277 3043 9309 3060
rect 9329 3043 9338 3063
rect 9277 3040 9338 3043
rect 9251 3033 9338 3040
rect 9397 3063 9434 3073
rect 9397 3043 9405 3063
rect 9425 3043 9434 3063
rect 9251 3032 9282 3033
rect 8885 2972 9226 2973
rect 8354 2940 8391 2971
rect 8567 2969 8603 2971
rect 8567 2940 8604 2969
rect 8810 2967 9226 2972
rect 8810 2947 8813 2967
rect 8833 2947 9226 2967
rect 9397 2964 9434 3043
rect 9464 3072 9495 3125
rect 9845 3123 9882 3124
rect 9844 3114 9883 3123
rect 9844 3096 9854 3114
rect 9872 3096 9883 3114
rect 9756 3079 9803 3080
rect 9844 3079 9883 3096
rect 9756 3075 9883 3079
rect 9514 3072 9551 3073
rect 9464 3063 9551 3072
rect 9464 3043 9522 3063
rect 9542 3043 9551 3063
rect 9464 3033 9551 3043
rect 9610 3063 9647 3073
rect 9610 3043 9618 3063
rect 9638 3043 9647 3063
rect 9464 3032 9495 3033
rect 9459 2964 9569 2977
rect 9610 2964 9647 3043
rect 9756 3046 9766 3075
rect 9795 3046 9883 3075
rect 9756 3040 9883 3046
rect 9756 3036 9803 3040
rect 9841 3026 9883 3040
rect 9841 3008 9852 3026
rect 9870 3008 9883 3026
rect 9841 3003 9883 3008
rect 9842 3000 9883 3003
rect 9842 2999 9879 3000
rect 9397 2962 9647 2964
rect 9397 2959 9498 2962
rect 9397 2940 9462 2959
rect 7806 2931 7841 2932
rect 7783 2926 7841 2931
rect 7783 2906 7786 2926
rect 7806 2912 7841 2926
rect 7861 2912 7870 2932
rect 7806 2904 7870 2912
rect 7832 2903 7870 2904
rect 7833 2902 7870 2903
rect 7936 2936 7972 2937
rect 8044 2936 8080 2937
rect 7936 2929 8080 2936
rect 7936 2928 7994 2929
rect 7936 2908 7944 2928
rect 7964 2910 7994 2928
rect 8023 2928 8080 2929
rect 8023 2910 8052 2928
rect 7964 2908 8052 2910
rect 8072 2908 8080 2928
rect 7936 2902 8080 2908
rect 8146 2932 8184 2940
rect 8252 2936 8288 2937
rect 8146 2912 8155 2932
rect 8175 2912 8184 2932
rect 8146 2903 8184 2912
rect 8203 2929 8288 2936
rect 8203 2909 8210 2929
rect 8231 2928 8288 2929
rect 8231 2909 8260 2928
rect 8203 2908 8260 2909
rect 8280 2908 8288 2928
rect 8146 2902 8183 2903
rect 8203 2902 8288 2908
rect 8354 2932 8392 2940
rect 8465 2936 8501 2937
rect 8354 2912 8363 2932
rect 8383 2912 8392 2932
rect 8354 2903 8392 2912
rect 8416 2928 8501 2936
rect 8416 2908 8473 2928
rect 8493 2908 8501 2928
rect 8354 2902 8391 2903
rect 8416 2902 8501 2908
rect 8567 2932 8605 2940
rect 8567 2912 8576 2932
rect 8596 2912 8605 2932
rect 9459 2932 9462 2940
rect 9491 2932 9498 2959
rect 9526 2935 9536 2962
rect 9565 2940 9647 2962
rect 9565 2935 9569 2940
rect 9526 2932 9569 2935
rect 9459 2918 9569 2932
rect 9835 2936 9882 2937
rect 9835 2927 9883 2936
rect 8567 2903 8605 2912
rect 9835 2909 9854 2927
rect 9872 2909 9883 2927
rect 9835 2907 9883 2909
rect 8567 2902 8604 2903
rect 7990 2881 8026 2902
rect 8416 2881 8447 2902
rect 7823 2877 7923 2881
rect 7823 2873 7885 2877
rect 7823 2847 7830 2873
rect 7856 2851 7885 2873
rect 7911 2851 7923 2877
rect 7856 2847 7923 2851
rect 7823 2844 7923 2847
rect 7991 2844 8026 2881
rect 8088 2878 8447 2881
rect 8088 2873 8310 2878
rect 8088 2849 8101 2873
rect 8125 2854 8310 2873
rect 8334 2854 8447 2878
rect 8125 2849 8447 2854
rect 8088 2845 8447 2849
rect 8514 2873 8663 2881
rect 8514 2853 8525 2873
rect 8545 2853 8663 2873
rect 8514 2846 8663 2853
rect 9196 2850 9234 2852
rect 9844 2850 9883 2907
rect 8514 2845 8555 2846
rect 7838 2792 7875 2793
rect 7934 2792 7971 2793
rect 7990 2792 8026 2844
rect 8045 2792 8082 2793
rect 7738 2783 7876 2792
rect 7738 2763 7847 2783
rect 7867 2763 7876 2783
rect 7738 2756 7876 2763
rect 7934 2783 8082 2792
rect 7934 2763 7943 2783
rect 7963 2763 8053 2783
rect 8073 2763 8082 2783
rect 7738 2754 7834 2756
rect 7934 2753 8082 2763
rect 8141 2783 8178 2793
rect 8253 2792 8290 2793
rect 8234 2790 8290 2792
rect 8141 2763 8149 2783
rect 8169 2763 8178 2783
rect 7990 2752 8026 2753
rect 7838 2693 7875 2694
rect 8141 2693 8178 2763
rect 8203 2783 8290 2790
rect 8203 2780 8261 2783
rect 8203 2760 8208 2780
rect 8229 2763 8261 2780
rect 8281 2763 8290 2783
rect 8229 2760 8290 2763
rect 8203 2753 8290 2760
rect 8349 2783 8386 2793
rect 8349 2763 8357 2783
rect 8377 2763 8386 2783
rect 8203 2752 8234 2753
rect 7837 2692 8178 2693
rect 7762 2687 8178 2692
rect 7762 2667 7765 2687
rect 7785 2667 8178 2687
rect 8349 2684 8386 2763
rect 8416 2792 8447 2845
rect 9196 2817 9882 2850
rect 8466 2792 8503 2793
rect 8416 2783 8503 2792
rect 8416 2763 8474 2783
rect 8494 2763 8503 2783
rect 8416 2753 8503 2763
rect 8562 2783 8599 2793
rect 8562 2763 8570 2783
rect 8590 2763 8599 2783
rect 8416 2752 8447 2753
rect 8411 2684 8521 2697
rect 8562 2684 8599 2763
rect 8349 2682 8599 2684
rect 8349 2679 8450 2682
rect 8349 2660 8414 2679
rect 7229 2647 7308 2655
rect 7140 2645 7308 2647
rect 6864 2638 7308 2645
rect 8411 2652 8414 2660
rect 8443 2652 8450 2679
rect 8478 2655 8488 2682
rect 8517 2660 8599 2682
rect 8788 2729 8956 2730
rect 9196 2729 9234 2817
rect 9495 2815 9542 2817
rect 9842 2793 9882 2817
rect 8788 2706 9234 2729
rect 9460 2760 9571 2774
rect 9460 2758 9502 2760
rect 9460 2738 9467 2758
rect 9486 2738 9502 2758
rect 9460 2730 9502 2738
rect 9530 2758 9571 2760
rect 9530 2738 9544 2758
rect 9563 2738 9571 2758
rect 9843 2749 9882 2793
rect 9530 2730 9571 2738
rect 9460 2724 9571 2730
rect 8788 2703 9232 2706
rect 8788 2701 8956 2703
rect 8517 2655 8521 2660
rect 8478 2652 8521 2655
rect 8411 2638 8521 2652
rect 6525 2618 6636 2624
rect 6864 2619 7234 2638
rect 7140 2618 7234 2619
rect 6525 2610 6566 2618
rect 6525 2590 6533 2610
rect 6552 2590 6566 2610
rect 6525 2588 6566 2590
rect 6594 2610 6636 2618
rect 6594 2590 6610 2610
rect 6629 2590 6636 2610
rect 7229 2609 7234 2618
rect 7282 2618 7308 2638
rect 7282 2609 7299 2618
rect 7229 2600 7299 2609
rect 6594 2588 6636 2590
rect 5973 2584 6009 2585
rect 5821 2554 5830 2574
rect 5850 2554 5858 2574
rect 5709 2545 5765 2547
rect 5709 2544 5746 2545
rect 5821 2544 5858 2554
rect 5917 2574 6065 2584
rect 6165 2581 6261 2583
rect 5917 2554 5926 2574
rect 5946 2554 6036 2574
rect 6056 2554 6065 2574
rect 5917 2545 6065 2554
rect 6123 2574 6261 2581
rect 6123 2554 6132 2574
rect 6152 2554 6261 2574
rect 6525 2573 6636 2588
rect 6123 2545 6261 2554
rect 5917 2544 5954 2545
rect 5973 2493 6009 2545
rect 6028 2544 6065 2545
rect 6124 2544 6161 2545
rect 5444 2491 5485 2492
rect 5336 2484 5485 2491
rect 4459 2482 4496 2483
rect 4409 2473 4496 2482
rect 4409 2453 4467 2473
rect 4487 2453 4496 2473
rect 4409 2443 4496 2453
rect 4555 2473 4592 2483
rect 4555 2453 4563 2473
rect 4583 2453 4592 2473
rect 5336 2464 5454 2484
rect 5474 2464 5485 2484
rect 5336 2456 5485 2464
rect 5552 2488 5911 2492
rect 5552 2483 5874 2488
rect 5552 2459 5665 2483
rect 5689 2464 5874 2483
rect 5898 2464 5911 2488
rect 5689 2459 5911 2464
rect 5552 2456 5911 2459
rect 5973 2456 6008 2493
rect 6076 2490 6176 2493
rect 6076 2486 6143 2490
rect 6076 2460 6088 2486
rect 6114 2464 6143 2486
rect 6169 2464 6176 2490
rect 6114 2460 6176 2464
rect 6076 2456 6176 2460
rect 4409 2442 4440 2443
rect 4404 2374 4514 2387
rect 4555 2374 4592 2453
rect 4789 2438 4826 2439
rect 4785 2429 4826 2438
rect 5552 2435 5583 2456
rect 5973 2435 6009 2456
rect 5395 2434 5432 2435
rect 5169 2431 5203 2432
rect 4785 2411 4798 2429
rect 4816 2411 4826 2429
rect 4785 2402 4826 2411
rect 5168 2422 5205 2431
rect 5168 2404 5177 2422
rect 5195 2404 5205 2422
rect 4785 2382 4825 2402
rect 5168 2394 5205 2404
rect 5394 2425 5432 2434
rect 5394 2405 5403 2425
rect 5423 2405 5432 2425
rect 5394 2397 5432 2405
rect 5498 2429 5583 2435
rect 5608 2434 5645 2435
rect 5498 2409 5506 2429
rect 5526 2409 5583 2429
rect 5498 2401 5583 2409
rect 5607 2425 5645 2434
rect 5607 2405 5616 2425
rect 5636 2405 5645 2425
rect 5498 2400 5534 2401
rect 5607 2397 5645 2405
rect 5711 2429 5796 2435
rect 5816 2434 5853 2435
rect 5711 2409 5719 2429
rect 5739 2428 5796 2429
rect 5739 2409 5768 2428
rect 5711 2408 5768 2409
rect 5789 2408 5796 2428
rect 5711 2401 5796 2408
rect 5815 2425 5853 2434
rect 5815 2405 5824 2425
rect 5844 2405 5853 2425
rect 5711 2400 5747 2401
rect 5815 2397 5853 2405
rect 5919 2429 6063 2435
rect 5919 2409 5927 2429
rect 5947 2428 6035 2429
rect 5947 2409 5978 2428
rect 5919 2408 5978 2409
rect 6003 2409 6035 2428
rect 6055 2409 6063 2429
rect 6003 2408 6063 2409
rect 5919 2401 6063 2408
rect 5919 2400 5955 2401
rect 6027 2400 6063 2401
rect 6129 2434 6166 2435
rect 6129 2433 6167 2434
rect 6129 2425 6193 2433
rect 6129 2405 6138 2425
rect 6158 2411 6193 2425
rect 6213 2411 6216 2431
rect 6158 2406 6216 2411
rect 6158 2405 6193 2406
rect 4342 2372 4592 2374
rect 4342 2369 4443 2372
rect 2860 2312 2924 2324
rect 3200 2320 3237 2347
rect 3408 2320 3445 2351
rect 3621 2349 3657 2351
rect 4342 2350 4407 2369
rect 3621 2320 3658 2349
rect 4404 2342 4407 2350
rect 4436 2342 4443 2369
rect 4471 2345 4481 2372
rect 4510 2350 4592 2372
rect 4700 2372 4825 2382
rect 4700 2353 4708 2372
rect 4733 2353 4825 2372
rect 4510 2345 4514 2350
rect 4700 2346 4825 2353
rect 4471 2342 4514 2345
rect 4404 2328 4514 2342
rect 2860 2311 2895 2312
rect 2837 2306 2895 2311
rect 2837 2286 2840 2306
rect 2860 2292 2895 2306
rect 2915 2292 2924 2312
rect 2860 2284 2924 2292
rect 2886 2283 2924 2284
rect 2887 2282 2924 2283
rect 2990 2316 3026 2317
rect 3098 2316 3134 2317
rect 2990 2308 3134 2316
rect 2990 2288 2998 2308
rect 3018 2288 3106 2308
rect 3126 2288 3134 2308
rect 2990 2282 3134 2288
rect 3200 2312 3238 2320
rect 3306 2316 3342 2317
rect 3200 2292 3209 2312
rect 3229 2292 3238 2312
rect 3200 2283 3238 2292
rect 3257 2309 3342 2316
rect 3257 2289 3264 2309
rect 3285 2308 3342 2309
rect 3285 2289 3314 2308
rect 3257 2288 3314 2289
rect 3334 2288 3342 2308
rect 3200 2282 3237 2283
rect 3257 2282 3342 2288
rect 3408 2312 3446 2320
rect 3519 2316 3555 2317
rect 3408 2292 3417 2312
rect 3437 2292 3446 2312
rect 3408 2283 3446 2292
rect 3470 2308 3555 2316
rect 3470 2288 3527 2308
rect 3547 2288 3555 2308
rect 3408 2282 3445 2283
rect 3470 2282 3555 2288
rect 3621 2312 3659 2320
rect 3621 2292 3630 2312
rect 3650 2292 3659 2312
rect 3621 2283 3659 2292
rect 4785 2298 4825 2346
rect 5169 2366 5203 2394
rect 5395 2368 5432 2397
rect 5396 2366 5432 2368
rect 5608 2366 5645 2397
rect 5169 2365 5341 2366
rect 5169 2333 5355 2365
rect 5396 2344 5645 2366
rect 5816 2365 5853 2397
rect 6129 2393 6193 2405
rect 6233 2367 6260 2545
rect 8788 2523 8815 2701
rect 8855 2663 8919 2675
rect 9195 2671 9232 2703
rect 9403 2702 9652 2724
rect 9403 2671 9440 2702
rect 9616 2700 9652 2702
rect 9616 2671 9653 2700
rect 8855 2662 8890 2663
rect 8832 2657 8890 2662
rect 8832 2637 8835 2657
rect 8855 2643 8890 2657
rect 8910 2643 8919 2663
rect 8855 2635 8919 2643
rect 8881 2634 8919 2635
rect 8882 2633 8919 2634
rect 8985 2667 9021 2668
rect 9093 2667 9129 2668
rect 8985 2662 9129 2667
rect 8985 2659 9047 2662
rect 8985 2639 8993 2659
rect 9013 2642 9047 2659
rect 9070 2659 9129 2662
rect 9070 2642 9101 2659
rect 9013 2639 9101 2642
rect 9121 2639 9129 2659
rect 8985 2633 9129 2639
rect 9195 2663 9233 2671
rect 9301 2667 9337 2668
rect 9195 2643 9204 2663
rect 9224 2643 9233 2663
rect 9195 2634 9233 2643
rect 9252 2660 9337 2667
rect 9252 2640 9259 2660
rect 9280 2659 9337 2660
rect 9280 2640 9309 2659
rect 9252 2639 9309 2640
rect 9329 2639 9337 2659
rect 9195 2633 9232 2634
rect 9252 2633 9337 2639
rect 9403 2663 9441 2671
rect 9514 2667 9550 2668
rect 9403 2643 9412 2663
rect 9432 2643 9441 2663
rect 9403 2634 9441 2643
rect 9465 2659 9550 2667
rect 9465 2639 9522 2659
rect 9542 2639 9550 2659
rect 9403 2633 9440 2634
rect 9465 2633 9550 2639
rect 9616 2663 9654 2671
rect 9616 2643 9625 2663
rect 9645 2643 9654 2663
rect 9616 2634 9654 2643
rect 9616 2633 9653 2634
rect 9039 2612 9075 2633
rect 9465 2612 9496 2633
rect 8872 2608 8972 2612
rect 8872 2604 8934 2608
rect 8872 2578 8879 2604
rect 8905 2582 8934 2604
rect 8960 2582 8972 2608
rect 8905 2578 8972 2582
rect 8872 2575 8972 2578
rect 9040 2575 9075 2612
rect 9137 2609 9496 2612
rect 9137 2604 9359 2609
rect 9137 2580 9150 2604
rect 9174 2585 9359 2604
rect 9383 2585 9496 2609
rect 9174 2580 9496 2585
rect 9137 2576 9496 2580
rect 9563 2604 9712 2612
rect 9563 2584 9574 2604
rect 9594 2584 9712 2604
rect 9563 2577 9712 2584
rect 9563 2576 9604 2577
rect 8887 2523 8924 2524
rect 8983 2523 9020 2524
rect 9039 2523 9075 2575
rect 9094 2523 9131 2524
rect 8787 2514 8925 2523
rect 8787 2494 8896 2514
rect 8916 2494 8925 2514
rect 8787 2487 8925 2494
rect 8983 2514 9131 2523
rect 8983 2494 8992 2514
rect 9012 2494 9102 2514
rect 9122 2494 9131 2514
rect 8787 2485 8883 2487
rect 8983 2484 9131 2494
rect 9190 2514 9227 2524
rect 9302 2523 9339 2524
rect 9283 2521 9339 2523
rect 9190 2494 9198 2514
rect 9218 2494 9227 2514
rect 9039 2483 9075 2484
rect 6416 2441 6526 2455
rect 6416 2438 6459 2441
rect 6416 2433 6420 2438
rect 6092 2365 6260 2367
rect 5816 2359 6260 2365
rect 5169 2301 5203 2333
rect 3621 2282 3658 2283
rect 3044 2261 3080 2282
rect 3470 2261 3501 2282
rect 4785 2280 4796 2298
rect 4814 2280 4825 2298
rect 4785 2272 4825 2280
rect 5165 2292 5203 2301
rect 5165 2274 5175 2292
rect 5193 2274 5203 2292
rect 4786 2271 4823 2272
rect 5165 2268 5203 2274
rect 5321 2270 5355 2333
rect 5477 2338 5588 2344
rect 5477 2330 5518 2338
rect 5477 2310 5485 2330
rect 5504 2310 5518 2330
rect 5477 2308 5518 2310
rect 5546 2330 5588 2338
rect 5546 2310 5562 2330
rect 5581 2310 5588 2330
rect 5546 2308 5588 2310
rect 5477 2293 5588 2308
rect 5815 2339 6260 2359
rect 5815 2270 5853 2339
rect 6092 2338 6260 2339
rect 6338 2411 6420 2433
rect 6449 2411 6459 2438
rect 6487 2414 6494 2441
rect 6523 2433 6526 2441
rect 8521 2450 8632 2465
rect 8521 2448 8563 2450
rect 6523 2414 6588 2433
rect 6487 2411 6588 2414
rect 6338 2409 6588 2411
rect 6338 2330 6375 2409
rect 6416 2396 6526 2409
rect 6490 2340 6521 2341
rect 6338 2310 6347 2330
rect 6367 2310 6375 2330
rect 6338 2300 6375 2310
rect 6434 2330 6521 2340
rect 6434 2310 6443 2330
rect 6463 2310 6521 2330
rect 6434 2301 6521 2310
rect 6434 2300 6471 2301
rect 5165 2264 5202 2268
rect 2877 2257 2977 2261
rect 2877 2253 2939 2257
rect 2877 2227 2884 2253
rect 2910 2231 2939 2253
rect 2965 2231 2977 2257
rect 2910 2227 2977 2231
rect 2877 2224 2977 2227
rect 3045 2224 3080 2261
rect 3142 2258 3501 2261
rect 3142 2253 3364 2258
rect 3142 2229 3155 2253
rect 3179 2234 3364 2253
rect 3388 2234 3501 2258
rect 3179 2229 3501 2234
rect 3142 2225 3501 2229
rect 3568 2253 3717 2261
rect 5321 2259 5853 2270
rect 3568 2233 3579 2253
rect 3599 2233 3717 2253
rect 5320 2243 5853 2259
rect 6490 2248 6521 2301
rect 6551 2330 6588 2409
rect 6759 2406 7152 2426
rect 7172 2406 7175 2426
rect 8254 2421 8295 2430
rect 6759 2401 7175 2406
rect 7849 2419 8017 2420
rect 8254 2419 8263 2421
rect 6759 2400 7100 2401
rect 6703 2340 6734 2341
rect 6551 2310 6560 2330
rect 6580 2310 6588 2330
rect 6551 2300 6588 2310
rect 6647 2333 6734 2340
rect 6647 2330 6708 2333
rect 6647 2310 6656 2330
rect 6676 2313 6708 2330
rect 6729 2313 6734 2333
rect 6676 2310 6734 2313
rect 6647 2303 6734 2310
rect 6759 2330 6796 2400
rect 7062 2399 7099 2400
rect 7849 2399 8263 2419
rect 8289 2399 8295 2421
rect 8521 2428 8528 2448
rect 8547 2428 8563 2448
rect 8521 2420 8563 2428
rect 8591 2448 8632 2450
rect 8591 2428 8605 2448
rect 8624 2428 8632 2448
rect 8591 2420 8632 2428
rect 8887 2424 8924 2425
rect 9190 2424 9227 2494
rect 9252 2514 9339 2521
rect 9252 2511 9310 2514
rect 9252 2491 9257 2511
rect 9278 2494 9310 2511
rect 9330 2494 9339 2514
rect 9278 2491 9339 2494
rect 9252 2484 9339 2491
rect 9398 2514 9435 2524
rect 9398 2494 9406 2514
rect 9426 2494 9435 2514
rect 9252 2483 9283 2484
rect 8886 2423 9227 2424
rect 8521 2414 8632 2420
rect 8811 2418 9227 2423
rect 7849 2393 8295 2399
rect 7849 2391 8017 2393
rect 6911 2340 6947 2341
rect 6759 2310 6768 2330
rect 6788 2310 6796 2330
rect 6647 2301 6703 2303
rect 6647 2300 6684 2301
rect 6759 2300 6796 2310
rect 6855 2330 7003 2340
rect 7103 2337 7199 2339
rect 6855 2310 6864 2330
rect 6884 2310 6974 2330
rect 6994 2310 7003 2330
rect 6855 2301 7003 2310
rect 7061 2330 7199 2337
rect 7061 2310 7070 2330
rect 7090 2310 7199 2330
rect 7061 2301 7199 2310
rect 6855 2300 6892 2301
rect 6911 2249 6947 2301
rect 6966 2300 7003 2301
rect 7062 2300 7099 2301
rect 6382 2247 6423 2248
rect 5320 2242 5834 2243
rect 3568 2226 3717 2233
rect 6274 2240 6423 2247
rect 4157 2230 4671 2231
rect 3568 2225 3609 2226
rect 3044 2189 3080 2224
rect 2892 2172 2929 2173
rect 2988 2172 3025 2173
rect 3044 2172 3051 2189
rect 2792 2163 2930 2172
rect 2792 2143 2901 2163
rect 2921 2143 2930 2163
rect 2792 2136 2930 2143
rect 2988 2163 3051 2172
rect 2988 2143 2997 2163
rect 3017 2148 3051 2163
rect 3072 2172 3080 2189
rect 3099 2172 3136 2173
rect 3072 2163 3136 2172
rect 3072 2148 3107 2163
rect 3017 2143 3107 2148
rect 3127 2143 3136 2163
rect 2792 2134 2888 2136
rect 2988 2133 3136 2143
rect 3195 2163 3232 2173
rect 3307 2172 3344 2173
rect 3288 2170 3344 2172
rect 3195 2143 3203 2163
rect 3223 2143 3232 2163
rect 3044 2132 3080 2133
rect 1974 2080 2142 2082
rect 1696 2074 2142 2080
rect 764 2050 1180 2055
rect 1359 2053 1470 2059
rect 764 2049 1105 2050
rect 708 1989 739 1990
rect 556 1959 565 1979
rect 585 1959 593 1979
rect 556 1949 593 1959
rect 652 1982 739 1989
rect 652 1979 713 1982
rect 652 1959 661 1979
rect 681 1962 713 1979
rect 734 1962 739 1982
rect 681 1959 739 1962
rect 652 1952 739 1959
rect 764 1979 801 2049
rect 1067 2048 1104 2049
rect 1359 2045 1400 2053
rect 1359 2025 1367 2045
rect 1386 2025 1400 2045
rect 1359 2023 1400 2025
rect 1428 2045 1470 2053
rect 1428 2025 1444 2045
rect 1463 2025 1470 2045
rect 1696 2052 1702 2074
rect 1728 2054 2142 2074
rect 2892 2073 2929 2074
rect 3195 2073 3232 2143
rect 3257 2163 3344 2170
rect 3257 2160 3315 2163
rect 3257 2140 3262 2160
rect 3283 2143 3315 2160
rect 3335 2143 3344 2163
rect 3283 2140 3344 2143
rect 3257 2133 3344 2140
rect 3403 2163 3440 2173
rect 3403 2143 3411 2163
rect 3431 2143 3440 2163
rect 3257 2132 3288 2133
rect 2891 2072 3232 2073
rect 1728 2052 1737 2054
rect 1974 2053 2142 2054
rect 2816 2071 3232 2072
rect 2816 2067 3192 2071
rect 1696 2043 1737 2052
rect 2816 2047 2819 2067
rect 2839 2054 3192 2067
rect 3224 2054 3232 2071
rect 2839 2047 3232 2054
rect 3403 2064 3440 2143
rect 3470 2172 3501 2225
rect 4138 2214 4671 2230
rect 6274 2220 6392 2240
rect 6412 2220 6423 2240
rect 4138 2203 4670 2214
rect 6274 2212 6423 2220
rect 6490 2244 6849 2248
rect 6490 2239 6812 2244
rect 6490 2215 6603 2239
rect 6627 2220 6812 2239
rect 6836 2220 6849 2244
rect 6627 2215 6849 2220
rect 6490 2212 6849 2215
rect 6911 2212 6946 2249
rect 7014 2246 7114 2249
rect 7014 2242 7081 2246
rect 7014 2216 7026 2242
rect 7052 2220 7081 2242
rect 7107 2220 7114 2246
rect 7052 2216 7114 2220
rect 7014 2212 7114 2216
rect 4789 2205 4826 2209
rect 3520 2172 3557 2173
rect 3470 2163 3557 2172
rect 3470 2143 3528 2163
rect 3548 2143 3557 2163
rect 3470 2133 3557 2143
rect 3616 2163 3653 2173
rect 3616 2143 3624 2163
rect 3644 2143 3653 2163
rect 3470 2132 3501 2133
rect 3465 2064 3575 2077
rect 3616 2064 3653 2143
rect 3403 2062 3653 2064
rect 3403 2059 3504 2062
rect 3403 2040 3468 2059
rect 1428 2023 1470 2025
rect 1359 2008 1470 2023
rect 3465 2032 3468 2040
rect 3497 2032 3504 2059
rect 3532 2035 3542 2062
rect 3571 2040 3653 2062
rect 3731 2134 3899 2135
rect 4138 2134 4176 2203
rect 3731 2114 4176 2134
rect 4403 2165 4514 2180
rect 4403 2163 4445 2165
rect 4403 2143 4410 2163
rect 4429 2143 4445 2163
rect 4403 2135 4445 2143
rect 4473 2163 4514 2165
rect 4473 2143 4487 2163
rect 4506 2143 4514 2163
rect 4473 2135 4514 2143
rect 4403 2129 4514 2135
rect 4636 2140 4670 2203
rect 4788 2199 4826 2205
rect 5168 2201 5205 2202
rect 4788 2181 4798 2199
rect 4816 2181 4826 2199
rect 4788 2172 4826 2181
rect 5166 2193 5206 2201
rect 5166 2175 5177 2193
rect 5195 2175 5206 2193
rect 6490 2191 6521 2212
rect 6911 2191 6947 2212
rect 6333 2190 6370 2191
rect 4788 2140 4822 2172
rect 3731 2108 4175 2114
rect 3731 2106 3899 2108
rect 3571 2035 3575 2040
rect 3532 2032 3575 2035
rect 3465 2018 3575 2032
rect 916 1989 952 1990
rect 764 1959 773 1979
rect 793 1959 801 1979
rect 652 1950 708 1952
rect 652 1949 689 1950
rect 764 1949 801 1959
rect 860 1979 1008 1989
rect 1108 1986 1204 1988
rect 860 1959 869 1979
rect 889 1959 979 1979
rect 999 1959 1008 1979
rect 860 1950 1008 1959
rect 1066 1979 1204 1986
rect 1066 1959 1075 1979
rect 1095 1959 1204 1979
rect 1066 1950 1204 1959
rect 860 1949 897 1950
rect 916 1898 952 1950
rect 971 1949 1008 1950
rect 1067 1949 1104 1950
rect 387 1896 428 1897
rect 279 1889 428 1896
rect 279 1869 397 1889
rect 417 1869 428 1889
rect 279 1861 428 1869
rect 495 1893 854 1897
rect 495 1888 817 1893
rect 495 1864 608 1888
rect 632 1869 817 1888
rect 841 1869 854 1893
rect 632 1864 854 1869
rect 495 1861 854 1864
rect 916 1861 951 1898
rect 1019 1895 1119 1898
rect 1019 1891 1086 1895
rect 1019 1865 1031 1891
rect 1057 1869 1086 1891
rect 1112 1869 1119 1895
rect 1057 1865 1119 1869
rect 1019 1861 1119 1865
rect 495 1840 526 1861
rect 916 1840 952 1861
rect 338 1839 375 1840
rect 337 1830 375 1839
rect 337 1810 346 1830
rect 366 1810 375 1830
rect 337 1802 375 1810
rect 441 1834 526 1840
rect 551 1839 588 1840
rect 441 1814 449 1834
rect 469 1814 526 1834
rect 441 1806 526 1814
rect 550 1830 588 1839
rect 550 1810 559 1830
rect 579 1810 588 1830
rect 441 1805 477 1806
rect 550 1802 588 1810
rect 654 1834 739 1840
rect 759 1839 796 1840
rect 654 1814 662 1834
rect 682 1833 739 1834
rect 682 1814 711 1833
rect 654 1813 711 1814
rect 732 1813 739 1833
rect 654 1806 739 1813
rect 758 1830 796 1839
rect 758 1810 767 1830
rect 787 1810 796 1830
rect 654 1805 690 1806
rect 758 1802 796 1810
rect 862 1834 1006 1840
rect 862 1814 870 1834
rect 890 1831 978 1834
rect 890 1814 921 1831
rect 862 1811 921 1814
rect 944 1814 978 1831
rect 998 1814 1006 1834
rect 944 1811 1006 1814
rect 862 1806 1006 1811
rect 862 1805 898 1806
rect 970 1805 1006 1806
rect 1072 1839 1109 1840
rect 1072 1838 1110 1839
rect 1072 1830 1136 1838
rect 1072 1810 1081 1830
rect 1101 1816 1136 1830
rect 1156 1816 1159 1836
rect 1101 1811 1159 1816
rect 1101 1810 1136 1811
rect 338 1773 375 1802
rect 339 1771 375 1773
rect 551 1771 588 1802
rect 339 1749 588 1771
rect 759 1770 796 1802
rect 1072 1798 1136 1810
rect 1176 1772 1203 1950
rect 3731 1928 3758 2106
rect 3798 2068 3862 2080
rect 4138 2076 4175 2108
rect 4346 2107 4595 2129
rect 4636 2108 4822 2140
rect 4650 2107 4822 2108
rect 4346 2076 4383 2107
rect 4559 2105 4595 2107
rect 4559 2076 4596 2105
rect 4788 2079 4822 2107
rect 5166 2127 5206 2175
rect 6332 2181 6370 2190
rect 6332 2161 6341 2181
rect 6361 2161 6370 2181
rect 6332 2153 6370 2161
rect 6436 2185 6521 2191
rect 6546 2190 6583 2191
rect 6436 2165 6444 2185
rect 6464 2165 6521 2185
rect 6436 2157 6521 2165
rect 6545 2181 6583 2190
rect 6545 2161 6554 2181
rect 6574 2161 6583 2181
rect 6436 2156 6472 2157
rect 6545 2153 6583 2161
rect 6649 2185 6734 2191
rect 6754 2190 6791 2191
rect 6649 2165 6657 2185
rect 6677 2184 6734 2185
rect 6677 2165 6706 2184
rect 6649 2164 6706 2165
rect 6727 2164 6734 2184
rect 6649 2157 6734 2164
rect 6753 2181 6791 2190
rect 6753 2161 6762 2181
rect 6782 2161 6791 2181
rect 6649 2156 6685 2157
rect 6753 2153 6791 2161
rect 6857 2185 7001 2191
rect 6857 2165 6865 2185
rect 6885 2168 6921 2185
rect 6941 2168 6973 2185
rect 6885 2165 6973 2168
rect 6993 2165 7001 2185
rect 6857 2157 7001 2165
rect 6857 2156 6893 2157
rect 6965 2156 7001 2157
rect 7067 2190 7104 2191
rect 7067 2189 7105 2190
rect 7067 2181 7131 2189
rect 7067 2161 7076 2181
rect 7096 2167 7131 2181
rect 7151 2167 7154 2187
rect 7096 2162 7154 2167
rect 7096 2161 7131 2162
rect 5477 2131 5587 2145
rect 5477 2128 5520 2131
rect 5166 2120 5291 2127
rect 5477 2123 5481 2128
rect 5166 2101 5258 2120
rect 5283 2101 5291 2120
rect 5166 2091 5291 2101
rect 5399 2101 5481 2123
rect 5510 2101 5520 2128
rect 5548 2104 5555 2131
rect 5584 2123 5587 2131
rect 6333 2124 6370 2153
rect 5584 2104 5649 2123
rect 6334 2122 6370 2124
rect 6546 2122 6583 2153
rect 6754 2126 6791 2153
rect 7067 2149 7131 2161
rect 5548 2101 5649 2104
rect 5399 2099 5649 2101
rect 3798 2067 3833 2068
rect 3775 2062 3833 2067
rect 3775 2042 3778 2062
rect 3798 2048 3833 2062
rect 3853 2048 3862 2068
rect 3798 2040 3862 2048
rect 3824 2039 3862 2040
rect 3825 2038 3862 2039
rect 3928 2072 3964 2073
rect 4036 2072 4072 2073
rect 3928 2065 4072 2072
rect 3928 2064 3988 2065
rect 3928 2044 3936 2064
rect 3956 2045 3988 2064
rect 4013 2064 4072 2065
rect 4013 2045 4044 2064
rect 3956 2044 4044 2045
rect 4064 2044 4072 2064
rect 3928 2038 4072 2044
rect 4138 2068 4176 2076
rect 4244 2072 4280 2073
rect 4138 2048 4147 2068
rect 4167 2048 4176 2068
rect 4138 2039 4176 2048
rect 4195 2065 4280 2072
rect 4195 2045 4202 2065
rect 4223 2064 4280 2065
rect 4223 2045 4252 2064
rect 4195 2044 4252 2045
rect 4272 2044 4280 2064
rect 4138 2038 4175 2039
rect 4195 2038 4280 2044
rect 4346 2068 4384 2076
rect 4457 2072 4493 2073
rect 4346 2048 4355 2068
rect 4375 2048 4384 2068
rect 4346 2039 4384 2048
rect 4408 2064 4493 2072
rect 4408 2044 4465 2064
rect 4485 2044 4493 2064
rect 4346 2038 4383 2039
rect 4408 2038 4493 2044
rect 4559 2068 4597 2076
rect 4559 2048 4568 2068
rect 4588 2048 4597 2068
rect 4559 2039 4597 2048
rect 4786 2069 4823 2079
rect 5166 2071 5206 2091
rect 4786 2051 4796 2069
rect 4814 2051 4823 2069
rect 4786 2042 4823 2051
rect 5165 2062 5206 2071
rect 5165 2044 5175 2062
rect 5193 2044 5206 2062
rect 4788 2041 4822 2042
rect 4559 2038 4596 2039
rect 3982 2017 4018 2038
rect 4408 2017 4439 2038
rect 5165 2035 5206 2044
rect 5165 2034 5202 2035
rect 5399 2020 5436 2099
rect 5477 2086 5587 2099
rect 5551 2030 5582 2031
rect 3815 2013 3915 2017
rect 3815 2009 3877 2013
rect 3815 1983 3822 2009
rect 3848 1987 3877 2009
rect 3903 1987 3915 2013
rect 3848 1983 3915 1987
rect 3815 1980 3915 1983
rect 3983 1980 4018 2017
rect 4080 2014 4439 2017
rect 4080 2009 4302 2014
rect 4080 1985 4093 2009
rect 4117 1990 4302 2009
rect 4326 1990 4439 2014
rect 4117 1985 4439 1990
rect 4080 1981 4439 1985
rect 4506 2009 4655 2017
rect 4506 1989 4517 2009
rect 4537 1989 4655 2009
rect 5399 2000 5408 2020
rect 5428 2000 5436 2020
rect 5399 1990 5436 2000
rect 5495 2020 5582 2030
rect 5495 2000 5504 2020
rect 5524 2000 5582 2020
rect 5495 1991 5582 2000
rect 5495 1990 5532 1991
rect 4506 1982 4655 1989
rect 4506 1981 4547 1982
rect 3830 1928 3867 1929
rect 3926 1928 3963 1929
rect 3982 1928 4018 1980
rect 4037 1928 4074 1929
rect 3730 1919 3868 1928
rect 3325 1898 3436 1913
rect 3325 1896 3367 1898
rect 2995 1875 3100 1877
rect 2653 1867 2821 1868
rect 2995 1867 3044 1875
rect 2653 1848 3044 1867
rect 3075 1848 3100 1875
rect 3325 1876 3332 1896
rect 3351 1876 3367 1896
rect 3325 1868 3367 1876
rect 3395 1896 3436 1898
rect 3395 1876 3409 1896
rect 3428 1876 3436 1896
rect 3730 1899 3839 1919
rect 3859 1899 3868 1919
rect 3730 1892 3868 1899
rect 3926 1919 4074 1928
rect 3926 1899 3935 1919
rect 3955 1899 4045 1919
rect 4065 1899 4074 1919
rect 3730 1890 3826 1892
rect 3926 1889 4074 1899
rect 4133 1919 4170 1929
rect 4245 1928 4282 1929
rect 4226 1926 4282 1928
rect 4133 1899 4141 1919
rect 4161 1899 4170 1919
rect 3982 1888 4018 1889
rect 3395 1868 3436 1876
rect 3325 1862 3436 1868
rect 2653 1841 3100 1848
rect 2653 1839 2821 1841
rect 1501 1808 1611 1822
rect 1501 1805 1544 1808
rect 1501 1800 1505 1805
rect 1035 1770 1203 1772
rect 759 1767 1203 1770
rect 420 1743 531 1749
rect 420 1735 461 1743
rect 109 1680 148 1724
rect 420 1715 428 1735
rect 447 1715 461 1735
rect 420 1713 461 1715
rect 489 1735 531 1743
rect 489 1715 505 1735
rect 524 1715 531 1735
rect 489 1713 531 1715
rect 420 1698 531 1713
rect 757 1744 1203 1767
rect 109 1656 149 1680
rect 449 1656 496 1658
rect 757 1656 795 1744
rect 1035 1743 1203 1744
rect 1423 1778 1505 1800
rect 1534 1778 1544 1805
rect 1572 1781 1579 1808
rect 1608 1800 1611 1808
rect 1608 1781 1673 1800
rect 1572 1778 1673 1781
rect 1423 1776 1673 1778
rect 1423 1697 1460 1776
rect 1501 1763 1611 1776
rect 1575 1707 1606 1708
rect 1423 1677 1432 1697
rect 1452 1677 1460 1697
rect 1423 1667 1460 1677
rect 1519 1697 1606 1707
rect 1519 1677 1528 1697
rect 1548 1677 1606 1697
rect 1519 1668 1606 1677
rect 1519 1667 1556 1668
rect 109 1623 795 1656
rect 109 1566 148 1623
rect 757 1621 795 1623
rect 1575 1615 1606 1668
rect 1636 1697 1673 1776
rect 1844 1789 2237 1793
rect 1844 1772 1863 1789
rect 1883 1773 2237 1789
rect 2257 1773 2260 1793
rect 1883 1772 2260 1773
rect 1844 1768 2260 1772
rect 1844 1767 2185 1768
rect 1788 1707 1819 1708
rect 1636 1677 1645 1697
rect 1665 1677 1673 1697
rect 1636 1667 1673 1677
rect 1732 1700 1819 1707
rect 1732 1697 1793 1700
rect 1732 1677 1741 1697
rect 1761 1680 1793 1697
rect 1814 1680 1819 1700
rect 1761 1677 1819 1680
rect 1732 1670 1819 1677
rect 1844 1697 1881 1767
rect 2147 1766 2184 1767
rect 1996 1707 2032 1708
rect 1844 1677 1853 1697
rect 1873 1677 1881 1697
rect 1732 1668 1788 1670
rect 1732 1667 1769 1668
rect 1844 1667 1881 1677
rect 1940 1697 2088 1707
rect 2256 1706 2285 1707
rect 2188 1704 2285 1706
rect 1940 1677 1949 1697
rect 1969 1693 2059 1697
rect 1969 1677 2002 1693
rect 1940 1668 2002 1677
rect 1940 1667 1977 1668
rect 1996 1655 2002 1668
rect 2025 1677 2059 1693
rect 2079 1677 2088 1697
rect 2025 1668 2088 1677
rect 2146 1697 2285 1704
rect 2146 1677 2155 1697
rect 2175 1677 2285 1697
rect 2146 1668 2285 1677
rect 2025 1655 2032 1668
rect 2051 1667 2088 1668
rect 2147 1667 2184 1668
rect 1996 1616 2032 1655
rect 1467 1614 1508 1615
rect 1359 1607 1508 1614
rect 1359 1587 1477 1607
rect 1497 1587 1508 1607
rect 1359 1579 1508 1587
rect 1575 1611 1934 1615
rect 1575 1606 1897 1611
rect 1575 1582 1688 1606
rect 1712 1587 1897 1606
rect 1921 1587 1934 1611
rect 1712 1582 1934 1587
rect 1575 1579 1934 1582
rect 1996 1579 2031 1616
rect 2099 1613 2199 1616
rect 2099 1609 2166 1613
rect 2099 1583 2111 1609
rect 2137 1587 2166 1609
rect 2192 1587 2199 1613
rect 2137 1583 2199 1587
rect 2099 1579 2199 1583
rect 109 1564 157 1566
rect 109 1546 120 1564
rect 138 1546 157 1564
rect 1575 1558 1606 1579
rect 1996 1558 2032 1579
rect 1418 1557 1455 1558
rect 109 1537 157 1546
rect 110 1536 157 1537
rect 423 1541 533 1555
rect 423 1538 466 1541
rect 423 1533 427 1538
rect 345 1511 427 1533
rect 456 1511 466 1538
rect 494 1514 501 1541
rect 530 1533 533 1541
rect 1417 1548 1455 1557
rect 530 1514 595 1533
rect 1417 1528 1426 1548
rect 1446 1528 1455 1548
rect 494 1511 595 1514
rect 345 1509 595 1511
rect 113 1473 150 1474
rect 109 1470 150 1473
rect 109 1465 151 1470
rect 109 1447 122 1465
rect 140 1447 151 1465
rect 109 1433 151 1447
rect 189 1433 236 1437
rect 109 1427 236 1433
rect 109 1398 197 1427
rect 226 1398 236 1427
rect 345 1430 382 1509
rect 423 1496 533 1509
rect 497 1440 528 1441
rect 345 1410 354 1430
rect 374 1410 382 1430
rect 345 1400 382 1410
rect 441 1430 528 1440
rect 441 1410 450 1430
rect 470 1410 528 1430
rect 441 1401 528 1410
rect 441 1400 478 1401
rect 109 1394 236 1398
rect 109 1377 148 1394
rect 189 1393 236 1394
rect 109 1359 120 1377
rect 138 1359 148 1377
rect 109 1350 148 1359
rect 110 1349 147 1350
rect 497 1348 528 1401
rect 558 1430 595 1509
rect 766 1506 1159 1526
rect 1179 1506 1182 1526
rect 1417 1520 1455 1528
rect 1521 1552 1606 1558
rect 1631 1557 1668 1558
rect 1521 1532 1529 1552
rect 1549 1532 1606 1552
rect 1521 1524 1606 1532
rect 1630 1548 1668 1557
rect 1630 1528 1639 1548
rect 1659 1528 1668 1548
rect 1521 1523 1557 1524
rect 1630 1520 1668 1528
rect 1734 1552 1819 1558
rect 1839 1557 1876 1558
rect 1734 1532 1742 1552
rect 1762 1551 1819 1552
rect 1762 1532 1791 1551
rect 1734 1531 1791 1532
rect 1812 1531 1819 1551
rect 1734 1524 1819 1531
rect 1838 1548 1876 1557
rect 1838 1528 1847 1548
rect 1867 1528 1876 1548
rect 1734 1523 1770 1524
rect 1838 1520 1876 1528
rect 1942 1552 2086 1558
rect 1942 1532 1950 1552
rect 1970 1532 2058 1552
rect 2078 1532 2086 1552
rect 1942 1524 2086 1532
rect 1942 1523 1978 1524
rect 2050 1523 2086 1524
rect 2152 1557 2189 1558
rect 2152 1556 2190 1557
rect 2152 1548 2216 1556
rect 2152 1528 2161 1548
rect 2181 1534 2216 1548
rect 2236 1534 2239 1554
rect 2181 1529 2239 1534
rect 2181 1528 2216 1529
rect 766 1501 1182 1506
rect 766 1500 1107 1501
rect 710 1440 741 1441
rect 558 1410 567 1430
rect 587 1410 595 1430
rect 558 1400 595 1410
rect 654 1433 741 1440
rect 654 1430 715 1433
rect 654 1410 663 1430
rect 683 1413 715 1430
rect 736 1413 741 1433
rect 683 1410 741 1413
rect 654 1403 741 1410
rect 766 1430 803 1500
rect 1069 1499 1106 1500
rect 1418 1491 1455 1520
rect 1419 1489 1455 1491
rect 1631 1489 1668 1520
rect 1419 1467 1668 1489
rect 1839 1488 1876 1520
rect 2152 1516 2216 1528
rect 2256 1490 2285 1668
rect 2653 1661 2680 1839
rect 2720 1801 2784 1813
rect 3060 1809 3097 1841
rect 3268 1840 3517 1862
rect 3268 1809 3305 1840
rect 3481 1838 3517 1840
rect 3481 1809 3518 1838
rect 3830 1829 3867 1830
rect 4133 1829 4170 1899
rect 4195 1919 4282 1926
rect 4195 1916 4253 1919
rect 4195 1896 4200 1916
rect 4221 1899 4253 1916
rect 4273 1899 4282 1919
rect 4221 1896 4282 1899
rect 4195 1889 4282 1896
rect 4341 1919 4378 1929
rect 4341 1899 4349 1919
rect 4369 1899 4378 1919
rect 4195 1888 4226 1889
rect 3829 1828 4170 1829
rect 3754 1823 4170 1828
rect 2720 1800 2755 1801
rect 2697 1795 2755 1800
rect 2697 1775 2700 1795
rect 2720 1781 2755 1795
rect 2775 1781 2784 1801
rect 2720 1773 2784 1781
rect 2746 1772 2784 1773
rect 2747 1771 2784 1772
rect 2850 1805 2886 1806
rect 2958 1805 2994 1806
rect 2850 1800 2994 1805
rect 2850 1797 2910 1800
rect 2850 1777 2858 1797
rect 2878 1779 2910 1797
rect 2937 1797 2994 1800
rect 2937 1779 2966 1797
rect 2878 1777 2966 1779
rect 2986 1777 2994 1797
rect 2850 1771 2994 1777
rect 3060 1801 3098 1809
rect 3166 1805 3202 1806
rect 3060 1781 3069 1801
rect 3089 1781 3098 1801
rect 3060 1772 3098 1781
rect 3117 1798 3202 1805
rect 3117 1778 3124 1798
rect 3145 1797 3202 1798
rect 3145 1778 3174 1797
rect 3117 1777 3174 1778
rect 3194 1777 3202 1797
rect 3060 1771 3097 1772
rect 3117 1771 3202 1777
rect 3268 1801 3306 1809
rect 3379 1805 3415 1806
rect 3268 1781 3277 1801
rect 3297 1781 3306 1801
rect 3268 1772 3306 1781
rect 3330 1797 3415 1805
rect 3330 1777 3387 1797
rect 3407 1777 3415 1797
rect 3268 1771 3305 1772
rect 3330 1771 3415 1777
rect 3481 1801 3519 1809
rect 3754 1803 3757 1823
rect 3777 1803 4170 1823
rect 4341 1820 4378 1899
rect 4408 1928 4439 1981
rect 4789 1979 4826 1980
rect 4788 1970 4827 1979
rect 4788 1952 4798 1970
rect 4816 1952 4827 1970
rect 5168 1968 5205 1972
rect 4700 1935 4747 1936
rect 4788 1935 4827 1952
rect 4700 1931 4827 1935
rect 4458 1928 4495 1929
rect 4408 1919 4495 1928
rect 4408 1899 4466 1919
rect 4486 1899 4495 1919
rect 4408 1889 4495 1899
rect 4554 1919 4591 1929
rect 4554 1899 4562 1919
rect 4582 1899 4591 1919
rect 4408 1888 4439 1889
rect 4403 1820 4513 1833
rect 4554 1820 4591 1899
rect 4700 1902 4710 1931
rect 4739 1902 4827 1931
rect 4700 1896 4827 1902
rect 4700 1892 4747 1896
rect 4785 1882 4827 1896
rect 4785 1864 4796 1882
rect 4814 1864 4827 1882
rect 4785 1859 4827 1864
rect 4786 1856 4827 1859
rect 5165 1963 5205 1968
rect 5165 1945 5177 1963
rect 5195 1945 5205 1963
rect 4786 1855 4823 1856
rect 4341 1818 4591 1820
rect 4341 1815 4442 1818
rect 3481 1781 3490 1801
rect 3510 1781 3519 1801
rect 4341 1796 4406 1815
rect 3481 1772 3519 1781
rect 4403 1788 4406 1796
rect 4435 1788 4442 1815
rect 4470 1791 4480 1818
rect 4509 1796 4591 1818
rect 4509 1791 4513 1796
rect 4470 1788 4513 1791
rect 4403 1774 4513 1788
rect 4779 1792 4826 1793
rect 4779 1783 4827 1792
rect 3481 1771 3518 1772
rect 2904 1750 2940 1771
rect 3330 1750 3361 1771
rect 4779 1765 4798 1783
rect 4816 1765 4827 1783
rect 4779 1763 4827 1765
rect 2737 1746 2837 1750
rect 2737 1742 2799 1746
rect 2737 1716 2744 1742
rect 2770 1720 2799 1742
rect 2825 1720 2837 1746
rect 2770 1716 2837 1720
rect 2737 1713 2837 1716
rect 2905 1713 2940 1750
rect 3002 1747 3361 1750
rect 3002 1742 3224 1747
rect 3002 1718 3015 1742
rect 3039 1723 3224 1742
rect 3248 1723 3361 1747
rect 3039 1718 3361 1723
rect 3002 1714 3361 1718
rect 3428 1742 3577 1750
rect 3428 1722 3439 1742
rect 3459 1722 3577 1742
rect 3428 1715 3577 1722
rect 3428 1714 3469 1715
rect 2752 1661 2789 1662
rect 2848 1661 2885 1662
rect 2904 1661 2940 1713
rect 2959 1661 2996 1662
rect 2652 1652 2790 1661
rect 2652 1632 2761 1652
rect 2781 1632 2790 1652
rect 2652 1625 2790 1632
rect 2848 1652 2996 1661
rect 2848 1632 2857 1652
rect 2877 1632 2967 1652
rect 2987 1632 2996 1652
rect 2652 1623 2748 1625
rect 2848 1622 2996 1632
rect 3055 1652 3092 1662
rect 3167 1661 3204 1662
rect 3148 1659 3204 1661
rect 3055 1632 3063 1652
rect 3083 1632 3092 1652
rect 2904 1621 2940 1622
rect 2752 1562 2789 1563
rect 3055 1562 3092 1632
rect 3117 1652 3204 1659
rect 3117 1649 3175 1652
rect 3117 1629 3122 1649
rect 3143 1632 3175 1649
rect 3195 1632 3204 1652
rect 3143 1629 3204 1632
rect 3117 1622 3204 1629
rect 3263 1652 3300 1662
rect 3263 1632 3271 1652
rect 3291 1632 3300 1652
rect 3117 1621 3148 1622
rect 2751 1561 3092 1562
rect 2676 1557 3092 1561
rect 2676 1556 3053 1557
rect 2676 1536 2679 1556
rect 2699 1540 3053 1556
rect 3073 1540 3092 1557
rect 2699 1536 3092 1540
rect 3263 1553 3300 1632
rect 3330 1661 3361 1714
rect 4141 1706 4179 1708
rect 4788 1706 4827 1763
rect 4141 1673 4827 1706
rect 3380 1661 3417 1662
rect 3330 1652 3417 1661
rect 3330 1632 3388 1652
rect 3408 1632 3417 1652
rect 3330 1622 3417 1632
rect 3476 1652 3513 1662
rect 3476 1632 3484 1652
rect 3504 1632 3513 1652
rect 3330 1621 3361 1622
rect 3325 1553 3435 1566
rect 3476 1553 3513 1632
rect 3263 1551 3513 1553
rect 3263 1548 3364 1551
rect 3263 1529 3328 1548
rect 3325 1521 3328 1529
rect 3357 1521 3364 1548
rect 3392 1524 3402 1551
rect 3431 1529 3513 1551
rect 3733 1585 3901 1586
rect 4141 1585 4179 1673
rect 4440 1671 4487 1673
rect 4787 1649 4827 1673
rect 3733 1562 4179 1585
rect 4405 1616 4516 1631
rect 4405 1614 4447 1616
rect 4405 1594 4412 1614
rect 4431 1594 4447 1614
rect 4405 1586 4447 1594
rect 4475 1614 4516 1616
rect 4475 1594 4489 1614
rect 4508 1594 4516 1614
rect 4788 1605 4827 1649
rect 4475 1586 4516 1594
rect 4405 1580 4516 1586
rect 3733 1559 4177 1562
rect 3733 1557 3901 1559
rect 3431 1524 3435 1529
rect 3392 1521 3435 1524
rect 3325 1507 3435 1521
rect 2115 1488 2285 1490
rect 1836 1481 2285 1488
rect 1500 1461 1611 1467
rect 1500 1453 1541 1461
rect 918 1440 954 1441
rect 766 1410 775 1430
rect 795 1410 803 1430
rect 654 1401 710 1403
rect 654 1400 691 1401
rect 766 1400 803 1410
rect 862 1430 1010 1440
rect 1110 1437 1206 1439
rect 862 1410 871 1430
rect 891 1410 981 1430
rect 1001 1410 1010 1430
rect 862 1401 1010 1410
rect 1068 1430 1206 1437
rect 1068 1410 1077 1430
rect 1097 1410 1206 1430
rect 1500 1433 1508 1453
rect 1527 1433 1541 1453
rect 1500 1431 1541 1433
rect 1569 1453 1611 1461
rect 1569 1433 1585 1453
rect 1604 1433 1611 1453
rect 1836 1454 1861 1481
rect 1892 1462 2285 1481
rect 1892 1454 1941 1462
rect 2115 1461 2285 1462
rect 1836 1452 1941 1454
rect 1569 1431 1611 1433
rect 1500 1416 1611 1431
rect 1068 1401 1206 1410
rect 862 1400 899 1401
rect 918 1349 954 1401
rect 973 1400 1010 1401
rect 1069 1400 1106 1401
rect 389 1347 430 1348
rect 281 1340 430 1347
rect 281 1320 399 1340
rect 419 1320 430 1340
rect 281 1312 430 1320
rect 497 1344 856 1348
rect 497 1339 819 1344
rect 497 1315 610 1339
rect 634 1320 819 1339
rect 843 1320 856 1344
rect 634 1315 856 1320
rect 497 1312 856 1315
rect 918 1312 953 1349
rect 1021 1346 1121 1349
rect 1021 1342 1088 1346
rect 1021 1316 1033 1342
rect 1059 1320 1088 1342
rect 1114 1320 1121 1346
rect 1059 1316 1121 1320
rect 1021 1312 1121 1316
rect 497 1291 528 1312
rect 918 1291 954 1312
rect 340 1290 377 1291
rect 114 1287 148 1288
rect 113 1278 150 1287
rect 113 1260 122 1278
rect 140 1260 150 1278
rect 113 1250 150 1260
rect 339 1281 377 1290
rect 339 1261 348 1281
rect 368 1261 377 1281
rect 339 1253 377 1261
rect 443 1285 528 1291
rect 553 1290 590 1291
rect 443 1265 451 1285
rect 471 1265 528 1285
rect 443 1257 528 1265
rect 552 1281 590 1290
rect 552 1261 561 1281
rect 581 1261 590 1281
rect 443 1256 479 1257
rect 552 1253 590 1261
rect 656 1285 741 1291
rect 761 1290 798 1291
rect 656 1265 664 1285
rect 684 1284 741 1285
rect 684 1265 713 1284
rect 656 1264 713 1265
rect 734 1264 741 1284
rect 656 1257 741 1264
rect 760 1281 798 1290
rect 760 1261 769 1281
rect 789 1261 798 1281
rect 656 1256 692 1257
rect 760 1253 798 1261
rect 864 1285 1008 1291
rect 864 1265 872 1285
rect 892 1284 980 1285
rect 892 1265 923 1284
rect 864 1264 923 1265
rect 948 1265 980 1284
rect 1000 1265 1008 1285
rect 948 1264 1008 1265
rect 864 1257 1008 1264
rect 864 1256 900 1257
rect 972 1256 1008 1257
rect 1074 1290 1111 1291
rect 1074 1289 1112 1290
rect 1074 1281 1138 1289
rect 1074 1261 1083 1281
rect 1103 1267 1138 1281
rect 1158 1267 1161 1287
rect 1103 1262 1161 1267
rect 1103 1261 1138 1262
rect 114 1222 148 1250
rect 340 1224 377 1253
rect 341 1222 377 1224
rect 553 1222 590 1253
rect 114 1221 286 1222
rect 114 1189 300 1221
rect 341 1200 590 1222
rect 761 1221 798 1253
rect 1074 1249 1138 1261
rect 1178 1223 1205 1401
rect 3733 1379 3760 1557
rect 3800 1519 3864 1531
rect 4140 1527 4177 1559
rect 4348 1558 4597 1580
rect 4348 1527 4385 1558
rect 4561 1556 4597 1558
rect 4561 1527 4598 1556
rect 3800 1518 3835 1519
rect 3777 1513 3835 1518
rect 3777 1493 3780 1513
rect 3800 1499 3835 1513
rect 3855 1499 3864 1519
rect 3800 1491 3864 1499
rect 3826 1490 3864 1491
rect 3827 1489 3864 1490
rect 3930 1523 3966 1524
rect 4038 1523 4074 1524
rect 3930 1518 4074 1523
rect 3930 1515 3992 1518
rect 3930 1495 3938 1515
rect 3958 1498 3992 1515
rect 4015 1515 4074 1518
rect 4015 1498 4046 1515
rect 3958 1495 4046 1498
rect 4066 1495 4074 1515
rect 3930 1489 4074 1495
rect 4140 1519 4178 1527
rect 4246 1523 4282 1524
rect 4140 1499 4149 1519
rect 4169 1499 4178 1519
rect 4140 1490 4178 1499
rect 4197 1516 4282 1523
rect 4197 1496 4204 1516
rect 4225 1515 4282 1516
rect 4225 1496 4254 1515
rect 4197 1495 4254 1496
rect 4274 1495 4282 1515
rect 4140 1489 4177 1490
rect 4197 1489 4282 1495
rect 4348 1519 4386 1527
rect 4459 1523 4495 1524
rect 4348 1499 4357 1519
rect 4377 1499 4386 1519
rect 4348 1490 4386 1499
rect 4410 1515 4495 1523
rect 4410 1495 4467 1515
rect 4487 1495 4495 1515
rect 4348 1489 4385 1490
rect 4410 1489 4495 1495
rect 4561 1519 4599 1527
rect 4561 1499 4570 1519
rect 4590 1499 4599 1519
rect 4561 1490 4599 1499
rect 4561 1489 4598 1490
rect 3984 1468 4020 1489
rect 4410 1468 4441 1489
rect 3817 1464 3917 1468
rect 3817 1460 3879 1464
rect 3817 1434 3824 1460
rect 3850 1438 3879 1460
rect 3905 1438 3917 1464
rect 3850 1434 3917 1438
rect 3817 1431 3917 1434
rect 3985 1431 4020 1468
rect 4082 1465 4441 1468
rect 4082 1460 4304 1465
rect 4082 1436 4095 1460
rect 4119 1441 4304 1460
rect 4328 1441 4441 1465
rect 4119 1436 4441 1441
rect 4082 1432 4441 1436
rect 4508 1460 4657 1468
rect 4508 1440 4519 1460
rect 4539 1440 4657 1460
rect 4508 1433 4657 1440
rect 4508 1432 4549 1433
rect 3832 1379 3869 1380
rect 3928 1379 3965 1380
rect 3984 1379 4020 1431
rect 4039 1379 4076 1380
rect 3732 1370 3870 1379
rect 3732 1350 3841 1370
rect 3861 1350 3870 1370
rect 3732 1343 3870 1350
rect 3928 1370 4076 1379
rect 3928 1350 3937 1370
rect 3957 1350 4047 1370
rect 4067 1350 4076 1370
rect 3732 1341 3828 1343
rect 3928 1340 4076 1350
rect 4135 1370 4172 1380
rect 4247 1379 4284 1380
rect 4228 1377 4284 1379
rect 4135 1350 4143 1370
rect 4163 1350 4172 1370
rect 3984 1339 4020 1340
rect 1361 1297 1471 1311
rect 1361 1294 1404 1297
rect 1361 1289 1365 1294
rect 1037 1221 1205 1223
rect 761 1215 1205 1221
rect 114 1157 148 1189
rect 110 1148 148 1157
rect 110 1130 120 1148
rect 138 1130 148 1148
rect 110 1124 148 1130
rect 266 1126 300 1189
rect 422 1194 533 1200
rect 422 1186 463 1194
rect 422 1166 430 1186
rect 449 1166 463 1186
rect 422 1164 463 1166
rect 491 1186 533 1194
rect 491 1166 507 1186
rect 526 1166 533 1186
rect 491 1164 533 1166
rect 422 1149 533 1164
rect 760 1195 1205 1215
rect 760 1126 798 1195
rect 1037 1194 1205 1195
rect 1283 1267 1365 1289
rect 1394 1267 1404 1294
rect 1432 1270 1439 1297
rect 1468 1289 1471 1297
rect 3466 1306 3577 1321
rect 3466 1304 3508 1306
rect 1468 1270 1533 1289
rect 1432 1267 1533 1270
rect 1283 1265 1533 1267
rect 1283 1186 1320 1265
rect 1361 1252 1471 1265
rect 1435 1196 1466 1197
rect 1283 1166 1292 1186
rect 1312 1166 1320 1186
rect 1283 1156 1320 1166
rect 1379 1186 1466 1196
rect 1379 1166 1388 1186
rect 1408 1166 1466 1186
rect 1379 1157 1466 1166
rect 1379 1156 1416 1157
rect 110 1120 147 1124
rect 266 1115 798 1126
rect 265 1099 798 1115
rect 1435 1104 1466 1157
rect 1496 1186 1533 1265
rect 1704 1275 2097 1282
rect 1704 1258 1712 1275
rect 1744 1262 2097 1275
rect 2117 1262 2120 1282
rect 3199 1277 3240 1286
rect 1744 1258 2120 1262
rect 1704 1257 2120 1258
rect 2794 1275 2962 1276
rect 3199 1275 3208 1277
rect 1704 1256 2045 1257
rect 1648 1196 1679 1197
rect 1496 1166 1505 1186
rect 1525 1166 1533 1186
rect 1496 1156 1533 1166
rect 1592 1189 1679 1196
rect 1592 1186 1653 1189
rect 1592 1166 1601 1186
rect 1621 1169 1653 1186
rect 1674 1169 1679 1189
rect 1621 1166 1679 1169
rect 1592 1159 1679 1166
rect 1704 1186 1741 1256
rect 2007 1255 2044 1256
rect 2794 1255 3208 1275
rect 3234 1255 3240 1277
rect 3466 1284 3473 1304
rect 3492 1284 3508 1304
rect 3466 1276 3508 1284
rect 3536 1304 3577 1306
rect 3536 1284 3550 1304
rect 3569 1284 3577 1304
rect 3536 1276 3577 1284
rect 3832 1280 3869 1281
rect 4135 1280 4172 1350
rect 4197 1370 4284 1377
rect 4197 1367 4255 1370
rect 4197 1347 4202 1367
rect 4223 1350 4255 1367
rect 4275 1350 4284 1370
rect 4223 1347 4284 1350
rect 4197 1340 4284 1347
rect 4343 1370 4380 1380
rect 4343 1350 4351 1370
rect 4371 1350 4380 1370
rect 4197 1339 4228 1340
rect 3831 1279 4172 1280
rect 3466 1270 3577 1276
rect 3756 1274 4172 1279
rect 2794 1249 3240 1255
rect 2794 1247 2962 1249
rect 1856 1196 1892 1197
rect 1704 1166 1713 1186
rect 1733 1166 1741 1186
rect 1592 1157 1648 1159
rect 1592 1156 1629 1157
rect 1704 1156 1741 1166
rect 1800 1186 1948 1196
rect 2048 1193 2144 1195
rect 1800 1166 1809 1186
rect 1829 1181 1919 1186
rect 1829 1166 1864 1181
rect 1800 1157 1864 1166
rect 1800 1156 1837 1157
rect 1856 1140 1864 1157
rect 1885 1166 1919 1181
rect 1939 1166 1948 1186
rect 1885 1157 1948 1166
rect 2006 1186 2144 1193
rect 2006 1166 2015 1186
rect 2035 1166 2144 1186
rect 2006 1157 2144 1166
rect 1885 1140 1892 1157
rect 1911 1156 1948 1157
rect 2007 1156 2044 1157
rect 1856 1105 1892 1140
rect 1327 1103 1368 1104
rect 265 1098 779 1099
rect 1219 1096 1368 1103
rect 1219 1076 1337 1096
rect 1357 1076 1368 1096
rect 1219 1068 1368 1076
rect 1435 1100 1794 1104
rect 1435 1095 1757 1100
rect 1435 1071 1548 1095
rect 1572 1076 1757 1095
rect 1781 1076 1794 1100
rect 1572 1071 1794 1076
rect 1435 1068 1794 1071
rect 1856 1068 1891 1105
rect 1959 1102 2059 1105
rect 1959 1098 2026 1102
rect 1959 1072 1971 1098
rect 1997 1076 2026 1098
rect 2052 1076 2059 1102
rect 1997 1072 2059 1076
rect 1959 1068 2059 1072
rect 113 1057 150 1058
rect 111 1049 151 1057
rect 111 1031 122 1049
rect 140 1031 151 1049
rect 1435 1047 1466 1068
rect 1856 1047 1892 1068
rect 1278 1046 1315 1047
rect 111 983 151 1031
rect 1277 1037 1315 1046
rect 1277 1017 1286 1037
rect 1306 1017 1315 1037
rect 1277 1009 1315 1017
rect 1381 1041 1466 1047
rect 1491 1046 1528 1047
rect 1381 1021 1389 1041
rect 1409 1021 1466 1041
rect 1381 1013 1466 1021
rect 1490 1037 1528 1046
rect 1490 1017 1499 1037
rect 1519 1017 1528 1037
rect 1381 1012 1417 1013
rect 1490 1009 1528 1017
rect 1594 1041 1679 1047
rect 1699 1046 1736 1047
rect 1594 1021 1602 1041
rect 1622 1040 1679 1041
rect 1622 1021 1651 1040
rect 1594 1020 1651 1021
rect 1672 1020 1679 1040
rect 1594 1013 1679 1020
rect 1698 1037 1736 1046
rect 1698 1017 1707 1037
rect 1727 1017 1736 1037
rect 1594 1012 1630 1013
rect 1698 1009 1736 1017
rect 1802 1041 1946 1047
rect 1802 1021 1810 1041
rect 1830 1021 1918 1041
rect 1938 1021 1946 1041
rect 1802 1013 1946 1021
rect 1802 1012 1838 1013
rect 1910 1012 1946 1013
rect 2012 1046 2049 1047
rect 2012 1045 2050 1046
rect 2012 1037 2076 1045
rect 2012 1017 2021 1037
rect 2041 1023 2076 1037
rect 2096 1023 2099 1043
rect 2041 1018 2099 1023
rect 2041 1017 2076 1018
rect 422 987 532 1001
rect 422 984 465 987
rect 111 976 236 983
rect 422 979 426 984
rect 111 957 203 976
rect 228 957 236 976
rect 111 947 236 957
rect 344 957 426 979
rect 455 957 465 984
rect 493 960 500 987
rect 529 979 532 987
rect 1278 980 1315 1009
rect 529 960 594 979
rect 1279 978 1315 980
rect 1491 978 1528 1009
rect 1699 982 1736 1009
rect 2012 1005 2076 1017
rect 493 957 594 960
rect 344 955 594 957
rect 111 927 151 947
rect 110 918 151 927
rect 110 900 120 918
rect 138 900 151 918
rect 110 891 151 900
rect 110 890 147 891
rect 344 876 381 955
rect 422 942 532 955
rect 496 886 527 887
rect 344 856 353 876
rect 373 856 381 876
rect 344 846 381 856
rect 440 876 527 886
rect 440 856 449 876
rect 469 856 527 876
rect 440 847 527 856
rect 440 846 477 847
rect 113 824 150 828
rect 110 819 150 824
rect 110 801 122 819
rect 140 801 150 819
rect 110 621 150 801
rect 496 794 527 847
rect 557 876 594 955
rect 765 952 1158 972
rect 1178 952 1181 972
rect 1279 956 1528 978
rect 1697 977 1738 982
rect 2116 979 2143 1157
rect 2794 1069 2821 1247
rect 3199 1244 3240 1249
rect 3409 1248 3658 1270
rect 3756 1254 3759 1274
rect 3779 1254 4172 1274
rect 4343 1271 4380 1350
rect 4410 1379 4441 1432
rect 4787 1425 4827 1605
rect 5165 1765 5205 1945
rect 5551 1938 5582 1991
rect 5612 2020 5649 2099
rect 5820 2096 6213 2116
rect 6233 2096 6236 2116
rect 6334 2100 6583 2122
rect 6752 2121 6793 2126
rect 7171 2123 7198 2301
rect 7849 2213 7876 2391
rect 8254 2388 8295 2393
rect 8464 2392 8713 2414
rect 8811 2398 8814 2418
rect 8834 2398 9227 2418
rect 9398 2415 9435 2494
rect 9465 2523 9496 2576
rect 9842 2569 9882 2749
rect 9842 2551 9852 2569
rect 9870 2551 9882 2569
rect 9842 2546 9882 2551
rect 9842 2542 9879 2546
rect 9515 2523 9552 2524
rect 9465 2514 9552 2523
rect 9465 2494 9523 2514
rect 9543 2494 9552 2514
rect 9465 2484 9552 2494
rect 9611 2514 9648 2524
rect 9611 2494 9619 2514
rect 9639 2494 9648 2514
rect 9465 2483 9496 2484
rect 9460 2415 9570 2428
rect 9611 2415 9648 2494
rect 9845 2479 9882 2480
rect 9841 2470 9882 2479
rect 9841 2452 9854 2470
rect 9872 2452 9882 2470
rect 9841 2443 9882 2452
rect 9841 2423 9881 2443
rect 9398 2413 9648 2415
rect 9398 2410 9499 2413
rect 7916 2353 7980 2365
rect 8256 2361 8293 2388
rect 8464 2361 8501 2392
rect 8677 2390 8713 2392
rect 9398 2391 9463 2410
rect 8677 2361 8714 2390
rect 9460 2383 9463 2391
rect 9492 2383 9499 2410
rect 9527 2386 9537 2413
rect 9566 2391 9648 2413
rect 9756 2413 9881 2423
rect 9756 2394 9764 2413
rect 9789 2394 9881 2413
rect 9566 2386 9570 2391
rect 9756 2387 9881 2394
rect 9527 2383 9570 2386
rect 9460 2369 9570 2383
rect 7916 2352 7951 2353
rect 7893 2347 7951 2352
rect 7893 2327 7896 2347
rect 7916 2333 7951 2347
rect 7971 2333 7980 2353
rect 7916 2325 7980 2333
rect 7942 2324 7980 2325
rect 7943 2323 7980 2324
rect 8046 2357 8082 2358
rect 8154 2357 8190 2358
rect 8046 2349 8190 2357
rect 8046 2329 8054 2349
rect 8074 2329 8162 2349
rect 8182 2329 8190 2349
rect 8046 2323 8190 2329
rect 8256 2353 8294 2361
rect 8362 2357 8398 2358
rect 8256 2333 8265 2353
rect 8285 2333 8294 2353
rect 8256 2324 8294 2333
rect 8313 2350 8398 2357
rect 8313 2330 8320 2350
rect 8341 2349 8398 2350
rect 8341 2330 8370 2349
rect 8313 2329 8370 2330
rect 8390 2329 8398 2349
rect 8256 2323 8293 2324
rect 8313 2323 8398 2329
rect 8464 2353 8502 2361
rect 8575 2357 8611 2358
rect 8464 2333 8473 2353
rect 8493 2333 8502 2353
rect 8464 2324 8502 2333
rect 8526 2349 8611 2357
rect 8526 2329 8583 2349
rect 8603 2329 8611 2349
rect 8464 2323 8501 2324
rect 8526 2323 8611 2329
rect 8677 2353 8715 2361
rect 8677 2333 8686 2353
rect 8706 2333 8715 2353
rect 8677 2324 8715 2333
rect 9841 2339 9881 2387
rect 8677 2323 8714 2324
rect 8100 2302 8136 2323
rect 8526 2302 8557 2323
rect 9841 2321 9852 2339
rect 9870 2321 9881 2339
rect 9841 2313 9881 2321
rect 9842 2312 9879 2313
rect 7933 2298 8033 2302
rect 7933 2294 7995 2298
rect 7933 2268 7940 2294
rect 7966 2272 7995 2294
rect 8021 2272 8033 2298
rect 7966 2268 8033 2272
rect 7933 2265 8033 2268
rect 8101 2265 8136 2302
rect 8198 2299 8557 2302
rect 8198 2294 8420 2299
rect 8198 2270 8211 2294
rect 8235 2275 8420 2294
rect 8444 2275 8557 2299
rect 8235 2270 8557 2275
rect 8198 2266 8557 2270
rect 8624 2294 8773 2302
rect 8624 2274 8635 2294
rect 8655 2274 8773 2294
rect 8624 2267 8773 2274
rect 9213 2271 9727 2272
rect 8624 2266 8665 2267
rect 8100 2230 8136 2265
rect 7948 2213 7985 2214
rect 8044 2213 8081 2214
rect 8100 2213 8107 2230
rect 7848 2204 7986 2213
rect 7848 2184 7957 2204
rect 7977 2184 7986 2204
rect 7848 2177 7986 2184
rect 8044 2204 8107 2213
rect 8044 2184 8053 2204
rect 8073 2189 8107 2204
rect 8128 2213 8136 2230
rect 8155 2213 8192 2214
rect 8128 2204 8192 2213
rect 8128 2189 8163 2204
rect 8073 2184 8163 2189
rect 8183 2184 8192 2204
rect 7848 2175 7944 2177
rect 8044 2174 8192 2184
rect 8251 2204 8288 2214
rect 8363 2213 8400 2214
rect 8344 2211 8400 2213
rect 8251 2184 8259 2204
rect 8279 2184 8288 2204
rect 8100 2173 8136 2174
rect 7030 2121 7198 2123
rect 6752 2115 7198 2121
rect 5820 2091 6236 2096
rect 6415 2094 6526 2100
rect 5820 2090 6161 2091
rect 5764 2030 5795 2031
rect 5612 2000 5621 2020
rect 5641 2000 5649 2020
rect 5612 1990 5649 2000
rect 5708 2023 5795 2030
rect 5708 2020 5769 2023
rect 5708 2000 5717 2020
rect 5737 2003 5769 2020
rect 5790 2003 5795 2023
rect 5737 2000 5795 2003
rect 5708 1993 5795 2000
rect 5820 2020 5857 2090
rect 6123 2089 6160 2090
rect 6415 2086 6456 2094
rect 6415 2066 6423 2086
rect 6442 2066 6456 2086
rect 6415 2064 6456 2066
rect 6484 2086 6526 2094
rect 6484 2066 6500 2086
rect 6519 2066 6526 2086
rect 6752 2093 6758 2115
rect 6784 2095 7198 2115
rect 7948 2114 7985 2115
rect 8251 2114 8288 2184
rect 8313 2204 8400 2211
rect 8313 2201 8371 2204
rect 8313 2181 8318 2201
rect 8339 2184 8371 2201
rect 8391 2184 8400 2204
rect 8339 2181 8400 2184
rect 8313 2174 8400 2181
rect 8459 2204 8496 2214
rect 8459 2184 8467 2204
rect 8487 2184 8496 2204
rect 8313 2173 8344 2174
rect 7947 2113 8288 2114
rect 6784 2093 6793 2095
rect 7030 2094 7198 2095
rect 7872 2112 8288 2113
rect 7872 2108 8248 2112
rect 6752 2084 6793 2093
rect 7872 2088 7875 2108
rect 7895 2095 8248 2108
rect 8280 2095 8288 2112
rect 7895 2088 8288 2095
rect 8459 2105 8496 2184
rect 8526 2213 8557 2266
rect 9194 2255 9727 2271
rect 9194 2244 9726 2255
rect 9845 2246 9882 2250
rect 8576 2213 8613 2214
rect 8526 2204 8613 2213
rect 8526 2184 8584 2204
rect 8604 2184 8613 2204
rect 8526 2174 8613 2184
rect 8672 2204 8709 2214
rect 8672 2184 8680 2204
rect 8700 2184 8709 2204
rect 8526 2173 8557 2174
rect 8521 2105 8631 2118
rect 8672 2105 8709 2184
rect 8459 2103 8709 2105
rect 8459 2100 8560 2103
rect 8459 2081 8524 2100
rect 6484 2064 6526 2066
rect 6415 2049 6526 2064
rect 8521 2073 8524 2081
rect 8553 2073 8560 2100
rect 8588 2076 8598 2103
rect 8627 2081 8709 2103
rect 8787 2175 8955 2176
rect 9194 2175 9232 2244
rect 8787 2155 9232 2175
rect 9459 2206 9570 2221
rect 9459 2204 9501 2206
rect 9459 2184 9466 2204
rect 9485 2184 9501 2204
rect 9459 2176 9501 2184
rect 9529 2204 9570 2206
rect 9529 2184 9543 2204
rect 9562 2184 9570 2204
rect 9529 2176 9570 2184
rect 9459 2170 9570 2176
rect 9692 2181 9726 2244
rect 9844 2240 9882 2246
rect 9844 2222 9854 2240
rect 9872 2222 9882 2240
rect 9844 2213 9882 2222
rect 9844 2181 9878 2213
rect 8787 2149 9231 2155
rect 8787 2147 8955 2149
rect 8627 2076 8631 2081
rect 8588 2073 8631 2076
rect 8521 2059 8631 2073
rect 5972 2030 6008 2031
rect 5820 2000 5829 2020
rect 5849 2000 5857 2020
rect 5708 1991 5764 1993
rect 5708 1990 5745 1991
rect 5820 1990 5857 2000
rect 5916 2020 6064 2030
rect 6164 2027 6260 2029
rect 5916 2000 5925 2020
rect 5945 2000 6035 2020
rect 6055 2000 6064 2020
rect 5916 1991 6064 2000
rect 6122 2020 6260 2027
rect 6122 2000 6131 2020
rect 6151 2000 6260 2020
rect 6122 1991 6260 2000
rect 5916 1990 5953 1991
rect 5972 1939 6008 1991
rect 6027 1990 6064 1991
rect 6123 1990 6160 1991
rect 5443 1937 5484 1938
rect 5335 1930 5484 1937
rect 5335 1910 5453 1930
rect 5473 1910 5484 1930
rect 5335 1902 5484 1910
rect 5551 1934 5910 1938
rect 5551 1929 5873 1934
rect 5551 1905 5664 1929
rect 5688 1910 5873 1929
rect 5897 1910 5910 1934
rect 5688 1905 5910 1910
rect 5551 1902 5910 1905
rect 5972 1902 6007 1939
rect 6075 1936 6175 1939
rect 6075 1932 6142 1936
rect 6075 1906 6087 1932
rect 6113 1910 6142 1932
rect 6168 1910 6175 1936
rect 6113 1906 6175 1910
rect 6075 1902 6175 1906
rect 5551 1881 5582 1902
rect 5972 1881 6008 1902
rect 5394 1880 5431 1881
rect 5393 1871 5431 1880
rect 5393 1851 5402 1871
rect 5422 1851 5431 1871
rect 5393 1843 5431 1851
rect 5497 1875 5582 1881
rect 5607 1880 5644 1881
rect 5497 1855 5505 1875
rect 5525 1855 5582 1875
rect 5497 1847 5582 1855
rect 5606 1871 5644 1880
rect 5606 1851 5615 1871
rect 5635 1851 5644 1871
rect 5497 1846 5533 1847
rect 5606 1843 5644 1851
rect 5710 1875 5795 1881
rect 5815 1880 5852 1881
rect 5710 1855 5718 1875
rect 5738 1874 5795 1875
rect 5738 1855 5767 1874
rect 5710 1854 5767 1855
rect 5788 1854 5795 1874
rect 5710 1847 5795 1854
rect 5814 1871 5852 1880
rect 5814 1851 5823 1871
rect 5843 1851 5852 1871
rect 5710 1846 5746 1847
rect 5814 1843 5852 1851
rect 5918 1875 6062 1881
rect 5918 1855 5926 1875
rect 5946 1872 6034 1875
rect 5946 1855 5977 1872
rect 5918 1852 5977 1855
rect 6000 1855 6034 1872
rect 6054 1855 6062 1875
rect 6000 1852 6062 1855
rect 5918 1847 6062 1852
rect 5918 1846 5954 1847
rect 6026 1846 6062 1847
rect 6128 1880 6165 1881
rect 6128 1879 6166 1880
rect 6128 1871 6192 1879
rect 6128 1851 6137 1871
rect 6157 1857 6192 1871
rect 6212 1857 6215 1877
rect 6157 1852 6215 1857
rect 6157 1851 6192 1852
rect 5394 1814 5431 1843
rect 5395 1812 5431 1814
rect 5607 1812 5644 1843
rect 5395 1790 5644 1812
rect 5815 1811 5852 1843
rect 6128 1839 6192 1851
rect 6232 1813 6259 1991
rect 8787 1969 8814 2147
rect 8854 2109 8918 2121
rect 9194 2117 9231 2149
rect 9402 2148 9651 2170
rect 9692 2149 9878 2181
rect 9706 2148 9878 2149
rect 9402 2117 9439 2148
rect 9615 2146 9651 2148
rect 9615 2117 9652 2146
rect 9844 2120 9878 2148
rect 8854 2108 8889 2109
rect 8831 2103 8889 2108
rect 8831 2083 8834 2103
rect 8854 2089 8889 2103
rect 8909 2089 8918 2109
rect 8854 2081 8918 2089
rect 8880 2080 8918 2081
rect 8881 2079 8918 2080
rect 8984 2113 9020 2114
rect 9092 2113 9128 2114
rect 8984 2106 9128 2113
rect 8984 2105 9044 2106
rect 8984 2085 8992 2105
rect 9012 2086 9044 2105
rect 9069 2105 9128 2106
rect 9069 2086 9100 2105
rect 9012 2085 9100 2086
rect 9120 2085 9128 2105
rect 8984 2079 9128 2085
rect 9194 2109 9232 2117
rect 9300 2113 9336 2114
rect 9194 2089 9203 2109
rect 9223 2089 9232 2109
rect 9194 2080 9232 2089
rect 9251 2106 9336 2113
rect 9251 2086 9258 2106
rect 9279 2105 9336 2106
rect 9279 2086 9308 2105
rect 9251 2085 9308 2086
rect 9328 2085 9336 2105
rect 9194 2079 9231 2080
rect 9251 2079 9336 2085
rect 9402 2109 9440 2117
rect 9513 2113 9549 2114
rect 9402 2089 9411 2109
rect 9431 2089 9440 2109
rect 9402 2080 9440 2089
rect 9464 2105 9549 2113
rect 9464 2085 9521 2105
rect 9541 2085 9549 2105
rect 9402 2079 9439 2080
rect 9464 2079 9549 2085
rect 9615 2109 9653 2117
rect 9615 2089 9624 2109
rect 9644 2089 9653 2109
rect 9615 2080 9653 2089
rect 9842 2110 9879 2120
rect 9842 2092 9852 2110
rect 9870 2092 9879 2110
rect 9842 2083 9879 2092
rect 9844 2082 9878 2083
rect 9615 2079 9652 2080
rect 9038 2058 9074 2079
rect 9464 2058 9495 2079
rect 8871 2054 8971 2058
rect 8871 2050 8933 2054
rect 8871 2024 8878 2050
rect 8904 2028 8933 2050
rect 8959 2028 8971 2054
rect 8904 2024 8971 2028
rect 8871 2021 8971 2024
rect 9039 2021 9074 2058
rect 9136 2055 9495 2058
rect 9136 2050 9358 2055
rect 9136 2026 9149 2050
rect 9173 2031 9358 2050
rect 9382 2031 9495 2055
rect 9173 2026 9495 2031
rect 9136 2022 9495 2026
rect 9562 2050 9711 2058
rect 9562 2030 9573 2050
rect 9593 2030 9711 2050
rect 9562 2023 9711 2030
rect 9562 2022 9603 2023
rect 8886 1969 8923 1970
rect 8982 1969 9019 1970
rect 9038 1969 9074 2021
rect 9093 1969 9130 1970
rect 8786 1960 8924 1969
rect 8381 1939 8492 1954
rect 8381 1937 8423 1939
rect 8051 1916 8156 1918
rect 7709 1908 7877 1909
rect 8051 1908 8100 1916
rect 7709 1889 8100 1908
rect 8131 1889 8156 1916
rect 8381 1917 8388 1937
rect 8407 1917 8423 1937
rect 8381 1909 8423 1917
rect 8451 1937 8492 1939
rect 8451 1917 8465 1937
rect 8484 1917 8492 1937
rect 8786 1940 8895 1960
rect 8915 1940 8924 1960
rect 8786 1933 8924 1940
rect 8982 1960 9130 1969
rect 8982 1940 8991 1960
rect 9011 1940 9101 1960
rect 9121 1940 9130 1960
rect 8786 1931 8882 1933
rect 8982 1930 9130 1940
rect 9189 1960 9226 1970
rect 9301 1969 9338 1970
rect 9282 1967 9338 1969
rect 9189 1940 9197 1960
rect 9217 1940 9226 1960
rect 9038 1929 9074 1930
rect 8451 1909 8492 1917
rect 8381 1903 8492 1909
rect 7709 1882 8156 1889
rect 7709 1880 7877 1882
rect 6557 1849 6667 1863
rect 6557 1846 6600 1849
rect 6557 1841 6561 1846
rect 6091 1811 6259 1813
rect 5815 1808 6259 1811
rect 5476 1784 5587 1790
rect 5476 1776 5517 1784
rect 5165 1721 5204 1765
rect 5476 1756 5484 1776
rect 5503 1756 5517 1776
rect 5476 1754 5517 1756
rect 5545 1776 5587 1784
rect 5545 1756 5561 1776
rect 5580 1756 5587 1776
rect 5545 1754 5587 1756
rect 5476 1739 5587 1754
rect 5813 1785 6259 1808
rect 5165 1697 5205 1721
rect 5505 1697 5552 1699
rect 5813 1697 5851 1785
rect 6091 1784 6259 1785
rect 6479 1819 6561 1841
rect 6590 1819 6600 1846
rect 6628 1822 6635 1849
rect 6664 1841 6667 1849
rect 6664 1822 6729 1841
rect 6628 1819 6729 1822
rect 6479 1817 6729 1819
rect 6479 1738 6516 1817
rect 6557 1804 6667 1817
rect 6631 1748 6662 1749
rect 6479 1718 6488 1738
rect 6508 1718 6516 1738
rect 6479 1708 6516 1718
rect 6575 1738 6662 1748
rect 6575 1718 6584 1738
rect 6604 1718 6662 1738
rect 6575 1709 6662 1718
rect 6575 1708 6612 1709
rect 5165 1664 5851 1697
rect 5165 1607 5204 1664
rect 5813 1662 5851 1664
rect 6631 1656 6662 1709
rect 6692 1738 6729 1817
rect 6900 1830 7293 1834
rect 6900 1813 6919 1830
rect 6939 1814 7293 1830
rect 7313 1814 7316 1834
rect 6939 1813 7316 1814
rect 6900 1809 7316 1813
rect 6900 1808 7241 1809
rect 6844 1748 6875 1749
rect 6692 1718 6701 1738
rect 6721 1718 6729 1738
rect 6692 1708 6729 1718
rect 6788 1741 6875 1748
rect 6788 1738 6849 1741
rect 6788 1718 6797 1738
rect 6817 1721 6849 1738
rect 6870 1721 6875 1741
rect 6817 1718 6875 1721
rect 6788 1711 6875 1718
rect 6900 1738 6937 1808
rect 7203 1807 7240 1808
rect 7052 1748 7088 1749
rect 6900 1718 6909 1738
rect 6929 1718 6937 1738
rect 6788 1709 6844 1711
rect 6788 1708 6825 1709
rect 6900 1708 6937 1718
rect 6996 1738 7144 1748
rect 7312 1747 7341 1748
rect 7244 1745 7341 1747
rect 6996 1718 7005 1738
rect 7025 1734 7115 1738
rect 7025 1718 7058 1734
rect 6996 1709 7058 1718
rect 6996 1708 7033 1709
rect 7052 1696 7058 1709
rect 7081 1718 7115 1734
rect 7135 1718 7144 1738
rect 7081 1709 7144 1718
rect 7202 1738 7341 1745
rect 7202 1718 7211 1738
rect 7231 1718 7341 1738
rect 7202 1709 7341 1718
rect 7081 1696 7088 1709
rect 7107 1708 7144 1709
rect 7203 1708 7240 1709
rect 7052 1657 7088 1696
rect 6523 1655 6564 1656
rect 6415 1648 6564 1655
rect 6415 1628 6533 1648
rect 6553 1628 6564 1648
rect 6415 1620 6564 1628
rect 6631 1652 6990 1656
rect 6631 1647 6953 1652
rect 6631 1623 6744 1647
rect 6768 1628 6953 1647
rect 6977 1628 6990 1652
rect 6768 1623 6990 1628
rect 6631 1620 6990 1623
rect 7052 1620 7087 1657
rect 7155 1654 7255 1657
rect 7155 1650 7222 1654
rect 7155 1624 7167 1650
rect 7193 1628 7222 1650
rect 7248 1628 7255 1654
rect 7193 1624 7255 1628
rect 7155 1620 7255 1624
rect 5165 1605 5213 1607
rect 5165 1587 5176 1605
rect 5194 1587 5213 1605
rect 6631 1599 6662 1620
rect 7052 1599 7088 1620
rect 6474 1598 6511 1599
rect 5165 1578 5213 1587
rect 5166 1577 5213 1578
rect 5479 1582 5589 1596
rect 5479 1579 5522 1582
rect 5479 1574 5483 1579
rect 5401 1552 5483 1574
rect 5512 1552 5522 1579
rect 5550 1555 5557 1582
rect 5586 1574 5589 1582
rect 6473 1589 6511 1598
rect 5586 1555 5651 1574
rect 6473 1569 6482 1589
rect 6502 1569 6511 1589
rect 5550 1552 5651 1555
rect 5401 1550 5651 1552
rect 5169 1514 5206 1515
rect 4787 1407 4797 1425
rect 4815 1407 4827 1425
rect 4787 1402 4827 1407
rect 5165 1511 5206 1514
rect 5165 1506 5207 1511
rect 5165 1488 5178 1506
rect 5196 1488 5207 1506
rect 5165 1474 5207 1488
rect 5245 1474 5292 1478
rect 5165 1468 5292 1474
rect 5165 1439 5253 1468
rect 5282 1439 5292 1468
rect 5401 1471 5438 1550
rect 5479 1537 5589 1550
rect 5553 1481 5584 1482
rect 5401 1451 5410 1471
rect 5430 1451 5438 1471
rect 5401 1441 5438 1451
rect 5497 1471 5584 1481
rect 5497 1451 5506 1471
rect 5526 1451 5584 1471
rect 5497 1442 5584 1451
rect 5497 1441 5534 1442
rect 5165 1435 5292 1439
rect 5165 1418 5204 1435
rect 5245 1434 5292 1435
rect 4787 1398 4824 1402
rect 5165 1400 5176 1418
rect 5194 1400 5204 1418
rect 5165 1391 5204 1400
rect 5166 1390 5203 1391
rect 5553 1389 5584 1442
rect 5614 1471 5651 1550
rect 5822 1547 6215 1567
rect 6235 1547 6238 1567
rect 6473 1561 6511 1569
rect 6577 1593 6662 1599
rect 6687 1598 6724 1599
rect 6577 1573 6585 1593
rect 6605 1573 6662 1593
rect 6577 1565 6662 1573
rect 6686 1589 6724 1598
rect 6686 1569 6695 1589
rect 6715 1569 6724 1589
rect 6577 1564 6613 1565
rect 6686 1561 6724 1569
rect 6790 1593 6875 1599
rect 6895 1598 6932 1599
rect 6790 1573 6798 1593
rect 6818 1592 6875 1593
rect 6818 1573 6847 1592
rect 6790 1572 6847 1573
rect 6868 1572 6875 1592
rect 6790 1565 6875 1572
rect 6894 1589 6932 1598
rect 6894 1569 6903 1589
rect 6923 1569 6932 1589
rect 6790 1564 6826 1565
rect 6894 1561 6932 1569
rect 6998 1593 7142 1599
rect 6998 1573 7006 1593
rect 7026 1573 7114 1593
rect 7134 1573 7142 1593
rect 6998 1565 7142 1573
rect 6998 1564 7034 1565
rect 7106 1564 7142 1565
rect 7208 1598 7245 1599
rect 7208 1597 7246 1598
rect 7208 1589 7272 1597
rect 7208 1569 7217 1589
rect 7237 1575 7272 1589
rect 7292 1575 7295 1595
rect 7237 1570 7295 1575
rect 7237 1569 7272 1570
rect 5822 1542 6238 1547
rect 5822 1541 6163 1542
rect 5766 1481 5797 1482
rect 5614 1451 5623 1471
rect 5643 1451 5651 1471
rect 5614 1441 5651 1451
rect 5710 1474 5797 1481
rect 5710 1471 5771 1474
rect 5710 1451 5719 1471
rect 5739 1454 5771 1471
rect 5792 1454 5797 1474
rect 5739 1451 5797 1454
rect 5710 1444 5797 1451
rect 5822 1471 5859 1541
rect 6125 1540 6162 1541
rect 6474 1532 6511 1561
rect 6475 1530 6511 1532
rect 6687 1530 6724 1561
rect 6475 1508 6724 1530
rect 6895 1529 6932 1561
rect 7208 1557 7272 1569
rect 7312 1531 7341 1709
rect 7709 1702 7736 1880
rect 7776 1842 7840 1854
rect 8116 1850 8153 1882
rect 8324 1881 8573 1903
rect 8324 1850 8361 1881
rect 8537 1879 8573 1881
rect 8537 1850 8574 1879
rect 8886 1870 8923 1871
rect 9189 1870 9226 1940
rect 9251 1960 9338 1967
rect 9251 1957 9309 1960
rect 9251 1937 9256 1957
rect 9277 1940 9309 1957
rect 9329 1940 9338 1960
rect 9277 1937 9338 1940
rect 9251 1930 9338 1937
rect 9397 1960 9434 1970
rect 9397 1940 9405 1960
rect 9425 1940 9434 1960
rect 9251 1929 9282 1930
rect 8885 1869 9226 1870
rect 8810 1864 9226 1869
rect 7776 1841 7811 1842
rect 7753 1836 7811 1841
rect 7753 1816 7756 1836
rect 7776 1822 7811 1836
rect 7831 1822 7840 1842
rect 7776 1814 7840 1822
rect 7802 1813 7840 1814
rect 7803 1812 7840 1813
rect 7906 1846 7942 1847
rect 8014 1846 8050 1847
rect 7906 1841 8050 1846
rect 7906 1838 7966 1841
rect 7906 1818 7914 1838
rect 7934 1820 7966 1838
rect 7993 1838 8050 1841
rect 7993 1820 8022 1838
rect 7934 1818 8022 1820
rect 8042 1818 8050 1838
rect 7906 1812 8050 1818
rect 8116 1842 8154 1850
rect 8222 1846 8258 1847
rect 8116 1822 8125 1842
rect 8145 1822 8154 1842
rect 8116 1813 8154 1822
rect 8173 1839 8258 1846
rect 8173 1819 8180 1839
rect 8201 1838 8258 1839
rect 8201 1819 8230 1838
rect 8173 1818 8230 1819
rect 8250 1818 8258 1838
rect 8116 1812 8153 1813
rect 8173 1812 8258 1818
rect 8324 1842 8362 1850
rect 8435 1846 8471 1847
rect 8324 1822 8333 1842
rect 8353 1822 8362 1842
rect 8324 1813 8362 1822
rect 8386 1838 8471 1846
rect 8386 1818 8443 1838
rect 8463 1818 8471 1838
rect 8324 1812 8361 1813
rect 8386 1812 8471 1818
rect 8537 1842 8575 1850
rect 8810 1844 8813 1864
rect 8833 1844 9226 1864
rect 9397 1861 9434 1940
rect 9464 1969 9495 2022
rect 9845 2020 9882 2021
rect 9844 2011 9883 2020
rect 9844 1993 9854 2011
rect 9872 1993 9883 2011
rect 9756 1976 9803 1977
rect 9844 1976 9883 1993
rect 9756 1972 9883 1976
rect 9514 1969 9551 1970
rect 9464 1960 9551 1969
rect 9464 1940 9522 1960
rect 9542 1940 9551 1960
rect 9464 1930 9551 1940
rect 9610 1960 9647 1970
rect 9610 1940 9618 1960
rect 9638 1940 9647 1960
rect 9464 1929 9495 1930
rect 9459 1861 9569 1874
rect 9610 1861 9647 1940
rect 9756 1943 9766 1972
rect 9795 1943 9883 1972
rect 9756 1937 9883 1943
rect 9756 1933 9803 1937
rect 9841 1923 9883 1937
rect 9841 1905 9852 1923
rect 9870 1905 9883 1923
rect 9841 1900 9883 1905
rect 9842 1897 9883 1900
rect 9842 1896 9879 1897
rect 9397 1859 9647 1861
rect 9397 1856 9498 1859
rect 8537 1822 8546 1842
rect 8566 1822 8575 1842
rect 9397 1837 9462 1856
rect 8537 1813 8575 1822
rect 9459 1829 9462 1837
rect 9491 1829 9498 1856
rect 9526 1832 9536 1859
rect 9565 1837 9647 1859
rect 9565 1832 9569 1837
rect 9526 1829 9569 1832
rect 9459 1815 9569 1829
rect 9835 1833 9882 1834
rect 9835 1824 9883 1833
rect 8537 1812 8574 1813
rect 7960 1791 7996 1812
rect 8386 1791 8417 1812
rect 9835 1806 9854 1824
rect 9872 1806 9883 1824
rect 9835 1804 9883 1806
rect 7793 1787 7893 1791
rect 7793 1783 7855 1787
rect 7793 1757 7800 1783
rect 7826 1761 7855 1783
rect 7881 1761 7893 1787
rect 7826 1757 7893 1761
rect 7793 1754 7893 1757
rect 7961 1754 7996 1791
rect 8058 1788 8417 1791
rect 8058 1783 8280 1788
rect 8058 1759 8071 1783
rect 8095 1764 8280 1783
rect 8304 1764 8417 1788
rect 8095 1759 8417 1764
rect 8058 1755 8417 1759
rect 8484 1783 8633 1791
rect 8484 1763 8495 1783
rect 8515 1763 8633 1783
rect 8484 1756 8633 1763
rect 8484 1755 8525 1756
rect 7808 1702 7845 1703
rect 7904 1702 7941 1703
rect 7960 1702 7996 1754
rect 8015 1702 8052 1703
rect 7708 1693 7846 1702
rect 7708 1673 7817 1693
rect 7837 1673 7846 1693
rect 7708 1666 7846 1673
rect 7904 1693 8052 1702
rect 7904 1673 7913 1693
rect 7933 1673 8023 1693
rect 8043 1673 8052 1693
rect 7708 1664 7804 1666
rect 7904 1663 8052 1673
rect 8111 1693 8148 1703
rect 8223 1702 8260 1703
rect 8204 1700 8260 1702
rect 8111 1673 8119 1693
rect 8139 1673 8148 1693
rect 7960 1662 7996 1663
rect 7808 1603 7845 1604
rect 8111 1603 8148 1673
rect 8173 1693 8260 1700
rect 8173 1690 8231 1693
rect 8173 1670 8178 1690
rect 8199 1673 8231 1690
rect 8251 1673 8260 1693
rect 8199 1670 8260 1673
rect 8173 1663 8260 1670
rect 8319 1693 8356 1703
rect 8319 1673 8327 1693
rect 8347 1673 8356 1693
rect 8173 1662 8204 1663
rect 7807 1602 8148 1603
rect 7732 1598 8148 1602
rect 7732 1597 8109 1598
rect 7732 1577 7735 1597
rect 7755 1581 8109 1597
rect 8129 1581 8148 1598
rect 7755 1577 8148 1581
rect 8319 1594 8356 1673
rect 8386 1702 8417 1755
rect 9197 1747 9235 1749
rect 9844 1747 9883 1804
rect 9197 1714 9883 1747
rect 8436 1702 8473 1703
rect 8386 1693 8473 1702
rect 8386 1673 8444 1693
rect 8464 1673 8473 1693
rect 8386 1663 8473 1673
rect 8532 1693 8569 1703
rect 8532 1673 8540 1693
rect 8560 1673 8569 1693
rect 8386 1662 8417 1663
rect 8381 1594 8491 1607
rect 8532 1594 8569 1673
rect 8319 1592 8569 1594
rect 8319 1589 8420 1592
rect 8319 1570 8384 1589
rect 8381 1562 8384 1570
rect 8413 1562 8420 1589
rect 8448 1565 8458 1592
rect 8487 1570 8569 1592
rect 8789 1626 8957 1627
rect 9197 1626 9235 1714
rect 9496 1712 9543 1714
rect 9843 1690 9883 1714
rect 8789 1603 9235 1626
rect 9461 1657 9572 1672
rect 9461 1655 9503 1657
rect 9461 1635 9468 1655
rect 9487 1635 9503 1655
rect 9461 1627 9503 1635
rect 9531 1655 9572 1657
rect 9531 1635 9545 1655
rect 9564 1635 9572 1655
rect 9844 1646 9883 1690
rect 9531 1627 9572 1635
rect 9461 1621 9572 1627
rect 8789 1600 9233 1603
rect 8789 1598 8957 1600
rect 8487 1565 8491 1570
rect 8448 1562 8491 1565
rect 8381 1548 8491 1562
rect 7171 1529 7341 1531
rect 6892 1522 7341 1529
rect 6556 1502 6667 1508
rect 6556 1494 6597 1502
rect 5974 1481 6010 1482
rect 5822 1451 5831 1471
rect 5851 1451 5859 1471
rect 5710 1442 5766 1444
rect 5710 1441 5747 1442
rect 5822 1441 5859 1451
rect 5918 1471 6066 1481
rect 6166 1478 6262 1480
rect 5918 1451 5927 1471
rect 5947 1451 6037 1471
rect 6057 1451 6066 1471
rect 5918 1442 6066 1451
rect 6124 1471 6262 1478
rect 6124 1451 6133 1471
rect 6153 1451 6262 1471
rect 6556 1474 6564 1494
rect 6583 1474 6597 1494
rect 6556 1472 6597 1474
rect 6625 1494 6667 1502
rect 6625 1474 6641 1494
rect 6660 1474 6667 1494
rect 6892 1495 6917 1522
rect 6948 1503 7341 1522
rect 6948 1495 6997 1503
rect 7171 1502 7341 1503
rect 6892 1493 6997 1495
rect 6625 1472 6667 1474
rect 6556 1457 6667 1472
rect 6124 1442 6262 1451
rect 5918 1441 5955 1442
rect 5974 1390 6010 1442
rect 6029 1441 6066 1442
rect 6125 1441 6162 1442
rect 5445 1388 5486 1389
rect 5337 1381 5486 1388
rect 4460 1379 4497 1380
rect 4410 1370 4497 1379
rect 4410 1350 4468 1370
rect 4488 1350 4497 1370
rect 4410 1340 4497 1350
rect 4556 1370 4593 1380
rect 4556 1350 4564 1370
rect 4584 1350 4593 1370
rect 5337 1361 5455 1381
rect 5475 1361 5486 1381
rect 5337 1353 5486 1361
rect 5553 1385 5912 1389
rect 5553 1380 5875 1385
rect 5553 1356 5666 1380
rect 5690 1361 5875 1380
rect 5899 1361 5912 1385
rect 5690 1356 5912 1361
rect 5553 1353 5912 1356
rect 5974 1353 6009 1390
rect 6077 1387 6177 1390
rect 6077 1383 6144 1387
rect 6077 1357 6089 1383
rect 6115 1361 6144 1383
rect 6170 1361 6177 1387
rect 6115 1357 6177 1361
rect 6077 1353 6177 1357
rect 4410 1339 4441 1340
rect 4405 1271 4515 1284
rect 4556 1271 4593 1350
rect 4790 1335 4827 1336
rect 4786 1326 4827 1335
rect 5553 1332 5584 1353
rect 5974 1332 6010 1353
rect 5396 1331 5433 1332
rect 5170 1328 5204 1329
rect 4786 1308 4799 1326
rect 4817 1308 4827 1326
rect 4786 1299 4827 1308
rect 5169 1319 5206 1328
rect 5169 1301 5178 1319
rect 5196 1301 5206 1319
rect 4786 1279 4826 1299
rect 5169 1291 5206 1301
rect 5395 1322 5433 1331
rect 5395 1302 5404 1322
rect 5424 1302 5433 1322
rect 5395 1294 5433 1302
rect 5499 1326 5584 1332
rect 5609 1331 5646 1332
rect 5499 1306 5507 1326
rect 5527 1306 5584 1326
rect 5499 1298 5584 1306
rect 5608 1322 5646 1331
rect 5608 1302 5617 1322
rect 5637 1302 5646 1322
rect 5499 1297 5535 1298
rect 5608 1294 5646 1302
rect 5712 1326 5797 1332
rect 5817 1331 5854 1332
rect 5712 1306 5720 1326
rect 5740 1325 5797 1326
rect 5740 1306 5769 1325
rect 5712 1305 5769 1306
rect 5790 1305 5797 1325
rect 5712 1298 5797 1305
rect 5816 1322 5854 1331
rect 5816 1302 5825 1322
rect 5845 1302 5854 1322
rect 5712 1297 5748 1298
rect 5816 1294 5854 1302
rect 5920 1326 6064 1332
rect 5920 1306 5928 1326
rect 5948 1325 6036 1326
rect 5948 1306 5979 1325
rect 5920 1305 5979 1306
rect 6004 1306 6036 1325
rect 6056 1306 6064 1326
rect 6004 1305 6064 1306
rect 5920 1298 6064 1305
rect 5920 1297 5956 1298
rect 6028 1297 6064 1298
rect 6130 1331 6167 1332
rect 6130 1330 6168 1331
rect 6130 1322 6194 1330
rect 6130 1302 6139 1322
rect 6159 1308 6194 1322
rect 6214 1308 6217 1328
rect 6159 1303 6217 1308
rect 6159 1302 6194 1303
rect 4343 1269 4593 1271
rect 4343 1266 4444 1269
rect 2861 1209 2925 1221
rect 3201 1217 3238 1244
rect 3409 1217 3446 1248
rect 3622 1246 3658 1248
rect 4343 1247 4408 1266
rect 3622 1217 3659 1246
rect 4405 1239 4408 1247
rect 4437 1239 4444 1266
rect 4472 1242 4482 1269
rect 4511 1247 4593 1269
rect 4701 1269 4826 1279
rect 4701 1250 4709 1269
rect 4734 1250 4826 1269
rect 4511 1242 4515 1247
rect 4701 1243 4826 1250
rect 4472 1239 4515 1242
rect 4405 1225 4515 1239
rect 2861 1208 2896 1209
rect 2838 1203 2896 1208
rect 2838 1183 2841 1203
rect 2861 1189 2896 1203
rect 2916 1189 2925 1209
rect 2861 1181 2925 1189
rect 2887 1180 2925 1181
rect 2888 1179 2925 1180
rect 2991 1213 3027 1214
rect 3099 1213 3135 1214
rect 2991 1205 3135 1213
rect 2991 1185 2999 1205
rect 3019 1202 3107 1205
rect 3019 1185 3051 1202
rect 3071 1185 3107 1202
rect 3127 1185 3135 1205
rect 2991 1179 3135 1185
rect 3201 1209 3239 1217
rect 3307 1213 3343 1214
rect 3201 1189 3210 1209
rect 3230 1189 3239 1209
rect 3201 1180 3239 1189
rect 3258 1206 3343 1213
rect 3258 1186 3265 1206
rect 3286 1205 3343 1206
rect 3286 1186 3315 1205
rect 3258 1185 3315 1186
rect 3335 1185 3343 1205
rect 3201 1179 3238 1180
rect 3258 1179 3343 1185
rect 3409 1209 3447 1217
rect 3520 1213 3556 1214
rect 3409 1189 3418 1209
rect 3438 1189 3447 1209
rect 3409 1180 3447 1189
rect 3471 1205 3556 1213
rect 3471 1185 3528 1205
rect 3548 1185 3556 1205
rect 3409 1179 3446 1180
rect 3471 1179 3556 1185
rect 3622 1209 3660 1217
rect 3622 1189 3631 1209
rect 3651 1189 3660 1209
rect 3622 1180 3660 1189
rect 4786 1195 4826 1243
rect 5170 1263 5204 1291
rect 5396 1265 5433 1294
rect 5397 1263 5433 1265
rect 5609 1263 5646 1294
rect 5170 1262 5342 1263
rect 5170 1230 5356 1262
rect 5397 1241 5646 1263
rect 5817 1262 5854 1294
rect 6130 1290 6194 1302
rect 6234 1264 6261 1442
rect 8789 1420 8816 1598
rect 8856 1560 8920 1572
rect 9196 1568 9233 1600
rect 9404 1599 9653 1621
rect 9404 1568 9441 1599
rect 9617 1597 9653 1599
rect 9617 1568 9654 1597
rect 8856 1559 8891 1560
rect 8833 1554 8891 1559
rect 8833 1534 8836 1554
rect 8856 1540 8891 1554
rect 8911 1540 8920 1560
rect 8856 1532 8920 1540
rect 8882 1531 8920 1532
rect 8883 1530 8920 1531
rect 8986 1564 9022 1565
rect 9094 1564 9130 1565
rect 8986 1559 9130 1564
rect 8986 1556 9048 1559
rect 8986 1536 8994 1556
rect 9014 1539 9048 1556
rect 9071 1556 9130 1559
rect 9071 1539 9102 1556
rect 9014 1536 9102 1539
rect 9122 1536 9130 1556
rect 8986 1530 9130 1536
rect 9196 1560 9234 1568
rect 9302 1564 9338 1565
rect 9196 1540 9205 1560
rect 9225 1540 9234 1560
rect 9196 1531 9234 1540
rect 9253 1557 9338 1564
rect 9253 1537 9260 1557
rect 9281 1556 9338 1557
rect 9281 1537 9310 1556
rect 9253 1536 9310 1537
rect 9330 1536 9338 1556
rect 9196 1530 9233 1531
rect 9253 1530 9338 1536
rect 9404 1560 9442 1568
rect 9515 1564 9551 1565
rect 9404 1540 9413 1560
rect 9433 1540 9442 1560
rect 9404 1531 9442 1540
rect 9466 1556 9551 1564
rect 9466 1536 9523 1556
rect 9543 1536 9551 1556
rect 9404 1530 9441 1531
rect 9466 1530 9551 1536
rect 9617 1560 9655 1568
rect 9617 1540 9626 1560
rect 9646 1540 9655 1560
rect 9617 1531 9655 1540
rect 9617 1530 9654 1531
rect 9040 1509 9076 1530
rect 9466 1509 9497 1530
rect 8873 1505 8973 1509
rect 8873 1501 8935 1505
rect 8873 1475 8880 1501
rect 8906 1479 8935 1501
rect 8961 1479 8973 1505
rect 8906 1475 8973 1479
rect 8873 1472 8973 1475
rect 9041 1472 9076 1509
rect 9138 1506 9497 1509
rect 9138 1501 9360 1506
rect 9138 1477 9151 1501
rect 9175 1482 9360 1501
rect 9384 1482 9497 1506
rect 9175 1477 9497 1482
rect 9138 1473 9497 1477
rect 9564 1501 9713 1509
rect 9564 1481 9575 1501
rect 9595 1481 9713 1501
rect 9564 1474 9713 1481
rect 9564 1473 9605 1474
rect 8888 1420 8925 1421
rect 8984 1420 9021 1421
rect 9040 1420 9076 1472
rect 9095 1420 9132 1421
rect 8788 1411 8926 1420
rect 8788 1391 8897 1411
rect 8917 1391 8926 1411
rect 8788 1384 8926 1391
rect 8984 1411 9132 1420
rect 8984 1391 8993 1411
rect 9013 1391 9103 1411
rect 9123 1391 9132 1411
rect 8788 1382 8884 1384
rect 8984 1381 9132 1391
rect 9191 1411 9228 1421
rect 9303 1420 9340 1421
rect 9284 1418 9340 1420
rect 9191 1391 9199 1411
rect 9219 1391 9228 1411
rect 9040 1380 9076 1381
rect 6417 1338 6527 1352
rect 6417 1335 6460 1338
rect 6417 1330 6421 1335
rect 6093 1262 6261 1264
rect 5817 1256 6261 1262
rect 5170 1198 5204 1230
rect 3622 1179 3659 1180
rect 3045 1158 3081 1179
rect 3471 1158 3502 1179
rect 4786 1177 4797 1195
rect 4815 1177 4826 1195
rect 4786 1169 4826 1177
rect 5166 1189 5204 1198
rect 5166 1171 5176 1189
rect 5194 1171 5204 1189
rect 4787 1168 4824 1169
rect 5166 1165 5204 1171
rect 5322 1167 5356 1230
rect 5478 1235 5589 1241
rect 5478 1227 5519 1235
rect 5478 1207 5486 1227
rect 5505 1207 5519 1227
rect 5478 1205 5519 1207
rect 5547 1227 5589 1235
rect 5547 1207 5563 1227
rect 5582 1207 5589 1227
rect 5547 1205 5589 1207
rect 5478 1190 5589 1205
rect 5816 1236 6261 1256
rect 5816 1167 5854 1236
rect 6093 1235 6261 1236
rect 6339 1308 6421 1330
rect 6450 1308 6460 1335
rect 6488 1311 6495 1338
rect 6524 1330 6527 1338
rect 8522 1347 8633 1362
rect 8522 1345 8564 1347
rect 6524 1311 6589 1330
rect 6488 1308 6589 1311
rect 6339 1306 6589 1308
rect 6339 1227 6376 1306
rect 6417 1293 6527 1306
rect 6491 1237 6522 1238
rect 6339 1207 6348 1227
rect 6368 1207 6376 1227
rect 6339 1197 6376 1207
rect 6435 1227 6522 1237
rect 6435 1207 6444 1227
rect 6464 1207 6522 1227
rect 6435 1198 6522 1207
rect 6435 1197 6472 1198
rect 5166 1161 5203 1165
rect 2878 1154 2978 1158
rect 2878 1150 2940 1154
rect 2878 1124 2885 1150
rect 2911 1128 2940 1150
rect 2966 1128 2978 1154
rect 2911 1124 2978 1128
rect 2878 1121 2978 1124
rect 3046 1121 3081 1158
rect 3143 1155 3502 1158
rect 3143 1150 3365 1155
rect 3143 1126 3156 1150
rect 3180 1131 3365 1150
rect 3389 1131 3502 1155
rect 3180 1126 3502 1131
rect 3143 1122 3502 1126
rect 3569 1150 3718 1158
rect 5322 1156 5854 1167
rect 3569 1130 3580 1150
rect 3600 1130 3718 1150
rect 5321 1140 5854 1156
rect 6491 1145 6522 1198
rect 6552 1227 6589 1306
rect 6760 1316 7153 1323
rect 6760 1299 6768 1316
rect 6800 1303 7153 1316
rect 7173 1303 7176 1323
rect 8255 1318 8296 1327
rect 6800 1299 7176 1303
rect 6760 1298 7176 1299
rect 7850 1316 8018 1317
rect 8255 1316 8264 1318
rect 6760 1297 7101 1298
rect 6704 1237 6735 1238
rect 6552 1207 6561 1227
rect 6581 1207 6589 1227
rect 6552 1197 6589 1207
rect 6648 1230 6735 1237
rect 6648 1227 6709 1230
rect 6648 1207 6657 1227
rect 6677 1210 6709 1227
rect 6730 1210 6735 1230
rect 6677 1207 6735 1210
rect 6648 1200 6735 1207
rect 6760 1227 6797 1297
rect 7063 1296 7100 1297
rect 7850 1296 8264 1316
rect 8290 1296 8296 1318
rect 8522 1325 8529 1345
rect 8548 1325 8564 1345
rect 8522 1317 8564 1325
rect 8592 1345 8633 1347
rect 8592 1325 8606 1345
rect 8625 1325 8633 1345
rect 8592 1317 8633 1325
rect 8888 1321 8925 1322
rect 9191 1321 9228 1391
rect 9253 1411 9340 1418
rect 9253 1408 9311 1411
rect 9253 1388 9258 1408
rect 9279 1391 9311 1408
rect 9331 1391 9340 1411
rect 9279 1388 9340 1391
rect 9253 1381 9340 1388
rect 9399 1411 9436 1421
rect 9399 1391 9407 1411
rect 9427 1391 9436 1411
rect 9253 1380 9284 1381
rect 8887 1320 9228 1321
rect 8522 1311 8633 1317
rect 8812 1315 9228 1320
rect 7850 1290 8296 1296
rect 7850 1288 8018 1290
rect 6912 1237 6948 1238
rect 6760 1207 6769 1227
rect 6789 1207 6797 1227
rect 6648 1198 6704 1200
rect 6648 1197 6685 1198
rect 6760 1197 6797 1207
rect 6856 1227 7004 1237
rect 7104 1234 7200 1236
rect 6856 1207 6865 1227
rect 6885 1222 6975 1227
rect 6885 1207 6920 1222
rect 6856 1198 6920 1207
rect 6856 1197 6893 1198
rect 6912 1181 6920 1198
rect 6941 1207 6975 1222
rect 6995 1207 7004 1227
rect 6941 1198 7004 1207
rect 7062 1227 7200 1234
rect 7062 1207 7071 1227
rect 7091 1207 7200 1227
rect 7062 1198 7200 1207
rect 6941 1181 6948 1198
rect 6967 1197 7004 1198
rect 7063 1197 7100 1198
rect 6912 1146 6948 1181
rect 6383 1144 6424 1145
rect 5321 1139 5835 1140
rect 3569 1123 3718 1130
rect 6275 1137 6424 1144
rect 4158 1127 4672 1128
rect 3569 1122 3610 1123
rect 2893 1069 2930 1070
rect 2989 1069 3026 1070
rect 3045 1069 3081 1121
rect 3100 1069 3137 1070
rect 2793 1060 2931 1069
rect 2793 1040 2902 1060
rect 2922 1040 2931 1060
rect 2793 1033 2931 1040
rect 2989 1060 3137 1069
rect 2989 1040 2998 1060
rect 3018 1040 3108 1060
rect 3128 1040 3137 1060
rect 2793 1031 2889 1033
rect 2989 1030 3137 1040
rect 3196 1060 3233 1070
rect 3308 1069 3345 1070
rect 3289 1067 3345 1069
rect 3196 1040 3204 1060
rect 3224 1040 3233 1060
rect 3045 1029 3081 1030
rect 1975 977 2143 979
rect 1697 971 2143 977
rect 765 947 1181 952
rect 1360 950 1471 956
rect 765 946 1106 947
rect 709 886 740 887
rect 557 856 566 876
rect 586 856 594 876
rect 557 846 594 856
rect 653 879 740 886
rect 653 876 714 879
rect 653 856 662 876
rect 682 859 714 876
rect 735 859 740 879
rect 682 856 740 859
rect 653 849 740 856
rect 765 876 802 946
rect 1068 945 1105 946
rect 1360 942 1401 950
rect 1360 922 1368 942
rect 1387 922 1401 942
rect 1360 920 1401 922
rect 1429 942 1471 950
rect 1429 922 1445 942
rect 1464 922 1471 942
rect 1697 949 1703 971
rect 1729 951 2143 971
rect 2893 970 2930 971
rect 3196 970 3233 1040
rect 3258 1060 3345 1067
rect 3258 1057 3316 1060
rect 3258 1037 3263 1057
rect 3284 1040 3316 1057
rect 3336 1040 3345 1060
rect 3284 1037 3345 1040
rect 3258 1030 3345 1037
rect 3404 1060 3441 1070
rect 3404 1040 3412 1060
rect 3432 1040 3441 1060
rect 3258 1029 3289 1030
rect 2892 969 3233 970
rect 1729 949 1738 951
rect 1975 950 2143 951
rect 2817 964 3233 969
rect 1697 940 1738 949
rect 2817 944 2820 964
rect 2840 944 3233 964
rect 3404 961 3441 1040
rect 3471 1069 3502 1122
rect 4139 1111 4672 1127
rect 6275 1117 6393 1137
rect 6413 1117 6424 1137
rect 4139 1100 4671 1111
rect 6275 1109 6424 1117
rect 6491 1141 6850 1145
rect 6491 1136 6813 1141
rect 6491 1112 6604 1136
rect 6628 1117 6813 1136
rect 6837 1117 6850 1141
rect 6628 1112 6850 1117
rect 6491 1109 6850 1112
rect 6912 1109 6947 1146
rect 7015 1143 7115 1146
rect 7015 1139 7082 1143
rect 7015 1113 7027 1139
rect 7053 1117 7082 1139
rect 7108 1117 7115 1143
rect 7053 1113 7115 1117
rect 7015 1109 7115 1113
rect 4790 1102 4827 1106
rect 3521 1069 3558 1070
rect 3471 1060 3558 1069
rect 3471 1040 3529 1060
rect 3549 1040 3558 1060
rect 3471 1030 3558 1040
rect 3617 1060 3654 1070
rect 3617 1040 3625 1060
rect 3645 1040 3654 1060
rect 3471 1029 3502 1030
rect 3466 961 3576 974
rect 3617 961 3654 1040
rect 3404 959 3654 961
rect 3404 956 3505 959
rect 3404 937 3469 956
rect 1429 920 1471 922
rect 1360 905 1471 920
rect 3466 929 3469 937
rect 3498 929 3505 956
rect 3533 932 3543 959
rect 3572 937 3654 959
rect 3732 1031 3900 1032
rect 4139 1031 4177 1100
rect 3732 1011 4177 1031
rect 4404 1062 4515 1077
rect 4404 1060 4446 1062
rect 4404 1040 4411 1060
rect 4430 1040 4446 1060
rect 4404 1032 4446 1040
rect 4474 1060 4515 1062
rect 4474 1040 4488 1060
rect 4507 1040 4515 1060
rect 4474 1032 4515 1040
rect 4404 1026 4515 1032
rect 4637 1037 4671 1100
rect 4789 1096 4827 1102
rect 5169 1098 5206 1099
rect 4789 1078 4799 1096
rect 4817 1078 4827 1096
rect 4789 1069 4827 1078
rect 5167 1090 5207 1098
rect 5167 1072 5178 1090
rect 5196 1072 5207 1090
rect 6491 1088 6522 1109
rect 6912 1088 6948 1109
rect 6334 1087 6371 1088
rect 4789 1037 4823 1069
rect 3732 1005 4176 1011
rect 3732 1003 3900 1005
rect 3572 932 3576 937
rect 3533 929 3576 932
rect 3466 915 3576 929
rect 917 886 953 887
rect 765 856 774 876
rect 794 856 802 876
rect 653 847 709 849
rect 653 846 690 847
rect 765 846 802 856
rect 861 876 1009 886
rect 1109 883 1205 885
rect 861 856 870 876
rect 890 856 980 876
rect 1000 856 1009 876
rect 861 847 1009 856
rect 1067 876 1205 883
rect 1067 856 1076 876
rect 1096 856 1205 876
rect 1067 847 1205 856
rect 861 846 898 847
rect 917 795 953 847
rect 972 846 1009 847
rect 1068 846 1105 847
rect 388 793 429 794
rect 280 786 429 793
rect 280 766 398 786
rect 418 766 429 786
rect 280 758 429 766
rect 496 790 855 794
rect 496 785 818 790
rect 496 761 609 785
rect 633 766 818 785
rect 842 766 855 790
rect 633 761 855 766
rect 496 758 855 761
rect 917 758 952 795
rect 1020 792 1120 795
rect 1020 788 1087 792
rect 1020 762 1032 788
rect 1058 766 1087 788
rect 1113 766 1120 792
rect 1058 762 1120 766
rect 1020 758 1120 762
rect 496 737 527 758
rect 917 737 953 758
rect 339 736 376 737
rect 338 727 376 736
rect 338 707 347 727
rect 367 707 376 727
rect 338 699 376 707
rect 442 731 527 737
rect 552 736 589 737
rect 442 711 450 731
rect 470 711 527 731
rect 442 703 527 711
rect 551 727 589 736
rect 551 707 560 727
rect 580 707 589 727
rect 442 702 478 703
rect 551 699 589 707
rect 655 731 740 737
rect 760 736 797 737
rect 655 711 663 731
rect 683 730 740 731
rect 683 711 712 730
rect 655 710 712 711
rect 733 710 740 730
rect 655 703 740 710
rect 759 727 797 736
rect 759 707 768 727
rect 788 707 797 727
rect 655 702 691 703
rect 759 699 797 707
rect 863 731 1007 737
rect 863 711 871 731
rect 891 728 979 731
rect 891 711 922 728
rect 863 708 922 711
rect 945 711 979 728
rect 999 711 1007 731
rect 945 708 1007 711
rect 863 703 1007 708
rect 863 702 899 703
rect 971 702 1007 703
rect 1073 736 1110 737
rect 1073 735 1111 736
rect 1073 727 1137 735
rect 1073 707 1082 727
rect 1102 713 1137 727
rect 1157 713 1160 733
rect 1102 708 1160 713
rect 1102 707 1137 708
rect 339 670 376 699
rect 340 668 376 670
rect 552 668 589 699
rect 340 646 589 668
rect 760 667 797 699
rect 1073 695 1137 707
rect 1177 669 1204 847
rect 3732 825 3759 1003
rect 3799 965 3863 977
rect 4139 973 4176 1005
rect 4347 1004 4596 1026
rect 4637 1005 4823 1037
rect 4651 1004 4823 1005
rect 4347 973 4384 1004
rect 4560 1002 4596 1004
rect 4560 973 4597 1002
rect 4789 976 4823 1004
rect 5167 1024 5207 1072
rect 6333 1078 6371 1087
rect 6333 1058 6342 1078
rect 6362 1058 6371 1078
rect 6333 1050 6371 1058
rect 6437 1082 6522 1088
rect 6547 1087 6584 1088
rect 6437 1062 6445 1082
rect 6465 1062 6522 1082
rect 6437 1054 6522 1062
rect 6546 1078 6584 1087
rect 6546 1058 6555 1078
rect 6575 1058 6584 1078
rect 6437 1053 6473 1054
rect 6546 1050 6584 1058
rect 6650 1082 6735 1088
rect 6755 1087 6792 1088
rect 6650 1062 6658 1082
rect 6678 1081 6735 1082
rect 6678 1062 6707 1081
rect 6650 1061 6707 1062
rect 6728 1061 6735 1081
rect 6650 1054 6735 1061
rect 6754 1078 6792 1087
rect 6754 1058 6763 1078
rect 6783 1058 6792 1078
rect 6650 1053 6686 1054
rect 6754 1050 6792 1058
rect 6858 1082 7002 1088
rect 6858 1062 6866 1082
rect 6886 1062 6974 1082
rect 6994 1062 7002 1082
rect 6858 1054 7002 1062
rect 6858 1053 6894 1054
rect 6966 1053 7002 1054
rect 7068 1087 7105 1088
rect 7068 1086 7106 1087
rect 7068 1078 7132 1086
rect 7068 1058 7077 1078
rect 7097 1064 7132 1078
rect 7152 1064 7155 1084
rect 7097 1059 7155 1064
rect 7097 1058 7132 1059
rect 5478 1028 5588 1042
rect 5478 1025 5521 1028
rect 5167 1017 5292 1024
rect 5478 1020 5482 1025
rect 5167 998 5259 1017
rect 5284 998 5292 1017
rect 5167 988 5292 998
rect 5400 998 5482 1020
rect 5511 998 5521 1025
rect 5549 1001 5556 1028
rect 5585 1020 5588 1028
rect 6334 1021 6371 1050
rect 5585 1001 5650 1020
rect 6335 1019 6371 1021
rect 6547 1019 6584 1050
rect 6755 1023 6792 1050
rect 7068 1046 7132 1058
rect 5549 998 5650 1001
rect 5400 996 5650 998
rect 3799 964 3834 965
rect 3776 959 3834 964
rect 3776 939 3779 959
rect 3799 945 3834 959
rect 3854 945 3863 965
rect 3799 937 3863 945
rect 3825 936 3863 937
rect 3826 935 3863 936
rect 3929 969 3965 970
rect 4037 969 4073 970
rect 3929 962 4073 969
rect 3929 961 3989 962
rect 3929 941 3937 961
rect 3957 942 3989 961
rect 4014 961 4073 962
rect 4014 942 4045 961
rect 3957 941 4045 942
rect 4065 941 4073 961
rect 3929 935 4073 941
rect 4139 965 4177 973
rect 4245 969 4281 970
rect 4139 945 4148 965
rect 4168 945 4177 965
rect 4139 936 4177 945
rect 4196 962 4281 969
rect 4196 942 4203 962
rect 4224 961 4281 962
rect 4224 942 4253 961
rect 4196 941 4253 942
rect 4273 941 4281 961
rect 4139 935 4176 936
rect 4196 935 4281 941
rect 4347 965 4385 973
rect 4458 969 4494 970
rect 4347 945 4356 965
rect 4376 945 4385 965
rect 4347 936 4385 945
rect 4409 961 4494 969
rect 4409 941 4466 961
rect 4486 941 4494 961
rect 4347 935 4384 936
rect 4409 935 4494 941
rect 4560 965 4598 973
rect 4560 945 4569 965
rect 4589 945 4598 965
rect 4560 936 4598 945
rect 4787 966 4824 976
rect 5167 968 5207 988
rect 4787 948 4797 966
rect 4815 948 4824 966
rect 4787 939 4824 948
rect 5166 959 5207 968
rect 5166 941 5176 959
rect 5194 941 5207 959
rect 4789 938 4823 939
rect 4560 935 4597 936
rect 3983 914 4019 935
rect 4409 914 4440 935
rect 5166 932 5207 941
rect 5166 931 5203 932
rect 5400 917 5437 996
rect 5478 983 5588 996
rect 5552 927 5583 928
rect 3816 910 3916 914
rect 3816 906 3878 910
rect 3816 880 3823 906
rect 3849 884 3878 906
rect 3904 884 3916 910
rect 3849 880 3916 884
rect 3816 877 3916 880
rect 3984 877 4019 914
rect 4081 911 4440 914
rect 4081 906 4303 911
rect 4081 882 4094 906
rect 4118 887 4303 906
rect 4327 887 4440 911
rect 4118 882 4440 887
rect 4081 878 4440 882
rect 4507 906 4656 914
rect 4507 886 4518 906
rect 4538 886 4656 906
rect 5400 897 5409 917
rect 5429 897 5437 917
rect 5400 887 5437 897
rect 5496 917 5583 927
rect 5496 897 5505 917
rect 5525 897 5583 917
rect 5496 888 5583 897
rect 5496 887 5533 888
rect 4507 879 4656 886
rect 4507 878 4548 879
rect 3831 825 3868 826
rect 3927 825 3964 826
rect 3983 825 4019 877
rect 4038 825 4075 826
rect 3731 816 3869 825
rect 3731 796 3840 816
rect 3860 796 3869 816
rect 3731 789 3869 796
rect 3927 816 4075 825
rect 3927 796 3936 816
rect 3956 796 4046 816
rect 4066 796 4075 816
rect 3731 787 3827 789
rect 3927 786 4075 796
rect 4134 816 4171 826
rect 4246 825 4283 826
rect 4227 823 4283 825
rect 4134 796 4142 816
rect 4162 796 4171 816
rect 3983 785 4019 786
rect 3831 726 3868 727
rect 4134 726 4171 796
rect 4196 816 4283 823
rect 4196 813 4254 816
rect 4196 793 4201 813
rect 4222 796 4254 813
rect 4274 796 4283 816
rect 4222 793 4283 796
rect 4196 786 4283 793
rect 4342 816 4379 826
rect 4342 796 4350 816
rect 4370 796 4379 816
rect 4196 785 4227 786
rect 3830 725 4171 726
rect 3755 720 4171 725
rect 3755 700 3758 720
rect 3778 700 4171 720
rect 4342 717 4379 796
rect 4409 825 4440 878
rect 4790 876 4827 877
rect 4789 867 4828 876
rect 4789 849 4799 867
rect 4817 849 4828 867
rect 5169 865 5206 869
rect 4701 832 4748 833
rect 4789 832 4828 849
rect 4701 828 4828 832
rect 4459 825 4496 826
rect 4409 816 4496 825
rect 4409 796 4467 816
rect 4487 796 4496 816
rect 4409 786 4496 796
rect 4555 816 4592 826
rect 4555 796 4563 816
rect 4583 796 4592 816
rect 4409 785 4440 786
rect 4404 717 4514 730
rect 4555 717 4592 796
rect 4701 799 4711 828
rect 4740 799 4828 828
rect 4701 793 4828 799
rect 4701 789 4748 793
rect 4786 779 4828 793
rect 4786 761 4797 779
rect 4815 761 4828 779
rect 4786 756 4828 761
rect 4787 753 4828 756
rect 5166 860 5206 865
rect 5166 842 5178 860
rect 5196 842 5206 860
rect 4787 752 4824 753
rect 4342 715 4592 717
rect 4342 712 4443 715
rect 4342 693 4407 712
rect 4404 685 4407 693
rect 4436 685 4443 712
rect 4471 688 4481 715
rect 4510 693 4592 715
rect 4510 688 4514 693
rect 4471 685 4514 688
rect 4404 671 4514 685
rect 4780 689 4827 690
rect 4780 680 4828 689
rect 1036 667 1204 669
rect 760 664 1204 667
rect 421 640 532 646
rect 421 632 462 640
rect 110 577 149 621
rect 421 612 429 632
rect 448 612 462 632
rect 421 610 462 612
rect 490 634 532 640
rect 758 641 1204 664
rect 4780 662 4799 680
rect 4817 662 4828 680
rect 4780 660 4828 662
rect 4789 641 4828 660
rect 5166 662 5206 842
rect 5552 835 5583 888
rect 5613 917 5650 996
rect 5821 993 6214 1013
rect 6234 993 6237 1013
rect 6335 997 6584 1019
rect 6753 1018 6794 1023
rect 7172 1020 7199 1198
rect 7850 1110 7877 1288
rect 8255 1285 8296 1290
rect 8465 1289 8714 1311
rect 8812 1295 8815 1315
rect 8835 1295 9228 1315
rect 9399 1312 9436 1391
rect 9466 1420 9497 1473
rect 9843 1466 9883 1646
rect 9843 1448 9853 1466
rect 9871 1448 9883 1466
rect 9843 1443 9883 1448
rect 9843 1439 9880 1443
rect 9516 1420 9553 1421
rect 9466 1411 9553 1420
rect 9466 1391 9524 1411
rect 9544 1391 9553 1411
rect 9466 1381 9553 1391
rect 9612 1411 9649 1421
rect 9612 1391 9620 1411
rect 9640 1391 9649 1411
rect 9466 1380 9497 1381
rect 9461 1312 9571 1325
rect 9612 1312 9649 1391
rect 9846 1376 9883 1377
rect 9842 1367 9883 1376
rect 9842 1349 9855 1367
rect 9873 1349 9883 1367
rect 9842 1340 9883 1349
rect 9842 1320 9882 1340
rect 9399 1310 9649 1312
rect 9399 1307 9500 1310
rect 7917 1250 7981 1262
rect 8257 1258 8294 1285
rect 8465 1258 8502 1289
rect 8678 1287 8714 1289
rect 9399 1288 9464 1307
rect 8678 1258 8715 1287
rect 9461 1280 9464 1288
rect 9493 1280 9500 1307
rect 9528 1283 9538 1310
rect 9567 1288 9649 1310
rect 9757 1310 9882 1320
rect 9757 1291 9765 1310
rect 9790 1291 9882 1310
rect 9567 1283 9571 1288
rect 9757 1284 9882 1291
rect 9528 1280 9571 1283
rect 9461 1266 9571 1280
rect 7917 1249 7952 1250
rect 7894 1244 7952 1249
rect 7894 1224 7897 1244
rect 7917 1230 7952 1244
rect 7972 1230 7981 1250
rect 7917 1222 7981 1230
rect 7943 1221 7981 1222
rect 7944 1220 7981 1221
rect 8047 1254 8083 1255
rect 8155 1254 8191 1255
rect 8047 1246 8191 1254
rect 8047 1226 8055 1246
rect 8075 1243 8163 1246
rect 8075 1226 8107 1243
rect 8127 1226 8163 1243
rect 8183 1226 8191 1246
rect 8047 1220 8191 1226
rect 8257 1250 8295 1258
rect 8363 1254 8399 1255
rect 8257 1230 8266 1250
rect 8286 1230 8295 1250
rect 8257 1221 8295 1230
rect 8314 1247 8399 1254
rect 8314 1227 8321 1247
rect 8342 1246 8399 1247
rect 8342 1227 8371 1246
rect 8314 1226 8371 1227
rect 8391 1226 8399 1246
rect 8257 1220 8294 1221
rect 8314 1220 8399 1226
rect 8465 1250 8503 1258
rect 8576 1254 8612 1255
rect 8465 1230 8474 1250
rect 8494 1230 8503 1250
rect 8465 1221 8503 1230
rect 8527 1246 8612 1254
rect 8527 1226 8584 1246
rect 8604 1226 8612 1246
rect 8465 1220 8502 1221
rect 8527 1220 8612 1226
rect 8678 1250 8716 1258
rect 8678 1230 8687 1250
rect 8707 1230 8716 1250
rect 8678 1221 8716 1230
rect 9842 1236 9882 1284
rect 8678 1220 8715 1221
rect 8101 1199 8137 1220
rect 8527 1199 8558 1220
rect 9842 1218 9853 1236
rect 9871 1218 9882 1236
rect 9842 1210 9882 1218
rect 9843 1209 9880 1210
rect 7934 1195 8034 1199
rect 7934 1191 7996 1195
rect 7934 1165 7941 1191
rect 7967 1169 7996 1191
rect 8022 1169 8034 1195
rect 7967 1165 8034 1169
rect 7934 1162 8034 1165
rect 8102 1162 8137 1199
rect 8199 1196 8558 1199
rect 8199 1191 8421 1196
rect 8199 1167 8212 1191
rect 8236 1172 8421 1191
rect 8445 1172 8558 1196
rect 8236 1167 8558 1172
rect 8199 1163 8558 1167
rect 8625 1191 8774 1199
rect 8625 1171 8636 1191
rect 8656 1171 8774 1191
rect 8625 1164 8774 1171
rect 9214 1168 9728 1169
rect 8625 1163 8666 1164
rect 7949 1110 7986 1111
rect 8045 1110 8082 1111
rect 8101 1110 8137 1162
rect 8156 1110 8193 1111
rect 7849 1101 7987 1110
rect 7849 1081 7958 1101
rect 7978 1081 7987 1101
rect 7849 1074 7987 1081
rect 8045 1101 8193 1110
rect 8045 1081 8054 1101
rect 8074 1081 8164 1101
rect 8184 1081 8193 1101
rect 7849 1072 7945 1074
rect 8045 1071 8193 1081
rect 8252 1101 8289 1111
rect 8364 1110 8401 1111
rect 8345 1108 8401 1110
rect 8252 1081 8260 1101
rect 8280 1081 8289 1101
rect 8101 1070 8137 1071
rect 7031 1018 7199 1020
rect 6753 1012 7199 1018
rect 5821 988 6237 993
rect 6416 991 6527 997
rect 5821 987 6162 988
rect 5765 927 5796 928
rect 5613 897 5622 917
rect 5642 897 5650 917
rect 5613 887 5650 897
rect 5709 920 5796 927
rect 5709 917 5770 920
rect 5709 897 5718 917
rect 5738 900 5770 917
rect 5791 900 5796 920
rect 5738 897 5796 900
rect 5709 890 5796 897
rect 5821 917 5858 987
rect 6124 986 6161 987
rect 6416 983 6457 991
rect 6416 963 6424 983
rect 6443 963 6457 983
rect 6416 961 6457 963
rect 6485 983 6527 991
rect 6485 963 6501 983
rect 6520 963 6527 983
rect 6753 990 6759 1012
rect 6785 992 7199 1012
rect 7949 1011 7986 1012
rect 8252 1011 8289 1081
rect 8314 1101 8401 1108
rect 8314 1098 8372 1101
rect 8314 1078 8319 1098
rect 8340 1081 8372 1098
rect 8392 1081 8401 1101
rect 8340 1078 8401 1081
rect 8314 1071 8401 1078
rect 8460 1101 8497 1111
rect 8460 1081 8468 1101
rect 8488 1081 8497 1101
rect 8314 1070 8345 1071
rect 7948 1010 8289 1011
rect 6785 990 6794 992
rect 7031 991 7199 992
rect 7873 1005 8289 1010
rect 6753 981 6794 990
rect 7873 985 7876 1005
rect 7896 985 8289 1005
rect 8460 1002 8497 1081
rect 8527 1110 8558 1163
rect 9195 1152 9728 1168
rect 9195 1141 9727 1152
rect 9846 1143 9883 1147
rect 8577 1110 8614 1111
rect 8527 1101 8614 1110
rect 8527 1081 8585 1101
rect 8605 1081 8614 1101
rect 8527 1071 8614 1081
rect 8673 1101 8710 1111
rect 8673 1081 8681 1101
rect 8701 1081 8710 1101
rect 8527 1070 8558 1071
rect 8522 1002 8632 1015
rect 8673 1002 8710 1081
rect 8460 1000 8710 1002
rect 8460 997 8561 1000
rect 8460 978 8525 997
rect 6485 961 6527 963
rect 6416 946 6527 961
rect 8522 970 8525 978
rect 8554 970 8561 997
rect 8589 973 8599 1000
rect 8628 978 8710 1000
rect 8788 1072 8956 1073
rect 9195 1072 9233 1141
rect 8788 1052 9233 1072
rect 9460 1103 9571 1118
rect 9460 1101 9502 1103
rect 9460 1081 9467 1101
rect 9486 1081 9502 1101
rect 9460 1073 9502 1081
rect 9530 1101 9571 1103
rect 9530 1081 9544 1101
rect 9563 1081 9571 1101
rect 9530 1073 9571 1081
rect 9460 1067 9571 1073
rect 9693 1078 9727 1141
rect 9845 1137 9883 1143
rect 9845 1119 9855 1137
rect 9873 1119 9883 1137
rect 9845 1110 9883 1119
rect 9845 1078 9879 1110
rect 8788 1046 9232 1052
rect 8788 1044 8956 1046
rect 8628 973 8632 978
rect 8589 970 8632 973
rect 8522 956 8632 970
rect 5973 927 6009 928
rect 5821 897 5830 917
rect 5850 897 5858 917
rect 5709 888 5765 890
rect 5709 887 5746 888
rect 5821 887 5858 897
rect 5917 917 6065 927
rect 6165 924 6261 926
rect 5917 897 5926 917
rect 5946 897 6036 917
rect 6056 897 6065 917
rect 5917 888 6065 897
rect 6123 917 6261 924
rect 6123 897 6132 917
rect 6152 897 6261 917
rect 6123 888 6261 897
rect 5917 887 5954 888
rect 5973 836 6009 888
rect 6028 887 6065 888
rect 6124 887 6161 888
rect 5444 834 5485 835
rect 5336 827 5485 834
rect 5336 807 5454 827
rect 5474 807 5485 827
rect 5336 799 5485 807
rect 5552 831 5911 835
rect 5552 826 5874 831
rect 5552 802 5665 826
rect 5689 807 5874 826
rect 5898 807 5911 831
rect 5689 802 5911 807
rect 5552 799 5911 802
rect 5973 799 6008 836
rect 6076 833 6176 836
rect 6076 829 6143 833
rect 6076 803 6088 829
rect 6114 807 6143 829
rect 6169 807 6176 833
rect 6114 803 6176 807
rect 6076 799 6176 803
rect 5552 778 5583 799
rect 5973 778 6009 799
rect 5395 777 5432 778
rect 5394 768 5432 777
rect 5394 748 5403 768
rect 5423 748 5432 768
rect 5394 740 5432 748
rect 5498 772 5583 778
rect 5608 777 5645 778
rect 5498 752 5506 772
rect 5526 752 5583 772
rect 5498 744 5583 752
rect 5607 768 5645 777
rect 5607 748 5616 768
rect 5636 748 5645 768
rect 5498 743 5534 744
rect 5607 740 5645 748
rect 5711 772 5796 778
rect 5816 777 5853 778
rect 5711 752 5719 772
rect 5739 771 5796 772
rect 5739 752 5768 771
rect 5711 751 5768 752
rect 5789 751 5796 771
rect 5711 744 5796 751
rect 5815 768 5853 777
rect 5815 748 5824 768
rect 5844 748 5853 768
rect 5711 743 5747 744
rect 5815 740 5853 748
rect 5919 772 6063 778
rect 5919 752 5927 772
rect 5947 769 6035 772
rect 5947 752 5978 769
rect 5919 749 5978 752
rect 6001 752 6035 769
rect 6055 752 6063 772
rect 6001 749 6063 752
rect 5919 744 6063 749
rect 5919 743 5955 744
rect 6027 743 6063 744
rect 6129 777 6166 778
rect 6129 776 6167 777
rect 6129 768 6193 776
rect 6129 748 6138 768
rect 6158 754 6193 768
rect 6213 754 6216 774
rect 6158 749 6216 754
rect 6158 748 6193 749
rect 5395 711 5432 740
rect 5396 709 5432 711
rect 5608 709 5645 740
rect 5396 687 5645 709
rect 5816 708 5853 740
rect 6129 736 6193 748
rect 6233 710 6260 888
rect 8788 866 8815 1044
rect 8855 1006 8919 1018
rect 9195 1014 9232 1046
rect 9403 1045 9652 1067
rect 9693 1046 9879 1078
rect 9707 1045 9879 1046
rect 9403 1014 9440 1045
rect 9616 1043 9652 1045
rect 9616 1014 9653 1043
rect 9845 1017 9879 1045
rect 8855 1005 8890 1006
rect 8832 1000 8890 1005
rect 8832 980 8835 1000
rect 8855 986 8890 1000
rect 8910 986 8919 1006
rect 8855 978 8919 986
rect 8881 977 8919 978
rect 8882 976 8919 977
rect 8985 1010 9021 1011
rect 9093 1010 9129 1011
rect 8985 1003 9129 1010
rect 8985 1002 9045 1003
rect 8985 982 8993 1002
rect 9013 983 9045 1002
rect 9070 1002 9129 1003
rect 9070 983 9101 1002
rect 9013 982 9101 983
rect 9121 982 9129 1002
rect 8985 976 9129 982
rect 9195 1006 9233 1014
rect 9301 1010 9337 1011
rect 9195 986 9204 1006
rect 9224 986 9233 1006
rect 9195 977 9233 986
rect 9252 1003 9337 1010
rect 9252 983 9259 1003
rect 9280 1002 9337 1003
rect 9280 983 9309 1002
rect 9252 982 9309 983
rect 9329 982 9337 1002
rect 9195 976 9232 977
rect 9252 976 9337 982
rect 9403 1006 9441 1014
rect 9514 1010 9550 1011
rect 9403 986 9412 1006
rect 9432 986 9441 1006
rect 9403 977 9441 986
rect 9465 1002 9550 1010
rect 9465 982 9522 1002
rect 9542 982 9550 1002
rect 9403 976 9440 977
rect 9465 976 9550 982
rect 9616 1006 9654 1014
rect 9616 986 9625 1006
rect 9645 986 9654 1006
rect 9616 977 9654 986
rect 9843 1007 9880 1017
rect 9843 989 9853 1007
rect 9871 989 9880 1007
rect 9843 980 9880 989
rect 9845 979 9879 980
rect 9616 976 9653 977
rect 9039 955 9075 976
rect 9465 955 9496 976
rect 8872 951 8972 955
rect 8872 947 8934 951
rect 8872 921 8879 947
rect 8905 925 8934 947
rect 8960 925 8972 951
rect 8905 921 8972 925
rect 8872 918 8972 921
rect 9040 918 9075 955
rect 9137 952 9496 955
rect 9137 947 9359 952
rect 9137 923 9150 947
rect 9174 928 9359 947
rect 9383 928 9496 952
rect 9174 923 9496 928
rect 9137 919 9496 923
rect 9563 947 9712 955
rect 9563 927 9574 947
rect 9594 927 9712 947
rect 9563 920 9712 927
rect 9563 919 9604 920
rect 8887 866 8924 867
rect 8983 866 9020 867
rect 9039 866 9075 918
rect 9094 866 9131 867
rect 8787 857 8925 866
rect 8787 837 8896 857
rect 8916 837 8925 857
rect 8787 830 8925 837
rect 8983 857 9131 866
rect 8983 837 8992 857
rect 9012 837 9102 857
rect 9122 837 9131 857
rect 8787 828 8883 830
rect 8983 827 9131 837
rect 9190 857 9227 867
rect 9302 866 9339 867
rect 9283 864 9339 866
rect 9190 837 9198 857
rect 9218 837 9227 857
rect 9039 826 9075 827
rect 8887 767 8924 768
rect 9190 767 9227 837
rect 9252 857 9339 864
rect 9252 854 9310 857
rect 9252 834 9257 854
rect 9278 837 9310 854
rect 9330 837 9339 857
rect 9278 834 9339 837
rect 9252 827 9339 834
rect 9398 857 9435 867
rect 9398 837 9406 857
rect 9426 837 9435 857
rect 9252 826 9283 827
rect 8886 766 9227 767
rect 8811 761 9227 766
rect 8811 741 8814 761
rect 8834 741 9227 761
rect 9398 758 9435 837
rect 9465 866 9496 919
rect 9846 917 9883 918
rect 9845 908 9884 917
rect 9845 890 9855 908
rect 9873 890 9884 908
rect 9757 873 9804 874
rect 9845 873 9884 890
rect 9757 869 9884 873
rect 9515 866 9552 867
rect 9465 857 9552 866
rect 9465 837 9523 857
rect 9543 837 9552 857
rect 9465 827 9552 837
rect 9611 857 9648 867
rect 9611 837 9619 857
rect 9639 837 9648 857
rect 9465 826 9496 827
rect 9460 758 9570 771
rect 9611 758 9648 837
rect 9757 840 9767 869
rect 9796 840 9884 869
rect 9757 834 9884 840
rect 9757 830 9804 834
rect 9842 820 9884 834
rect 9842 802 9853 820
rect 9871 802 9884 820
rect 9842 797 9884 802
rect 9843 794 9884 797
rect 9843 793 9880 794
rect 9398 756 9648 758
rect 9398 753 9499 756
rect 9398 734 9463 753
rect 9460 726 9463 734
rect 9492 726 9499 753
rect 9527 729 9537 756
rect 9566 734 9648 756
rect 9566 729 9570 734
rect 9527 726 9570 729
rect 9460 712 9570 726
rect 9836 730 9883 731
rect 9836 721 9884 730
rect 6092 708 6260 710
rect 5816 705 6260 708
rect 5477 681 5588 687
rect 5477 673 5518 681
rect 490 632 531 634
rect 490 612 506 632
rect 525 612 531 632
rect 490 610 531 612
rect 421 595 531 610
rect 110 553 150 577
rect 758 567 796 641
rect 1036 640 1204 641
rect 718 553 797 567
rect 110 552 400 553
rect 566 552 797 553
rect 110 550 797 552
rect 110 529 757 550
rect 786 529 797 550
rect 110 520 797 529
rect 4787 554 4831 641
rect 5166 618 5205 662
rect 5477 653 5485 673
rect 5504 653 5518 673
rect 5477 651 5518 653
rect 5546 675 5588 681
rect 5814 682 6260 705
rect 9836 703 9855 721
rect 9873 703 9884 721
rect 9836 701 9884 703
rect 9845 682 9884 701
rect 5546 673 5587 675
rect 5546 653 5562 673
rect 5581 653 5587 673
rect 5546 651 5587 653
rect 5477 636 5587 651
rect 5166 594 5206 618
rect 5814 608 5852 682
rect 6092 681 6260 682
rect 5774 594 5853 608
rect 5166 593 5456 594
rect 5622 593 5853 594
rect 5166 591 5853 593
rect 5166 570 5813 591
rect 5842 570 5853 591
rect 5166 561 5853 570
rect 9843 595 9887 682
rect 9843 574 9848 595
rect 9877 574 9887 595
rect 9843 561 9887 574
rect 4787 533 4792 554
rect 4821 533 4831 554
rect 5774 551 5853 561
rect 4787 520 4831 533
rect 718 510 797 520
rect 6725 469 6835 483
rect 6725 466 6768 469
rect 6725 461 6729 466
rect 1669 428 1779 442
rect 1669 425 1712 428
rect 1669 420 1673 425
rect 1591 398 1673 420
rect 1702 398 1712 425
rect 1740 401 1747 428
rect 1776 420 1779 428
rect 6647 439 6729 461
rect 6758 439 6768 466
rect 6796 442 6803 469
rect 6832 461 6835 469
rect 6832 442 6897 461
rect 6796 439 6897 442
rect 6647 437 6897 439
rect 1776 401 1841 420
rect 1740 398 1841 401
rect 1591 396 1841 398
rect 1591 317 1628 396
rect 1669 383 1779 396
rect 1743 327 1774 328
rect 1591 297 1600 317
rect 1620 297 1628 317
rect 1591 287 1628 297
rect 1687 317 1774 327
rect 1687 297 1696 317
rect 1716 297 1774 317
rect 1687 288 1774 297
rect 1687 287 1724 288
rect 1743 235 1774 288
rect 1804 317 1841 396
rect 2012 393 2405 413
rect 2425 393 2428 413
rect 4619 408 4729 422
rect 4619 405 4662 408
rect 4619 400 4623 405
rect 2012 388 2428 393
rect 2012 387 2353 388
rect 1956 327 1987 328
rect 1804 297 1813 317
rect 1833 297 1841 317
rect 1804 287 1841 297
rect 1900 320 1987 327
rect 1900 317 1961 320
rect 1900 297 1909 317
rect 1929 300 1961 317
rect 1982 300 1987 320
rect 1929 297 1987 300
rect 1900 290 1987 297
rect 2012 317 2049 387
rect 2315 386 2352 387
rect 4541 378 4623 400
rect 4652 378 4662 405
rect 4690 381 4697 408
rect 4726 400 4729 408
rect 4726 381 4791 400
rect 4690 378 4791 381
rect 4541 376 4791 378
rect 2164 327 2200 328
rect 2012 297 2021 317
rect 2041 297 2049 317
rect 1900 288 1956 290
rect 1900 287 1937 288
rect 2012 287 2049 297
rect 2108 317 2256 327
rect 2356 324 2452 326
rect 2108 297 2117 317
rect 2137 297 2227 317
rect 2247 297 2256 317
rect 2108 288 2256 297
rect 2314 317 2452 324
rect 2314 297 2323 317
rect 2343 297 2452 317
rect 2314 288 2452 297
rect 4541 297 4578 376
rect 4619 363 4729 376
rect 4693 307 4724 308
rect 2108 287 2145 288
rect 2164 236 2200 288
rect 2219 287 2256 288
rect 2315 287 2352 288
rect 1635 234 1676 235
rect 1527 227 1676 234
rect 1527 207 1645 227
rect 1665 207 1676 227
rect 1527 199 1676 207
rect 1743 231 2102 235
rect 1743 226 2065 231
rect 1743 202 1856 226
rect 1880 207 2065 226
rect 2089 207 2102 231
rect 1880 202 2102 207
rect 1743 199 2102 202
rect 2164 199 2199 236
rect 2267 233 2367 236
rect 2267 229 2334 233
rect 2267 203 2279 229
rect 2305 207 2334 229
rect 2360 207 2367 233
rect 2305 203 2367 207
rect 2267 199 2367 203
rect 1743 178 1774 199
rect 2164 178 2200 199
rect 1586 177 1623 178
rect 1585 168 1623 177
rect 1585 148 1594 168
rect 1614 148 1623 168
rect 1585 140 1623 148
rect 1689 172 1774 178
rect 1799 177 1836 178
rect 1689 152 1697 172
rect 1717 152 1774 172
rect 1689 144 1774 152
rect 1798 168 1836 177
rect 1798 148 1807 168
rect 1827 148 1836 168
rect 1689 143 1725 144
rect 1798 140 1836 148
rect 1902 172 1987 178
rect 2007 177 2044 178
rect 1902 152 1910 172
rect 1930 171 1987 172
rect 1930 152 1959 171
rect 1902 151 1959 152
rect 1980 151 1987 171
rect 1902 144 1987 151
rect 2006 168 2044 177
rect 2006 148 2015 168
rect 2035 148 2044 168
rect 1902 143 1938 144
rect 2006 140 2044 148
rect 2110 172 2254 178
rect 2110 152 2118 172
rect 2138 170 2226 172
rect 2138 152 2165 170
rect 2110 150 2165 152
rect 2199 152 2226 170
rect 2246 152 2254 172
rect 2199 150 2254 152
rect 2110 144 2254 150
rect 2110 143 2146 144
rect 2218 143 2254 144
rect 2320 177 2357 178
rect 2320 176 2358 177
rect 2320 168 2384 176
rect 2320 148 2329 168
rect 2349 154 2384 168
rect 2404 154 2407 174
rect 2349 149 2407 154
rect 2349 148 2384 149
rect 1586 111 1623 140
rect 1587 109 1623 111
rect 1799 109 1836 140
rect 1587 87 1836 109
rect 2007 108 2044 140
rect 2320 136 2384 148
rect 2424 119 2451 288
rect 4541 277 4550 297
rect 4570 277 4578 297
rect 4541 267 4578 277
rect 4637 297 4724 307
rect 4637 277 4646 297
rect 4666 277 4724 297
rect 4637 268 4724 277
rect 4637 267 4674 268
rect 4693 215 4724 268
rect 4754 297 4791 376
rect 4962 373 5355 393
rect 5375 373 5378 393
rect 4962 368 5378 373
rect 4962 367 5303 368
rect 4906 307 4937 308
rect 4754 277 4763 297
rect 4783 277 4791 297
rect 4754 267 4791 277
rect 4850 300 4937 307
rect 4850 297 4911 300
rect 4850 277 4859 297
rect 4879 280 4911 297
rect 4932 280 4937 300
rect 4879 277 4937 280
rect 4850 270 4937 277
rect 4962 297 4999 367
rect 5265 366 5302 367
rect 6647 358 6684 437
rect 6725 424 6835 437
rect 6799 368 6830 369
rect 6647 338 6656 358
rect 6676 338 6684 358
rect 6647 328 6684 338
rect 6743 358 6830 368
rect 6743 338 6752 358
rect 6772 338 6830 358
rect 6743 329 6830 338
rect 6743 328 6780 329
rect 5114 307 5150 308
rect 4962 277 4971 297
rect 4991 277 4999 297
rect 4850 268 4906 270
rect 4850 267 4887 268
rect 4962 267 4999 277
rect 5058 297 5206 307
rect 5306 304 5402 306
rect 5058 277 5067 297
rect 5087 277 5177 297
rect 5197 277 5206 297
rect 5058 268 5206 277
rect 5264 297 5402 304
rect 5264 277 5273 297
rect 5293 277 5402 297
rect 5264 268 5402 277
rect 6799 276 6830 329
rect 6860 358 6897 437
rect 7068 434 7461 454
rect 7481 434 7484 454
rect 7068 429 7484 434
rect 7068 428 7409 429
rect 7012 368 7043 369
rect 6860 338 6869 358
rect 6889 338 6897 358
rect 6860 328 6897 338
rect 6956 361 7043 368
rect 6956 358 7017 361
rect 6956 338 6965 358
rect 6985 341 7017 358
rect 7038 341 7043 361
rect 6985 338 7043 341
rect 6956 331 7043 338
rect 7068 358 7105 428
rect 7371 427 7408 428
rect 7220 368 7256 369
rect 7068 338 7077 358
rect 7097 338 7105 358
rect 6956 329 7012 331
rect 6956 328 6993 329
rect 7068 328 7105 338
rect 7164 358 7312 368
rect 7412 365 7508 367
rect 7164 338 7173 358
rect 7193 338 7283 358
rect 7303 338 7312 358
rect 7164 329 7312 338
rect 7370 358 7508 365
rect 7370 338 7379 358
rect 7399 338 7508 358
rect 7370 329 7508 338
rect 7164 328 7201 329
rect 7220 277 7256 329
rect 7275 328 7312 329
rect 7371 328 7408 329
rect 6691 275 6732 276
rect 6583 268 6732 275
rect 5058 267 5095 268
rect 5114 216 5150 268
rect 5169 267 5206 268
rect 5265 267 5302 268
rect 4585 214 4626 215
rect 4477 207 4626 214
rect 4477 187 4595 207
rect 4615 187 4626 207
rect 4477 179 4626 187
rect 4693 211 5052 215
rect 4693 206 5015 211
rect 4693 182 4806 206
rect 4830 187 5015 206
rect 5039 187 5052 211
rect 4830 182 5052 187
rect 4693 179 5052 182
rect 5114 179 5149 216
rect 5217 213 5317 216
rect 5217 209 5284 213
rect 5217 183 5229 209
rect 5255 187 5284 209
rect 5310 187 5317 213
rect 5255 183 5317 187
rect 5217 179 5317 183
rect 4693 158 4724 179
rect 5114 158 5150 179
rect 4536 157 4573 158
rect 4535 148 4573 157
rect 4535 128 4544 148
rect 4564 128 4573 148
rect 4535 120 4573 128
rect 4639 152 4724 158
rect 4749 157 4786 158
rect 4639 132 4647 152
rect 4667 132 4724 152
rect 4639 124 4724 132
rect 4748 148 4786 157
rect 4748 128 4757 148
rect 4777 128 4786 148
rect 4639 123 4675 124
rect 4748 120 4786 128
rect 4852 152 4937 158
rect 4957 157 4994 158
rect 4852 132 4860 152
rect 4880 151 4937 152
rect 4880 132 4909 151
rect 4852 131 4909 132
rect 4930 131 4937 151
rect 4852 124 4937 131
rect 4956 148 4994 157
rect 4956 128 4965 148
rect 4985 128 4994 148
rect 4852 123 4888 124
rect 4956 120 4994 128
rect 5060 152 5204 158
rect 5060 132 5068 152
rect 5088 132 5176 152
rect 5196 132 5204 152
rect 5060 124 5204 132
rect 5060 123 5096 124
rect 5168 123 5204 124
rect 5270 157 5307 158
rect 5270 156 5308 157
rect 5270 148 5334 156
rect 5270 128 5279 148
rect 5299 134 5334 148
rect 5354 134 5357 154
rect 5299 129 5357 134
rect 5299 128 5334 129
rect 2397 113 2525 119
rect 2397 110 2486 113
rect 2283 108 2486 110
rect 2007 92 2486 108
rect 2513 92 2525 113
rect 1668 81 1779 87
rect 2007 82 2525 92
rect 4536 91 4573 120
rect 2283 81 2525 82
rect 1668 73 1709 81
rect 1668 53 1676 73
rect 1695 53 1709 73
rect 1668 51 1709 53
rect 1737 73 1779 81
rect 2397 79 2525 81
rect 4537 89 4573 91
rect 4749 89 4786 120
rect 1737 53 1753 73
rect 1772 53 1779 73
rect 4537 67 4786 89
rect 4957 88 4994 120
rect 5270 116 5334 128
rect 5374 108 5401 268
rect 6583 248 6701 268
rect 6721 248 6732 268
rect 6583 240 6732 248
rect 6799 272 7158 276
rect 6799 267 7121 272
rect 6799 243 6912 267
rect 6936 248 7121 267
rect 7145 248 7158 272
rect 6936 243 7158 248
rect 6799 240 7158 243
rect 7220 240 7255 277
rect 7323 274 7423 277
rect 7323 270 7390 274
rect 7323 244 7335 270
rect 7361 248 7390 270
rect 7416 248 7423 274
rect 7361 244 7423 248
rect 7323 240 7423 244
rect 6799 219 6830 240
rect 7220 219 7256 240
rect 6642 218 6679 219
rect 6641 209 6679 218
rect 6641 189 6650 209
rect 6670 189 6679 209
rect 6641 181 6679 189
rect 6745 213 6830 219
rect 6855 218 6892 219
rect 6745 193 6753 213
rect 6773 193 6830 213
rect 6745 185 6830 193
rect 6854 209 6892 218
rect 6854 189 6863 209
rect 6883 189 6892 209
rect 6745 184 6781 185
rect 6854 181 6892 189
rect 6958 213 7043 219
rect 7063 218 7100 219
rect 6958 193 6966 213
rect 6986 212 7043 213
rect 6986 193 7015 212
rect 6958 192 7015 193
rect 7036 192 7043 212
rect 6958 185 7043 192
rect 7062 209 7100 218
rect 7062 189 7071 209
rect 7091 189 7100 209
rect 6958 184 6994 185
rect 7062 181 7100 189
rect 7166 213 7310 219
rect 7166 193 7174 213
rect 7194 211 7282 213
rect 7194 193 7221 211
rect 7166 191 7221 193
rect 7255 193 7282 211
rect 7302 193 7310 213
rect 7255 191 7310 193
rect 7166 185 7310 191
rect 7166 184 7202 185
rect 7274 184 7310 185
rect 7376 218 7413 219
rect 7376 217 7414 218
rect 7376 209 7440 217
rect 7376 189 7385 209
rect 7405 195 7440 209
rect 7460 195 7463 215
rect 7405 190 7463 195
rect 7405 189 7440 190
rect 6642 152 6679 181
rect 6643 150 6679 152
rect 6855 150 6892 181
rect 6643 128 6892 150
rect 7063 149 7100 181
rect 7376 177 7440 189
rect 7480 160 7507 329
rect 7453 154 7581 160
rect 7453 151 7542 154
rect 7339 149 7542 151
rect 7063 133 7542 149
rect 7569 133 7581 154
rect 6724 122 6835 128
rect 7063 123 7581 133
rect 7339 122 7581 123
rect 6724 114 6765 122
rect 5370 94 5493 108
rect 5370 90 5422 94
rect 5233 88 5422 90
rect 4957 68 5422 88
rect 5481 68 5493 94
rect 6724 94 6732 114
rect 6751 94 6765 114
rect 6724 92 6765 94
rect 6793 114 6835 122
rect 7453 120 7581 122
rect 6793 94 6809 114
rect 6828 94 6835 114
rect 6793 92 6835 94
rect 6724 77 6835 92
rect 1737 51 1779 53
rect 1668 36 1779 51
rect 4618 61 4729 67
rect 4957 62 5493 68
rect 5233 61 5493 62
rect 4618 53 4659 61
rect 4618 33 4626 53
rect 4645 33 4659 53
rect 4618 31 4659 33
rect 4687 53 4729 61
rect 5361 59 5493 61
rect 5404 57 5493 59
rect 4687 33 4703 53
rect 4722 33 4729 53
rect 4687 31 4729 33
rect 4618 16 4729 31
<< viali >>
rect 4408 9315 4427 9335
rect 4485 9315 4504 9335
rect 423 9232 452 9259
rect 497 9235 526 9262
rect 193 9119 222 9148
rect 1155 9227 1175 9247
rect 711 9134 732 9154
rect 1084 9041 1110 9067
rect 709 8985 730 9005
rect 919 8985 944 9005
rect 1134 8988 1154 9008
rect 3776 9214 3796 9234
rect 3988 9219 4011 9239
rect 4200 9217 4221 9237
rect 3820 9155 3846 9181
rect 426 8887 445 8907
rect 503 8887 522 8907
rect 1361 8988 1390 9015
rect 1435 8991 1464 9018
rect 2093 8983 2113 9003
rect 1649 8890 1670 8910
rect 3204 8976 3230 8998
rect 3469 9005 3488 9025
rect 3546 9005 3565 9025
rect 4198 9068 4219 9088
rect 2022 8797 2048 8823
rect 1647 8741 1668 8761
rect 1862 8745 1882 8762
rect 2072 8744 2092 8764
rect 199 8678 224 8697
rect 422 8678 451 8705
rect 496 8681 525 8708
rect 1154 8673 1174 8693
rect 3755 8975 3775 8995
rect 9464 9356 9483 9376
rect 9541 9356 9560 9376
rect 5479 9273 5508 9300
rect 5553 9276 5582 9303
rect 5249 9160 5278 9189
rect 6211 9268 6231 9288
rect 5767 9175 5788 9195
rect 6140 9082 6166 9108
rect 5765 9026 5786 9046
rect 5975 9026 6000 9046
rect 6190 9029 6210 9049
rect 4404 8960 4433 8987
rect 4478 8963 4507 8990
rect 4705 8971 4730 8990
rect 2837 8904 2857 8924
rect 3261 8907 3282 8927
rect 8832 9255 8852 9275
rect 9044 9260 9067 9280
rect 9256 9258 9277 9278
rect 8876 9196 8902 9222
rect 5482 8928 5501 8948
rect 5559 8928 5578 8948
rect 6417 9029 6446 9056
rect 6491 9032 6520 9059
rect 2881 8845 2907 8871
rect 7149 9024 7169 9044
rect 6705 8931 6726 8951
rect 8260 9017 8286 9039
rect 8525 9046 8544 9066
rect 8602 9046 8621 9066
rect 9254 9109 9275 9129
rect 3048 8766 3069 8807
rect 710 8580 731 8600
rect 1364 8643 1383 8663
rect 1441 8643 1460 8663
rect 1699 8670 1725 8692
rect 3259 8758 3280 8778
rect 2816 8665 2836 8685
rect 3189 8672 3221 8689
rect 7078 8838 7104 8864
rect 3465 8650 3494 8677
rect 3539 8653 3568 8680
rect 4407 8761 4426 8781
rect 4484 8761 4503 8781
rect 1083 8487 1109 8513
rect 708 8431 729 8451
rect 918 8429 941 8449
rect 1133 8434 1153 8454
rect 6703 8782 6724 8802
rect 6918 8786 6938 8803
rect 7128 8785 7148 8805
rect 5255 8719 5280 8738
rect 5478 8719 5507 8746
rect 5552 8722 5581 8749
rect 3775 8660 3795 8680
rect 3985 8663 4010 8683
rect 4199 8663 4220 8683
rect 3819 8601 3845 8627
rect 3041 8466 3072 8493
rect 3329 8494 3348 8514
rect 3406 8494 3425 8514
rect 425 8333 444 8353
rect 502 8333 521 8353
rect 1502 8396 1531 8423
rect 1576 8399 1605 8426
rect 1860 8390 1880 8407
rect 2234 8391 2254 8411
rect 1790 8298 1811 8318
rect 2163 8205 2189 8231
rect 424 8129 453 8156
rect 498 8132 527 8159
rect 194 8016 223 8045
rect 1156 8124 1176 8144
rect 1788 8149 1809 8169
rect 1996 8147 2023 8168
rect 2213 8152 2233 8172
rect 712 8031 733 8051
rect 4197 8514 4218 8534
rect 2697 8393 2717 8413
rect 3121 8396 3142 8416
rect 3754 8421 3774 8441
rect 4707 8520 4736 8549
rect 4403 8406 4432 8433
rect 4477 8409 4506 8436
rect 2741 8334 2767 8360
rect 2908 8254 2931 8292
rect 3119 8247 3140 8267
rect 2676 8154 2696 8174
rect 3050 8158 3070 8175
rect 3325 8139 3354 8166
rect 3399 8142 3428 8169
rect 4409 8212 4428 8232
rect 4486 8212 4505 8232
rect 1505 8051 1524 8071
rect 1582 8051 1601 8071
rect 1858 8072 1889 8099
rect 1085 7938 1111 7964
rect 710 7882 731 7902
rect 920 7882 945 7902
rect 1135 7885 1155 7905
rect 3777 8111 3797 8131
rect 3989 8116 4012 8136
rect 4201 8114 4222 8134
rect 3821 8052 3847 8078
rect 427 7784 446 7804
rect 504 7784 523 7804
rect 1362 7885 1391 7912
rect 1436 7888 1465 7915
rect 1709 7876 1741 7893
rect 2094 7880 2114 7900
rect 1650 7787 1671 7807
rect 3205 7873 3231 7895
rect 3470 7902 3489 7922
rect 3547 7902 3566 7922
rect 4199 7965 4220 7985
rect 1861 7758 1882 7799
rect 2023 7694 2049 7720
rect 1648 7638 1669 7658
rect 2073 7641 2093 7661
rect 200 7575 225 7594
rect 423 7575 452 7602
rect 497 7578 526 7605
rect 1155 7570 1175 7590
rect 3756 7872 3776 7892
rect 6210 8714 6230 8734
rect 8811 9016 8831 9036
rect 9460 9001 9489 9028
rect 9534 9004 9563 9031
rect 9761 9012 9786 9031
rect 7893 8945 7913 8965
rect 8317 8948 8338 8968
rect 7937 8886 7963 8912
rect 8104 8807 8125 8848
rect 5766 8621 5787 8641
rect 6420 8684 6439 8704
rect 6497 8684 6516 8704
rect 6755 8711 6781 8733
rect 8315 8799 8336 8819
rect 7872 8706 7892 8726
rect 8245 8713 8277 8730
rect 8521 8691 8550 8718
rect 8595 8694 8624 8721
rect 9463 8802 9482 8822
rect 9540 8802 9559 8822
rect 6139 8528 6165 8554
rect 5764 8472 5785 8492
rect 5974 8470 5997 8490
rect 6189 8475 6209 8495
rect 8831 8701 8851 8721
rect 9041 8704 9066 8724
rect 9255 8704 9276 8724
rect 8875 8642 8901 8668
rect 8097 8507 8128 8534
rect 8385 8535 8404 8555
rect 8462 8535 8481 8555
rect 5481 8374 5500 8394
rect 5558 8374 5577 8394
rect 6558 8437 6587 8464
rect 6632 8440 6661 8467
rect 6916 8431 6936 8448
rect 7290 8432 7310 8452
rect 6846 8339 6867 8359
rect 7219 8246 7245 8272
rect 5480 8170 5509 8197
rect 5554 8173 5583 8200
rect 5250 8057 5279 8086
rect 6212 8165 6232 8185
rect 6844 8190 6865 8210
rect 7052 8188 7079 8209
rect 7269 8193 7289 8213
rect 5768 8072 5789 8092
rect 9253 8555 9274 8575
rect 7753 8434 7773 8454
rect 8177 8437 8198 8457
rect 8810 8462 8830 8482
rect 9763 8561 9792 8590
rect 9459 8447 9488 8474
rect 9533 8450 9562 8477
rect 7797 8375 7823 8401
rect 7964 8295 7987 8333
rect 8175 8288 8196 8308
rect 7732 8195 7752 8215
rect 8106 8199 8126 8216
rect 8381 8180 8410 8207
rect 8455 8183 8484 8210
rect 9465 8253 9484 8273
rect 9542 8253 9561 8273
rect 6561 8092 6580 8112
rect 6638 8092 6657 8112
rect 6914 8113 6945 8140
rect 6141 7979 6167 8005
rect 5766 7923 5787 7943
rect 5976 7923 6001 7943
rect 6191 7926 6211 7946
rect 4405 7857 4434 7884
rect 4479 7860 4508 7887
rect 4706 7868 4731 7887
rect 2838 7801 2858 7821
rect 3048 7803 3068 7820
rect 3262 7804 3283 7824
rect 8833 8152 8853 8172
rect 9045 8157 9068 8177
rect 9257 8155 9278 8175
rect 8877 8093 8903 8119
rect 5483 7825 5502 7845
rect 5560 7825 5579 7845
rect 6418 7926 6447 7953
rect 6492 7929 6521 7956
rect 2882 7742 2908 7768
rect 6765 7917 6797 7934
rect 7150 7921 7170 7941
rect 6706 7828 6727 7848
rect 8261 7914 8287 7936
rect 8526 7943 8545 7963
rect 8603 7943 8622 7963
rect 9255 8006 9276 8026
rect 6917 7799 6938 7840
rect 711 7477 732 7497
rect 1365 7540 1384 7560
rect 1442 7540 1461 7560
rect 1700 7567 1726 7589
rect 3260 7655 3281 7675
rect 2817 7562 2837 7582
rect 7079 7735 7105 7761
rect 3466 7547 3495 7574
rect 3540 7550 3569 7577
rect 4408 7658 4427 7678
rect 4485 7658 4504 7678
rect 1084 7384 1110 7410
rect 709 7328 730 7348
rect 919 7326 942 7346
rect 1134 7331 1154 7351
rect 6704 7679 6725 7699
rect 7129 7682 7149 7702
rect 5256 7616 5281 7635
rect 5479 7616 5508 7643
rect 5553 7619 5582 7646
rect 3776 7557 3796 7577
rect 3986 7560 4011 7580
rect 4200 7560 4221 7580
rect 3820 7498 3846 7524
rect 2707 7350 2755 7379
rect 3360 7378 3379 7398
rect 3437 7378 3456 7398
rect 426 7230 445 7250
rect 503 7230 522 7250
rect 1472 7306 1501 7333
rect 1546 7309 1575 7336
rect 2204 7301 2224 7321
rect 1760 7208 1781 7228
rect 2133 7115 2159 7141
rect 424 7026 453 7053
rect 498 7029 527 7056
rect 1758 7059 1779 7079
rect 1966 7059 1995 7078
rect 2183 7062 2203 7082
rect 194 6913 223 6942
rect 1156 7021 1176 7041
rect 712 6928 733 6948
rect 4198 7411 4219 7431
rect 3755 7318 3775 7338
rect 4708 7417 4737 7446
rect 2728 7277 2748 7297
rect 3152 7280 3173 7300
rect 4404 7303 4433 7330
rect 4478 7306 4507 7333
rect 2772 7218 2798 7244
rect 6211 7611 6231 7631
rect 8812 7913 8832 7933
rect 9461 7898 9490 7925
rect 9535 7901 9564 7928
rect 9762 7909 9787 7928
rect 7894 7842 7914 7862
rect 8104 7844 8124 7861
rect 8318 7845 8339 7865
rect 7938 7783 7964 7809
rect 5767 7518 5788 7538
rect 6421 7581 6440 7601
rect 6498 7581 6517 7601
rect 6756 7608 6782 7630
rect 8316 7696 8337 7716
rect 7873 7603 7893 7623
rect 8522 7588 8551 7615
rect 8596 7591 8625 7618
rect 9464 7699 9483 7719
rect 9541 7699 9560 7719
rect 6140 7425 6166 7451
rect 5765 7369 5786 7389
rect 5975 7367 5998 7387
rect 6190 7372 6210 7392
rect 8832 7598 8852 7618
rect 9042 7601 9067 7621
rect 9256 7601 9277 7621
rect 8876 7539 8902 7565
rect 7763 7391 7811 7420
rect 8416 7419 8435 7439
rect 8493 7419 8512 7439
rect 5482 7271 5501 7291
rect 5559 7271 5578 7291
rect 2937 7143 2964 7175
rect 3150 7131 3171 7151
rect 2707 7040 2727 7058
rect 3097 7036 3118 7056
rect 3356 7023 3385 7050
rect 3430 7026 3459 7053
rect 6528 7347 6557 7374
rect 6602 7350 6631 7377
rect 7260 7342 7280 7362
rect 6816 7249 6837 7269
rect 4409 7109 4428 7129
rect 4486 7109 4505 7129
rect 1475 6961 1494 6981
rect 1552 6961 1571 6981
rect 1085 6835 1111 6861
rect 710 6779 731 6799
rect 920 6779 945 6799
rect 1135 6782 1155 6802
rect 3777 7008 3797 7028
rect 3989 7013 4012 7033
rect 4201 7011 4222 7031
rect 3821 6949 3847 6975
rect 2176 6840 2224 6869
rect 427 6681 446 6701
rect 504 6681 523 6701
rect 1362 6782 1391 6809
rect 1436 6785 1465 6812
rect 2094 6777 2114 6797
rect 1650 6684 1671 6704
rect 3205 6770 3231 6792
rect 3470 6799 3489 6819
rect 3547 6799 3566 6819
rect 4199 6862 4220 6882
rect 2023 6591 2049 6617
rect 1648 6535 1669 6555
rect 1863 6539 1883 6556
rect 2073 6538 2093 6558
rect 200 6472 225 6491
rect 423 6472 452 6499
rect 497 6475 526 6502
rect 1155 6467 1175 6487
rect 3756 6769 3776 6789
rect 7189 7156 7215 7182
rect 5480 7067 5509 7094
rect 5554 7070 5583 7097
rect 6814 7100 6835 7120
rect 7022 7100 7051 7119
rect 7239 7103 7259 7123
rect 5250 6954 5279 6983
rect 6212 7062 6232 7082
rect 5768 6969 5789 6989
rect 9254 7452 9275 7472
rect 8811 7359 8831 7379
rect 9764 7458 9793 7487
rect 7784 7318 7804 7338
rect 8208 7321 8229 7341
rect 9460 7344 9489 7371
rect 9534 7347 9563 7374
rect 7828 7259 7854 7285
rect 7993 7184 8020 7216
rect 8206 7172 8227 7192
rect 7763 7081 7783 7099
rect 8153 7077 8174 7097
rect 8412 7064 8441 7091
rect 8486 7067 8515 7094
rect 9465 7150 9484 7170
rect 9542 7150 9561 7170
rect 6531 7002 6550 7022
rect 6608 7002 6627 7022
rect 6141 6876 6167 6902
rect 5766 6820 5787 6840
rect 5976 6820 6001 6840
rect 6191 6823 6211 6843
rect 4405 6754 4434 6781
rect 4479 6757 4508 6784
rect 4706 6765 4731 6784
rect 2838 6698 2858 6718
rect 3262 6701 3283 6721
rect 8833 7049 8853 7069
rect 9045 7054 9068 7074
rect 9257 7052 9278 7072
rect 8877 6990 8903 7016
rect 7232 6881 7280 6910
rect 5483 6722 5502 6742
rect 5560 6722 5579 6742
rect 6418 6823 6447 6850
rect 6492 6826 6521 6853
rect 2882 6639 2908 6665
rect 7150 6818 7170 6838
rect 6706 6725 6727 6745
rect 8261 6811 8287 6833
rect 8526 6840 8545 6860
rect 8603 6840 8622 6860
rect 9255 6903 9276 6923
rect 3049 6560 3070 6601
rect 711 6374 732 6394
rect 1365 6437 1384 6457
rect 1442 6437 1461 6457
rect 1700 6464 1726 6486
rect 3260 6552 3281 6572
rect 2817 6459 2837 6479
rect 3190 6466 3222 6483
rect 7079 6632 7105 6658
rect 3466 6444 3495 6471
rect 3540 6447 3569 6474
rect 4408 6555 4427 6575
rect 4485 6555 4504 6575
rect 1084 6281 1110 6307
rect 709 6225 730 6245
rect 919 6223 942 6243
rect 1134 6228 1154 6248
rect 6704 6576 6725 6596
rect 6919 6580 6939 6597
rect 7129 6579 7149 6599
rect 5256 6513 5281 6532
rect 5479 6513 5508 6540
rect 5553 6516 5582 6543
rect 3776 6454 3796 6474
rect 3986 6457 4011 6477
rect 4200 6457 4221 6477
rect 3820 6395 3846 6421
rect 3042 6260 3073 6287
rect 3330 6288 3349 6308
rect 3407 6288 3426 6308
rect 426 6127 445 6147
rect 503 6127 522 6147
rect 1503 6190 1532 6217
rect 1577 6193 1606 6220
rect 1861 6184 1881 6201
rect 2235 6185 2255 6205
rect 1791 6092 1812 6112
rect 2000 6067 2023 6105
rect 2164 5999 2190 6025
rect 425 5923 454 5950
rect 499 5926 528 5953
rect 195 5810 224 5839
rect 1157 5918 1177 5938
rect 1789 5943 1810 5963
rect 2214 5946 2234 5966
rect 713 5825 734 5845
rect 4198 6308 4219 6328
rect 2698 6187 2718 6207
rect 2908 6191 2935 6212
rect 3122 6190 3143 6210
rect 3755 6215 3775 6235
rect 4708 6314 4737 6343
rect 4404 6200 4433 6227
rect 4478 6203 4507 6230
rect 2742 6128 2768 6154
rect 3120 6041 3141 6061
rect 2677 5948 2697 5968
rect 3051 5952 3071 5969
rect 3326 5933 3355 5960
rect 3400 5936 3429 5963
rect 4410 6006 4429 6026
rect 4487 6006 4506 6026
rect 1506 5845 1525 5865
rect 1583 5845 1602 5865
rect 1859 5866 1890 5893
rect 1086 5732 1112 5758
rect 711 5676 732 5696
rect 921 5676 946 5696
rect 1136 5679 1156 5699
rect 3778 5905 3798 5925
rect 3990 5910 4013 5930
rect 4202 5908 4223 5928
rect 3822 5846 3848 5872
rect 428 5578 447 5598
rect 505 5578 524 5598
rect 1363 5679 1392 5706
rect 1437 5682 1466 5709
rect 1710 5670 1742 5687
rect 2095 5674 2115 5694
rect 1651 5581 1672 5601
rect 3206 5667 3232 5689
rect 3471 5696 3490 5716
rect 3548 5696 3567 5716
rect 4200 5759 4221 5779
rect 1862 5552 1883 5593
rect 2024 5488 2050 5514
rect 1649 5432 1670 5452
rect 2074 5435 2094 5455
rect 201 5369 226 5388
rect 424 5369 453 5396
rect 498 5372 527 5399
rect 1156 5364 1176 5384
rect 3757 5666 3777 5686
rect 6211 6508 6231 6528
rect 8812 6810 8832 6830
rect 9461 6795 9490 6822
rect 9535 6798 9564 6825
rect 9762 6806 9787 6825
rect 7894 6739 7914 6759
rect 8318 6742 8339 6762
rect 7938 6680 7964 6706
rect 8105 6601 8126 6642
rect 5767 6415 5788 6435
rect 6421 6478 6440 6498
rect 6498 6478 6517 6498
rect 6756 6505 6782 6527
rect 8316 6593 8337 6613
rect 7873 6500 7893 6520
rect 8246 6507 8278 6524
rect 8522 6485 8551 6512
rect 8596 6488 8625 6515
rect 9464 6596 9483 6616
rect 9541 6596 9560 6616
rect 6140 6322 6166 6348
rect 5765 6266 5786 6286
rect 5975 6264 5998 6284
rect 6190 6269 6210 6289
rect 8832 6495 8852 6515
rect 9042 6498 9067 6518
rect 9256 6498 9277 6518
rect 8876 6436 8902 6462
rect 8098 6301 8129 6328
rect 8386 6329 8405 6349
rect 8463 6329 8482 6349
rect 5482 6168 5501 6188
rect 5559 6168 5578 6188
rect 6559 6231 6588 6258
rect 6633 6234 6662 6261
rect 6917 6225 6937 6242
rect 7291 6226 7311 6246
rect 6847 6133 6868 6153
rect 7056 6108 7079 6146
rect 7220 6040 7246 6066
rect 5481 5964 5510 5991
rect 5555 5967 5584 5994
rect 5251 5851 5280 5880
rect 6213 5959 6233 5979
rect 6845 5984 6866 6004
rect 7270 5987 7290 6007
rect 5769 5866 5790 5886
rect 9254 6349 9275 6369
rect 7754 6228 7774 6248
rect 7964 6232 7991 6253
rect 8178 6231 8199 6251
rect 8811 6256 8831 6276
rect 9764 6355 9793 6384
rect 9460 6241 9489 6268
rect 9534 6244 9563 6271
rect 7798 6169 7824 6195
rect 8176 6082 8197 6102
rect 7733 5989 7753 6009
rect 8107 5993 8127 6010
rect 8382 5974 8411 6001
rect 8456 5977 8485 6004
rect 9466 6047 9485 6067
rect 9543 6047 9562 6067
rect 6562 5886 6581 5906
rect 6639 5886 6658 5906
rect 6915 5907 6946 5934
rect 6142 5773 6168 5799
rect 5767 5717 5788 5737
rect 5977 5717 6002 5737
rect 6192 5720 6212 5740
rect 4406 5651 4435 5678
rect 4480 5654 4509 5681
rect 4707 5662 4732 5681
rect 2839 5595 2859 5615
rect 3049 5597 3069 5614
rect 3263 5598 3284 5618
rect 8834 5946 8854 5966
rect 9046 5951 9069 5971
rect 9258 5949 9279 5969
rect 8878 5887 8904 5913
rect 5484 5619 5503 5639
rect 5561 5619 5580 5639
rect 6419 5720 6448 5747
rect 6493 5723 6522 5750
rect 2883 5536 2909 5562
rect 6766 5711 6798 5728
rect 7151 5715 7171 5735
rect 6707 5622 6728 5642
rect 8262 5708 8288 5730
rect 8527 5737 8546 5757
rect 8604 5737 8623 5757
rect 9256 5800 9277 5820
rect 6918 5593 6939 5634
rect 712 5271 733 5291
rect 1366 5334 1385 5354
rect 1443 5334 1462 5354
rect 1701 5361 1727 5383
rect 3261 5449 3282 5469
rect 2818 5356 2838 5376
rect 7080 5529 7106 5555
rect 3467 5341 3496 5368
rect 3541 5344 3570 5371
rect 4409 5452 4428 5472
rect 4486 5452 4505 5472
rect 2567 5283 2594 5323
rect 1085 5178 1111 5204
rect 710 5122 731 5142
rect 920 5120 943 5140
rect 1135 5125 1155 5145
rect 6705 5473 6726 5493
rect 7130 5476 7150 5496
rect 5257 5410 5282 5429
rect 5480 5410 5509 5437
rect 5554 5413 5583 5440
rect 3777 5351 3797 5371
rect 3987 5354 4012 5374
rect 4201 5354 4222 5374
rect 3821 5292 3847 5318
rect 3362 5166 3381 5186
rect 3439 5166 3458 5186
rect 427 5024 446 5044
rect 504 5024 523 5044
rect 1472 5106 1501 5133
rect 1546 5109 1575 5136
rect 2204 5101 2224 5121
rect 1760 5008 1781 5028
rect 2133 4915 2159 4941
rect 425 4820 454 4847
rect 499 4823 528 4850
rect 1758 4859 1779 4879
rect 1966 4858 1992 4882
rect 2183 4862 2203 4882
rect 195 4707 224 4736
rect 1157 4815 1177 4835
rect 713 4722 734 4742
rect 4199 5205 4220 5225
rect 3756 5112 3776 5132
rect 4709 5211 4738 5240
rect 2730 5065 2750 5085
rect 2937 5068 2962 5088
rect 3154 5068 3175 5088
rect 4405 5097 4434 5124
rect 4479 5100 4508 5127
rect 2774 5006 2800 5032
rect 6212 5405 6232 5425
rect 8813 5707 8833 5727
rect 9462 5692 9491 5719
rect 9536 5695 9565 5722
rect 9763 5703 9788 5722
rect 7895 5636 7915 5656
rect 8105 5638 8125 5655
rect 8319 5639 8340 5659
rect 7939 5577 7965 5603
rect 5768 5312 5789 5332
rect 6422 5375 6441 5395
rect 6499 5375 6518 5395
rect 6757 5402 6783 5424
rect 8317 5490 8338 5510
rect 7874 5397 7894 5417
rect 8523 5382 8552 5409
rect 8597 5385 8626 5412
rect 9465 5493 9484 5513
rect 9542 5493 9561 5513
rect 7623 5324 7650 5364
rect 6141 5219 6167 5245
rect 5766 5163 5787 5183
rect 5976 5161 5999 5181
rect 6191 5166 6211 5186
rect 8833 5392 8853 5412
rect 9043 5395 9068 5415
rect 9257 5395 9278 5415
rect 8877 5333 8903 5359
rect 8418 5207 8437 5227
rect 8495 5207 8514 5227
rect 3152 4919 3173 4939
rect 2709 4826 2729 4846
rect 5483 5065 5502 5085
rect 5560 5065 5579 5085
rect 6528 5147 6557 5174
rect 6602 5150 6631 5177
rect 3358 4811 3387 4838
rect 3432 4814 3461 4841
rect 4410 4903 4429 4923
rect 4487 4903 4506 4923
rect 7260 5142 7280 5162
rect 6816 5049 6837 5069
rect 1475 4761 1494 4781
rect 1552 4761 1571 4781
rect 1086 4629 1112 4655
rect 711 4573 732 4593
rect 921 4573 946 4593
rect 1136 4576 1156 4596
rect 3778 4802 3798 4822
rect 3990 4807 4013 4827
rect 4202 4805 4223 4825
rect 3822 4743 3848 4769
rect 2339 4624 2366 4664
rect 428 4475 447 4495
rect 505 4475 524 4495
rect 1363 4576 1392 4603
rect 1437 4579 1466 4606
rect 2095 4571 2115 4591
rect 1651 4478 1672 4498
rect 3206 4564 3232 4586
rect 3471 4593 3490 4613
rect 3548 4593 3567 4613
rect 4200 4656 4221 4676
rect 2024 4385 2050 4411
rect 1649 4329 1670 4349
rect 1864 4333 1884 4350
rect 2074 4332 2094 4352
rect 201 4266 226 4285
rect 424 4266 453 4293
rect 498 4269 527 4296
rect 1156 4261 1176 4281
rect 3757 4563 3777 4583
rect 7189 4956 7215 4982
rect 5481 4861 5510 4888
rect 5555 4864 5584 4891
rect 6814 4900 6835 4920
rect 7022 4899 7048 4923
rect 7239 4903 7259 4923
rect 5251 4748 5280 4777
rect 6213 4856 6233 4876
rect 5769 4763 5790 4783
rect 9255 5246 9276 5266
rect 8812 5153 8832 5173
rect 9765 5252 9794 5281
rect 7786 5106 7806 5126
rect 7993 5109 8018 5129
rect 8210 5109 8231 5129
rect 9461 5138 9490 5165
rect 9535 5141 9564 5168
rect 7830 5047 7856 5073
rect 8208 4960 8229 4980
rect 7765 4867 7785 4887
rect 8414 4852 8443 4879
rect 8488 4855 8517 4882
rect 9466 4944 9485 4964
rect 9543 4944 9562 4964
rect 6531 4802 6550 4822
rect 6608 4802 6627 4822
rect 6142 4670 6168 4696
rect 5767 4614 5788 4634
rect 5977 4614 6002 4634
rect 6192 4617 6212 4637
rect 4406 4548 4435 4575
rect 4480 4551 4509 4578
rect 4707 4559 4732 4578
rect 2839 4492 2859 4512
rect 3263 4495 3284 4515
rect 8834 4843 8854 4863
rect 9046 4848 9069 4868
rect 9258 4846 9279 4866
rect 8878 4784 8904 4810
rect 7395 4665 7422 4705
rect 5484 4516 5503 4536
rect 5561 4516 5580 4536
rect 6419 4617 6448 4644
rect 6493 4620 6522 4647
rect 2883 4433 2909 4459
rect 7151 4612 7171 4632
rect 6707 4519 6728 4539
rect 8262 4605 8288 4627
rect 8527 4634 8546 4654
rect 8604 4634 8623 4654
rect 9256 4697 9277 4717
rect 3050 4354 3071 4395
rect 712 4168 733 4188
rect 1366 4231 1385 4251
rect 1443 4231 1462 4251
rect 1701 4258 1727 4280
rect 3261 4346 3282 4366
rect 2818 4253 2838 4273
rect 3191 4260 3223 4277
rect 7080 4426 7106 4452
rect 3467 4238 3496 4265
rect 3541 4241 3570 4268
rect 4409 4349 4428 4369
rect 4486 4349 4505 4369
rect 1085 4075 1111 4101
rect 710 4019 731 4039
rect 920 4017 943 4037
rect 1135 4022 1155 4042
rect 6705 4370 6726 4390
rect 6920 4374 6940 4391
rect 7130 4373 7150 4393
rect 5257 4307 5282 4326
rect 5480 4307 5509 4334
rect 5554 4310 5583 4337
rect 3777 4248 3797 4268
rect 3987 4251 4012 4271
rect 4201 4251 4222 4271
rect 3821 4189 3847 4215
rect 3043 4054 3074 4081
rect 3331 4082 3350 4102
rect 3408 4082 3427 4102
rect 427 3921 446 3941
rect 504 3921 523 3941
rect 1504 3984 1533 4011
rect 1578 3987 1607 4014
rect 1862 3978 1882 3995
rect 2236 3979 2256 3999
rect 1792 3886 1813 3906
rect 2165 3793 2191 3819
rect 426 3717 455 3744
rect 500 3720 529 3747
rect 196 3604 225 3633
rect 1158 3712 1178 3732
rect 1790 3737 1811 3757
rect 1998 3735 2025 3756
rect 2215 3740 2235 3760
rect 714 3619 735 3639
rect 4199 4102 4220 4122
rect 2699 3981 2719 4001
rect 3123 3984 3144 4004
rect 3756 4009 3776 4029
rect 4709 4108 4738 4137
rect 4405 3994 4434 4021
rect 4479 3997 4508 4024
rect 2743 3922 2769 3948
rect 2910 3842 2933 3880
rect 3121 3835 3142 3855
rect 2678 3742 2698 3762
rect 3052 3746 3072 3763
rect 3327 3727 3356 3754
rect 3401 3730 3430 3757
rect 4411 3800 4430 3820
rect 4488 3800 4507 3820
rect 1507 3639 1526 3659
rect 1584 3639 1603 3659
rect 1860 3660 1891 3687
rect 1087 3526 1113 3552
rect 712 3470 733 3490
rect 922 3470 947 3490
rect 1137 3473 1157 3493
rect 3779 3699 3799 3719
rect 3991 3704 4014 3724
rect 4203 3702 4224 3722
rect 3823 3640 3849 3666
rect 429 3372 448 3392
rect 506 3372 525 3392
rect 1364 3473 1393 3500
rect 1438 3476 1467 3503
rect 1711 3464 1743 3481
rect 2096 3468 2116 3488
rect 1652 3375 1673 3395
rect 3207 3461 3233 3483
rect 3472 3490 3491 3510
rect 3549 3490 3568 3510
rect 4201 3553 4222 3573
rect 1863 3346 1884 3387
rect 2025 3282 2051 3308
rect 1650 3226 1671 3246
rect 2075 3229 2095 3249
rect 202 3163 227 3182
rect 425 3163 454 3190
rect 499 3166 528 3193
rect 1157 3158 1177 3178
rect 3758 3460 3778 3480
rect 6212 4302 6232 4322
rect 8813 4604 8833 4624
rect 9462 4589 9491 4616
rect 9536 4592 9565 4619
rect 9763 4600 9788 4619
rect 7895 4533 7915 4553
rect 8319 4536 8340 4556
rect 7939 4474 7965 4500
rect 8106 4395 8127 4436
rect 5768 4209 5789 4229
rect 6422 4272 6441 4292
rect 6499 4272 6518 4292
rect 6757 4299 6783 4321
rect 8317 4387 8338 4407
rect 7874 4294 7894 4314
rect 8247 4301 8279 4318
rect 8523 4279 8552 4306
rect 8597 4282 8626 4309
rect 9465 4390 9484 4410
rect 9542 4390 9561 4410
rect 6141 4116 6167 4142
rect 5766 4060 5787 4080
rect 5976 4058 5999 4078
rect 6191 4063 6211 4083
rect 8833 4289 8853 4309
rect 9043 4292 9068 4312
rect 9257 4292 9278 4312
rect 8877 4230 8903 4256
rect 8099 4095 8130 4122
rect 8387 4123 8406 4143
rect 8464 4123 8483 4143
rect 5483 3962 5502 3982
rect 5560 3962 5579 3982
rect 6560 4025 6589 4052
rect 6634 4028 6663 4055
rect 6918 4019 6938 4036
rect 7292 4020 7312 4040
rect 6848 3927 6869 3947
rect 7221 3834 7247 3860
rect 5482 3758 5511 3785
rect 5556 3761 5585 3788
rect 5252 3645 5281 3674
rect 6214 3753 6234 3773
rect 6846 3778 6867 3798
rect 7054 3776 7081 3797
rect 7271 3781 7291 3801
rect 5770 3660 5791 3680
rect 9255 4143 9276 4163
rect 7755 4022 7775 4042
rect 8179 4025 8200 4045
rect 8812 4050 8832 4070
rect 9765 4149 9794 4178
rect 9461 4035 9490 4062
rect 9535 4038 9564 4065
rect 7799 3963 7825 3989
rect 7966 3883 7989 3921
rect 8177 3876 8198 3896
rect 7734 3783 7754 3803
rect 8108 3787 8128 3804
rect 8383 3768 8412 3795
rect 8457 3771 8486 3798
rect 9467 3841 9486 3861
rect 9544 3841 9563 3861
rect 6563 3680 6582 3700
rect 6640 3680 6659 3700
rect 6916 3701 6947 3728
rect 6143 3567 6169 3593
rect 5768 3511 5789 3531
rect 5978 3511 6003 3531
rect 6193 3514 6213 3534
rect 4407 3445 4436 3472
rect 4481 3448 4510 3475
rect 4708 3456 4733 3475
rect 2840 3389 2860 3409
rect 3050 3391 3070 3408
rect 3264 3392 3285 3412
rect 8835 3740 8855 3760
rect 9047 3745 9070 3765
rect 9259 3743 9280 3763
rect 8879 3681 8905 3707
rect 5485 3413 5504 3433
rect 5562 3413 5581 3433
rect 6420 3514 6449 3541
rect 6494 3517 6523 3544
rect 2884 3330 2910 3356
rect 6767 3505 6799 3522
rect 7152 3509 7172 3529
rect 6708 3416 6729 3436
rect 8263 3502 8289 3524
rect 8528 3531 8547 3551
rect 8605 3531 8624 3551
rect 9257 3594 9278 3614
rect 6919 3387 6940 3428
rect 713 3065 734 3085
rect 1367 3128 1386 3148
rect 1444 3128 1463 3148
rect 1702 3155 1728 3177
rect 3262 3243 3283 3263
rect 2819 3150 2839 3170
rect 7081 3323 7107 3349
rect 3468 3135 3497 3162
rect 3542 3138 3571 3165
rect 4410 3246 4429 3266
rect 4487 3246 4506 3266
rect 2709 3078 2757 3107
rect 1086 2972 1112 2998
rect 711 2916 732 2936
rect 921 2914 944 2934
rect 1136 2919 1156 2939
rect 6706 3267 6727 3287
rect 7131 3270 7151 3290
rect 5258 3204 5283 3223
rect 5481 3204 5510 3231
rect 5555 3207 5584 3234
rect 3778 3145 3798 3165
rect 3988 3148 4013 3168
rect 4202 3148 4223 3168
rect 3822 3086 3848 3112
rect 3362 2966 3381 2986
rect 3439 2966 3458 2986
rect 428 2818 447 2838
rect 505 2818 524 2838
rect 1474 2894 1503 2921
rect 1548 2897 1577 2924
rect 1815 2891 1836 2911
rect 2206 2889 2226 2907
rect 1762 2796 1783 2816
rect 1969 2772 1996 2804
rect 2135 2703 2161 2729
rect 426 2614 455 2641
rect 500 2617 529 2644
rect 1760 2647 1781 2667
rect 2185 2650 2205 2670
rect 196 2501 225 2530
rect 1158 2609 1178 2629
rect 714 2516 735 2536
rect 4200 2999 4221 3019
rect 3757 2906 3777 2926
rect 4710 3005 4739 3034
rect 2730 2865 2750 2885
rect 2938 2869 2967 2888
rect 3154 2868 3175 2888
rect 4406 2891 4435 2918
rect 4480 2894 4509 2921
rect 2774 2806 2800 2832
rect 6213 3199 6233 3219
rect 8814 3501 8834 3521
rect 9463 3486 9492 3513
rect 9537 3489 9566 3516
rect 9764 3497 9789 3516
rect 7896 3430 7916 3450
rect 8106 3432 8126 3449
rect 8320 3433 8341 3453
rect 7940 3371 7966 3397
rect 5769 3106 5790 3126
rect 6423 3169 6442 3189
rect 6500 3169 6519 3189
rect 6758 3196 6784 3218
rect 8318 3284 8339 3304
rect 7875 3191 7895 3211
rect 8524 3176 8553 3203
rect 8598 3179 8627 3206
rect 9466 3287 9485 3307
rect 9543 3287 9562 3307
rect 7765 3119 7813 3148
rect 6142 3013 6168 3039
rect 5767 2957 5788 2977
rect 5977 2955 6000 2975
rect 6192 2960 6212 2980
rect 8834 3186 8854 3206
rect 9044 3189 9069 3209
rect 9258 3189 9279 3209
rect 8878 3127 8904 3153
rect 8418 3007 8437 3027
rect 8495 3007 8514 3027
rect 5484 2859 5503 2879
rect 5561 2859 5580 2879
rect 3152 2719 3173 2739
rect 2709 2626 2729 2646
rect 3358 2611 3387 2638
rect 3432 2614 3461 2641
rect 6530 2935 6559 2962
rect 6604 2938 6633 2965
rect 6871 2932 6892 2952
rect 7262 2930 7282 2948
rect 6818 2837 6839 2857
rect 7025 2813 7052 2845
rect 4411 2697 4430 2717
rect 4488 2697 4507 2717
rect 1477 2549 1496 2569
rect 1554 2549 1573 2569
rect 2178 2568 2226 2597
rect 1087 2423 1113 2449
rect 712 2367 733 2387
rect 922 2367 947 2387
rect 1137 2370 1157 2390
rect 3779 2596 3799 2616
rect 3991 2601 4014 2621
rect 4203 2599 4224 2619
rect 3823 2537 3849 2563
rect 429 2269 448 2289
rect 506 2269 525 2289
rect 1364 2370 1393 2397
rect 1438 2373 1467 2400
rect 2096 2365 2116 2385
rect 1652 2272 1673 2292
rect 3207 2358 3233 2380
rect 3472 2387 3491 2407
rect 3549 2387 3568 2407
rect 4201 2450 4222 2470
rect 2025 2179 2051 2205
rect 1650 2123 1671 2143
rect 1865 2127 1885 2144
rect 2075 2126 2095 2146
rect 202 2060 227 2079
rect 425 2060 454 2087
rect 499 2063 528 2090
rect 1157 2055 1177 2075
rect 3758 2357 3778 2377
rect 7191 2744 7217 2770
rect 5482 2655 5511 2682
rect 5556 2658 5585 2685
rect 6816 2688 6837 2708
rect 7241 2691 7261 2711
rect 5252 2542 5281 2571
rect 6214 2650 6234 2670
rect 5770 2557 5791 2577
rect 9256 3040 9277 3060
rect 8813 2947 8833 2967
rect 9766 3046 9795 3075
rect 7786 2906 7806 2926
rect 7994 2910 8023 2929
rect 8210 2909 8231 2929
rect 9462 2932 9491 2959
rect 9536 2935 9565 2962
rect 7830 2847 7856 2873
rect 8208 2760 8229 2780
rect 7765 2667 7785 2687
rect 8414 2652 8443 2679
rect 8488 2655 8517 2682
rect 9467 2738 9486 2758
rect 9544 2738 9563 2758
rect 6533 2590 6552 2610
rect 6610 2590 6629 2610
rect 7234 2609 7282 2638
rect 6143 2464 6169 2490
rect 5768 2408 5789 2428
rect 5978 2408 6003 2428
rect 6193 2411 6213 2431
rect 4407 2342 4436 2369
rect 4481 2345 4510 2372
rect 4708 2353 4733 2372
rect 2840 2286 2860 2306
rect 3264 2289 3285 2309
rect 8835 2637 8855 2657
rect 9047 2642 9070 2662
rect 9259 2640 9280 2660
rect 8879 2578 8905 2604
rect 5485 2310 5504 2330
rect 5562 2310 5581 2330
rect 6420 2411 6449 2438
rect 6494 2414 6523 2441
rect 2884 2227 2910 2253
rect 7152 2406 7172 2426
rect 6708 2313 6729 2333
rect 8263 2399 8289 2421
rect 8528 2428 8547 2448
rect 8605 2428 8624 2448
rect 9257 2491 9278 2511
rect 3051 2148 3072 2189
rect 713 1962 734 1982
rect 1367 2025 1386 2045
rect 1444 2025 1463 2045
rect 1702 2052 1728 2074
rect 3262 2140 3283 2160
rect 2819 2047 2839 2067
rect 3192 2054 3224 2071
rect 7081 2220 7107 2246
rect 3468 2032 3497 2059
rect 3542 2035 3571 2062
rect 4410 2143 4429 2163
rect 4487 2143 4506 2163
rect 1086 1869 1112 1895
rect 711 1813 732 1833
rect 921 1811 944 1831
rect 1136 1816 1156 1836
rect 6706 2164 6727 2184
rect 6921 2168 6941 2185
rect 7131 2167 7151 2187
rect 5258 2101 5283 2120
rect 5481 2101 5510 2128
rect 5555 2104 5584 2131
rect 3778 2042 3798 2062
rect 3988 2045 4013 2065
rect 4202 2045 4223 2065
rect 3822 1983 3848 2009
rect 3044 1848 3075 1875
rect 3332 1876 3351 1896
rect 3409 1876 3428 1896
rect 428 1715 447 1735
rect 505 1715 524 1735
rect 1505 1778 1534 1805
rect 1579 1781 1608 1808
rect 1863 1772 1883 1789
rect 2237 1773 2257 1793
rect 1793 1680 1814 1700
rect 2002 1655 2025 1693
rect 2166 1587 2192 1613
rect 427 1511 456 1538
rect 501 1514 530 1541
rect 197 1398 226 1427
rect 1159 1506 1179 1526
rect 1791 1531 1812 1551
rect 2216 1534 2236 1554
rect 715 1413 736 1433
rect 4200 1896 4221 1916
rect 2700 1775 2720 1795
rect 2910 1779 2937 1800
rect 3124 1778 3145 1798
rect 3757 1803 3777 1823
rect 4710 1902 4739 1931
rect 4406 1788 4435 1815
rect 4480 1791 4509 1818
rect 2744 1716 2770 1742
rect 3122 1629 3143 1649
rect 2679 1536 2699 1556
rect 3053 1540 3073 1557
rect 3328 1521 3357 1548
rect 3402 1524 3431 1551
rect 4412 1594 4431 1614
rect 4489 1594 4508 1614
rect 1508 1433 1527 1453
rect 1585 1433 1604 1453
rect 1861 1454 1892 1481
rect 1088 1320 1114 1346
rect 713 1264 734 1284
rect 923 1264 948 1284
rect 1138 1267 1158 1287
rect 3780 1493 3800 1513
rect 3992 1498 4015 1518
rect 4204 1496 4225 1516
rect 3824 1434 3850 1460
rect 430 1166 449 1186
rect 507 1166 526 1186
rect 1365 1267 1394 1294
rect 1439 1270 1468 1297
rect 1712 1258 1744 1275
rect 2097 1262 2117 1282
rect 1653 1169 1674 1189
rect 3208 1255 3234 1277
rect 3473 1284 3492 1304
rect 3550 1284 3569 1304
rect 4202 1347 4223 1367
rect 1864 1140 1885 1181
rect 2026 1076 2052 1102
rect 1651 1020 1672 1040
rect 2076 1023 2096 1043
rect 203 957 228 976
rect 426 957 455 984
rect 500 960 529 987
rect 1158 952 1178 972
rect 3759 1254 3779 1274
rect 6213 2096 6233 2116
rect 8814 2398 8834 2418
rect 9463 2383 9492 2410
rect 9537 2386 9566 2413
rect 9764 2394 9789 2413
rect 7896 2327 7916 2347
rect 8320 2330 8341 2350
rect 7940 2268 7966 2294
rect 8107 2189 8128 2230
rect 5769 2003 5790 2023
rect 6423 2066 6442 2086
rect 6500 2066 6519 2086
rect 6758 2093 6784 2115
rect 8318 2181 8339 2201
rect 7875 2088 7895 2108
rect 8248 2095 8280 2112
rect 8524 2073 8553 2100
rect 8598 2076 8627 2103
rect 9466 2184 9485 2204
rect 9543 2184 9562 2204
rect 6142 1910 6168 1936
rect 5767 1854 5788 1874
rect 5977 1852 6000 1872
rect 6192 1857 6212 1877
rect 8834 2083 8854 2103
rect 9044 2086 9069 2106
rect 9258 2086 9279 2106
rect 8878 2024 8904 2050
rect 8100 1889 8131 1916
rect 8388 1917 8407 1937
rect 8465 1917 8484 1937
rect 5484 1756 5503 1776
rect 5561 1756 5580 1776
rect 6561 1819 6590 1846
rect 6635 1822 6664 1849
rect 6919 1813 6939 1830
rect 7293 1814 7313 1834
rect 6849 1721 6870 1741
rect 7058 1696 7081 1734
rect 7222 1628 7248 1654
rect 5483 1552 5512 1579
rect 5557 1555 5586 1582
rect 5253 1439 5282 1468
rect 6215 1547 6235 1567
rect 6847 1572 6868 1592
rect 7272 1575 7292 1595
rect 5771 1454 5792 1474
rect 9256 1937 9277 1957
rect 7756 1816 7776 1836
rect 7966 1820 7993 1841
rect 8180 1819 8201 1839
rect 8813 1844 8833 1864
rect 9766 1943 9795 1972
rect 9462 1829 9491 1856
rect 9536 1832 9565 1859
rect 7800 1757 7826 1783
rect 8178 1670 8199 1690
rect 7735 1577 7755 1597
rect 8109 1581 8129 1598
rect 8384 1562 8413 1589
rect 8458 1565 8487 1592
rect 9468 1635 9487 1655
rect 9545 1635 9564 1655
rect 6564 1474 6583 1494
rect 6641 1474 6660 1494
rect 6917 1495 6948 1522
rect 6144 1361 6170 1387
rect 5769 1305 5790 1325
rect 5979 1305 6004 1325
rect 6194 1308 6214 1328
rect 4408 1239 4437 1266
rect 4482 1242 4511 1269
rect 4709 1250 4734 1269
rect 2841 1183 2861 1203
rect 3051 1185 3071 1202
rect 3265 1186 3286 1206
rect 8836 1534 8856 1554
rect 9048 1539 9071 1559
rect 9260 1537 9281 1557
rect 8880 1475 8906 1501
rect 5486 1207 5505 1227
rect 5563 1207 5582 1227
rect 6421 1308 6450 1335
rect 6495 1311 6524 1338
rect 2885 1124 2911 1150
rect 6768 1299 6800 1316
rect 7153 1303 7173 1323
rect 6709 1210 6730 1230
rect 8264 1296 8290 1318
rect 8529 1325 8548 1345
rect 8606 1325 8625 1345
rect 9258 1388 9279 1408
rect 6920 1181 6941 1222
rect 714 859 735 879
rect 1368 922 1387 942
rect 1445 922 1464 942
rect 1703 949 1729 971
rect 3263 1037 3284 1057
rect 2820 944 2840 964
rect 7082 1117 7108 1143
rect 3469 929 3498 956
rect 3543 932 3572 959
rect 4411 1040 4430 1060
rect 4488 1040 4507 1060
rect 1087 766 1113 792
rect 712 710 733 730
rect 922 708 945 728
rect 1137 713 1157 733
rect 6707 1061 6728 1081
rect 7132 1064 7152 1084
rect 5259 998 5284 1017
rect 5482 998 5511 1025
rect 5556 1001 5585 1028
rect 3779 939 3799 959
rect 3989 942 4014 962
rect 4203 942 4224 962
rect 3823 880 3849 906
rect 4201 793 4222 813
rect 3758 700 3778 720
rect 4711 799 4740 828
rect 4407 685 4436 712
rect 4481 688 4510 715
rect 429 612 448 632
rect 6214 993 6234 1013
rect 8815 1295 8835 1315
rect 9464 1280 9493 1307
rect 9538 1283 9567 1310
rect 9765 1291 9790 1310
rect 7897 1224 7917 1244
rect 8107 1226 8127 1243
rect 8321 1227 8342 1247
rect 7941 1165 7967 1191
rect 5770 900 5791 920
rect 6424 963 6443 983
rect 6501 963 6520 983
rect 6759 990 6785 1012
rect 8319 1078 8340 1098
rect 7876 985 7896 1005
rect 8525 970 8554 997
rect 8599 973 8628 1000
rect 9467 1081 9486 1101
rect 9544 1081 9563 1101
rect 6143 807 6169 833
rect 5768 751 5789 771
rect 5978 749 6001 769
rect 6193 754 6213 774
rect 8835 980 8855 1000
rect 9045 983 9070 1003
rect 9259 983 9280 1003
rect 8879 921 8905 947
rect 9257 834 9278 854
rect 8814 741 8834 761
rect 9767 840 9796 869
rect 9463 726 9492 753
rect 9537 729 9566 756
rect 506 612 525 632
rect 757 529 786 550
rect 5485 653 5504 673
rect 5562 653 5581 673
rect 5813 570 5842 591
rect 9848 574 9877 595
rect 4792 533 4821 554
rect 1673 398 1702 425
rect 1747 401 1776 428
rect 6729 439 6758 466
rect 6803 442 6832 469
rect 2405 393 2425 413
rect 1961 300 1982 320
rect 4623 378 4652 405
rect 4697 381 4726 408
rect 2334 207 2360 233
rect 1959 151 1980 171
rect 2165 150 2199 170
rect 2384 154 2404 174
rect 5355 373 5375 393
rect 4911 280 4932 300
rect 7461 434 7481 454
rect 7017 341 7038 361
rect 5284 187 5310 213
rect 4909 131 4930 151
rect 5334 134 5354 154
rect 2486 92 2513 113
rect 1676 53 1695 73
rect 1753 53 1772 73
rect 7390 248 7416 274
rect 7015 192 7036 212
rect 7221 191 7255 211
rect 7440 195 7460 215
rect 7542 133 7569 154
rect 5422 68 5481 94
rect 6732 94 6751 114
rect 6809 94 6828 114
rect 4626 33 4645 53
rect 4703 33 4722 53
<< metal1 >>
rect 8775 9394 9077 9396
rect 6206 9371 6241 9373
rect 5242 9368 6241 9371
rect 3719 9353 4021 9355
rect 1150 9330 1185 9332
rect 186 9327 1185 9330
rect 185 9303 1185 9327
rect 185 9148 233 9303
rect 419 9262 529 9276
rect 419 9259 497 9262
rect 419 9232 423 9259
rect 452 9235 497 9259
rect 526 9235 529 9262
rect 1150 9252 1185 9303
rect 452 9232 529 9235
rect 419 9217 529 9232
rect 1148 9247 1185 9252
rect 1148 9227 1155 9247
rect 1175 9227 1185 9247
rect 1148 9220 1185 9227
rect 3658 9324 4021 9353
rect 3658 9322 3719 9324
rect 1148 9219 1183 9220
rect 185 9119 193 9148
rect 222 9119 233 9148
rect 185 9114 233 9119
rect 704 9154 736 9161
rect 704 9134 711 9154
rect 732 9134 736 9154
rect 704 9069 736 9134
rect 1074 9069 1114 9070
rect 704 9067 1116 9069
rect 704 9041 1084 9067
rect 1110 9041 1116 9067
rect 704 9033 1116 9041
rect 704 9005 736 9033
rect 1149 9013 1183 9219
rect 3200 9102 3237 9104
rect 3658 9102 3691 9322
rect 3979 9243 4021 9324
rect 4401 9335 4512 9352
rect 4401 9315 4408 9335
rect 4427 9315 4485 9335
rect 4504 9315 4512 9335
rect 4401 9293 4512 9315
rect 5241 9344 6241 9368
rect 3768 9241 3803 9242
rect 2087 9086 2121 9087
rect 1218 9051 2122 9086
rect 3200 9073 3691 9102
rect 704 8985 709 9005
rect 730 8985 736 9005
rect 704 8978 736 8985
rect 911 9005 950 9011
rect 911 8985 919 9005
rect 944 8985 950 9005
rect 911 8978 950 8985
rect 1127 9008 1183 9013
rect 1127 8988 1134 9008
rect 1154 8988 1183 9008
rect 1127 8981 1183 8988
rect 1127 8980 1162 8981
rect 919 8932 950 8978
rect 418 8907 529 8929
rect 418 8887 426 8907
rect 445 8887 503 8907
rect 522 8887 529 8907
rect 918 8915 950 8932
rect 1219 8915 1256 9051
rect 1357 9018 1467 9032
rect 1357 9015 1435 9018
rect 1357 8988 1361 9015
rect 1390 8991 1435 9015
rect 1464 8991 1467 9018
rect 2087 9008 2121 9051
rect 1390 8988 1467 8991
rect 1357 8973 1467 8988
rect 2086 9003 2121 9008
rect 3200 9007 3237 9073
rect 3658 9072 3691 9073
rect 3747 9234 3803 9241
rect 3747 9214 3776 9234
rect 3796 9214 3803 9234
rect 3747 9209 3803 9214
rect 3977 9239 4021 9243
rect 3977 9219 3988 9239
rect 4011 9219 4021 9239
rect 3977 9212 4021 9219
rect 4194 9237 4226 9244
rect 4194 9217 4200 9237
rect 4221 9217 4226 9237
rect 3977 9210 4020 9212
rect 2086 8983 2093 9003
rect 2113 8983 2121 9003
rect 2086 8975 2121 8983
rect 918 8902 1256 8915
rect 418 8870 529 8887
rect 919 8883 1256 8902
rect 1198 8882 1256 8883
rect 1642 8910 1674 8917
rect 1642 8890 1649 8910
rect 1670 8890 1674 8910
rect 1642 8825 1674 8890
rect 2012 8825 2052 8826
rect 1642 8823 2054 8825
rect 1642 8797 2022 8823
rect 2048 8797 2054 8823
rect 1642 8789 2054 8797
rect 188 8750 1184 8776
rect 1642 8761 1674 8789
rect 190 8697 232 8750
rect 190 8678 199 8697
rect 224 8678 232 8697
rect 190 8668 232 8678
rect 418 8708 528 8722
rect 418 8705 496 8708
rect 418 8678 422 8705
rect 451 8681 496 8705
rect 525 8681 528 8708
rect 1148 8698 1182 8750
rect 1642 8741 1647 8761
rect 1668 8741 1674 8761
rect 1642 8734 1674 8741
rect 1852 8762 1890 8772
rect 2087 8769 2121 8975
rect 3195 8998 3237 9007
rect 3195 8976 3204 8998
rect 3230 8976 3237 8998
rect 3462 9025 3573 9042
rect 3462 9005 3469 9025
rect 3488 9005 3546 9025
rect 3565 9005 3573 9025
rect 3462 8983 3573 9005
rect 3747 9003 3781 9209
rect 4194 9189 4226 9217
rect 3814 9181 4226 9189
rect 3814 9155 3820 9181
rect 3846 9155 4226 9181
rect 5241 9189 5289 9344
rect 5475 9303 5585 9317
rect 5475 9300 5553 9303
rect 5475 9273 5479 9300
rect 5508 9276 5553 9300
rect 5582 9276 5585 9303
rect 6206 9293 6241 9344
rect 5508 9273 5585 9276
rect 5475 9258 5585 9273
rect 6204 9288 6241 9293
rect 6204 9268 6211 9288
rect 6231 9268 6241 9288
rect 6204 9261 6241 9268
rect 8714 9365 9077 9394
rect 8714 9363 8775 9365
rect 6204 9260 6239 9261
rect 5241 9160 5249 9189
rect 5278 9160 5289 9189
rect 5241 9155 5289 9160
rect 5760 9195 5792 9202
rect 5760 9175 5767 9195
rect 5788 9175 5792 9195
rect 3814 9153 4226 9155
rect 3816 9152 3856 9153
rect 4194 9088 4226 9153
rect 4194 9068 4198 9088
rect 4219 9068 4226 9088
rect 4194 9061 4226 9068
rect 5760 9110 5792 9175
rect 6130 9110 6170 9111
rect 5760 9108 6172 9110
rect 5760 9082 6140 9108
rect 6166 9082 6172 9108
rect 5760 9074 6172 9082
rect 5760 9046 5792 9074
rect 6205 9054 6239 9260
rect 8256 9143 8293 9145
rect 8714 9143 8747 9363
rect 9035 9284 9077 9365
rect 9457 9376 9568 9393
rect 9457 9356 9464 9376
rect 9483 9356 9541 9376
rect 9560 9356 9568 9376
rect 9457 9334 9568 9356
rect 8824 9282 8859 9283
rect 7143 9127 7177 9128
rect 6274 9092 7178 9127
rect 8256 9114 8747 9143
rect 5760 9026 5765 9046
rect 5786 9026 5792 9046
rect 5760 9019 5792 9026
rect 5967 9046 6006 9052
rect 5967 9026 5975 9046
rect 6000 9026 6006 9046
rect 5967 9019 6006 9026
rect 6183 9049 6239 9054
rect 6183 9029 6190 9049
rect 6210 9029 6239 9049
rect 6183 9022 6239 9029
rect 6183 9021 6218 9022
rect 3747 8995 3782 9003
rect 3195 8966 3237 8976
rect 3747 8975 3755 8995
rect 3775 8975 3782 8995
rect 3747 8970 3782 8975
rect 4401 8990 4511 9005
rect 4401 8987 4478 8990
rect 3195 8965 3236 8966
rect 2829 8931 2864 8932
rect 1852 8745 1862 8762
rect 1882 8745 1890 8762
rect 1693 8702 1734 8703
rect 451 8678 528 8681
rect 418 8663 528 8678
rect 1147 8693 1182 8698
rect 1147 8673 1154 8693
rect 1174 8673 1182 8693
rect 1692 8692 1734 8702
rect 1147 8665 1182 8673
rect 703 8600 735 8607
rect 703 8580 710 8600
rect 731 8580 735 8600
rect 703 8515 735 8580
rect 1073 8515 1113 8516
rect 703 8513 1115 8515
rect 703 8487 1083 8513
rect 1109 8487 1115 8513
rect 703 8479 1115 8487
rect 703 8451 735 8479
rect 1148 8459 1182 8665
rect 1356 8663 1467 8685
rect 1356 8643 1364 8663
rect 1383 8643 1441 8663
rect 1460 8643 1467 8663
rect 1356 8626 1467 8643
rect 1692 8670 1699 8692
rect 1725 8670 1734 8692
rect 1692 8661 1734 8670
rect 909 8456 952 8458
rect 703 8431 708 8451
rect 729 8431 735 8451
rect 703 8424 735 8431
rect 908 8449 952 8456
rect 908 8429 918 8449
rect 941 8429 952 8449
rect 908 8425 952 8429
rect 1126 8454 1182 8459
rect 1126 8434 1133 8454
rect 1153 8434 1182 8454
rect 1126 8427 1182 8434
rect 1238 8595 1271 8596
rect 1692 8595 1729 8661
rect 1238 8566 1729 8595
rect 1126 8426 1161 8427
rect 417 8353 528 8375
rect 417 8333 425 8353
rect 444 8333 502 8353
rect 521 8333 528 8353
rect 417 8316 528 8333
rect 908 8344 950 8425
rect 1238 8346 1271 8566
rect 1692 8564 1729 8566
rect 1498 8426 1608 8440
rect 1498 8423 1576 8426
rect 1498 8396 1502 8423
rect 1531 8399 1576 8423
rect 1605 8399 1608 8426
rect 1531 8396 1608 8399
rect 1498 8381 1608 8396
rect 1852 8407 1890 8745
rect 2065 8764 2121 8769
rect 2065 8744 2072 8764
rect 2092 8744 2121 8764
rect 2065 8737 2121 8744
rect 2808 8924 2864 8931
rect 2808 8904 2837 8924
rect 2857 8904 2864 8924
rect 2808 8899 2864 8904
rect 3255 8927 3287 8934
rect 3255 8907 3261 8927
rect 3282 8907 3287 8927
rect 3747 8918 3781 8970
rect 4401 8960 4404 8987
rect 4433 8963 4478 8987
rect 4507 8963 4511 8990
rect 4433 8960 4511 8963
rect 4401 8946 4511 8960
rect 4697 8990 4739 9000
rect 4697 8971 4705 8990
rect 4730 8971 4739 8990
rect 5975 8973 6006 9019
rect 4697 8918 4739 8971
rect 5474 8948 5585 8970
rect 5474 8928 5482 8948
rect 5501 8928 5559 8948
rect 5578 8928 5585 8948
rect 5974 8956 6006 8973
rect 6275 8956 6312 9092
rect 6413 9059 6523 9073
rect 6413 9056 6491 9059
rect 6413 9029 6417 9056
rect 6446 9032 6491 9056
rect 6520 9032 6523 9059
rect 7143 9049 7177 9092
rect 6446 9029 6523 9032
rect 6413 9014 6523 9029
rect 7142 9044 7177 9049
rect 8256 9048 8293 9114
rect 8714 9113 8747 9114
rect 8803 9275 8859 9282
rect 8803 9255 8832 9275
rect 8852 9255 8859 9275
rect 8803 9250 8859 9255
rect 9033 9280 9077 9284
rect 9033 9260 9044 9280
rect 9067 9260 9077 9280
rect 9033 9253 9077 9260
rect 9250 9278 9282 9285
rect 9250 9258 9256 9278
rect 9277 9258 9282 9278
rect 9033 9251 9076 9253
rect 7142 9024 7149 9044
rect 7169 9024 7177 9044
rect 7142 9016 7177 9024
rect 5974 8943 6312 8956
rect 2065 8736 2100 8737
rect 2808 8693 2842 8899
rect 3255 8879 3287 8907
rect 3745 8892 4741 8918
rect 5474 8911 5585 8928
rect 5975 8924 6312 8943
rect 6254 8923 6312 8924
rect 6698 8951 6730 8958
rect 6698 8931 6705 8951
rect 6726 8931 6730 8951
rect 2875 8871 3287 8879
rect 2875 8845 2881 8871
rect 2907 8845 3287 8871
rect 2875 8843 3287 8845
rect 2877 8842 2917 8843
rect 3037 8807 3076 8822
rect 3037 8766 3048 8807
rect 3069 8766 3076 8807
rect 2807 8685 2843 8693
rect 2807 8665 2816 8685
rect 2836 8665 2843 8685
rect 2807 8664 2843 8665
rect 2807 8653 2841 8664
rect 3037 8493 3076 8766
rect 3255 8778 3287 8843
rect 6698 8866 6730 8931
rect 7068 8866 7108 8867
rect 6698 8864 7110 8866
rect 6698 8838 7078 8864
rect 7104 8838 7110 8864
rect 6698 8830 7110 8838
rect 3255 8758 3259 8778
rect 3280 8758 3287 8778
rect 3255 8751 3287 8758
rect 3673 8785 3731 8786
rect 3673 8766 4010 8785
rect 4400 8781 4511 8798
rect 5244 8791 6240 8817
rect 6698 8802 6730 8830
rect 3673 8753 4011 8766
rect 3177 8689 3230 8692
rect 3177 8672 3189 8689
rect 3221 8672 3230 8689
rect 3177 8664 3230 8672
rect 3176 8617 3230 8664
rect 3462 8680 3572 8695
rect 3462 8677 3539 8680
rect 3462 8650 3465 8677
rect 3494 8653 3539 8677
rect 3568 8653 3572 8680
rect 3494 8650 3572 8653
rect 3462 8636 3572 8650
rect 3673 8617 3710 8753
rect 3979 8736 4011 8753
rect 4400 8761 4407 8781
rect 4426 8761 4484 8781
rect 4503 8761 4511 8781
rect 4400 8739 4511 8761
rect 5246 8738 5288 8791
rect 3979 8690 4010 8736
rect 5246 8719 5255 8738
rect 5280 8719 5288 8738
rect 5246 8709 5288 8719
rect 5474 8749 5584 8763
rect 5474 8746 5552 8749
rect 5474 8719 5478 8746
rect 5507 8722 5552 8746
rect 5581 8722 5584 8749
rect 6204 8739 6238 8791
rect 6698 8782 6703 8802
rect 6724 8782 6730 8802
rect 6698 8775 6730 8782
rect 6908 8803 6946 8813
rect 7143 8810 7177 9016
rect 8251 9039 8293 9048
rect 8251 9017 8260 9039
rect 8286 9017 8293 9039
rect 8518 9066 8629 9083
rect 8518 9046 8525 9066
rect 8544 9046 8602 9066
rect 8621 9046 8629 9066
rect 8518 9024 8629 9046
rect 8803 9044 8837 9250
rect 9250 9230 9282 9258
rect 8870 9222 9282 9230
rect 8870 9196 8876 9222
rect 8902 9196 9282 9222
rect 8870 9194 9282 9196
rect 8872 9193 8912 9194
rect 9250 9129 9282 9194
rect 9250 9109 9254 9129
rect 9275 9109 9282 9129
rect 9250 9102 9282 9109
rect 8803 9036 8838 9044
rect 8251 9007 8293 9017
rect 8803 9016 8811 9036
rect 8831 9016 8838 9036
rect 8803 9011 8838 9016
rect 9457 9031 9567 9046
rect 9457 9028 9534 9031
rect 8251 9006 8292 9007
rect 7885 8972 7920 8973
rect 6908 8786 6918 8803
rect 6938 8786 6946 8803
rect 6749 8743 6790 8744
rect 5507 8719 5584 8722
rect 5474 8704 5584 8719
rect 6203 8734 6238 8739
rect 6203 8714 6210 8734
rect 6230 8714 6238 8734
rect 6748 8733 6790 8743
rect 6203 8706 6238 8714
rect 3767 8687 3802 8688
rect 3746 8680 3802 8687
rect 3746 8660 3775 8680
rect 3795 8660 3802 8680
rect 3746 8655 3802 8660
rect 3979 8683 4018 8690
rect 3979 8663 3985 8683
rect 4010 8663 4018 8683
rect 3979 8657 4018 8663
rect 4193 8683 4225 8690
rect 4193 8663 4199 8683
rect 4220 8663 4225 8683
rect 3176 8582 3711 8617
rect 3176 8578 3229 8582
rect 3037 8466 3041 8493
rect 3072 8466 3076 8493
rect 3322 8514 3433 8531
rect 3322 8494 3329 8514
rect 3348 8494 3406 8514
rect 3425 8494 3433 8514
rect 3322 8472 3433 8494
rect 3037 8459 3076 8466
rect 3746 8449 3780 8655
rect 4193 8635 4225 8663
rect 3813 8627 4225 8635
rect 3813 8601 3819 8627
rect 3845 8601 4225 8627
rect 3813 8599 4225 8601
rect 3815 8598 3855 8599
rect 4193 8534 4225 8599
rect 5759 8641 5791 8648
rect 5759 8621 5766 8641
rect 5787 8621 5791 8641
rect 5759 8556 5791 8621
rect 6129 8556 6169 8557
rect 5759 8554 6171 8556
rect 4193 8514 4197 8534
rect 4218 8514 4225 8534
rect 4193 8507 4225 8514
rect 4696 8549 4744 8554
rect 4696 8520 4707 8549
rect 4736 8520 4744 8549
rect 3746 8448 3781 8449
rect 3744 8441 3781 8448
rect 2689 8420 2724 8421
rect 2230 8416 2262 8417
rect 1852 8390 1860 8407
rect 1880 8390 1890 8407
rect 1852 8384 1890 8390
rect 2227 8411 2262 8416
rect 2227 8391 2234 8411
rect 2254 8391 2262 8411
rect 2227 8383 2262 8391
rect 1210 8344 1271 8346
rect 908 8315 1271 8344
rect 1783 8318 1815 8325
rect 908 8313 1210 8315
rect 1783 8298 1790 8318
rect 1811 8298 1815 8318
rect 1783 8233 1815 8298
rect 2153 8233 2193 8234
rect 1783 8231 2195 8233
rect 1151 8227 1186 8229
rect 187 8224 1186 8227
rect 186 8200 1186 8224
rect 186 8045 234 8200
rect 420 8159 530 8173
rect 420 8156 498 8159
rect 420 8129 424 8156
rect 453 8132 498 8156
rect 527 8132 530 8159
rect 1151 8149 1186 8200
rect 453 8129 530 8132
rect 420 8114 530 8129
rect 1149 8144 1186 8149
rect 1149 8124 1156 8144
rect 1176 8124 1186 8144
rect 1783 8205 2163 8231
rect 2189 8205 2195 8231
rect 1783 8197 2195 8205
rect 1783 8169 1815 8197
rect 1783 8149 1788 8169
rect 1809 8149 1815 8169
rect 1783 8142 1815 8149
rect 1989 8168 2031 8179
rect 2228 8177 2262 8383
rect 2666 8413 2724 8420
rect 2666 8393 2697 8413
rect 2717 8393 2724 8413
rect 2666 8388 2724 8393
rect 3115 8416 3147 8423
rect 3115 8396 3121 8416
rect 3142 8396 3147 8416
rect 2666 8240 2702 8388
rect 3115 8368 3147 8396
rect 2735 8360 3147 8368
rect 2735 8334 2741 8360
rect 2767 8334 3147 8360
rect 3744 8421 3754 8441
rect 3774 8421 3781 8441
rect 3744 8416 3781 8421
rect 4400 8436 4510 8451
rect 4400 8433 4477 8436
rect 3744 8365 3779 8416
rect 4400 8406 4403 8433
rect 4432 8409 4477 8433
rect 4506 8409 4510 8436
rect 4432 8406 4510 8409
rect 4400 8392 4510 8406
rect 4696 8365 4744 8520
rect 5759 8528 6139 8554
rect 6165 8528 6171 8554
rect 5759 8520 6171 8528
rect 5759 8492 5791 8520
rect 6204 8500 6238 8706
rect 6412 8704 6523 8726
rect 6412 8684 6420 8704
rect 6439 8684 6497 8704
rect 6516 8684 6523 8704
rect 6412 8667 6523 8684
rect 6748 8711 6755 8733
rect 6781 8711 6790 8733
rect 6748 8702 6790 8711
rect 5965 8497 6008 8499
rect 5759 8472 5764 8492
rect 5785 8472 5791 8492
rect 5759 8465 5791 8472
rect 5964 8490 6008 8497
rect 5964 8470 5974 8490
rect 5997 8470 6008 8490
rect 5964 8466 6008 8470
rect 6182 8495 6238 8500
rect 6182 8475 6189 8495
rect 6209 8475 6238 8495
rect 6182 8468 6238 8475
rect 6294 8636 6327 8637
rect 6748 8636 6785 8702
rect 6294 8607 6785 8636
rect 6182 8467 6217 8468
rect 3744 8341 4744 8365
rect 5473 8394 5584 8416
rect 5473 8374 5481 8394
rect 5500 8374 5558 8394
rect 5577 8374 5584 8394
rect 5473 8357 5584 8374
rect 5964 8385 6006 8466
rect 6294 8387 6327 8607
rect 6748 8605 6785 8607
rect 6554 8467 6664 8481
rect 6554 8464 6632 8467
rect 6554 8437 6558 8464
rect 6587 8440 6632 8464
rect 6661 8440 6664 8467
rect 6587 8437 6664 8440
rect 6554 8422 6664 8437
rect 6908 8448 6946 8786
rect 7121 8805 7177 8810
rect 7121 8785 7128 8805
rect 7148 8785 7177 8805
rect 7121 8778 7177 8785
rect 7864 8965 7920 8972
rect 7864 8945 7893 8965
rect 7913 8945 7920 8965
rect 7864 8940 7920 8945
rect 8311 8968 8343 8975
rect 8311 8948 8317 8968
rect 8338 8948 8343 8968
rect 8803 8959 8837 9011
rect 9457 9001 9460 9028
rect 9489 9004 9534 9028
rect 9563 9004 9567 9031
rect 9489 9001 9567 9004
rect 9457 8987 9567 9001
rect 9753 9031 9795 9041
rect 9753 9012 9761 9031
rect 9786 9012 9795 9031
rect 9753 8959 9795 9012
rect 7121 8777 7156 8778
rect 7864 8734 7898 8940
rect 8311 8920 8343 8948
rect 8801 8933 9797 8959
rect 7931 8912 8343 8920
rect 7931 8886 7937 8912
rect 7963 8886 8343 8912
rect 7931 8884 8343 8886
rect 7933 8883 7973 8884
rect 8093 8848 8132 8863
rect 8093 8807 8104 8848
rect 8125 8807 8132 8848
rect 7863 8726 7899 8734
rect 7863 8706 7872 8726
rect 7892 8706 7899 8726
rect 7863 8705 7899 8706
rect 7863 8694 7897 8705
rect 8093 8534 8132 8807
rect 8311 8819 8343 8884
rect 8311 8799 8315 8819
rect 8336 8799 8343 8819
rect 8311 8792 8343 8799
rect 8729 8826 8787 8827
rect 8729 8807 9066 8826
rect 9456 8822 9567 8839
rect 8729 8794 9067 8807
rect 8233 8730 8286 8733
rect 8233 8713 8245 8730
rect 8277 8713 8286 8730
rect 8233 8705 8286 8713
rect 8232 8658 8286 8705
rect 8518 8721 8628 8736
rect 8518 8718 8595 8721
rect 8518 8691 8521 8718
rect 8550 8694 8595 8718
rect 8624 8694 8628 8721
rect 8550 8691 8628 8694
rect 8518 8677 8628 8691
rect 8729 8658 8766 8794
rect 9035 8777 9067 8794
rect 9456 8802 9463 8822
rect 9482 8802 9540 8822
rect 9559 8802 9567 8822
rect 9456 8780 9567 8802
rect 9035 8731 9066 8777
rect 8823 8728 8858 8729
rect 8802 8721 8858 8728
rect 8802 8701 8831 8721
rect 8851 8701 8858 8721
rect 8802 8696 8858 8701
rect 9035 8724 9074 8731
rect 9035 8704 9041 8724
rect 9066 8704 9074 8724
rect 9035 8698 9074 8704
rect 9249 8724 9281 8731
rect 9249 8704 9255 8724
rect 9276 8704 9281 8724
rect 8232 8623 8767 8658
rect 8232 8619 8285 8623
rect 8093 8507 8097 8534
rect 8128 8507 8132 8534
rect 8378 8555 8489 8572
rect 8378 8535 8385 8555
rect 8404 8535 8462 8555
rect 8481 8535 8489 8555
rect 8378 8513 8489 8535
rect 8093 8500 8132 8507
rect 8802 8490 8836 8696
rect 9249 8676 9281 8704
rect 8869 8668 9281 8676
rect 8869 8642 8875 8668
rect 8901 8642 9281 8668
rect 8869 8640 9281 8642
rect 8871 8639 8911 8640
rect 9249 8575 9281 8640
rect 9249 8555 9253 8575
rect 9274 8555 9281 8575
rect 9249 8548 9281 8555
rect 9752 8590 9800 8595
rect 9752 8561 9763 8590
rect 9792 8561 9800 8590
rect 8802 8489 8837 8490
rect 8800 8482 8837 8489
rect 7745 8461 7780 8462
rect 7286 8457 7318 8458
rect 6908 8431 6916 8448
rect 6936 8431 6946 8448
rect 6908 8425 6946 8431
rect 7283 8452 7318 8457
rect 7283 8432 7290 8452
rect 7310 8432 7318 8452
rect 7283 8424 7318 8432
rect 6266 8385 6327 8387
rect 5964 8356 6327 8385
rect 6839 8359 6871 8366
rect 5964 8354 6266 8356
rect 3744 8338 4743 8341
rect 6839 8339 6846 8359
rect 6867 8339 6871 8359
rect 3744 8336 3779 8338
rect 2735 8332 3147 8334
rect 2737 8331 2777 8332
rect 1989 8147 1996 8168
rect 2023 8147 2031 8168
rect 1149 8117 1186 8124
rect 1149 8116 1184 8117
rect 186 8016 194 8045
rect 223 8016 234 8045
rect 186 8011 234 8016
rect 705 8051 737 8058
rect 705 8031 712 8051
rect 733 8031 737 8051
rect 705 7966 737 8031
rect 1075 7966 1115 7967
rect 705 7964 1117 7966
rect 705 7938 1085 7964
rect 1111 7938 1117 7964
rect 705 7930 1117 7938
rect 705 7902 737 7930
rect 1150 7910 1184 8116
rect 1854 8099 1893 8106
rect 1497 8071 1608 8093
rect 1497 8051 1505 8071
rect 1524 8051 1582 8071
rect 1601 8051 1608 8071
rect 1497 8034 1608 8051
rect 1854 8072 1858 8099
rect 1889 8072 1893 8099
rect 1701 7983 1754 7987
rect 1219 7948 1754 7983
rect 705 7882 710 7902
rect 731 7882 737 7902
rect 705 7875 737 7882
rect 912 7902 951 7908
rect 912 7882 920 7902
rect 945 7882 951 7902
rect 912 7875 951 7882
rect 1128 7905 1184 7910
rect 1128 7885 1135 7905
rect 1155 7885 1184 7905
rect 1128 7878 1184 7885
rect 1128 7877 1163 7878
rect 920 7829 951 7875
rect 419 7804 530 7826
rect 419 7784 427 7804
rect 446 7784 504 7804
rect 523 7784 530 7804
rect 919 7812 951 7829
rect 1220 7812 1257 7948
rect 1358 7915 1468 7929
rect 1358 7912 1436 7915
rect 1358 7885 1362 7912
rect 1391 7888 1436 7912
rect 1465 7888 1468 7915
rect 1391 7885 1468 7888
rect 1358 7870 1468 7885
rect 1700 7901 1754 7948
rect 1700 7893 1753 7901
rect 1700 7876 1709 7893
rect 1741 7876 1753 7893
rect 1700 7873 1753 7876
rect 919 7799 1257 7812
rect 419 7767 530 7784
rect 920 7780 1257 7799
rect 1199 7779 1257 7780
rect 1643 7807 1675 7814
rect 1643 7787 1650 7807
rect 1671 7787 1675 7807
rect 1643 7722 1675 7787
rect 1854 7799 1893 8072
rect 1989 7976 2031 8147
rect 2206 8172 2262 8177
rect 2206 8152 2213 8172
rect 2233 8152 2262 8172
rect 2206 8145 2262 8152
rect 2669 8182 2702 8240
rect 2899 8292 2937 8302
rect 2899 8254 2908 8292
rect 2931 8254 2937 8292
rect 2669 8174 2703 8182
rect 2669 8154 2676 8174
rect 2696 8154 2703 8174
rect 2669 8149 2703 8154
rect 2669 8148 2700 8149
rect 2206 8144 2241 8145
rect 2899 8118 2937 8254
rect 3115 8267 3147 8332
rect 6839 8274 6871 8339
rect 7209 8274 7249 8275
rect 6839 8272 7251 8274
rect 6207 8268 6242 8270
rect 3115 8247 3119 8267
rect 3140 8247 3147 8267
rect 5243 8265 6242 8268
rect 3720 8250 4022 8252
rect 3115 8240 3147 8247
rect 3659 8221 4022 8250
rect 3659 8219 3720 8221
rect 3040 8175 3078 8181
rect 3040 8158 3050 8175
rect 3070 8158 3078 8175
rect 1989 7942 2233 7976
rect 2899 7964 2943 8118
rect 2736 7962 2943 7964
rect 2196 7934 2233 7942
rect 2089 7901 2123 7912
rect 2087 7900 2123 7901
rect 2087 7880 2094 7900
rect 2114 7880 2123 7900
rect 2087 7872 2123 7880
rect 1854 7758 1861 7799
rect 1882 7758 1893 7799
rect 1854 7743 1893 7758
rect 2013 7722 2053 7723
rect 1643 7720 2055 7722
rect 1643 7694 2023 7720
rect 2049 7694 2055 7720
rect 1643 7686 2055 7694
rect 189 7647 1185 7673
rect 1643 7658 1675 7686
rect 2088 7666 2122 7872
rect 191 7594 233 7647
rect 191 7575 200 7594
rect 225 7575 233 7594
rect 191 7565 233 7575
rect 419 7605 529 7619
rect 419 7602 497 7605
rect 419 7575 423 7602
rect 452 7578 497 7602
rect 526 7578 529 7605
rect 1149 7595 1183 7647
rect 1643 7638 1648 7658
rect 1669 7638 1675 7658
rect 1643 7631 1675 7638
rect 2066 7661 2122 7666
rect 2066 7641 2073 7661
rect 2093 7641 2122 7661
rect 2066 7634 2122 7641
rect 2066 7633 2101 7634
rect 1694 7599 1735 7600
rect 452 7575 529 7578
rect 419 7560 529 7575
rect 1148 7590 1183 7595
rect 1148 7570 1155 7590
rect 1175 7570 1183 7590
rect 1693 7589 1735 7599
rect 1148 7562 1183 7570
rect 704 7497 736 7504
rect 704 7477 711 7497
rect 732 7477 736 7497
rect 704 7412 736 7477
rect 1074 7412 1114 7413
rect 704 7410 1116 7412
rect 704 7384 1084 7410
rect 1110 7384 1116 7410
rect 704 7376 1116 7384
rect 704 7348 736 7376
rect 1149 7356 1183 7562
rect 1357 7560 1468 7582
rect 1357 7540 1365 7560
rect 1384 7540 1442 7560
rect 1461 7540 1468 7560
rect 1357 7523 1468 7540
rect 1693 7567 1700 7589
rect 1726 7567 1735 7589
rect 1693 7558 1735 7567
rect 910 7353 953 7355
rect 704 7328 709 7348
rect 730 7328 736 7348
rect 704 7321 736 7328
rect 909 7346 953 7353
rect 909 7326 919 7346
rect 942 7326 953 7346
rect 909 7322 953 7326
rect 1127 7351 1183 7356
rect 1127 7331 1134 7351
rect 1154 7331 1183 7351
rect 1127 7324 1183 7331
rect 1239 7492 1272 7493
rect 1693 7492 1730 7558
rect 1239 7463 1730 7492
rect 1127 7323 1162 7324
rect 418 7250 529 7272
rect 418 7230 426 7250
rect 445 7230 503 7250
rect 522 7230 529 7250
rect 418 7214 529 7230
rect 909 7241 951 7322
rect 1239 7243 1272 7463
rect 1693 7461 1730 7463
rect 1468 7336 1578 7350
rect 1468 7333 1546 7336
rect 1468 7306 1472 7333
rect 1501 7309 1546 7333
rect 1575 7309 1578 7336
rect 1501 7306 1578 7309
rect 1468 7291 1578 7306
rect 2196 7321 2234 7934
rect 2712 7929 2943 7962
rect 2712 7388 2762 7929
rect 2899 7925 2943 7929
rect 2830 7828 2865 7829
rect 2809 7821 2865 7828
rect 2809 7801 2838 7821
rect 2858 7801 2865 7821
rect 2809 7796 2865 7801
rect 3040 7820 3078 8158
rect 3322 8169 3432 8184
rect 3322 8166 3399 8169
rect 3322 8139 3325 8166
rect 3354 8142 3399 8166
rect 3428 8142 3432 8169
rect 3354 8139 3432 8142
rect 3322 8125 3432 8139
rect 3201 7999 3238 8001
rect 3659 7999 3692 8219
rect 3980 8140 4022 8221
rect 4402 8232 4513 8249
rect 4402 8212 4409 8232
rect 4428 8212 4486 8232
rect 4505 8212 4513 8232
rect 4402 8190 4513 8212
rect 5242 8241 6242 8265
rect 3769 8138 3804 8139
rect 3201 7970 3692 7999
rect 3201 7904 3238 7970
rect 3659 7969 3692 7970
rect 3748 8131 3804 8138
rect 3748 8111 3777 8131
rect 3797 8111 3804 8131
rect 3748 8106 3804 8111
rect 3978 8136 4022 8140
rect 3978 8116 3989 8136
rect 4012 8116 4022 8136
rect 3978 8109 4022 8116
rect 4195 8134 4227 8141
rect 4195 8114 4201 8134
rect 4222 8114 4227 8134
rect 3978 8107 4021 8109
rect 3196 7895 3238 7904
rect 3196 7873 3205 7895
rect 3231 7873 3238 7895
rect 3463 7922 3574 7939
rect 3463 7902 3470 7922
rect 3489 7902 3547 7922
rect 3566 7902 3574 7922
rect 3463 7880 3574 7902
rect 3748 7900 3782 8106
rect 4195 8086 4227 8114
rect 3815 8078 4227 8086
rect 3815 8052 3821 8078
rect 3847 8052 4227 8078
rect 5242 8086 5290 8241
rect 5476 8200 5586 8214
rect 5476 8197 5554 8200
rect 5476 8170 5480 8197
rect 5509 8173 5554 8197
rect 5583 8173 5586 8200
rect 6207 8190 6242 8241
rect 5509 8170 5586 8173
rect 5476 8155 5586 8170
rect 6205 8185 6242 8190
rect 6205 8165 6212 8185
rect 6232 8165 6242 8185
rect 6839 8246 7219 8272
rect 7245 8246 7251 8272
rect 6839 8238 7251 8246
rect 6839 8210 6871 8238
rect 6839 8190 6844 8210
rect 6865 8190 6871 8210
rect 6839 8183 6871 8190
rect 7045 8209 7087 8220
rect 7284 8218 7318 8424
rect 7722 8454 7780 8461
rect 7722 8434 7753 8454
rect 7773 8434 7780 8454
rect 7722 8429 7780 8434
rect 8171 8457 8203 8464
rect 8171 8437 8177 8457
rect 8198 8437 8203 8457
rect 7722 8281 7758 8429
rect 8171 8409 8203 8437
rect 7791 8401 8203 8409
rect 7791 8375 7797 8401
rect 7823 8375 8203 8401
rect 8800 8462 8810 8482
rect 8830 8462 8837 8482
rect 8800 8457 8837 8462
rect 9456 8477 9566 8492
rect 9456 8474 9533 8477
rect 8800 8406 8835 8457
rect 9456 8447 9459 8474
rect 9488 8450 9533 8474
rect 9562 8450 9566 8477
rect 9488 8447 9566 8450
rect 9456 8433 9566 8447
rect 9752 8406 9800 8561
rect 8800 8382 9800 8406
rect 8800 8379 9799 8382
rect 8800 8377 8835 8379
rect 7791 8373 8203 8375
rect 7793 8372 7833 8373
rect 7045 8188 7052 8209
rect 7079 8188 7087 8209
rect 6205 8158 6242 8165
rect 6205 8157 6240 8158
rect 5242 8057 5250 8086
rect 5279 8057 5290 8086
rect 5242 8052 5290 8057
rect 5761 8092 5793 8099
rect 5761 8072 5768 8092
rect 5789 8072 5793 8092
rect 3815 8050 4227 8052
rect 3817 8049 3857 8050
rect 4195 7985 4227 8050
rect 4195 7965 4199 7985
rect 4220 7965 4227 7985
rect 4195 7958 4227 7965
rect 5761 8007 5793 8072
rect 6131 8007 6171 8008
rect 5761 8005 6173 8007
rect 5761 7979 6141 8005
rect 6167 7979 6173 8005
rect 5761 7971 6173 7979
rect 5761 7943 5793 7971
rect 6206 7951 6240 8157
rect 6910 8140 6949 8147
rect 6553 8112 6664 8134
rect 6553 8092 6561 8112
rect 6580 8092 6638 8112
rect 6657 8092 6664 8112
rect 6553 8075 6664 8092
rect 6910 8113 6914 8140
rect 6945 8113 6949 8140
rect 6757 8024 6810 8028
rect 6275 7989 6810 8024
rect 5761 7923 5766 7943
rect 5787 7923 5793 7943
rect 5761 7916 5793 7923
rect 5968 7943 6007 7949
rect 5968 7923 5976 7943
rect 6001 7923 6007 7943
rect 5968 7916 6007 7923
rect 6184 7946 6240 7951
rect 6184 7926 6191 7946
rect 6211 7926 6240 7946
rect 6184 7919 6240 7926
rect 6184 7918 6219 7919
rect 3748 7892 3783 7900
rect 3196 7863 3238 7873
rect 3748 7872 3756 7892
rect 3776 7872 3783 7892
rect 3748 7867 3783 7872
rect 4402 7887 4512 7902
rect 4402 7884 4479 7887
rect 3196 7862 3237 7863
rect 3040 7803 3048 7820
rect 3068 7803 3078 7820
rect 2809 7590 2843 7796
rect 3040 7793 3078 7803
rect 3256 7824 3288 7831
rect 3256 7804 3262 7824
rect 3283 7804 3288 7824
rect 3748 7815 3782 7867
rect 4402 7857 4405 7884
rect 4434 7860 4479 7884
rect 4508 7860 4512 7887
rect 4434 7857 4512 7860
rect 4402 7843 4512 7857
rect 4698 7887 4740 7897
rect 4698 7868 4706 7887
rect 4731 7868 4740 7887
rect 5976 7870 6007 7916
rect 4698 7815 4740 7868
rect 5475 7845 5586 7867
rect 5475 7825 5483 7845
rect 5502 7825 5560 7845
rect 5579 7825 5586 7845
rect 5975 7853 6007 7870
rect 6276 7853 6313 7989
rect 6414 7956 6524 7970
rect 6414 7953 6492 7956
rect 6414 7926 6418 7953
rect 6447 7929 6492 7953
rect 6521 7929 6524 7956
rect 6447 7926 6524 7929
rect 6414 7911 6524 7926
rect 6756 7942 6810 7989
rect 6756 7934 6809 7942
rect 6756 7917 6765 7934
rect 6797 7917 6809 7934
rect 6756 7914 6809 7917
rect 5975 7840 6313 7853
rect 3256 7776 3288 7804
rect 3746 7789 4742 7815
rect 5475 7808 5586 7825
rect 5976 7821 6313 7840
rect 6255 7820 6313 7821
rect 6699 7848 6731 7855
rect 6699 7828 6706 7848
rect 6727 7828 6731 7848
rect 2876 7768 3288 7776
rect 2876 7742 2882 7768
rect 2908 7742 3288 7768
rect 2876 7740 3288 7742
rect 2878 7739 2918 7740
rect 3256 7675 3288 7740
rect 6699 7763 6731 7828
rect 6910 7840 6949 8113
rect 7045 8017 7087 8188
rect 7262 8213 7318 8218
rect 7262 8193 7269 8213
rect 7289 8193 7318 8213
rect 7262 8186 7318 8193
rect 7725 8223 7758 8281
rect 7955 8333 7993 8343
rect 7955 8295 7964 8333
rect 7987 8295 7993 8333
rect 7725 8215 7759 8223
rect 7725 8195 7732 8215
rect 7752 8195 7759 8215
rect 7725 8190 7759 8195
rect 7725 8189 7756 8190
rect 7262 8185 7297 8186
rect 7955 8159 7993 8295
rect 8171 8308 8203 8373
rect 8171 8288 8175 8308
rect 8196 8288 8203 8308
rect 8776 8291 9078 8293
rect 8171 8281 8203 8288
rect 8715 8262 9078 8291
rect 8715 8260 8776 8262
rect 8096 8216 8134 8222
rect 8096 8199 8106 8216
rect 8126 8199 8134 8216
rect 7045 7983 7289 8017
rect 7955 8005 7999 8159
rect 7792 8003 7999 8005
rect 7252 7975 7289 7983
rect 7145 7942 7179 7953
rect 7143 7941 7179 7942
rect 7143 7921 7150 7941
rect 7170 7921 7179 7941
rect 7143 7913 7179 7921
rect 6910 7799 6917 7840
rect 6938 7799 6949 7840
rect 6910 7784 6949 7799
rect 7069 7763 7109 7764
rect 6699 7761 7111 7763
rect 6699 7735 7079 7761
rect 7105 7735 7111 7761
rect 6699 7727 7111 7735
rect 3256 7655 3260 7675
rect 3281 7655 3288 7675
rect 3256 7648 3288 7655
rect 3674 7682 3732 7683
rect 3674 7663 4011 7682
rect 4401 7678 4512 7695
rect 5245 7688 6241 7714
rect 6699 7699 6731 7727
rect 7144 7707 7178 7913
rect 3674 7650 4012 7663
rect 2809 7582 2844 7590
rect 2809 7562 2817 7582
rect 2837 7562 2844 7582
rect 2809 7557 2844 7562
rect 3463 7577 3573 7592
rect 3463 7574 3540 7577
rect 2809 7514 2843 7557
rect 3463 7547 3466 7574
rect 3495 7550 3540 7574
rect 3569 7550 3573 7577
rect 3495 7547 3573 7550
rect 3463 7533 3573 7547
rect 3674 7514 3711 7650
rect 3980 7633 4012 7650
rect 4401 7658 4408 7678
rect 4427 7658 4485 7678
rect 4504 7658 4512 7678
rect 4401 7636 4512 7658
rect 5247 7635 5289 7688
rect 3980 7587 4011 7633
rect 5247 7616 5256 7635
rect 5281 7616 5289 7635
rect 5247 7606 5289 7616
rect 5475 7646 5585 7660
rect 5475 7643 5553 7646
rect 5475 7616 5479 7643
rect 5508 7619 5553 7643
rect 5582 7619 5585 7646
rect 6205 7636 6239 7688
rect 6699 7679 6704 7699
rect 6725 7679 6731 7699
rect 6699 7672 6731 7679
rect 7122 7702 7178 7707
rect 7122 7682 7129 7702
rect 7149 7682 7178 7702
rect 7122 7675 7178 7682
rect 7122 7674 7157 7675
rect 6750 7640 6791 7641
rect 5508 7616 5585 7619
rect 5475 7601 5585 7616
rect 6204 7631 6239 7636
rect 6204 7611 6211 7631
rect 6231 7611 6239 7631
rect 6749 7630 6791 7640
rect 6204 7603 6239 7611
rect 3768 7584 3803 7585
rect 3747 7577 3803 7584
rect 3747 7557 3776 7577
rect 3796 7557 3803 7577
rect 3747 7552 3803 7557
rect 3980 7580 4019 7587
rect 3980 7560 3986 7580
rect 4011 7560 4019 7580
rect 3980 7554 4019 7560
rect 4194 7580 4226 7587
rect 4194 7560 4200 7580
rect 4221 7560 4226 7580
rect 2808 7479 3712 7514
rect 2809 7478 2843 7479
rect 2690 7379 2762 7388
rect 2690 7350 2707 7379
rect 2755 7350 2762 7379
rect 3353 7398 3464 7415
rect 3353 7378 3360 7398
rect 3379 7378 3437 7398
rect 3456 7378 3464 7398
rect 3353 7356 3464 7378
rect 2690 7343 2762 7350
rect 3747 7346 3781 7552
rect 4194 7532 4226 7560
rect 3814 7524 4226 7532
rect 3814 7498 3820 7524
rect 3846 7498 4226 7524
rect 3814 7496 4226 7498
rect 3816 7495 3856 7496
rect 4194 7431 4226 7496
rect 5760 7538 5792 7545
rect 5760 7518 5767 7538
rect 5788 7518 5792 7538
rect 5760 7453 5792 7518
rect 6130 7453 6170 7454
rect 5760 7451 6172 7453
rect 4194 7411 4198 7431
rect 4219 7411 4226 7431
rect 4194 7404 4226 7411
rect 4697 7446 4745 7451
rect 4697 7417 4708 7446
rect 4737 7417 4745 7446
rect 3747 7345 3782 7346
rect 2690 7333 2760 7343
rect 3745 7338 3782 7345
rect 2196 7301 2204 7321
rect 2224 7301 2234 7321
rect 3745 7318 3755 7338
rect 3775 7318 3782 7338
rect 3745 7313 3782 7318
rect 4401 7333 4511 7348
rect 4401 7330 4478 7333
rect 2720 7304 2755 7305
rect 2196 7294 2234 7301
rect 2699 7297 2755 7304
rect 2197 7293 2232 7294
rect 1211 7241 1272 7243
rect 909 7212 1272 7241
rect 1753 7228 1785 7235
rect 909 7210 1211 7212
rect 1753 7208 1760 7228
rect 1781 7208 1785 7228
rect 1753 7143 1785 7208
rect 2123 7143 2163 7144
rect 1753 7141 2165 7143
rect 1151 7124 1186 7126
rect 187 7121 1186 7124
rect 186 7097 1186 7121
rect 186 6942 234 7097
rect 420 7056 530 7070
rect 420 7053 498 7056
rect 420 7026 424 7053
rect 453 7029 498 7053
rect 527 7029 530 7056
rect 1151 7046 1186 7097
rect 1753 7115 2133 7141
rect 2159 7115 2165 7141
rect 1753 7107 2165 7115
rect 1753 7079 1785 7107
rect 1753 7059 1758 7079
rect 1779 7059 1785 7079
rect 1753 7052 1785 7059
rect 1959 7078 2004 7090
rect 2198 7087 2232 7293
rect 1959 7059 1966 7078
rect 1995 7059 2004 7078
rect 453 7026 530 7029
rect 420 7011 530 7026
rect 1149 7041 1186 7046
rect 1149 7021 1156 7041
rect 1176 7021 1186 7041
rect 1149 7014 1186 7021
rect 1149 7013 1184 7014
rect 186 6913 194 6942
rect 223 6913 234 6942
rect 186 6908 234 6913
rect 705 6948 737 6955
rect 705 6928 712 6948
rect 733 6928 737 6948
rect 705 6863 737 6928
rect 1075 6863 1115 6864
rect 705 6861 1117 6863
rect 705 6835 1085 6861
rect 1111 6835 1117 6861
rect 705 6827 1117 6835
rect 705 6799 737 6827
rect 1150 6807 1184 7013
rect 1467 6981 1578 7003
rect 1467 6961 1475 6981
rect 1494 6961 1552 6981
rect 1571 6961 1578 6981
rect 1467 6944 1578 6961
rect 1959 6976 2004 7059
rect 2176 7082 2232 7087
rect 2176 7062 2183 7082
rect 2203 7062 2232 7082
rect 2699 7277 2728 7297
rect 2748 7277 2755 7297
rect 2699 7272 2755 7277
rect 3146 7300 3178 7307
rect 3146 7280 3152 7300
rect 3173 7280 3178 7300
rect 2699 7066 2733 7272
rect 3146 7252 3178 7280
rect 2766 7244 3178 7252
rect 2766 7218 2772 7244
rect 2798 7218 3178 7244
rect 3745 7262 3780 7313
rect 4401 7303 4404 7330
rect 4433 7306 4478 7330
rect 4507 7306 4511 7333
rect 4433 7303 4511 7306
rect 4401 7289 4511 7303
rect 4697 7262 4745 7417
rect 5760 7425 6140 7451
rect 6166 7425 6172 7451
rect 5760 7417 6172 7425
rect 5760 7389 5792 7417
rect 6205 7397 6239 7603
rect 6413 7601 6524 7623
rect 6413 7581 6421 7601
rect 6440 7581 6498 7601
rect 6517 7581 6524 7601
rect 6413 7564 6524 7581
rect 6749 7608 6756 7630
rect 6782 7608 6791 7630
rect 6749 7599 6791 7608
rect 5966 7394 6009 7396
rect 5760 7369 5765 7389
rect 5786 7369 5792 7389
rect 5760 7362 5792 7369
rect 5965 7387 6009 7394
rect 5965 7367 5975 7387
rect 5998 7367 6009 7387
rect 5965 7363 6009 7367
rect 6183 7392 6239 7397
rect 6183 7372 6190 7392
rect 6210 7372 6239 7392
rect 6183 7365 6239 7372
rect 6295 7533 6328 7534
rect 6749 7533 6786 7599
rect 6295 7504 6786 7533
rect 6183 7364 6218 7365
rect 3745 7238 4745 7262
rect 5474 7291 5585 7313
rect 5474 7271 5482 7291
rect 5501 7271 5559 7291
rect 5578 7271 5585 7291
rect 5474 7255 5585 7271
rect 5965 7282 6007 7363
rect 6295 7284 6328 7504
rect 6749 7502 6786 7504
rect 6524 7377 6634 7391
rect 6524 7374 6602 7377
rect 6524 7347 6528 7374
rect 6557 7350 6602 7374
rect 6631 7350 6634 7377
rect 6557 7347 6634 7350
rect 6524 7332 6634 7347
rect 7252 7362 7290 7975
rect 7768 7970 7999 8003
rect 7768 7429 7818 7970
rect 7955 7966 7999 7970
rect 7886 7869 7921 7870
rect 7865 7862 7921 7869
rect 7865 7842 7894 7862
rect 7914 7842 7921 7862
rect 7865 7837 7921 7842
rect 8096 7861 8134 8199
rect 8378 8210 8488 8225
rect 8378 8207 8455 8210
rect 8378 8180 8381 8207
rect 8410 8183 8455 8207
rect 8484 8183 8488 8210
rect 8410 8180 8488 8183
rect 8378 8166 8488 8180
rect 8257 8040 8294 8042
rect 8715 8040 8748 8260
rect 9036 8181 9078 8262
rect 9458 8273 9569 8290
rect 9458 8253 9465 8273
rect 9484 8253 9542 8273
rect 9561 8253 9569 8273
rect 9458 8231 9569 8253
rect 8825 8179 8860 8180
rect 8257 8011 8748 8040
rect 8257 7945 8294 8011
rect 8715 8010 8748 8011
rect 8804 8172 8860 8179
rect 8804 8152 8833 8172
rect 8853 8152 8860 8172
rect 8804 8147 8860 8152
rect 9034 8177 9078 8181
rect 9034 8157 9045 8177
rect 9068 8157 9078 8177
rect 9034 8150 9078 8157
rect 9251 8175 9283 8182
rect 9251 8155 9257 8175
rect 9278 8155 9283 8175
rect 9034 8148 9077 8150
rect 8252 7936 8294 7945
rect 8252 7914 8261 7936
rect 8287 7914 8294 7936
rect 8519 7963 8630 7980
rect 8519 7943 8526 7963
rect 8545 7943 8603 7963
rect 8622 7943 8630 7963
rect 8519 7921 8630 7943
rect 8804 7941 8838 8147
rect 9251 8127 9283 8155
rect 8871 8119 9283 8127
rect 8871 8093 8877 8119
rect 8903 8093 9283 8119
rect 8871 8091 9283 8093
rect 8873 8090 8913 8091
rect 9251 8026 9283 8091
rect 9251 8006 9255 8026
rect 9276 8006 9283 8026
rect 9251 7999 9283 8006
rect 8804 7933 8839 7941
rect 8252 7904 8294 7914
rect 8804 7913 8812 7933
rect 8832 7913 8839 7933
rect 8804 7908 8839 7913
rect 9458 7928 9568 7943
rect 9458 7925 9535 7928
rect 8252 7903 8293 7904
rect 8096 7844 8104 7861
rect 8124 7844 8134 7861
rect 7865 7631 7899 7837
rect 8096 7834 8134 7844
rect 8312 7865 8344 7872
rect 8312 7845 8318 7865
rect 8339 7845 8344 7865
rect 8804 7856 8838 7908
rect 9458 7898 9461 7925
rect 9490 7901 9535 7925
rect 9564 7901 9568 7928
rect 9490 7898 9568 7901
rect 9458 7884 9568 7898
rect 9754 7928 9796 7938
rect 9754 7909 9762 7928
rect 9787 7909 9796 7928
rect 9754 7856 9796 7909
rect 8312 7817 8344 7845
rect 8802 7830 9798 7856
rect 7932 7809 8344 7817
rect 7932 7783 7938 7809
rect 7964 7783 8344 7809
rect 7932 7781 8344 7783
rect 7934 7780 7974 7781
rect 8312 7716 8344 7781
rect 8312 7696 8316 7716
rect 8337 7696 8344 7716
rect 8312 7689 8344 7696
rect 8730 7723 8788 7724
rect 8730 7704 9067 7723
rect 9457 7719 9568 7736
rect 8730 7691 9068 7704
rect 7865 7623 7900 7631
rect 7865 7603 7873 7623
rect 7893 7603 7900 7623
rect 7865 7598 7900 7603
rect 8519 7618 8629 7633
rect 8519 7615 8596 7618
rect 7865 7555 7899 7598
rect 8519 7588 8522 7615
rect 8551 7591 8596 7615
rect 8625 7591 8629 7618
rect 8551 7588 8629 7591
rect 8519 7574 8629 7588
rect 8730 7555 8767 7691
rect 9036 7674 9068 7691
rect 9457 7699 9464 7719
rect 9483 7699 9541 7719
rect 9560 7699 9568 7719
rect 9457 7677 9568 7699
rect 9036 7628 9067 7674
rect 8824 7625 8859 7626
rect 8803 7618 8859 7625
rect 8803 7598 8832 7618
rect 8852 7598 8859 7618
rect 8803 7593 8859 7598
rect 9036 7621 9075 7628
rect 9036 7601 9042 7621
rect 9067 7601 9075 7621
rect 9036 7595 9075 7601
rect 9250 7621 9282 7628
rect 9250 7601 9256 7621
rect 9277 7601 9282 7621
rect 7864 7520 8768 7555
rect 7865 7519 7899 7520
rect 7746 7420 7818 7429
rect 7746 7391 7763 7420
rect 7811 7391 7818 7420
rect 8409 7439 8520 7456
rect 8409 7419 8416 7439
rect 8435 7419 8493 7439
rect 8512 7419 8520 7439
rect 8409 7397 8520 7419
rect 7746 7384 7818 7391
rect 8803 7387 8837 7593
rect 9250 7573 9282 7601
rect 8870 7565 9282 7573
rect 8870 7539 8876 7565
rect 8902 7539 9282 7565
rect 8870 7537 9282 7539
rect 8872 7536 8912 7537
rect 9250 7472 9282 7537
rect 9250 7452 9254 7472
rect 9275 7452 9282 7472
rect 9250 7445 9282 7452
rect 9753 7487 9801 7492
rect 9753 7458 9764 7487
rect 9793 7458 9801 7487
rect 8803 7386 8838 7387
rect 7746 7374 7816 7384
rect 8801 7379 8838 7386
rect 7252 7342 7260 7362
rect 7280 7342 7290 7362
rect 8801 7359 8811 7379
rect 8831 7359 8838 7379
rect 8801 7354 8838 7359
rect 9457 7374 9567 7389
rect 9457 7371 9534 7374
rect 7776 7345 7811 7346
rect 7252 7335 7290 7342
rect 7755 7338 7811 7345
rect 7253 7334 7288 7335
rect 6267 7282 6328 7284
rect 5965 7253 6328 7282
rect 6809 7269 6841 7276
rect 5965 7251 6267 7253
rect 6809 7249 6816 7269
rect 6837 7249 6841 7269
rect 3745 7235 4744 7238
rect 3745 7233 3780 7235
rect 2766 7216 3178 7218
rect 2768 7215 2808 7216
rect 2934 7175 2969 7193
rect 2934 7143 2937 7175
rect 2964 7143 2969 7175
rect 2699 7065 2734 7066
rect 2176 7055 2232 7062
rect 2697 7058 2735 7065
rect 2176 7054 2211 7055
rect 2697 7054 2707 7058
rect 2691 7040 2707 7054
rect 2727 7054 2735 7058
rect 2727 7040 2741 7054
rect 2691 7033 2741 7040
rect 2324 6976 2374 6978
rect 1959 6942 2374 6976
rect 2088 6880 2122 6881
rect 1219 6845 2123 6880
rect 2171 6869 2239 6880
rect 2171 6848 2176 6869
rect 705 6779 710 6799
rect 731 6779 737 6799
rect 705 6772 737 6779
rect 912 6799 951 6805
rect 912 6779 920 6799
rect 945 6779 951 6799
rect 912 6772 951 6779
rect 1128 6802 1184 6807
rect 1128 6782 1135 6802
rect 1155 6782 1184 6802
rect 1128 6775 1184 6782
rect 1128 6774 1163 6775
rect 920 6726 951 6772
rect 419 6701 530 6723
rect 419 6681 427 6701
rect 446 6681 504 6701
rect 523 6681 530 6701
rect 919 6709 951 6726
rect 1220 6709 1257 6845
rect 1358 6812 1468 6826
rect 1358 6809 1436 6812
rect 1358 6782 1362 6809
rect 1391 6785 1436 6809
rect 1465 6785 1468 6812
rect 2088 6802 2122 6845
rect 1391 6782 1468 6785
rect 1358 6767 1468 6782
rect 2087 6797 2122 6802
rect 2087 6777 2094 6797
rect 2114 6777 2122 6797
rect 2087 6769 2122 6777
rect 919 6696 1257 6709
rect 419 6664 530 6681
rect 920 6677 1257 6696
rect 1199 6676 1257 6677
rect 1643 6704 1675 6711
rect 1643 6684 1650 6704
rect 1671 6684 1675 6704
rect 1643 6619 1675 6684
rect 2013 6619 2053 6620
rect 1643 6617 2055 6619
rect 1643 6591 2023 6617
rect 2049 6591 2055 6617
rect 1643 6583 2055 6591
rect 189 6544 1185 6570
rect 1643 6555 1675 6583
rect 191 6491 233 6544
rect 191 6472 200 6491
rect 225 6472 233 6491
rect 191 6462 233 6472
rect 419 6502 529 6516
rect 419 6499 497 6502
rect 419 6472 423 6499
rect 452 6475 497 6499
rect 526 6475 529 6502
rect 1149 6492 1183 6544
rect 1643 6535 1648 6555
rect 1669 6535 1675 6555
rect 1643 6528 1675 6535
rect 1853 6556 1891 6566
rect 2088 6563 2122 6769
rect 1853 6539 1863 6556
rect 1883 6539 1891 6556
rect 1694 6496 1735 6497
rect 452 6472 529 6475
rect 419 6457 529 6472
rect 1148 6487 1183 6492
rect 1148 6467 1155 6487
rect 1175 6467 1183 6487
rect 1693 6486 1735 6496
rect 1148 6459 1183 6467
rect 704 6394 736 6401
rect 704 6374 711 6394
rect 732 6374 736 6394
rect 704 6309 736 6374
rect 1074 6309 1114 6310
rect 704 6307 1116 6309
rect 704 6281 1084 6307
rect 1110 6281 1116 6307
rect 704 6273 1116 6281
rect 704 6245 736 6273
rect 1149 6253 1183 6459
rect 1357 6457 1468 6479
rect 1357 6437 1365 6457
rect 1384 6437 1442 6457
rect 1461 6437 1468 6457
rect 1357 6420 1468 6437
rect 1693 6464 1700 6486
rect 1726 6464 1735 6486
rect 1693 6455 1735 6464
rect 910 6250 953 6252
rect 704 6225 709 6245
rect 730 6225 736 6245
rect 704 6218 736 6225
rect 909 6243 953 6250
rect 909 6223 919 6243
rect 942 6223 953 6243
rect 909 6219 953 6223
rect 1127 6248 1183 6253
rect 1127 6228 1134 6248
rect 1154 6228 1183 6248
rect 1127 6221 1183 6228
rect 1239 6389 1272 6390
rect 1693 6389 1730 6455
rect 1239 6360 1730 6389
rect 1127 6220 1162 6221
rect 418 6147 529 6169
rect 418 6127 426 6147
rect 445 6127 503 6147
rect 522 6127 529 6147
rect 418 6110 529 6127
rect 909 6138 951 6219
rect 1239 6140 1272 6360
rect 1693 6358 1730 6360
rect 1499 6220 1609 6234
rect 1499 6217 1577 6220
rect 1499 6190 1503 6217
rect 1532 6193 1577 6217
rect 1606 6193 1609 6220
rect 1532 6190 1609 6193
rect 1499 6175 1609 6190
rect 1853 6201 1891 6539
rect 2066 6558 2122 6563
rect 2066 6538 2073 6558
rect 2093 6538 2122 6558
rect 2066 6531 2122 6538
rect 2169 6840 2176 6848
rect 2224 6840 2239 6869
rect 2169 6831 2239 6840
rect 2066 6530 2101 6531
rect 1988 6430 2032 6434
rect 2169 6430 2219 6831
rect 2324 6814 2374 6942
rect 2557 6955 2667 6957
rect 2934 6955 2969 7143
rect 3146 7151 3178 7216
rect 6809 7184 6841 7249
rect 7179 7184 7219 7185
rect 6809 7182 7221 7184
rect 6207 7165 6242 7167
rect 5243 7162 6242 7165
rect 3146 7131 3150 7151
rect 3171 7131 3178 7151
rect 3720 7147 4022 7149
rect 3146 7124 3178 7131
rect 3659 7118 4022 7147
rect 3659 7116 3720 7118
rect 2557 6925 2969 6955
rect 2557 6900 2601 6925
rect 2640 6922 2969 6925
rect 3088 7056 3122 7062
rect 3088 7036 3097 7056
rect 3118 7036 3122 7056
rect 1988 6397 2219 6430
rect 1988 6395 2195 6397
rect 1988 6241 2032 6395
rect 1853 6184 1861 6201
rect 1881 6184 1891 6201
rect 1853 6178 1891 6184
rect 1211 6138 1272 6140
rect 909 6109 1272 6138
rect 1784 6112 1816 6119
rect 909 6107 1211 6109
rect 1784 6092 1791 6112
rect 1812 6092 1816 6112
rect 1784 6027 1816 6092
rect 1994 6105 2032 6241
rect 2231 6210 2262 6211
rect 2228 6205 2262 6210
rect 2228 6185 2235 6205
rect 2255 6185 2262 6205
rect 2228 6177 2262 6185
rect 1994 6067 2000 6105
rect 2023 6067 2032 6105
rect 1994 6057 2032 6067
rect 2229 6119 2262 6177
rect 2154 6027 2194 6028
rect 1784 6025 2196 6027
rect 1152 6021 1187 6023
rect 188 6018 1187 6021
rect 187 5994 1187 6018
rect 187 5839 235 5994
rect 421 5953 531 5967
rect 421 5950 499 5953
rect 421 5923 425 5950
rect 454 5926 499 5950
rect 528 5926 531 5953
rect 1152 5943 1187 5994
rect 454 5923 531 5926
rect 421 5908 531 5923
rect 1150 5938 1187 5943
rect 1150 5918 1157 5938
rect 1177 5918 1187 5938
rect 1784 5999 2164 6025
rect 2190 5999 2196 6025
rect 1784 5991 2196 5999
rect 1784 5963 1816 5991
rect 2229 5971 2265 6119
rect 1784 5943 1789 5963
rect 1810 5943 1816 5963
rect 1784 5936 1816 5943
rect 2207 5966 2265 5971
rect 2207 5946 2214 5966
rect 2234 5946 2265 5966
rect 2207 5939 2265 5946
rect 2207 5938 2242 5939
rect 1150 5911 1187 5918
rect 1150 5910 1185 5911
rect 187 5810 195 5839
rect 224 5810 235 5839
rect 187 5805 235 5810
rect 706 5845 738 5852
rect 706 5825 713 5845
rect 734 5825 738 5845
rect 706 5760 738 5825
rect 1076 5760 1116 5761
rect 706 5758 1118 5760
rect 706 5732 1086 5758
rect 1112 5732 1118 5758
rect 706 5724 1118 5732
rect 706 5696 738 5724
rect 1151 5704 1185 5910
rect 1855 5893 1894 5900
rect 1498 5865 1609 5887
rect 1498 5845 1506 5865
rect 1525 5845 1583 5865
rect 1602 5845 1609 5865
rect 1498 5828 1609 5845
rect 1855 5866 1859 5893
rect 1890 5866 1894 5893
rect 1702 5777 1755 5781
rect 1220 5742 1755 5777
rect 706 5676 711 5696
rect 732 5676 738 5696
rect 706 5669 738 5676
rect 913 5696 952 5702
rect 913 5676 921 5696
rect 946 5676 952 5696
rect 913 5669 952 5676
rect 1129 5699 1185 5704
rect 1129 5679 1136 5699
rect 1156 5679 1185 5699
rect 1129 5672 1185 5679
rect 1129 5671 1164 5672
rect 921 5623 952 5669
rect 420 5598 531 5620
rect 420 5578 428 5598
rect 447 5578 505 5598
rect 524 5578 531 5598
rect 920 5606 952 5623
rect 1221 5606 1258 5742
rect 1359 5709 1469 5723
rect 1359 5706 1437 5709
rect 1359 5679 1363 5706
rect 1392 5682 1437 5706
rect 1466 5682 1469 5709
rect 1392 5679 1469 5682
rect 1359 5664 1469 5679
rect 1701 5695 1755 5742
rect 1701 5687 1754 5695
rect 1701 5670 1710 5687
rect 1742 5670 1754 5687
rect 1701 5667 1754 5670
rect 920 5593 1258 5606
rect 420 5561 531 5578
rect 921 5574 1258 5593
rect 1200 5573 1258 5574
rect 1644 5601 1676 5608
rect 1644 5581 1651 5601
rect 1672 5581 1676 5601
rect 1644 5516 1676 5581
rect 1855 5593 1894 5866
rect 2090 5695 2124 5706
rect 2088 5694 2124 5695
rect 2088 5674 2095 5694
rect 2115 5674 2124 5694
rect 2088 5666 2124 5674
rect 1855 5552 1862 5593
rect 1883 5552 1894 5593
rect 1855 5537 1894 5552
rect 2014 5516 2054 5517
rect 1644 5514 2056 5516
rect 1644 5488 2024 5514
rect 2050 5488 2056 5514
rect 1644 5480 2056 5488
rect 190 5441 1186 5467
rect 1644 5452 1676 5480
rect 2089 5460 2123 5666
rect 192 5388 234 5441
rect 192 5369 201 5388
rect 226 5369 234 5388
rect 192 5359 234 5369
rect 420 5399 530 5413
rect 420 5396 498 5399
rect 420 5369 424 5396
rect 453 5372 498 5396
rect 527 5372 530 5399
rect 1150 5389 1184 5441
rect 1644 5432 1649 5452
rect 1670 5432 1676 5452
rect 1644 5425 1676 5432
rect 2067 5455 2123 5460
rect 2067 5435 2074 5455
rect 2094 5435 2123 5455
rect 2067 5428 2123 5435
rect 2067 5427 2102 5428
rect 1695 5393 1736 5394
rect 453 5369 530 5372
rect 420 5354 530 5369
rect 1149 5384 1184 5389
rect 1149 5364 1156 5384
rect 1176 5364 1184 5384
rect 1694 5383 1736 5393
rect 1149 5356 1184 5364
rect 705 5291 737 5298
rect 705 5271 712 5291
rect 733 5271 737 5291
rect 705 5206 737 5271
rect 1075 5206 1115 5207
rect 705 5204 1117 5206
rect 705 5178 1085 5204
rect 1111 5178 1117 5204
rect 705 5170 1117 5178
rect 705 5142 737 5170
rect 1150 5150 1184 5356
rect 1358 5354 1469 5376
rect 1358 5334 1366 5354
rect 1385 5334 1443 5354
rect 1462 5334 1469 5354
rect 1358 5317 1469 5334
rect 1694 5361 1701 5383
rect 1727 5361 1736 5383
rect 1694 5352 1736 5361
rect 911 5147 954 5149
rect 705 5122 710 5142
rect 731 5122 737 5142
rect 705 5115 737 5122
rect 910 5140 954 5147
rect 910 5120 920 5140
rect 943 5120 954 5140
rect 910 5116 954 5120
rect 1128 5145 1184 5150
rect 1128 5125 1135 5145
rect 1155 5125 1184 5145
rect 1128 5118 1184 5125
rect 1240 5286 1273 5287
rect 1694 5286 1731 5352
rect 2326 5329 2372 6814
rect 1240 5257 1731 5286
rect 1128 5117 1163 5118
rect 419 5044 530 5066
rect 419 5024 427 5044
rect 446 5024 504 5044
rect 523 5024 530 5044
rect 419 5007 530 5024
rect 910 5035 952 5116
rect 1240 5037 1273 5257
rect 1694 5255 1731 5257
rect 2324 5305 2372 5329
rect 2554 5323 2601 6900
rect 3088 6857 3122 7036
rect 3353 7053 3463 7068
rect 3353 7050 3430 7053
rect 3353 7023 3356 7050
rect 3385 7026 3430 7050
rect 3459 7026 3463 7053
rect 3385 7023 3463 7026
rect 3353 7009 3463 7023
rect 2697 6832 3122 6857
rect 3201 6896 3238 6898
rect 3659 6896 3692 7116
rect 3980 7037 4022 7118
rect 4402 7129 4513 7145
rect 4402 7109 4409 7129
rect 4428 7109 4486 7129
rect 4505 7109 4513 7129
rect 4402 7087 4513 7109
rect 5242 7138 6242 7162
rect 3769 7035 3804 7036
rect 3201 6867 3692 6896
rect 2697 6816 3121 6832
rect 2697 6425 2735 6816
rect 3201 6801 3238 6867
rect 3659 6866 3692 6867
rect 3748 7028 3804 7035
rect 3748 7008 3777 7028
rect 3797 7008 3804 7028
rect 3748 7003 3804 7008
rect 3978 7033 4022 7037
rect 3978 7013 3989 7033
rect 4012 7013 4022 7033
rect 3978 7006 4022 7013
rect 4195 7031 4227 7038
rect 4195 7011 4201 7031
rect 4222 7011 4227 7031
rect 3978 7004 4021 7006
rect 3196 6792 3238 6801
rect 3196 6770 3205 6792
rect 3231 6770 3238 6792
rect 3463 6819 3574 6836
rect 3463 6799 3470 6819
rect 3489 6799 3547 6819
rect 3566 6799 3574 6819
rect 3463 6777 3574 6799
rect 3748 6797 3782 7003
rect 4195 6983 4227 7011
rect 3815 6975 4227 6983
rect 3815 6949 3821 6975
rect 3847 6949 4227 6975
rect 5242 6983 5290 7138
rect 5476 7097 5586 7111
rect 5476 7094 5554 7097
rect 5476 7067 5480 7094
rect 5509 7070 5554 7094
rect 5583 7070 5586 7097
rect 6207 7087 6242 7138
rect 6809 7156 7189 7182
rect 7215 7156 7221 7182
rect 6809 7148 7221 7156
rect 6809 7120 6841 7148
rect 6809 7100 6814 7120
rect 6835 7100 6841 7120
rect 6809 7093 6841 7100
rect 7015 7119 7060 7131
rect 7254 7128 7288 7334
rect 7015 7100 7022 7119
rect 7051 7100 7060 7119
rect 5509 7067 5586 7070
rect 5476 7052 5586 7067
rect 6205 7082 6242 7087
rect 6205 7062 6212 7082
rect 6232 7062 6242 7082
rect 6205 7055 6242 7062
rect 6205 7054 6240 7055
rect 5242 6954 5250 6983
rect 5279 6954 5290 6983
rect 5242 6949 5290 6954
rect 5761 6989 5793 6996
rect 5761 6969 5768 6989
rect 5789 6969 5793 6989
rect 3815 6947 4227 6949
rect 3817 6946 3857 6947
rect 4195 6882 4227 6947
rect 4195 6862 4199 6882
rect 4220 6862 4227 6882
rect 4195 6855 4227 6862
rect 5761 6904 5793 6969
rect 6131 6904 6171 6905
rect 5761 6902 6173 6904
rect 5761 6876 6141 6902
rect 6167 6876 6173 6902
rect 5761 6868 6173 6876
rect 5761 6840 5793 6868
rect 6206 6848 6240 7054
rect 6523 7022 6634 7044
rect 6523 7002 6531 7022
rect 6550 7002 6608 7022
rect 6627 7002 6634 7022
rect 6523 6985 6634 7002
rect 7015 7017 7060 7100
rect 7232 7123 7288 7128
rect 7232 7103 7239 7123
rect 7259 7103 7288 7123
rect 7755 7318 7784 7338
rect 7804 7318 7811 7338
rect 7755 7313 7811 7318
rect 8202 7341 8234 7348
rect 8202 7321 8208 7341
rect 8229 7321 8234 7341
rect 7755 7107 7789 7313
rect 8202 7293 8234 7321
rect 7822 7285 8234 7293
rect 7822 7259 7828 7285
rect 7854 7259 8234 7285
rect 8801 7303 8836 7354
rect 9457 7344 9460 7371
rect 9489 7347 9534 7371
rect 9563 7347 9567 7374
rect 9489 7344 9567 7347
rect 9457 7330 9567 7344
rect 9753 7303 9801 7458
rect 8801 7279 9801 7303
rect 8801 7276 9800 7279
rect 8801 7274 8836 7276
rect 7822 7257 8234 7259
rect 7824 7256 7864 7257
rect 7990 7216 8025 7234
rect 7990 7184 7993 7216
rect 8020 7184 8025 7216
rect 7755 7106 7790 7107
rect 7232 7096 7288 7103
rect 7753 7099 7791 7106
rect 7232 7095 7267 7096
rect 7753 7095 7763 7099
rect 7747 7081 7763 7095
rect 7783 7095 7791 7099
rect 7783 7081 7797 7095
rect 7747 7074 7797 7081
rect 7380 7017 7430 7019
rect 7015 6983 7430 7017
rect 7144 6921 7178 6922
rect 6275 6886 7179 6921
rect 7227 6910 7295 6921
rect 7227 6889 7232 6910
rect 5761 6820 5766 6840
rect 5787 6820 5793 6840
rect 5761 6813 5793 6820
rect 5968 6840 6007 6846
rect 5968 6820 5976 6840
rect 6001 6820 6007 6840
rect 5968 6813 6007 6820
rect 6184 6843 6240 6848
rect 6184 6823 6191 6843
rect 6211 6823 6240 6843
rect 6184 6816 6240 6823
rect 6184 6815 6219 6816
rect 3748 6789 3783 6797
rect 3196 6760 3238 6770
rect 3748 6769 3756 6789
rect 3776 6769 3783 6789
rect 3748 6764 3783 6769
rect 4402 6784 4512 6799
rect 4402 6781 4479 6784
rect 3196 6759 3237 6760
rect 2830 6725 2865 6726
rect 2809 6718 2865 6725
rect 2809 6698 2838 6718
rect 2858 6698 2865 6718
rect 2809 6693 2865 6698
rect 3256 6721 3288 6728
rect 3256 6701 3262 6721
rect 3283 6701 3288 6721
rect 3748 6712 3782 6764
rect 4402 6754 4405 6781
rect 4434 6757 4479 6781
rect 4508 6757 4512 6784
rect 4434 6754 4512 6757
rect 4402 6740 4512 6754
rect 4698 6784 4740 6794
rect 4698 6765 4706 6784
rect 4731 6765 4740 6784
rect 5976 6767 6007 6813
rect 4698 6712 4740 6765
rect 5475 6742 5586 6764
rect 5475 6722 5483 6742
rect 5502 6722 5560 6742
rect 5579 6722 5586 6742
rect 5975 6750 6007 6767
rect 6276 6750 6313 6886
rect 6414 6853 6524 6867
rect 6414 6850 6492 6853
rect 6414 6823 6418 6850
rect 6447 6826 6492 6850
rect 6521 6826 6524 6853
rect 7144 6843 7178 6886
rect 6447 6823 6524 6826
rect 6414 6808 6524 6823
rect 7143 6838 7178 6843
rect 7143 6818 7150 6838
rect 7170 6818 7178 6838
rect 7143 6810 7178 6818
rect 5975 6737 6313 6750
rect 2809 6487 2843 6693
rect 3256 6673 3288 6701
rect 3746 6686 4742 6712
rect 5475 6705 5586 6722
rect 5976 6718 6313 6737
rect 6255 6717 6313 6718
rect 6699 6745 6731 6752
rect 6699 6725 6706 6745
rect 6727 6725 6731 6745
rect 2876 6665 3288 6673
rect 2876 6639 2882 6665
rect 2908 6639 3288 6665
rect 2876 6637 3288 6639
rect 2878 6636 2918 6637
rect 3038 6601 3077 6616
rect 3038 6560 3049 6601
rect 3070 6560 3077 6601
rect 2808 6479 2844 6487
rect 2808 6459 2817 6479
rect 2837 6459 2844 6479
rect 2808 6458 2844 6459
rect 2808 6447 2842 6458
rect 2698 6417 2735 6425
rect 2698 6383 2942 6417
rect 2690 6214 2725 6215
rect 2669 6207 2725 6214
rect 2669 6187 2698 6207
rect 2718 6187 2725 6207
rect 2669 6182 2725 6187
rect 2900 6212 2942 6383
rect 3038 6287 3077 6560
rect 3256 6572 3288 6637
rect 6699 6660 6731 6725
rect 7069 6660 7109 6661
rect 6699 6658 7111 6660
rect 6699 6632 7079 6658
rect 7105 6632 7111 6658
rect 6699 6624 7111 6632
rect 3256 6552 3260 6572
rect 3281 6552 3288 6572
rect 3256 6545 3288 6552
rect 3674 6579 3732 6580
rect 3674 6560 4011 6579
rect 4401 6575 4512 6592
rect 5245 6585 6241 6611
rect 6699 6596 6731 6624
rect 3674 6547 4012 6560
rect 3178 6483 3231 6486
rect 3178 6466 3190 6483
rect 3222 6466 3231 6483
rect 3178 6458 3231 6466
rect 3177 6411 3231 6458
rect 3463 6474 3573 6489
rect 3463 6471 3540 6474
rect 3463 6444 3466 6471
rect 3495 6447 3540 6471
rect 3569 6447 3573 6474
rect 3495 6444 3573 6447
rect 3463 6430 3573 6444
rect 3674 6411 3711 6547
rect 3980 6530 4012 6547
rect 4401 6555 4408 6575
rect 4427 6555 4485 6575
rect 4504 6555 4512 6575
rect 4401 6533 4512 6555
rect 5247 6532 5289 6585
rect 3980 6484 4011 6530
rect 5247 6513 5256 6532
rect 5281 6513 5289 6532
rect 5247 6503 5289 6513
rect 5475 6543 5585 6557
rect 5475 6540 5553 6543
rect 5475 6513 5479 6540
rect 5508 6516 5553 6540
rect 5582 6516 5585 6543
rect 6205 6533 6239 6585
rect 6699 6576 6704 6596
rect 6725 6576 6731 6596
rect 6699 6569 6731 6576
rect 6909 6597 6947 6607
rect 7144 6604 7178 6810
rect 6909 6580 6919 6597
rect 6939 6580 6947 6597
rect 6750 6537 6791 6538
rect 5508 6513 5585 6516
rect 5475 6498 5585 6513
rect 6204 6528 6239 6533
rect 6204 6508 6211 6528
rect 6231 6508 6239 6528
rect 6749 6527 6791 6537
rect 6204 6500 6239 6508
rect 3768 6481 3803 6482
rect 3747 6474 3803 6481
rect 3747 6454 3776 6474
rect 3796 6454 3803 6474
rect 3747 6449 3803 6454
rect 3980 6477 4019 6484
rect 3980 6457 3986 6477
rect 4011 6457 4019 6477
rect 3980 6451 4019 6457
rect 4194 6477 4226 6484
rect 4194 6457 4200 6477
rect 4221 6457 4226 6477
rect 3177 6376 3712 6411
rect 3177 6372 3230 6376
rect 3038 6260 3042 6287
rect 3073 6260 3077 6287
rect 3323 6308 3434 6325
rect 3323 6288 3330 6308
rect 3349 6288 3407 6308
rect 3426 6288 3434 6308
rect 3323 6266 3434 6288
rect 3038 6253 3077 6260
rect 3747 6243 3781 6449
rect 4194 6429 4226 6457
rect 3814 6421 4226 6429
rect 3814 6395 3820 6421
rect 3846 6395 4226 6421
rect 3814 6393 4226 6395
rect 3816 6392 3856 6393
rect 4194 6328 4226 6393
rect 5760 6435 5792 6442
rect 5760 6415 5767 6435
rect 5788 6415 5792 6435
rect 5760 6350 5792 6415
rect 6130 6350 6170 6351
rect 5760 6348 6172 6350
rect 4194 6308 4198 6328
rect 4219 6308 4226 6328
rect 4194 6301 4226 6308
rect 4697 6343 4745 6348
rect 4697 6314 4708 6343
rect 4737 6314 4745 6343
rect 3747 6242 3782 6243
rect 3745 6235 3782 6242
rect 2900 6191 2908 6212
rect 2935 6191 2942 6212
rect 2669 5976 2703 6182
rect 2900 6180 2942 6191
rect 3116 6210 3148 6217
rect 3116 6190 3122 6210
rect 3143 6190 3148 6210
rect 3116 6162 3148 6190
rect 2736 6154 3148 6162
rect 2736 6128 2742 6154
rect 2768 6128 3148 6154
rect 3745 6215 3755 6235
rect 3775 6215 3782 6235
rect 3745 6210 3782 6215
rect 4401 6230 4511 6245
rect 4401 6227 4478 6230
rect 3745 6159 3780 6210
rect 4401 6200 4404 6227
rect 4433 6203 4478 6227
rect 4507 6203 4511 6230
rect 4433 6200 4511 6203
rect 4401 6186 4511 6200
rect 4697 6159 4745 6314
rect 5760 6322 6140 6348
rect 6166 6322 6172 6348
rect 5760 6314 6172 6322
rect 5760 6286 5792 6314
rect 6205 6294 6239 6500
rect 6413 6498 6524 6520
rect 6413 6478 6421 6498
rect 6440 6478 6498 6498
rect 6517 6478 6524 6498
rect 6413 6461 6524 6478
rect 6749 6505 6756 6527
rect 6782 6505 6791 6527
rect 6749 6496 6791 6505
rect 5966 6291 6009 6293
rect 5760 6266 5765 6286
rect 5786 6266 5792 6286
rect 5760 6259 5792 6266
rect 5965 6284 6009 6291
rect 5965 6264 5975 6284
rect 5998 6264 6009 6284
rect 5965 6260 6009 6264
rect 6183 6289 6239 6294
rect 6183 6269 6190 6289
rect 6210 6269 6239 6289
rect 6183 6262 6239 6269
rect 6295 6430 6328 6431
rect 6749 6430 6786 6496
rect 6295 6401 6786 6430
rect 6183 6261 6218 6262
rect 3745 6135 4745 6159
rect 5474 6188 5585 6210
rect 5474 6168 5482 6188
rect 5501 6168 5559 6188
rect 5578 6168 5585 6188
rect 5474 6151 5585 6168
rect 5965 6179 6007 6260
rect 6295 6181 6328 6401
rect 6749 6399 6786 6401
rect 6555 6261 6665 6275
rect 6555 6258 6633 6261
rect 6555 6231 6559 6258
rect 6588 6234 6633 6258
rect 6662 6234 6665 6261
rect 6588 6231 6665 6234
rect 6555 6216 6665 6231
rect 6909 6242 6947 6580
rect 7122 6599 7178 6604
rect 7122 6579 7129 6599
rect 7149 6579 7178 6599
rect 7122 6572 7178 6579
rect 7225 6881 7232 6889
rect 7280 6881 7295 6910
rect 7225 6872 7295 6881
rect 7122 6571 7157 6572
rect 7044 6471 7088 6475
rect 7225 6471 7275 6872
rect 7380 6855 7430 6983
rect 7613 6996 7723 6998
rect 7990 6996 8025 7184
rect 8202 7192 8234 7257
rect 8202 7172 8206 7192
rect 8227 7172 8234 7192
rect 8776 7188 9078 7190
rect 8202 7165 8234 7172
rect 8715 7159 9078 7188
rect 8715 7157 8776 7159
rect 7613 6966 8025 6996
rect 7613 6941 7657 6966
rect 7696 6963 8025 6966
rect 8144 7097 8178 7103
rect 8144 7077 8153 7097
rect 8174 7077 8178 7097
rect 7044 6438 7275 6471
rect 7044 6436 7251 6438
rect 7044 6282 7088 6436
rect 6909 6225 6917 6242
rect 6937 6225 6947 6242
rect 6909 6219 6947 6225
rect 6267 6179 6328 6181
rect 5965 6150 6328 6179
rect 6840 6153 6872 6160
rect 5965 6148 6267 6150
rect 3745 6132 4744 6135
rect 6840 6133 6847 6153
rect 6868 6133 6872 6153
rect 3745 6130 3780 6132
rect 2736 6126 3148 6128
rect 2738 6125 2778 6126
rect 3116 6061 3148 6126
rect 6840 6068 6872 6133
rect 7050 6146 7088 6282
rect 7287 6251 7318 6252
rect 7284 6246 7318 6251
rect 7284 6226 7291 6246
rect 7311 6226 7318 6246
rect 7284 6218 7318 6226
rect 7050 6108 7056 6146
rect 7079 6108 7088 6146
rect 7050 6098 7088 6108
rect 7285 6160 7318 6218
rect 7210 6068 7250 6069
rect 6840 6066 7252 6068
rect 6208 6062 6243 6064
rect 3116 6041 3120 6061
rect 3141 6041 3148 6061
rect 5244 6059 6243 6062
rect 3721 6044 4023 6046
rect 3116 6034 3148 6041
rect 3660 6015 4023 6044
rect 3660 6013 3721 6015
rect 2669 5968 2704 5976
rect 2669 5948 2677 5968
rect 2697 5948 2704 5968
rect 2669 5943 2704 5948
rect 3041 5969 3079 5975
rect 3041 5952 3051 5969
rect 3071 5952 3079 5969
rect 2669 5942 2701 5943
rect 2831 5622 2866 5623
rect 1468 5136 1578 5150
rect 1468 5133 1546 5136
rect 1468 5106 1472 5133
rect 1501 5109 1546 5133
rect 1575 5109 1578 5136
rect 2324 5127 2371 5305
rect 2554 5283 2567 5323
rect 2594 5283 2601 5323
rect 2810 5615 2866 5622
rect 2810 5595 2839 5615
rect 2859 5595 2866 5615
rect 2810 5590 2866 5595
rect 3041 5614 3079 5952
rect 3323 5963 3433 5978
rect 3323 5960 3400 5963
rect 3323 5933 3326 5960
rect 3355 5936 3400 5960
rect 3429 5936 3433 5963
rect 3355 5933 3433 5936
rect 3323 5919 3433 5933
rect 3202 5793 3239 5795
rect 3660 5793 3693 6013
rect 3981 5934 4023 6015
rect 4403 6026 4514 6043
rect 4403 6006 4410 6026
rect 4429 6006 4487 6026
rect 4506 6006 4514 6026
rect 4403 5984 4514 6006
rect 5243 6035 6243 6059
rect 3770 5932 3805 5933
rect 3202 5764 3693 5793
rect 3202 5698 3239 5764
rect 3660 5763 3693 5764
rect 3749 5925 3805 5932
rect 3749 5905 3778 5925
rect 3798 5905 3805 5925
rect 3749 5900 3805 5905
rect 3979 5930 4023 5934
rect 3979 5910 3990 5930
rect 4013 5910 4023 5930
rect 3979 5903 4023 5910
rect 4196 5928 4228 5935
rect 4196 5908 4202 5928
rect 4223 5908 4228 5928
rect 3979 5901 4022 5903
rect 3197 5689 3239 5698
rect 3197 5667 3206 5689
rect 3232 5667 3239 5689
rect 3464 5716 3575 5733
rect 3464 5696 3471 5716
rect 3490 5696 3548 5716
rect 3567 5696 3575 5716
rect 3464 5674 3575 5696
rect 3749 5694 3783 5900
rect 4196 5880 4228 5908
rect 3816 5872 4228 5880
rect 3816 5846 3822 5872
rect 3848 5846 4228 5872
rect 5243 5880 5291 6035
rect 5477 5994 5587 6008
rect 5477 5991 5555 5994
rect 5477 5964 5481 5991
rect 5510 5967 5555 5991
rect 5584 5967 5587 5994
rect 6208 5984 6243 6035
rect 5510 5964 5587 5967
rect 5477 5949 5587 5964
rect 6206 5979 6243 5984
rect 6206 5959 6213 5979
rect 6233 5959 6243 5979
rect 6840 6040 7220 6066
rect 7246 6040 7252 6066
rect 6840 6032 7252 6040
rect 6840 6004 6872 6032
rect 7285 6012 7321 6160
rect 6840 5984 6845 6004
rect 6866 5984 6872 6004
rect 6840 5977 6872 5984
rect 7263 6007 7321 6012
rect 7263 5987 7270 6007
rect 7290 5987 7321 6007
rect 7263 5980 7321 5987
rect 7263 5979 7298 5980
rect 6206 5952 6243 5959
rect 6206 5951 6241 5952
rect 5243 5851 5251 5880
rect 5280 5851 5291 5880
rect 5243 5846 5291 5851
rect 5762 5886 5794 5893
rect 5762 5866 5769 5886
rect 5790 5866 5794 5886
rect 3816 5844 4228 5846
rect 3818 5843 3858 5844
rect 4196 5779 4228 5844
rect 4196 5759 4200 5779
rect 4221 5759 4228 5779
rect 4196 5752 4228 5759
rect 5762 5801 5794 5866
rect 6132 5801 6172 5802
rect 5762 5799 6174 5801
rect 5762 5773 6142 5799
rect 6168 5773 6174 5799
rect 5762 5765 6174 5773
rect 5762 5737 5794 5765
rect 6207 5745 6241 5951
rect 6911 5934 6950 5941
rect 6554 5906 6665 5928
rect 6554 5886 6562 5906
rect 6581 5886 6639 5906
rect 6658 5886 6665 5906
rect 6554 5869 6665 5886
rect 6911 5907 6915 5934
rect 6946 5907 6950 5934
rect 6758 5818 6811 5822
rect 6276 5783 6811 5818
rect 5762 5717 5767 5737
rect 5788 5717 5794 5737
rect 5762 5710 5794 5717
rect 5969 5737 6008 5743
rect 5969 5717 5977 5737
rect 6002 5717 6008 5737
rect 5969 5710 6008 5717
rect 6185 5740 6241 5745
rect 6185 5720 6192 5740
rect 6212 5720 6241 5740
rect 6185 5713 6241 5720
rect 6185 5712 6220 5713
rect 3749 5686 3784 5694
rect 3197 5657 3239 5667
rect 3749 5666 3757 5686
rect 3777 5666 3784 5686
rect 3749 5661 3784 5666
rect 4403 5681 4513 5696
rect 4403 5678 4480 5681
rect 3197 5656 3238 5657
rect 3041 5597 3049 5614
rect 3069 5597 3079 5614
rect 2810 5384 2844 5590
rect 3041 5587 3079 5597
rect 3257 5618 3289 5625
rect 3257 5598 3263 5618
rect 3284 5598 3289 5618
rect 3749 5609 3783 5661
rect 4403 5651 4406 5678
rect 4435 5654 4480 5678
rect 4509 5654 4513 5681
rect 4435 5651 4513 5654
rect 4403 5637 4513 5651
rect 4699 5681 4741 5691
rect 4699 5662 4707 5681
rect 4732 5662 4741 5681
rect 5977 5664 6008 5710
rect 4699 5609 4741 5662
rect 5476 5639 5587 5661
rect 5476 5619 5484 5639
rect 5503 5619 5561 5639
rect 5580 5619 5587 5639
rect 5976 5647 6008 5664
rect 6277 5647 6314 5783
rect 6415 5750 6525 5764
rect 6415 5747 6493 5750
rect 6415 5720 6419 5747
rect 6448 5723 6493 5747
rect 6522 5723 6525 5750
rect 6448 5720 6525 5723
rect 6415 5705 6525 5720
rect 6757 5736 6811 5783
rect 6757 5728 6810 5736
rect 6757 5711 6766 5728
rect 6798 5711 6810 5728
rect 6757 5708 6810 5711
rect 5976 5634 6314 5647
rect 3257 5570 3289 5598
rect 3747 5583 4743 5609
rect 5476 5602 5587 5619
rect 5977 5615 6314 5634
rect 6256 5614 6314 5615
rect 6700 5642 6732 5649
rect 6700 5622 6707 5642
rect 6728 5622 6732 5642
rect 2877 5562 3289 5570
rect 2877 5536 2883 5562
rect 2909 5536 3289 5562
rect 2877 5534 3289 5536
rect 2879 5533 2919 5534
rect 3257 5469 3289 5534
rect 6700 5557 6732 5622
rect 6911 5634 6950 5907
rect 7146 5736 7180 5747
rect 7144 5735 7180 5736
rect 7144 5715 7151 5735
rect 7171 5715 7180 5735
rect 7144 5707 7180 5715
rect 6911 5593 6918 5634
rect 6939 5593 6950 5634
rect 6911 5578 6950 5593
rect 7070 5557 7110 5558
rect 6700 5555 7112 5557
rect 6700 5529 7080 5555
rect 7106 5529 7112 5555
rect 6700 5521 7112 5529
rect 3257 5449 3261 5469
rect 3282 5449 3289 5469
rect 3257 5442 3289 5449
rect 3675 5476 3733 5477
rect 3675 5457 4012 5476
rect 4402 5472 4513 5489
rect 5246 5482 6242 5508
rect 6700 5493 6732 5521
rect 7145 5501 7179 5707
rect 3675 5444 4013 5457
rect 2810 5376 2845 5384
rect 2810 5356 2818 5376
rect 2838 5356 2845 5376
rect 2810 5351 2845 5356
rect 3464 5371 3574 5386
rect 3464 5368 3541 5371
rect 2810 5308 2844 5351
rect 3464 5341 3467 5368
rect 3496 5344 3541 5368
rect 3570 5344 3574 5371
rect 3496 5341 3574 5344
rect 3464 5327 3574 5341
rect 3675 5308 3712 5444
rect 3981 5427 4013 5444
rect 4402 5452 4409 5472
rect 4428 5452 4486 5472
rect 4505 5452 4513 5472
rect 4402 5430 4513 5452
rect 5248 5429 5290 5482
rect 3981 5381 4012 5427
rect 5248 5410 5257 5429
rect 5282 5410 5290 5429
rect 5248 5400 5290 5410
rect 5476 5440 5586 5454
rect 5476 5437 5554 5440
rect 5476 5410 5480 5437
rect 5509 5413 5554 5437
rect 5583 5413 5586 5440
rect 6206 5430 6240 5482
rect 6700 5473 6705 5493
rect 6726 5473 6732 5493
rect 6700 5466 6732 5473
rect 7123 5496 7179 5501
rect 7123 5476 7130 5496
rect 7150 5476 7179 5496
rect 7123 5469 7179 5476
rect 7123 5468 7158 5469
rect 6751 5434 6792 5435
rect 5509 5410 5586 5413
rect 5476 5395 5586 5410
rect 6205 5425 6240 5430
rect 6205 5405 6212 5425
rect 6232 5405 6240 5425
rect 6750 5424 6792 5434
rect 6205 5397 6240 5405
rect 3769 5378 3804 5379
rect 3748 5371 3804 5378
rect 3748 5351 3777 5371
rect 3797 5351 3804 5371
rect 3748 5346 3804 5351
rect 3981 5374 4020 5381
rect 3981 5354 3987 5374
rect 4012 5354 4020 5374
rect 3981 5348 4020 5354
rect 4195 5374 4227 5381
rect 4195 5354 4201 5374
rect 4222 5354 4227 5374
rect 2554 5265 2601 5283
rect 2809 5273 3713 5308
rect 2810 5272 2844 5273
rect 2471 5206 2523 5211
rect 2926 5206 2971 5208
rect 2471 5191 2971 5206
rect 2471 5138 2485 5191
rect 2516 5167 2971 5191
rect 2516 5166 2541 5167
rect 2516 5138 2523 5166
rect 1501 5106 1578 5109
rect 1468 5091 1578 5106
rect 2193 5121 2374 5127
rect 2193 5101 2204 5121
rect 2224 5101 2374 5121
rect 2471 5114 2523 5138
rect 2193 5095 2374 5101
rect 2197 5093 2232 5095
rect 1212 5035 1273 5037
rect 910 5006 1273 5035
rect 1753 5028 1785 5035
rect 1753 5008 1760 5028
rect 1781 5008 1785 5028
rect 910 5004 1212 5006
rect 1753 4943 1785 5008
rect 2123 4943 2163 4944
rect 1753 4941 2165 4943
rect 1152 4918 1187 4920
rect 188 4915 1187 4918
rect 187 4891 1187 4915
rect 187 4736 235 4891
rect 421 4850 531 4864
rect 421 4847 499 4850
rect 421 4820 425 4847
rect 454 4823 499 4847
rect 528 4823 531 4850
rect 1152 4840 1187 4891
rect 1753 4915 2133 4941
rect 2159 4915 2165 4941
rect 1753 4907 2165 4915
rect 1753 4879 1785 4907
rect 2198 4887 2232 5093
rect 2722 5092 2757 5093
rect 1753 4859 1758 4879
rect 1779 4859 1785 4879
rect 1753 4852 1785 4859
rect 1955 4882 2000 4887
rect 1955 4858 1966 4882
rect 1992 4858 2000 4882
rect 1955 4847 2000 4858
rect 2176 4882 2232 4887
rect 2176 4862 2183 4882
rect 2203 4862 2232 4882
rect 2176 4855 2232 4862
rect 2701 5085 2757 5092
rect 2701 5065 2730 5085
rect 2750 5065 2757 5085
rect 2701 5060 2757 5065
rect 2926 5088 2971 5167
rect 3355 5186 3466 5203
rect 3355 5166 3362 5186
rect 3381 5166 3439 5186
rect 3458 5166 3466 5186
rect 3355 5144 3466 5166
rect 3748 5140 3782 5346
rect 4195 5326 4227 5354
rect 3815 5318 4227 5326
rect 3815 5292 3821 5318
rect 3847 5292 4227 5318
rect 3815 5290 4227 5292
rect 3817 5289 3857 5290
rect 4195 5225 4227 5290
rect 5761 5332 5793 5339
rect 5761 5312 5768 5332
rect 5789 5312 5793 5332
rect 5761 5247 5793 5312
rect 6131 5247 6171 5248
rect 5761 5245 6173 5247
rect 4195 5205 4199 5225
rect 4220 5205 4227 5225
rect 4195 5198 4227 5205
rect 4698 5240 4746 5245
rect 4698 5211 4709 5240
rect 4738 5211 4746 5240
rect 3748 5139 3783 5140
rect 3746 5132 3783 5139
rect 3746 5112 3756 5132
rect 3776 5112 3783 5132
rect 3746 5107 3783 5112
rect 4402 5127 4512 5142
rect 4402 5124 4479 5127
rect 2926 5068 2937 5088
rect 2962 5068 2971 5088
rect 2926 5064 2971 5068
rect 3148 5088 3180 5095
rect 3148 5068 3154 5088
rect 3175 5068 3180 5088
rect 2176 4854 2211 4855
rect 2701 4854 2735 5060
rect 3148 5040 3180 5068
rect 2768 5032 3180 5040
rect 2768 5006 2774 5032
rect 2800 5006 3180 5032
rect 3746 5056 3781 5107
rect 4402 5097 4405 5124
rect 4434 5100 4479 5124
rect 4508 5100 4512 5127
rect 4434 5097 4512 5100
rect 4402 5083 4512 5097
rect 4698 5056 4746 5211
rect 5761 5219 6141 5245
rect 6167 5219 6173 5245
rect 5761 5211 6173 5219
rect 5761 5183 5793 5211
rect 6206 5191 6240 5397
rect 6414 5395 6525 5417
rect 6414 5375 6422 5395
rect 6441 5375 6499 5395
rect 6518 5375 6525 5395
rect 6414 5358 6525 5375
rect 6750 5402 6757 5424
rect 6783 5402 6792 5424
rect 6750 5393 6792 5402
rect 5967 5188 6010 5190
rect 5761 5163 5766 5183
rect 5787 5163 5793 5183
rect 5761 5156 5793 5163
rect 5966 5181 6010 5188
rect 5966 5161 5976 5181
rect 5999 5161 6010 5181
rect 5966 5157 6010 5161
rect 6184 5186 6240 5191
rect 6184 5166 6191 5186
rect 6211 5166 6240 5186
rect 6184 5159 6240 5166
rect 6296 5327 6329 5328
rect 6750 5327 6787 5393
rect 7382 5370 7428 6855
rect 6296 5298 6787 5327
rect 6184 5158 6219 5159
rect 3746 5032 4746 5056
rect 5475 5085 5586 5107
rect 5475 5065 5483 5085
rect 5502 5065 5560 5085
rect 5579 5065 5586 5085
rect 5475 5048 5586 5065
rect 5966 5076 6008 5157
rect 6296 5078 6329 5298
rect 6750 5296 6787 5298
rect 7380 5346 7428 5370
rect 7610 5364 7657 6941
rect 8144 6898 8178 7077
rect 8409 7094 8519 7109
rect 8409 7091 8486 7094
rect 8409 7064 8412 7091
rect 8441 7067 8486 7091
rect 8515 7067 8519 7094
rect 8441 7064 8519 7067
rect 8409 7050 8519 7064
rect 7753 6873 8178 6898
rect 8257 6937 8294 6939
rect 8715 6937 8748 7157
rect 9036 7078 9078 7159
rect 9458 7170 9569 7186
rect 9458 7150 9465 7170
rect 9484 7150 9542 7170
rect 9561 7150 9569 7170
rect 9458 7128 9569 7150
rect 8825 7076 8860 7077
rect 8257 6908 8748 6937
rect 7753 6857 8177 6873
rect 7753 6466 7791 6857
rect 8257 6842 8294 6908
rect 8715 6907 8748 6908
rect 8804 7069 8860 7076
rect 8804 7049 8833 7069
rect 8853 7049 8860 7069
rect 8804 7044 8860 7049
rect 9034 7074 9078 7078
rect 9034 7054 9045 7074
rect 9068 7054 9078 7074
rect 9034 7047 9078 7054
rect 9251 7072 9283 7079
rect 9251 7052 9257 7072
rect 9278 7052 9283 7072
rect 9034 7045 9077 7047
rect 8252 6833 8294 6842
rect 8252 6811 8261 6833
rect 8287 6811 8294 6833
rect 8519 6860 8630 6877
rect 8519 6840 8526 6860
rect 8545 6840 8603 6860
rect 8622 6840 8630 6860
rect 8519 6818 8630 6840
rect 8804 6838 8838 7044
rect 9251 7024 9283 7052
rect 8871 7016 9283 7024
rect 8871 6990 8877 7016
rect 8903 6990 9283 7016
rect 8871 6988 9283 6990
rect 8873 6987 8913 6988
rect 9251 6923 9283 6988
rect 9251 6903 9255 6923
rect 9276 6903 9283 6923
rect 9251 6896 9283 6903
rect 8804 6830 8839 6838
rect 8252 6801 8294 6811
rect 8804 6810 8812 6830
rect 8832 6810 8839 6830
rect 8804 6805 8839 6810
rect 9458 6825 9568 6840
rect 9458 6822 9535 6825
rect 8252 6800 8293 6801
rect 7886 6766 7921 6767
rect 7865 6759 7921 6766
rect 7865 6739 7894 6759
rect 7914 6739 7921 6759
rect 7865 6734 7921 6739
rect 8312 6762 8344 6769
rect 8312 6742 8318 6762
rect 8339 6742 8344 6762
rect 8804 6753 8838 6805
rect 9458 6795 9461 6822
rect 9490 6798 9535 6822
rect 9564 6798 9568 6825
rect 9490 6795 9568 6798
rect 9458 6781 9568 6795
rect 9754 6825 9796 6835
rect 9754 6806 9762 6825
rect 9787 6806 9796 6825
rect 9754 6753 9796 6806
rect 7865 6528 7899 6734
rect 8312 6714 8344 6742
rect 8802 6727 9798 6753
rect 7932 6706 8344 6714
rect 7932 6680 7938 6706
rect 7964 6680 8344 6706
rect 7932 6678 8344 6680
rect 7934 6677 7974 6678
rect 8094 6642 8133 6657
rect 8094 6601 8105 6642
rect 8126 6601 8133 6642
rect 7864 6520 7900 6528
rect 7864 6500 7873 6520
rect 7893 6500 7900 6520
rect 7864 6499 7900 6500
rect 7864 6488 7898 6499
rect 7754 6458 7791 6466
rect 7754 6424 7998 6458
rect 7746 6255 7781 6256
rect 7725 6248 7781 6255
rect 7725 6228 7754 6248
rect 7774 6228 7781 6248
rect 7725 6223 7781 6228
rect 7956 6253 7998 6424
rect 8094 6328 8133 6601
rect 8312 6613 8344 6678
rect 8312 6593 8316 6613
rect 8337 6593 8344 6613
rect 8312 6586 8344 6593
rect 8730 6620 8788 6621
rect 8730 6601 9067 6620
rect 9457 6616 9568 6633
rect 8730 6588 9068 6601
rect 8234 6524 8287 6527
rect 8234 6507 8246 6524
rect 8278 6507 8287 6524
rect 8234 6499 8287 6507
rect 8233 6452 8287 6499
rect 8519 6515 8629 6530
rect 8519 6512 8596 6515
rect 8519 6485 8522 6512
rect 8551 6488 8596 6512
rect 8625 6488 8629 6515
rect 8551 6485 8629 6488
rect 8519 6471 8629 6485
rect 8730 6452 8767 6588
rect 9036 6571 9068 6588
rect 9457 6596 9464 6616
rect 9483 6596 9541 6616
rect 9560 6596 9568 6616
rect 9457 6574 9568 6596
rect 9036 6525 9067 6571
rect 8824 6522 8859 6523
rect 8803 6515 8859 6522
rect 8803 6495 8832 6515
rect 8852 6495 8859 6515
rect 8803 6490 8859 6495
rect 9036 6518 9075 6525
rect 9036 6498 9042 6518
rect 9067 6498 9075 6518
rect 9036 6492 9075 6498
rect 9250 6518 9282 6525
rect 9250 6498 9256 6518
rect 9277 6498 9282 6518
rect 8233 6417 8768 6452
rect 8233 6413 8286 6417
rect 8094 6301 8098 6328
rect 8129 6301 8133 6328
rect 8379 6349 8490 6366
rect 8379 6329 8386 6349
rect 8405 6329 8463 6349
rect 8482 6329 8490 6349
rect 8379 6307 8490 6329
rect 8094 6294 8133 6301
rect 8803 6284 8837 6490
rect 9250 6470 9282 6498
rect 8870 6462 9282 6470
rect 8870 6436 8876 6462
rect 8902 6436 9282 6462
rect 8870 6434 9282 6436
rect 8872 6433 8912 6434
rect 9250 6369 9282 6434
rect 9250 6349 9254 6369
rect 9275 6349 9282 6369
rect 9250 6342 9282 6349
rect 9753 6384 9801 6389
rect 9753 6355 9764 6384
rect 9793 6355 9801 6384
rect 8803 6283 8838 6284
rect 8801 6276 8838 6283
rect 7956 6232 7964 6253
rect 7991 6232 7998 6253
rect 7725 6017 7759 6223
rect 7956 6221 7998 6232
rect 8172 6251 8204 6258
rect 8172 6231 8178 6251
rect 8199 6231 8204 6251
rect 8172 6203 8204 6231
rect 7792 6195 8204 6203
rect 7792 6169 7798 6195
rect 7824 6169 8204 6195
rect 8801 6256 8811 6276
rect 8831 6256 8838 6276
rect 8801 6251 8838 6256
rect 9457 6271 9567 6286
rect 9457 6268 9534 6271
rect 8801 6200 8836 6251
rect 9457 6241 9460 6268
rect 9489 6244 9534 6268
rect 9563 6244 9567 6271
rect 9489 6241 9567 6244
rect 9457 6227 9567 6241
rect 9753 6200 9801 6355
rect 8801 6176 9801 6200
rect 8801 6173 9800 6176
rect 8801 6171 8836 6173
rect 7792 6167 8204 6169
rect 7794 6166 7834 6167
rect 8172 6102 8204 6167
rect 8172 6082 8176 6102
rect 8197 6082 8204 6102
rect 8777 6085 9079 6087
rect 8172 6075 8204 6082
rect 8716 6056 9079 6085
rect 8716 6054 8777 6056
rect 7725 6009 7760 6017
rect 7725 5989 7733 6009
rect 7753 5989 7760 6009
rect 7725 5984 7760 5989
rect 8097 6010 8135 6016
rect 8097 5993 8107 6010
rect 8127 5993 8135 6010
rect 7725 5983 7757 5984
rect 7887 5663 7922 5664
rect 6524 5177 6634 5191
rect 6524 5174 6602 5177
rect 6524 5147 6528 5174
rect 6557 5150 6602 5174
rect 6631 5150 6634 5177
rect 7380 5168 7427 5346
rect 7610 5324 7623 5364
rect 7650 5324 7657 5364
rect 7866 5656 7922 5663
rect 7866 5636 7895 5656
rect 7915 5636 7922 5656
rect 7866 5631 7922 5636
rect 8097 5655 8135 5993
rect 8379 6004 8489 6019
rect 8379 6001 8456 6004
rect 8379 5974 8382 6001
rect 8411 5977 8456 6001
rect 8485 5977 8489 6004
rect 8411 5974 8489 5977
rect 8379 5960 8489 5974
rect 8258 5834 8295 5836
rect 8716 5834 8749 6054
rect 9037 5975 9079 6056
rect 9459 6067 9570 6084
rect 9459 6047 9466 6067
rect 9485 6047 9543 6067
rect 9562 6047 9570 6067
rect 9459 6025 9570 6047
rect 8826 5973 8861 5974
rect 8258 5805 8749 5834
rect 8258 5739 8295 5805
rect 8716 5804 8749 5805
rect 8805 5966 8861 5973
rect 8805 5946 8834 5966
rect 8854 5946 8861 5966
rect 8805 5941 8861 5946
rect 9035 5971 9079 5975
rect 9035 5951 9046 5971
rect 9069 5951 9079 5971
rect 9035 5944 9079 5951
rect 9252 5969 9284 5976
rect 9252 5949 9258 5969
rect 9279 5949 9284 5969
rect 9035 5942 9078 5944
rect 8253 5730 8295 5739
rect 8253 5708 8262 5730
rect 8288 5708 8295 5730
rect 8520 5757 8631 5774
rect 8520 5737 8527 5757
rect 8546 5737 8604 5757
rect 8623 5737 8631 5757
rect 8520 5715 8631 5737
rect 8805 5735 8839 5941
rect 9252 5921 9284 5949
rect 8872 5913 9284 5921
rect 8872 5887 8878 5913
rect 8904 5887 9284 5913
rect 8872 5885 9284 5887
rect 8874 5884 8914 5885
rect 9252 5820 9284 5885
rect 9252 5800 9256 5820
rect 9277 5800 9284 5820
rect 9252 5793 9284 5800
rect 8805 5727 8840 5735
rect 8253 5698 8295 5708
rect 8805 5707 8813 5727
rect 8833 5707 8840 5727
rect 8805 5702 8840 5707
rect 9459 5722 9569 5737
rect 9459 5719 9536 5722
rect 8253 5697 8294 5698
rect 8097 5638 8105 5655
rect 8125 5638 8135 5655
rect 7866 5425 7900 5631
rect 8097 5628 8135 5638
rect 8313 5659 8345 5666
rect 8313 5639 8319 5659
rect 8340 5639 8345 5659
rect 8805 5650 8839 5702
rect 9459 5692 9462 5719
rect 9491 5695 9536 5719
rect 9565 5695 9569 5722
rect 9491 5692 9569 5695
rect 9459 5678 9569 5692
rect 9755 5722 9797 5732
rect 9755 5703 9763 5722
rect 9788 5703 9797 5722
rect 9755 5650 9797 5703
rect 8313 5611 8345 5639
rect 8803 5624 9799 5650
rect 7933 5603 8345 5611
rect 7933 5577 7939 5603
rect 7965 5577 8345 5603
rect 7933 5575 8345 5577
rect 7935 5574 7975 5575
rect 8313 5510 8345 5575
rect 8313 5490 8317 5510
rect 8338 5490 8345 5510
rect 8313 5483 8345 5490
rect 8731 5517 8789 5518
rect 8731 5498 9068 5517
rect 9458 5513 9569 5530
rect 8731 5485 9069 5498
rect 7866 5417 7901 5425
rect 7866 5397 7874 5417
rect 7894 5397 7901 5417
rect 7866 5392 7901 5397
rect 8520 5412 8630 5427
rect 8520 5409 8597 5412
rect 7866 5349 7900 5392
rect 8520 5382 8523 5409
rect 8552 5385 8597 5409
rect 8626 5385 8630 5412
rect 8552 5382 8630 5385
rect 8520 5368 8630 5382
rect 8731 5349 8768 5485
rect 9037 5468 9069 5485
rect 9458 5493 9465 5513
rect 9484 5493 9542 5513
rect 9561 5493 9569 5513
rect 9458 5471 9569 5493
rect 9037 5422 9068 5468
rect 8825 5419 8860 5420
rect 8804 5412 8860 5419
rect 8804 5392 8833 5412
rect 8853 5392 8860 5412
rect 8804 5387 8860 5392
rect 9037 5415 9076 5422
rect 9037 5395 9043 5415
rect 9068 5395 9076 5415
rect 9037 5389 9076 5395
rect 9251 5415 9283 5422
rect 9251 5395 9257 5415
rect 9278 5395 9283 5415
rect 7610 5306 7657 5324
rect 7865 5314 8769 5349
rect 7866 5313 7900 5314
rect 7527 5247 7579 5252
rect 7982 5247 8027 5249
rect 7527 5232 8027 5247
rect 7527 5179 7541 5232
rect 7572 5208 8027 5232
rect 7572 5207 7597 5208
rect 7572 5179 7579 5207
rect 6557 5147 6634 5150
rect 6524 5132 6634 5147
rect 7249 5162 7430 5168
rect 7249 5142 7260 5162
rect 7280 5142 7430 5162
rect 7527 5155 7579 5179
rect 7249 5136 7430 5142
rect 7253 5134 7288 5136
rect 6268 5076 6329 5078
rect 5966 5047 6329 5076
rect 6809 5069 6841 5076
rect 6809 5049 6816 5069
rect 6837 5049 6841 5069
rect 5966 5045 6268 5047
rect 3746 5029 4745 5032
rect 3746 5027 3781 5029
rect 2768 5004 3180 5006
rect 2770 5003 2810 5004
rect 3148 4939 3180 5004
rect 6809 4984 6841 5049
rect 7179 4984 7219 4985
rect 6809 4982 7221 4984
rect 6208 4959 6243 4961
rect 5244 4956 6243 4959
rect 3721 4941 4023 4943
rect 3148 4919 3152 4939
rect 3173 4919 3180 4939
rect 3148 4912 3180 4919
rect 3660 4912 4023 4941
rect 3660 4910 3721 4912
rect 2701 4852 2736 4854
rect 454 4820 531 4823
rect 421 4805 531 4820
rect 1150 4835 1187 4840
rect 1150 4815 1157 4835
rect 1177 4815 1187 4835
rect 1150 4808 1187 4815
rect 1956 4813 1994 4847
rect 2559 4846 2740 4852
rect 2559 4826 2709 4846
rect 2729 4826 2740 4846
rect 2559 4820 2740 4826
rect 3355 4841 3465 4856
rect 3355 4838 3432 4841
rect 2392 4813 2442 4817
rect 1150 4807 1185 4808
rect 187 4707 195 4736
rect 224 4707 235 4736
rect 187 4702 235 4707
rect 706 4742 738 4749
rect 706 4722 713 4742
rect 734 4722 738 4742
rect 706 4657 738 4722
rect 1076 4657 1116 4658
rect 706 4655 1118 4657
rect 706 4629 1086 4655
rect 1112 4629 1118 4655
rect 706 4621 1118 4629
rect 706 4593 738 4621
rect 1151 4601 1185 4807
rect 1956 4803 2442 4813
rect 1467 4781 1578 4803
rect 1467 4761 1475 4781
rect 1494 4761 1552 4781
rect 1571 4761 1578 4781
rect 1956 4771 2405 4803
rect 1467 4744 1578 4761
rect 2392 4750 2405 4771
rect 2436 4750 2442 4803
rect 2392 4733 2442 4750
rect 2089 4674 2123 4675
rect 1220 4639 2124 4674
rect 2332 4664 2379 4682
rect 706 4573 711 4593
rect 732 4573 738 4593
rect 706 4566 738 4573
rect 913 4593 952 4599
rect 913 4573 921 4593
rect 946 4573 952 4593
rect 913 4566 952 4573
rect 1129 4596 1185 4601
rect 1129 4576 1136 4596
rect 1156 4576 1185 4596
rect 1129 4569 1185 4576
rect 1129 4568 1164 4569
rect 921 4520 952 4566
rect 420 4495 531 4517
rect 420 4475 428 4495
rect 447 4475 505 4495
rect 524 4475 531 4495
rect 920 4503 952 4520
rect 1221 4503 1258 4639
rect 1359 4606 1469 4620
rect 1359 4603 1437 4606
rect 1359 4576 1363 4603
rect 1392 4579 1437 4603
rect 1466 4579 1469 4606
rect 2089 4596 2123 4639
rect 1392 4576 1469 4579
rect 1359 4561 1469 4576
rect 2088 4591 2123 4596
rect 2088 4571 2095 4591
rect 2115 4571 2123 4591
rect 2088 4563 2123 4571
rect 920 4490 1258 4503
rect 420 4458 531 4475
rect 921 4471 1258 4490
rect 1200 4470 1258 4471
rect 1644 4498 1676 4505
rect 1644 4478 1651 4498
rect 1672 4478 1676 4498
rect 1644 4413 1676 4478
rect 2014 4413 2054 4414
rect 1644 4411 2056 4413
rect 1644 4385 2024 4411
rect 2050 4385 2056 4411
rect 1644 4377 2056 4385
rect 190 4338 1186 4364
rect 1644 4349 1676 4377
rect 192 4285 234 4338
rect 192 4266 201 4285
rect 226 4266 234 4285
rect 192 4256 234 4266
rect 420 4296 530 4310
rect 420 4293 498 4296
rect 420 4266 424 4293
rect 453 4269 498 4293
rect 527 4269 530 4296
rect 1150 4286 1184 4338
rect 1644 4329 1649 4349
rect 1670 4329 1676 4349
rect 1644 4322 1676 4329
rect 1854 4350 1892 4360
rect 2089 4357 2123 4563
rect 1854 4333 1864 4350
rect 1884 4333 1892 4350
rect 1695 4290 1736 4291
rect 453 4266 530 4269
rect 420 4251 530 4266
rect 1149 4281 1184 4286
rect 1149 4261 1156 4281
rect 1176 4261 1184 4281
rect 1694 4280 1736 4290
rect 1149 4253 1184 4261
rect 705 4188 737 4195
rect 705 4168 712 4188
rect 733 4168 737 4188
rect 705 4103 737 4168
rect 1075 4103 1115 4104
rect 705 4101 1117 4103
rect 705 4075 1085 4101
rect 1111 4075 1117 4101
rect 705 4067 1117 4075
rect 705 4039 737 4067
rect 1150 4047 1184 4253
rect 1358 4251 1469 4273
rect 1358 4231 1366 4251
rect 1385 4231 1443 4251
rect 1462 4231 1469 4251
rect 1358 4214 1469 4231
rect 1694 4258 1701 4280
rect 1727 4258 1736 4280
rect 1694 4249 1736 4258
rect 911 4044 954 4046
rect 705 4019 710 4039
rect 731 4019 737 4039
rect 705 4012 737 4019
rect 910 4037 954 4044
rect 910 4017 920 4037
rect 943 4017 954 4037
rect 910 4013 954 4017
rect 1128 4042 1184 4047
rect 1128 4022 1135 4042
rect 1155 4022 1184 4042
rect 1128 4015 1184 4022
rect 1240 4183 1273 4184
rect 1694 4183 1731 4249
rect 1240 4154 1731 4183
rect 1128 4014 1163 4015
rect 419 3941 530 3963
rect 419 3921 427 3941
rect 446 3921 504 3941
rect 523 3921 530 3941
rect 419 3904 530 3921
rect 910 3932 952 4013
rect 1240 3934 1273 4154
rect 1694 4152 1731 4154
rect 1500 4014 1610 4028
rect 1500 4011 1578 4014
rect 1500 3984 1504 4011
rect 1533 3987 1578 4011
rect 1607 3987 1610 4014
rect 1533 3984 1610 3987
rect 1500 3969 1610 3984
rect 1854 3995 1892 4333
rect 2067 4352 2123 4357
rect 2067 4332 2074 4352
rect 2094 4332 2123 4352
rect 2067 4325 2123 4332
rect 2332 4624 2339 4664
rect 2366 4624 2379 4664
rect 2562 4642 2609 4820
rect 3355 4811 3358 4838
rect 3387 4814 3432 4838
rect 3461 4814 3465 4841
rect 3387 4811 3465 4814
rect 3355 4797 3465 4811
rect 2067 4324 2102 4325
rect 2232 4004 2264 4005
rect 1854 3978 1862 3995
rect 1882 3978 1892 3995
rect 1854 3972 1892 3978
rect 2229 3999 2264 4004
rect 2229 3979 2236 3999
rect 2256 3979 2264 3999
rect 2229 3971 2264 3979
rect 1212 3932 1273 3934
rect 910 3903 1273 3932
rect 1785 3906 1817 3913
rect 910 3901 1212 3903
rect 1785 3886 1792 3906
rect 1813 3886 1817 3906
rect 1785 3821 1817 3886
rect 2155 3821 2195 3822
rect 1785 3819 2197 3821
rect 1153 3815 1188 3817
rect 189 3812 1188 3815
rect 188 3788 1188 3812
rect 188 3633 236 3788
rect 422 3747 532 3761
rect 422 3744 500 3747
rect 422 3717 426 3744
rect 455 3720 500 3744
rect 529 3720 532 3747
rect 1153 3737 1188 3788
rect 455 3717 532 3720
rect 422 3702 532 3717
rect 1151 3732 1188 3737
rect 1151 3712 1158 3732
rect 1178 3712 1188 3732
rect 1785 3793 2165 3819
rect 2191 3793 2197 3819
rect 1785 3785 2197 3793
rect 1785 3757 1817 3785
rect 1785 3737 1790 3757
rect 1811 3737 1817 3757
rect 1785 3730 1817 3737
rect 1991 3756 2033 3767
rect 2230 3765 2264 3971
rect 1991 3735 1998 3756
rect 2025 3735 2033 3756
rect 1151 3705 1188 3712
rect 1151 3704 1186 3705
rect 188 3604 196 3633
rect 225 3604 236 3633
rect 188 3599 236 3604
rect 707 3639 739 3646
rect 707 3619 714 3639
rect 735 3619 739 3639
rect 707 3554 739 3619
rect 1077 3554 1117 3555
rect 707 3552 1119 3554
rect 707 3526 1087 3552
rect 1113 3526 1119 3552
rect 707 3518 1119 3526
rect 707 3490 739 3518
rect 1152 3498 1186 3704
rect 1856 3687 1895 3694
rect 1499 3659 1610 3681
rect 1499 3639 1507 3659
rect 1526 3639 1584 3659
rect 1603 3639 1610 3659
rect 1499 3622 1610 3639
rect 1856 3660 1860 3687
rect 1891 3660 1895 3687
rect 1703 3571 1756 3575
rect 1221 3536 1756 3571
rect 707 3470 712 3490
rect 733 3470 739 3490
rect 707 3463 739 3470
rect 914 3490 953 3496
rect 914 3470 922 3490
rect 947 3470 953 3490
rect 914 3463 953 3470
rect 1130 3493 1186 3498
rect 1130 3473 1137 3493
rect 1157 3473 1186 3493
rect 1130 3466 1186 3473
rect 1130 3465 1165 3466
rect 922 3417 953 3463
rect 421 3392 532 3414
rect 421 3372 429 3392
rect 448 3372 506 3392
rect 525 3372 532 3392
rect 921 3400 953 3417
rect 1222 3400 1259 3536
rect 1360 3503 1470 3517
rect 1360 3500 1438 3503
rect 1360 3473 1364 3500
rect 1393 3476 1438 3500
rect 1467 3476 1470 3503
rect 1393 3473 1470 3476
rect 1360 3458 1470 3473
rect 1702 3489 1756 3536
rect 1702 3481 1755 3489
rect 1702 3464 1711 3481
rect 1743 3464 1755 3481
rect 1702 3461 1755 3464
rect 921 3387 1259 3400
rect 421 3355 532 3372
rect 922 3368 1259 3387
rect 1201 3367 1259 3368
rect 1645 3395 1677 3402
rect 1645 3375 1652 3395
rect 1673 3375 1677 3395
rect 1645 3310 1677 3375
rect 1856 3387 1895 3660
rect 1991 3564 2033 3735
rect 2208 3760 2264 3765
rect 2208 3740 2215 3760
rect 2235 3740 2264 3760
rect 2208 3733 2264 3740
rect 2208 3732 2243 3733
rect 1991 3530 2235 3564
rect 2198 3522 2235 3530
rect 2091 3489 2125 3500
rect 2089 3488 2125 3489
rect 2089 3468 2096 3488
rect 2116 3468 2125 3488
rect 2089 3460 2125 3468
rect 1856 3346 1863 3387
rect 1884 3346 1895 3387
rect 1856 3331 1895 3346
rect 2015 3310 2055 3311
rect 1645 3308 2057 3310
rect 1645 3282 2025 3308
rect 2051 3282 2057 3308
rect 1645 3274 2057 3282
rect 191 3235 1187 3261
rect 1645 3246 1677 3274
rect 2090 3254 2124 3460
rect 193 3182 235 3235
rect 193 3163 202 3182
rect 227 3163 235 3182
rect 193 3153 235 3163
rect 421 3193 531 3207
rect 421 3190 499 3193
rect 421 3163 425 3190
rect 454 3166 499 3190
rect 528 3166 531 3193
rect 1151 3183 1185 3235
rect 1645 3226 1650 3246
rect 1671 3226 1677 3246
rect 1645 3219 1677 3226
rect 2068 3249 2124 3254
rect 2068 3229 2075 3249
rect 2095 3229 2124 3249
rect 2068 3222 2124 3229
rect 2068 3221 2103 3222
rect 1696 3187 1737 3188
rect 454 3163 531 3166
rect 421 3148 531 3163
rect 1150 3178 1185 3183
rect 1150 3158 1157 3178
rect 1177 3158 1185 3178
rect 1695 3177 1737 3187
rect 1150 3150 1185 3158
rect 706 3085 738 3092
rect 706 3065 713 3085
rect 734 3065 738 3085
rect 706 3000 738 3065
rect 1076 3000 1116 3001
rect 706 2998 1118 3000
rect 706 2972 1086 2998
rect 1112 2972 1118 2998
rect 706 2964 1118 2972
rect 706 2936 738 2964
rect 1151 2944 1185 3150
rect 1359 3148 1470 3170
rect 1359 3128 1367 3148
rect 1386 3128 1444 3148
rect 1463 3128 1470 3148
rect 1359 3111 1470 3128
rect 1695 3155 1702 3177
rect 1728 3155 1737 3177
rect 1695 3146 1737 3155
rect 912 2941 955 2943
rect 706 2916 711 2936
rect 732 2916 738 2936
rect 706 2909 738 2916
rect 911 2934 955 2941
rect 911 2914 921 2934
rect 944 2914 955 2934
rect 911 2910 955 2914
rect 1129 2939 1185 2944
rect 1129 2919 1136 2939
rect 1156 2919 1185 2939
rect 1129 2912 1185 2919
rect 1241 3080 1274 3081
rect 1695 3080 1732 3146
rect 2198 3131 2236 3522
rect 1812 3115 2236 3131
rect 1241 3051 1732 3080
rect 1129 2911 1164 2912
rect 420 2838 531 2860
rect 420 2818 428 2838
rect 447 2818 505 2838
rect 524 2818 531 2838
rect 420 2802 531 2818
rect 911 2829 953 2910
rect 1241 2831 1274 3051
rect 1695 3049 1732 3051
rect 1811 3090 2236 3115
rect 1470 2924 1580 2938
rect 1470 2921 1548 2924
rect 1470 2894 1474 2921
rect 1503 2897 1548 2921
rect 1577 2897 1580 2924
rect 1503 2894 1580 2897
rect 1470 2879 1580 2894
rect 1811 2911 1845 3090
rect 2332 3047 2379 4624
rect 2561 4618 2609 4642
rect 3202 4690 3239 4692
rect 3660 4690 3693 4910
rect 3981 4831 4023 4912
rect 4403 4923 4514 4940
rect 4403 4903 4410 4923
rect 4429 4903 4487 4923
rect 4506 4903 4514 4923
rect 4403 4881 4514 4903
rect 5243 4932 6243 4956
rect 3770 4829 3805 4830
rect 3202 4661 3693 4690
rect 2561 3133 2607 4618
rect 3202 4595 3239 4661
rect 3660 4660 3693 4661
rect 3749 4822 3805 4829
rect 3749 4802 3778 4822
rect 3798 4802 3805 4822
rect 3749 4797 3805 4802
rect 3979 4827 4023 4831
rect 3979 4807 3990 4827
rect 4013 4807 4023 4827
rect 3979 4800 4023 4807
rect 4196 4825 4228 4832
rect 4196 4805 4202 4825
rect 4223 4805 4228 4825
rect 3979 4798 4022 4800
rect 3197 4586 3239 4595
rect 3197 4564 3206 4586
rect 3232 4564 3239 4586
rect 3464 4613 3575 4630
rect 3464 4593 3471 4613
rect 3490 4593 3548 4613
rect 3567 4593 3575 4613
rect 3464 4571 3575 4593
rect 3749 4591 3783 4797
rect 4196 4777 4228 4805
rect 3816 4769 4228 4777
rect 3816 4743 3822 4769
rect 3848 4743 4228 4769
rect 5243 4777 5291 4932
rect 5477 4891 5587 4905
rect 5477 4888 5555 4891
rect 5477 4861 5481 4888
rect 5510 4864 5555 4888
rect 5584 4864 5587 4891
rect 6208 4881 6243 4932
rect 6809 4956 7189 4982
rect 7215 4956 7221 4982
rect 6809 4948 7221 4956
rect 6809 4920 6841 4948
rect 7254 4928 7288 5134
rect 7778 5133 7813 5134
rect 6809 4900 6814 4920
rect 6835 4900 6841 4920
rect 6809 4893 6841 4900
rect 7011 4923 7056 4928
rect 7011 4899 7022 4923
rect 7048 4899 7056 4923
rect 7011 4888 7056 4899
rect 7232 4923 7288 4928
rect 7232 4903 7239 4923
rect 7259 4903 7288 4923
rect 7232 4896 7288 4903
rect 7757 5126 7813 5133
rect 7757 5106 7786 5126
rect 7806 5106 7813 5126
rect 7757 5101 7813 5106
rect 7982 5129 8027 5208
rect 8411 5227 8522 5244
rect 8411 5207 8418 5227
rect 8437 5207 8495 5227
rect 8514 5207 8522 5227
rect 8411 5185 8522 5207
rect 8804 5181 8838 5387
rect 9251 5367 9283 5395
rect 8871 5359 9283 5367
rect 8871 5333 8877 5359
rect 8903 5333 9283 5359
rect 8871 5331 9283 5333
rect 8873 5330 8913 5331
rect 9251 5266 9283 5331
rect 9251 5246 9255 5266
rect 9276 5246 9283 5266
rect 9251 5239 9283 5246
rect 9754 5281 9802 5286
rect 9754 5252 9765 5281
rect 9794 5252 9802 5281
rect 8804 5180 8839 5181
rect 8802 5173 8839 5180
rect 8802 5153 8812 5173
rect 8832 5153 8839 5173
rect 8802 5148 8839 5153
rect 9458 5168 9568 5183
rect 9458 5165 9535 5168
rect 7982 5109 7993 5129
rect 8018 5109 8027 5129
rect 7982 5105 8027 5109
rect 8204 5129 8236 5136
rect 8204 5109 8210 5129
rect 8231 5109 8236 5129
rect 7232 4895 7267 4896
rect 7757 4895 7791 5101
rect 8204 5081 8236 5109
rect 7824 5073 8236 5081
rect 7824 5047 7830 5073
rect 7856 5047 8236 5073
rect 8802 5097 8837 5148
rect 9458 5138 9461 5165
rect 9490 5141 9535 5165
rect 9564 5141 9568 5168
rect 9490 5138 9568 5141
rect 9458 5124 9568 5138
rect 9754 5097 9802 5252
rect 8802 5073 9802 5097
rect 8802 5070 9801 5073
rect 8802 5068 8837 5070
rect 7824 5045 8236 5047
rect 7826 5044 7866 5045
rect 8204 4980 8236 5045
rect 8777 4982 9079 4984
rect 8204 4960 8208 4980
rect 8229 4960 8236 4980
rect 8204 4953 8236 4960
rect 8716 4953 9079 4982
rect 8716 4951 8777 4953
rect 7757 4893 7792 4895
rect 5510 4861 5587 4864
rect 5477 4846 5587 4861
rect 6206 4876 6243 4881
rect 6206 4856 6213 4876
rect 6233 4856 6243 4876
rect 6206 4849 6243 4856
rect 7012 4854 7050 4888
rect 7615 4887 7796 4893
rect 7615 4867 7765 4887
rect 7785 4867 7796 4887
rect 7615 4861 7796 4867
rect 8411 4882 8521 4897
rect 8411 4879 8488 4882
rect 7448 4854 7498 4858
rect 6206 4848 6241 4849
rect 5243 4748 5251 4777
rect 5280 4748 5291 4777
rect 5243 4743 5291 4748
rect 5762 4783 5794 4790
rect 5762 4763 5769 4783
rect 5790 4763 5794 4783
rect 3816 4741 4228 4743
rect 3818 4740 3858 4741
rect 4196 4676 4228 4741
rect 4196 4656 4200 4676
rect 4221 4656 4228 4676
rect 4196 4649 4228 4656
rect 5762 4698 5794 4763
rect 6132 4698 6172 4699
rect 5762 4696 6174 4698
rect 5762 4670 6142 4696
rect 6168 4670 6174 4696
rect 5762 4662 6174 4670
rect 5762 4634 5794 4662
rect 6207 4642 6241 4848
rect 7012 4844 7498 4854
rect 6523 4822 6634 4844
rect 6523 4802 6531 4822
rect 6550 4802 6608 4822
rect 6627 4802 6634 4822
rect 7012 4812 7461 4844
rect 6523 4785 6634 4802
rect 7448 4791 7461 4812
rect 7492 4791 7498 4844
rect 7448 4774 7498 4791
rect 7145 4715 7179 4716
rect 6276 4680 7180 4715
rect 7388 4705 7435 4723
rect 5762 4614 5767 4634
rect 5788 4614 5794 4634
rect 5762 4607 5794 4614
rect 5969 4634 6008 4640
rect 5969 4614 5977 4634
rect 6002 4614 6008 4634
rect 5969 4607 6008 4614
rect 6185 4637 6241 4642
rect 6185 4617 6192 4637
rect 6212 4617 6241 4637
rect 6185 4610 6241 4617
rect 6185 4609 6220 4610
rect 3749 4583 3784 4591
rect 3197 4554 3239 4564
rect 3749 4563 3757 4583
rect 3777 4563 3784 4583
rect 3749 4558 3784 4563
rect 4403 4578 4513 4593
rect 4403 4575 4480 4578
rect 3197 4553 3238 4554
rect 2831 4519 2866 4520
rect 2810 4512 2866 4519
rect 2810 4492 2839 4512
rect 2859 4492 2866 4512
rect 2810 4487 2866 4492
rect 3257 4515 3289 4522
rect 3257 4495 3263 4515
rect 3284 4495 3289 4515
rect 3749 4506 3783 4558
rect 4403 4548 4406 4575
rect 4435 4551 4480 4575
rect 4509 4551 4513 4578
rect 4435 4548 4513 4551
rect 4403 4534 4513 4548
rect 4699 4578 4741 4588
rect 4699 4559 4707 4578
rect 4732 4559 4741 4578
rect 5977 4561 6008 4607
rect 4699 4506 4741 4559
rect 5476 4536 5587 4558
rect 5476 4516 5484 4536
rect 5503 4516 5561 4536
rect 5580 4516 5587 4536
rect 5976 4544 6008 4561
rect 6277 4544 6314 4680
rect 6415 4647 6525 4661
rect 6415 4644 6493 4647
rect 6415 4617 6419 4644
rect 6448 4620 6493 4644
rect 6522 4620 6525 4647
rect 7145 4637 7179 4680
rect 6448 4617 6525 4620
rect 6415 4602 6525 4617
rect 7144 4632 7179 4637
rect 7144 4612 7151 4632
rect 7171 4612 7179 4632
rect 7144 4604 7179 4612
rect 5976 4531 6314 4544
rect 2810 4281 2844 4487
rect 3257 4467 3289 4495
rect 3747 4480 4743 4506
rect 5476 4499 5587 4516
rect 5977 4512 6314 4531
rect 6256 4511 6314 4512
rect 6700 4539 6732 4546
rect 6700 4519 6707 4539
rect 6728 4519 6732 4539
rect 2877 4459 3289 4467
rect 2877 4433 2883 4459
rect 2909 4433 3289 4459
rect 2877 4431 3289 4433
rect 2879 4430 2919 4431
rect 3039 4395 3078 4410
rect 3039 4354 3050 4395
rect 3071 4354 3078 4395
rect 2809 4273 2845 4281
rect 2809 4253 2818 4273
rect 2838 4253 2845 4273
rect 2809 4252 2845 4253
rect 2809 4241 2843 4252
rect 3039 4081 3078 4354
rect 3257 4366 3289 4431
rect 6700 4454 6732 4519
rect 7070 4454 7110 4455
rect 6700 4452 7112 4454
rect 6700 4426 7080 4452
rect 7106 4426 7112 4452
rect 6700 4418 7112 4426
rect 3257 4346 3261 4366
rect 3282 4346 3289 4366
rect 3257 4339 3289 4346
rect 3675 4373 3733 4374
rect 3675 4354 4012 4373
rect 4402 4369 4513 4386
rect 5246 4379 6242 4405
rect 6700 4390 6732 4418
rect 3675 4341 4013 4354
rect 3179 4277 3232 4280
rect 3179 4260 3191 4277
rect 3223 4260 3232 4277
rect 3179 4252 3232 4260
rect 3178 4205 3232 4252
rect 3464 4268 3574 4283
rect 3464 4265 3541 4268
rect 3464 4238 3467 4265
rect 3496 4241 3541 4265
rect 3570 4241 3574 4268
rect 3496 4238 3574 4241
rect 3464 4224 3574 4238
rect 3675 4205 3712 4341
rect 3981 4324 4013 4341
rect 4402 4349 4409 4369
rect 4428 4349 4486 4369
rect 4505 4349 4513 4369
rect 4402 4327 4513 4349
rect 5248 4326 5290 4379
rect 3981 4278 4012 4324
rect 5248 4307 5257 4326
rect 5282 4307 5290 4326
rect 5248 4297 5290 4307
rect 5476 4337 5586 4351
rect 5476 4334 5554 4337
rect 5476 4307 5480 4334
rect 5509 4310 5554 4334
rect 5583 4310 5586 4337
rect 6206 4327 6240 4379
rect 6700 4370 6705 4390
rect 6726 4370 6732 4390
rect 6700 4363 6732 4370
rect 6910 4391 6948 4401
rect 7145 4398 7179 4604
rect 6910 4374 6920 4391
rect 6940 4374 6948 4391
rect 6751 4331 6792 4332
rect 5509 4307 5586 4310
rect 5476 4292 5586 4307
rect 6205 4322 6240 4327
rect 6205 4302 6212 4322
rect 6232 4302 6240 4322
rect 6750 4321 6792 4331
rect 6205 4294 6240 4302
rect 3769 4275 3804 4276
rect 3748 4268 3804 4275
rect 3748 4248 3777 4268
rect 3797 4248 3804 4268
rect 3748 4243 3804 4248
rect 3981 4271 4020 4278
rect 3981 4251 3987 4271
rect 4012 4251 4020 4271
rect 3981 4245 4020 4251
rect 4195 4271 4227 4278
rect 4195 4251 4201 4271
rect 4222 4251 4227 4271
rect 3178 4170 3713 4205
rect 3178 4166 3231 4170
rect 3039 4054 3043 4081
rect 3074 4054 3078 4081
rect 3324 4102 3435 4119
rect 3324 4082 3331 4102
rect 3350 4082 3408 4102
rect 3427 4082 3435 4102
rect 3324 4060 3435 4082
rect 3039 4047 3078 4054
rect 3748 4037 3782 4243
rect 4195 4223 4227 4251
rect 3815 4215 4227 4223
rect 3815 4189 3821 4215
rect 3847 4189 4227 4215
rect 3815 4187 4227 4189
rect 3817 4186 3857 4187
rect 4195 4122 4227 4187
rect 5761 4229 5793 4236
rect 5761 4209 5768 4229
rect 5789 4209 5793 4229
rect 5761 4144 5793 4209
rect 6131 4144 6171 4145
rect 5761 4142 6173 4144
rect 4195 4102 4199 4122
rect 4220 4102 4227 4122
rect 4195 4095 4227 4102
rect 4698 4137 4746 4142
rect 4698 4108 4709 4137
rect 4738 4108 4746 4137
rect 3748 4036 3783 4037
rect 3746 4029 3783 4036
rect 2691 4008 2726 4009
rect 2668 4001 2726 4008
rect 2668 3981 2699 4001
rect 2719 3981 2726 4001
rect 2668 3976 2726 3981
rect 3117 4004 3149 4011
rect 3117 3984 3123 4004
rect 3144 3984 3149 4004
rect 2668 3828 2704 3976
rect 3117 3956 3149 3984
rect 2737 3948 3149 3956
rect 2737 3922 2743 3948
rect 2769 3922 3149 3948
rect 3746 4009 3756 4029
rect 3776 4009 3783 4029
rect 3746 4004 3783 4009
rect 4402 4024 4512 4039
rect 4402 4021 4479 4024
rect 3746 3953 3781 4004
rect 4402 3994 4405 4021
rect 4434 3997 4479 4021
rect 4508 3997 4512 4024
rect 4434 3994 4512 3997
rect 4402 3980 4512 3994
rect 4698 3953 4746 4108
rect 5761 4116 6141 4142
rect 6167 4116 6173 4142
rect 5761 4108 6173 4116
rect 5761 4080 5793 4108
rect 6206 4088 6240 4294
rect 6414 4292 6525 4314
rect 6414 4272 6422 4292
rect 6441 4272 6499 4292
rect 6518 4272 6525 4292
rect 6414 4255 6525 4272
rect 6750 4299 6757 4321
rect 6783 4299 6792 4321
rect 6750 4290 6792 4299
rect 5967 4085 6010 4087
rect 5761 4060 5766 4080
rect 5787 4060 5793 4080
rect 5761 4053 5793 4060
rect 5966 4078 6010 4085
rect 5966 4058 5976 4078
rect 5999 4058 6010 4078
rect 5966 4054 6010 4058
rect 6184 4083 6240 4088
rect 6184 4063 6191 4083
rect 6211 4063 6240 4083
rect 6184 4056 6240 4063
rect 6296 4224 6329 4225
rect 6750 4224 6787 4290
rect 6296 4195 6787 4224
rect 6184 4055 6219 4056
rect 3746 3929 4746 3953
rect 5475 3982 5586 4004
rect 5475 3962 5483 3982
rect 5502 3962 5560 3982
rect 5579 3962 5586 3982
rect 5475 3945 5586 3962
rect 5966 3973 6008 4054
rect 6296 3975 6329 4195
rect 6750 4193 6787 4195
rect 6556 4055 6666 4069
rect 6556 4052 6634 4055
rect 6556 4025 6560 4052
rect 6589 4028 6634 4052
rect 6663 4028 6666 4055
rect 6589 4025 6666 4028
rect 6556 4010 6666 4025
rect 6910 4036 6948 4374
rect 7123 4393 7179 4398
rect 7123 4373 7130 4393
rect 7150 4373 7179 4393
rect 7123 4366 7179 4373
rect 7388 4665 7395 4705
rect 7422 4665 7435 4705
rect 7618 4683 7665 4861
rect 8411 4852 8414 4879
rect 8443 4855 8488 4879
rect 8517 4855 8521 4882
rect 8443 4852 8521 4855
rect 8411 4838 8521 4852
rect 7123 4365 7158 4366
rect 7288 4045 7320 4046
rect 6910 4019 6918 4036
rect 6938 4019 6948 4036
rect 6910 4013 6948 4019
rect 7285 4040 7320 4045
rect 7285 4020 7292 4040
rect 7312 4020 7320 4040
rect 7285 4012 7320 4020
rect 6268 3973 6329 3975
rect 5966 3944 6329 3973
rect 6841 3947 6873 3954
rect 5966 3942 6268 3944
rect 3746 3926 4745 3929
rect 6841 3927 6848 3947
rect 6869 3927 6873 3947
rect 3746 3924 3781 3926
rect 2737 3920 3149 3922
rect 2739 3919 2779 3920
rect 2671 3770 2704 3828
rect 2901 3880 2939 3890
rect 2901 3842 2910 3880
rect 2933 3842 2939 3880
rect 2671 3762 2705 3770
rect 2671 3742 2678 3762
rect 2698 3742 2705 3762
rect 2671 3737 2705 3742
rect 2671 3736 2702 3737
rect 2901 3706 2939 3842
rect 3117 3855 3149 3920
rect 6841 3862 6873 3927
rect 7211 3862 7251 3863
rect 6841 3860 7253 3862
rect 6209 3856 6244 3858
rect 3117 3835 3121 3855
rect 3142 3835 3149 3855
rect 5245 3853 6244 3856
rect 3722 3838 4024 3840
rect 3117 3828 3149 3835
rect 3661 3809 4024 3838
rect 3661 3807 3722 3809
rect 3042 3763 3080 3769
rect 3042 3746 3052 3763
rect 3072 3746 3080 3763
rect 2901 3552 2945 3706
rect 2738 3550 2945 3552
rect 2714 3517 2945 3550
rect 1811 2891 1815 2911
rect 1836 2891 1845 2911
rect 1811 2885 1845 2891
rect 1964 3022 2293 3025
rect 2332 3022 2376 3047
rect 1964 2992 2376 3022
rect 1213 2829 1274 2831
rect 911 2800 1274 2829
rect 1755 2816 1787 2823
rect 911 2798 1213 2800
rect 1755 2796 1762 2816
rect 1783 2796 1787 2816
rect 1755 2731 1787 2796
rect 1964 2804 1999 2992
rect 2266 2990 2376 2992
rect 2559 3005 2609 3133
rect 2714 3116 2764 3517
rect 2901 3513 2945 3517
rect 2832 3416 2867 3417
rect 2694 3107 2764 3116
rect 2694 3078 2709 3107
rect 2757 3099 2764 3107
rect 2811 3409 2867 3416
rect 2811 3389 2840 3409
rect 2860 3389 2867 3409
rect 2811 3384 2867 3389
rect 3042 3408 3080 3746
rect 3324 3757 3434 3772
rect 3324 3754 3401 3757
rect 3324 3727 3327 3754
rect 3356 3730 3401 3754
rect 3430 3730 3434 3757
rect 3356 3727 3434 3730
rect 3324 3713 3434 3727
rect 3203 3587 3240 3589
rect 3661 3587 3694 3807
rect 3982 3728 4024 3809
rect 4404 3820 4515 3837
rect 4404 3800 4411 3820
rect 4430 3800 4488 3820
rect 4507 3800 4515 3820
rect 4404 3778 4515 3800
rect 5244 3829 6244 3853
rect 3771 3726 3806 3727
rect 3203 3558 3694 3587
rect 3203 3492 3240 3558
rect 3661 3557 3694 3558
rect 3750 3719 3806 3726
rect 3750 3699 3779 3719
rect 3799 3699 3806 3719
rect 3750 3694 3806 3699
rect 3980 3724 4024 3728
rect 3980 3704 3991 3724
rect 4014 3704 4024 3724
rect 3980 3697 4024 3704
rect 4197 3722 4229 3729
rect 4197 3702 4203 3722
rect 4224 3702 4229 3722
rect 3980 3695 4023 3697
rect 3198 3483 3240 3492
rect 3198 3461 3207 3483
rect 3233 3461 3240 3483
rect 3465 3510 3576 3527
rect 3465 3490 3472 3510
rect 3491 3490 3549 3510
rect 3568 3490 3576 3510
rect 3465 3468 3576 3490
rect 3750 3488 3784 3694
rect 4197 3674 4229 3702
rect 3817 3666 4229 3674
rect 3817 3640 3823 3666
rect 3849 3640 4229 3666
rect 5244 3674 5292 3829
rect 5478 3788 5588 3802
rect 5478 3785 5556 3788
rect 5478 3758 5482 3785
rect 5511 3761 5556 3785
rect 5585 3761 5588 3788
rect 6209 3778 6244 3829
rect 5511 3758 5588 3761
rect 5478 3743 5588 3758
rect 6207 3773 6244 3778
rect 6207 3753 6214 3773
rect 6234 3753 6244 3773
rect 6841 3834 7221 3860
rect 7247 3834 7253 3860
rect 6841 3826 7253 3834
rect 6841 3798 6873 3826
rect 6841 3778 6846 3798
rect 6867 3778 6873 3798
rect 6841 3771 6873 3778
rect 7047 3797 7089 3808
rect 7286 3806 7320 4012
rect 7047 3776 7054 3797
rect 7081 3776 7089 3797
rect 6207 3746 6244 3753
rect 6207 3745 6242 3746
rect 5244 3645 5252 3674
rect 5281 3645 5292 3674
rect 5244 3640 5292 3645
rect 5763 3680 5795 3687
rect 5763 3660 5770 3680
rect 5791 3660 5795 3680
rect 3817 3638 4229 3640
rect 3819 3637 3859 3638
rect 4197 3573 4229 3638
rect 4197 3553 4201 3573
rect 4222 3553 4229 3573
rect 4197 3546 4229 3553
rect 5763 3595 5795 3660
rect 6133 3595 6173 3596
rect 5763 3593 6175 3595
rect 5763 3567 6143 3593
rect 6169 3567 6175 3593
rect 5763 3559 6175 3567
rect 5763 3531 5795 3559
rect 6208 3539 6242 3745
rect 6912 3728 6951 3735
rect 6555 3700 6666 3722
rect 6555 3680 6563 3700
rect 6582 3680 6640 3700
rect 6659 3680 6666 3700
rect 6555 3663 6666 3680
rect 6912 3701 6916 3728
rect 6947 3701 6951 3728
rect 6759 3612 6812 3616
rect 6277 3577 6812 3612
rect 5763 3511 5768 3531
rect 5789 3511 5795 3531
rect 5763 3504 5795 3511
rect 5970 3531 6009 3537
rect 5970 3511 5978 3531
rect 6003 3511 6009 3531
rect 5970 3504 6009 3511
rect 6186 3534 6242 3539
rect 6186 3514 6193 3534
rect 6213 3514 6242 3534
rect 6186 3507 6242 3514
rect 6186 3506 6221 3507
rect 3750 3480 3785 3488
rect 3198 3451 3240 3461
rect 3750 3460 3758 3480
rect 3778 3460 3785 3480
rect 3750 3455 3785 3460
rect 4404 3475 4514 3490
rect 4404 3472 4481 3475
rect 3198 3450 3239 3451
rect 3042 3391 3050 3408
rect 3070 3391 3080 3408
rect 2811 3178 2845 3384
rect 3042 3381 3080 3391
rect 3258 3412 3290 3419
rect 3258 3392 3264 3412
rect 3285 3392 3290 3412
rect 3750 3403 3784 3455
rect 4404 3445 4407 3472
rect 4436 3448 4481 3472
rect 4510 3448 4514 3475
rect 4436 3445 4514 3448
rect 4404 3431 4514 3445
rect 4700 3475 4742 3485
rect 4700 3456 4708 3475
rect 4733 3456 4742 3475
rect 5978 3458 6009 3504
rect 4700 3403 4742 3456
rect 5477 3433 5588 3455
rect 5477 3413 5485 3433
rect 5504 3413 5562 3433
rect 5581 3413 5588 3433
rect 5977 3441 6009 3458
rect 6278 3441 6315 3577
rect 6416 3544 6526 3558
rect 6416 3541 6494 3544
rect 6416 3514 6420 3541
rect 6449 3517 6494 3541
rect 6523 3517 6526 3544
rect 6449 3514 6526 3517
rect 6416 3499 6526 3514
rect 6758 3530 6812 3577
rect 6758 3522 6811 3530
rect 6758 3505 6767 3522
rect 6799 3505 6811 3522
rect 6758 3502 6811 3505
rect 5977 3428 6315 3441
rect 3258 3364 3290 3392
rect 3748 3377 4744 3403
rect 5477 3396 5588 3413
rect 5978 3409 6315 3428
rect 6257 3408 6315 3409
rect 6701 3436 6733 3443
rect 6701 3416 6708 3436
rect 6729 3416 6733 3436
rect 2878 3356 3290 3364
rect 2878 3330 2884 3356
rect 2910 3330 3290 3356
rect 2878 3328 3290 3330
rect 2880 3327 2920 3328
rect 3258 3263 3290 3328
rect 6701 3351 6733 3416
rect 6912 3428 6951 3701
rect 7047 3605 7089 3776
rect 7264 3801 7320 3806
rect 7264 3781 7271 3801
rect 7291 3781 7320 3801
rect 7264 3774 7320 3781
rect 7264 3773 7299 3774
rect 7047 3571 7291 3605
rect 7254 3563 7291 3571
rect 7147 3530 7181 3541
rect 7145 3529 7181 3530
rect 7145 3509 7152 3529
rect 7172 3509 7181 3529
rect 7145 3501 7181 3509
rect 6912 3387 6919 3428
rect 6940 3387 6951 3428
rect 6912 3372 6951 3387
rect 7071 3351 7111 3352
rect 6701 3349 7113 3351
rect 6701 3323 7081 3349
rect 7107 3323 7113 3349
rect 6701 3315 7113 3323
rect 3258 3243 3262 3263
rect 3283 3243 3290 3263
rect 3258 3236 3290 3243
rect 3676 3270 3734 3271
rect 3676 3251 4013 3270
rect 4403 3266 4514 3283
rect 5247 3276 6243 3302
rect 6701 3287 6733 3315
rect 7146 3295 7180 3501
rect 3676 3238 4014 3251
rect 2811 3170 2846 3178
rect 2811 3150 2819 3170
rect 2839 3150 2846 3170
rect 2811 3145 2846 3150
rect 3465 3165 3575 3180
rect 3465 3162 3542 3165
rect 2811 3102 2845 3145
rect 3465 3135 3468 3162
rect 3497 3138 3542 3162
rect 3571 3138 3575 3165
rect 3497 3135 3575 3138
rect 3465 3121 3575 3135
rect 3676 3102 3713 3238
rect 3982 3221 4014 3238
rect 4403 3246 4410 3266
rect 4429 3246 4487 3266
rect 4506 3246 4514 3266
rect 4403 3224 4514 3246
rect 5249 3223 5291 3276
rect 3982 3175 4013 3221
rect 5249 3204 5258 3223
rect 5283 3204 5291 3223
rect 5249 3194 5291 3204
rect 5477 3234 5587 3248
rect 5477 3231 5555 3234
rect 5477 3204 5481 3231
rect 5510 3207 5555 3231
rect 5584 3207 5587 3234
rect 6207 3224 6241 3276
rect 6701 3267 6706 3287
rect 6727 3267 6733 3287
rect 6701 3260 6733 3267
rect 7124 3290 7180 3295
rect 7124 3270 7131 3290
rect 7151 3270 7180 3290
rect 7124 3263 7180 3270
rect 7124 3262 7159 3263
rect 6752 3228 6793 3229
rect 5510 3204 5587 3207
rect 5477 3189 5587 3204
rect 6206 3219 6241 3224
rect 6206 3199 6213 3219
rect 6233 3199 6241 3219
rect 6751 3218 6793 3228
rect 6206 3191 6241 3199
rect 3770 3172 3805 3173
rect 3749 3165 3805 3172
rect 3749 3145 3778 3165
rect 3798 3145 3805 3165
rect 3749 3140 3805 3145
rect 3982 3168 4021 3175
rect 3982 3148 3988 3168
rect 4013 3148 4021 3168
rect 3982 3142 4021 3148
rect 4196 3168 4228 3175
rect 4196 3148 4202 3168
rect 4223 3148 4228 3168
rect 2757 3078 2762 3099
rect 2694 3067 2762 3078
rect 2810 3067 3714 3102
rect 2811 3066 2845 3067
rect 2559 2971 2974 3005
rect 2559 2969 2609 2971
rect 2192 2907 2242 2914
rect 2192 2893 2206 2907
rect 2198 2889 2206 2893
rect 2226 2893 2242 2907
rect 2226 2889 2236 2893
rect 2722 2892 2757 2893
rect 2198 2882 2236 2889
rect 2701 2885 2757 2892
rect 2199 2881 2234 2882
rect 1964 2772 1969 2804
rect 1996 2772 1999 2804
rect 1964 2754 1999 2772
rect 2125 2731 2165 2732
rect 1755 2729 2167 2731
rect 1153 2712 1188 2714
rect 189 2709 1188 2712
rect 188 2685 1188 2709
rect 188 2530 236 2685
rect 422 2644 532 2658
rect 422 2641 500 2644
rect 422 2614 426 2641
rect 455 2617 500 2641
rect 529 2617 532 2644
rect 1153 2634 1188 2685
rect 1755 2703 2135 2729
rect 2161 2703 2167 2729
rect 1755 2695 2167 2703
rect 1755 2667 1787 2695
rect 2200 2675 2234 2881
rect 1755 2647 1760 2667
rect 1781 2647 1787 2667
rect 1755 2640 1787 2647
rect 2178 2670 2234 2675
rect 2178 2650 2185 2670
rect 2205 2650 2234 2670
rect 2701 2865 2730 2885
rect 2750 2865 2757 2885
rect 2701 2860 2757 2865
rect 2929 2888 2974 2971
rect 3355 2986 3466 3003
rect 3355 2966 3362 2986
rect 3381 2966 3439 2986
rect 3458 2966 3466 2986
rect 3355 2944 3466 2966
rect 3749 2934 3783 3140
rect 4196 3120 4228 3148
rect 3816 3112 4228 3120
rect 3816 3086 3822 3112
rect 3848 3086 4228 3112
rect 3816 3084 4228 3086
rect 3818 3083 3858 3084
rect 4196 3019 4228 3084
rect 5762 3126 5794 3133
rect 5762 3106 5769 3126
rect 5790 3106 5794 3126
rect 5762 3041 5794 3106
rect 6132 3041 6172 3042
rect 5762 3039 6174 3041
rect 4196 2999 4200 3019
rect 4221 2999 4228 3019
rect 4196 2992 4228 2999
rect 4699 3034 4747 3039
rect 4699 3005 4710 3034
rect 4739 3005 4747 3034
rect 3749 2933 3784 2934
rect 3747 2926 3784 2933
rect 3747 2906 3757 2926
rect 3777 2906 3784 2926
rect 3747 2901 3784 2906
rect 4403 2921 4513 2936
rect 4403 2918 4480 2921
rect 2929 2869 2938 2888
rect 2967 2869 2974 2888
rect 2701 2654 2735 2860
rect 2929 2857 2974 2869
rect 3148 2888 3180 2895
rect 3148 2868 3154 2888
rect 3175 2868 3180 2888
rect 3148 2840 3180 2868
rect 2768 2832 3180 2840
rect 2768 2806 2774 2832
rect 2800 2806 3180 2832
rect 3747 2850 3782 2901
rect 4403 2891 4406 2918
rect 4435 2894 4480 2918
rect 4509 2894 4513 2921
rect 4435 2891 4513 2894
rect 4403 2877 4513 2891
rect 4699 2850 4747 3005
rect 5762 3013 6142 3039
rect 6168 3013 6174 3039
rect 5762 3005 6174 3013
rect 5762 2977 5794 3005
rect 6207 2985 6241 3191
rect 6415 3189 6526 3211
rect 6415 3169 6423 3189
rect 6442 3169 6500 3189
rect 6519 3169 6526 3189
rect 6415 3152 6526 3169
rect 6751 3196 6758 3218
rect 6784 3196 6793 3218
rect 6751 3187 6793 3196
rect 5968 2982 6011 2984
rect 5762 2957 5767 2977
rect 5788 2957 5794 2977
rect 5762 2950 5794 2957
rect 5967 2975 6011 2982
rect 5967 2955 5977 2975
rect 6000 2955 6011 2975
rect 5967 2951 6011 2955
rect 6185 2980 6241 2985
rect 6185 2960 6192 2980
rect 6212 2960 6241 2980
rect 6185 2953 6241 2960
rect 6297 3121 6330 3122
rect 6751 3121 6788 3187
rect 7254 3172 7292 3563
rect 6868 3156 7292 3172
rect 6297 3092 6788 3121
rect 6185 2952 6220 2953
rect 3747 2826 4747 2850
rect 5476 2879 5587 2901
rect 5476 2859 5484 2879
rect 5503 2859 5561 2879
rect 5580 2859 5587 2879
rect 5476 2843 5587 2859
rect 5967 2870 6009 2951
rect 6297 2872 6330 3092
rect 6751 3090 6788 3092
rect 6867 3131 7292 3156
rect 6526 2965 6636 2979
rect 6526 2962 6604 2965
rect 6526 2935 6530 2962
rect 6559 2938 6604 2962
rect 6633 2938 6636 2965
rect 6559 2935 6636 2938
rect 6526 2920 6636 2935
rect 6867 2952 6901 3131
rect 7388 3088 7435 4665
rect 7617 4659 7665 4683
rect 8258 4731 8295 4733
rect 8716 4731 8749 4951
rect 9037 4872 9079 4953
rect 9459 4964 9570 4981
rect 9459 4944 9466 4964
rect 9485 4944 9543 4964
rect 9562 4944 9570 4964
rect 9459 4922 9570 4944
rect 8826 4870 8861 4871
rect 8258 4702 8749 4731
rect 7617 3174 7663 4659
rect 8258 4636 8295 4702
rect 8716 4701 8749 4702
rect 8805 4863 8861 4870
rect 8805 4843 8834 4863
rect 8854 4843 8861 4863
rect 8805 4838 8861 4843
rect 9035 4868 9079 4872
rect 9035 4848 9046 4868
rect 9069 4848 9079 4868
rect 9035 4841 9079 4848
rect 9252 4866 9284 4873
rect 9252 4846 9258 4866
rect 9279 4846 9284 4866
rect 9035 4839 9078 4841
rect 8253 4627 8295 4636
rect 8253 4605 8262 4627
rect 8288 4605 8295 4627
rect 8520 4654 8631 4671
rect 8520 4634 8527 4654
rect 8546 4634 8604 4654
rect 8623 4634 8631 4654
rect 8520 4612 8631 4634
rect 8805 4632 8839 4838
rect 9252 4818 9284 4846
rect 8872 4810 9284 4818
rect 8872 4784 8878 4810
rect 8904 4784 9284 4810
rect 8872 4782 9284 4784
rect 8874 4781 8914 4782
rect 9252 4717 9284 4782
rect 9252 4697 9256 4717
rect 9277 4697 9284 4717
rect 9252 4690 9284 4697
rect 8805 4624 8840 4632
rect 8253 4595 8295 4605
rect 8805 4604 8813 4624
rect 8833 4604 8840 4624
rect 8805 4599 8840 4604
rect 9459 4619 9569 4634
rect 9459 4616 9536 4619
rect 8253 4594 8294 4595
rect 7887 4560 7922 4561
rect 7866 4553 7922 4560
rect 7866 4533 7895 4553
rect 7915 4533 7922 4553
rect 7866 4528 7922 4533
rect 8313 4556 8345 4563
rect 8313 4536 8319 4556
rect 8340 4536 8345 4556
rect 8805 4547 8839 4599
rect 9459 4589 9462 4616
rect 9491 4592 9536 4616
rect 9565 4592 9569 4619
rect 9491 4589 9569 4592
rect 9459 4575 9569 4589
rect 9755 4619 9797 4629
rect 9755 4600 9763 4619
rect 9788 4600 9797 4619
rect 9755 4547 9797 4600
rect 7866 4322 7900 4528
rect 8313 4508 8345 4536
rect 8803 4521 9799 4547
rect 7933 4500 8345 4508
rect 7933 4474 7939 4500
rect 7965 4474 8345 4500
rect 7933 4472 8345 4474
rect 7935 4471 7975 4472
rect 8095 4436 8134 4451
rect 8095 4395 8106 4436
rect 8127 4395 8134 4436
rect 7865 4314 7901 4322
rect 7865 4294 7874 4314
rect 7894 4294 7901 4314
rect 7865 4293 7901 4294
rect 7865 4282 7899 4293
rect 8095 4122 8134 4395
rect 8313 4407 8345 4472
rect 8313 4387 8317 4407
rect 8338 4387 8345 4407
rect 8313 4380 8345 4387
rect 8731 4414 8789 4415
rect 8731 4395 9068 4414
rect 9458 4410 9569 4427
rect 8731 4382 9069 4395
rect 8235 4318 8288 4321
rect 8235 4301 8247 4318
rect 8279 4301 8288 4318
rect 8235 4293 8288 4301
rect 8234 4246 8288 4293
rect 8520 4309 8630 4324
rect 8520 4306 8597 4309
rect 8520 4279 8523 4306
rect 8552 4282 8597 4306
rect 8626 4282 8630 4309
rect 8552 4279 8630 4282
rect 8520 4265 8630 4279
rect 8731 4246 8768 4382
rect 9037 4365 9069 4382
rect 9458 4390 9465 4410
rect 9484 4390 9542 4410
rect 9561 4390 9569 4410
rect 9458 4368 9569 4390
rect 9037 4319 9068 4365
rect 8825 4316 8860 4317
rect 8804 4309 8860 4316
rect 8804 4289 8833 4309
rect 8853 4289 8860 4309
rect 8804 4284 8860 4289
rect 9037 4312 9076 4319
rect 9037 4292 9043 4312
rect 9068 4292 9076 4312
rect 9037 4286 9076 4292
rect 9251 4312 9283 4319
rect 9251 4292 9257 4312
rect 9278 4292 9283 4312
rect 8234 4211 8769 4246
rect 8234 4207 8287 4211
rect 8095 4095 8099 4122
rect 8130 4095 8134 4122
rect 8380 4143 8491 4160
rect 8380 4123 8387 4143
rect 8406 4123 8464 4143
rect 8483 4123 8491 4143
rect 8380 4101 8491 4123
rect 8095 4088 8134 4095
rect 8804 4078 8838 4284
rect 9251 4264 9283 4292
rect 8871 4256 9283 4264
rect 8871 4230 8877 4256
rect 8903 4230 9283 4256
rect 8871 4228 9283 4230
rect 8873 4227 8913 4228
rect 9251 4163 9283 4228
rect 9251 4143 9255 4163
rect 9276 4143 9283 4163
rect 9251 4136 9283 4143
rect 9754 4178 9802 4183
rect 9754 4149 9765 4178
rect 9794 4149 9802 4178
rect 8804 4077 8839 4078
rect 8802 4070 8839 4077
rect 7747 4049 7782 4050
rect 7724 4042 7782 4049
rect 7724 4022 7755 4042
rect 7775 4022 7782 4042
rect 7724 4017 7782 4022
rect 8173 4045 8205 4052
rect 8173 4025 8179 4045
rect 8200 4025 8205 4045
rect 7724 3869 7760 4017
rect 8173 3997 8205 4025
rect 7793 3989 8205 3997
rect 7793 3963 7799 3989
rect 7825 3963 8205 3989
rect 8802 4050 8812 4070
rect 8832 4050 8839 4070
rect 8802 4045 8839 4050
rect 9458 4065 9568 4080
rect 9458 4062 9535 4065
rect 8802 3994 8837 4045
rect 9458 4035 9461 4062
rect 9490 4038 9535 4062
rect 9564 4038 9568 4065
rect 9490 4035 9568 4038
rect 9458 4021 9568 4035
rect 9754 3994 9802 4149
rect 8802 3970 9802 3994
rect 8802 3967 9801 3970
rect 8802 3965 8837 3967
rect 7793 3961 8205 3963
rect 7795 3960 7835 3961
rect 7727 3811 7760 3869
rect 7957 3921 7995 3931
rect 7957 3883 7966 3921
rect 7989 3883 7995 3921
rect 7727 3803 7761 3811
rect 7727 3783 7734 3803
rect 7754 3783 7761 3803
rect 7727 3778 7761 3783
rect 7727 3777 7758 3778
rect 7957 3747 7995 3883
rect 8173 3896 8205 3961
rect 8173 3876 8177 3896
rect 8198 3876 8205 3896
rect 8778 3879 9080 3881
rect 8173 3869 8205 3876
rect 8717 3850 9080 3879
rect 8717 3848 8778 3850
rect 8098 3804 8136 3810
rect 8098 3787 8108 3804
rect 8128 3787 8136 3804
rect 7957 3593 8001 3747
rect 7794 3591 8001 3593
rect 7770 3558 8001 3591
rect 6867 2932 6871 2952
rect 6892 2932 6901 2952
rect 6867 2926 6901 2932
rect 7020 3063 7349 3066
rect 7388 3063 7432 3088
rect 7020 3033 7432 3063
rect 6269 2870 6330 2872
rect 5967 2841 6330 2870
rect 6811 2857 6843 2864
rect 5967 2839 6269 2841
rect 6811 2837 6818 2857
rect 6839 2837 6843 2857
rect 3747 2823 4746 2826
rect 3747 2821 3782 2823
rect 2768 2804 3180 2806
rect 2770 2803 2810 2804
rect 3148 2739 3180 2804
rect 6811 2772 6843 2837
rect 7020 2845 7055 3033
rect 7322 3031 7432 3033
rect 7615 3046 7665 3174
rect 7770 3157 7820 3558
rect 7957 3554 8001 3558
rect 7888 3457 7923 3458
rect 7750 3148 7820 3157
rect 7750 3119 7765 3148
rect 7813 3140 7820 3148
rect 7867 3450 7923 3457
rect 7867 3430 7896 3450
rect 7916 3430 7923 3450
rect 7867 3425 7923 3430
rect 8098 3449 8136 3787
rect 8380 3798 8490 3813
rect 8380 3795 8457 3798
rect 8380 3768 8383 3795
rect 8412 3771 8457 3795
rect 8486 3771 8490 3798
rect 8412 3768 8490 3771
rect 8380 3754 8490 3768
rect 8259 3628 8296 3630
rect 8717 3628 8750 3848
rect 9038 3769 9080 3850
rect 9460 3861 9571 3878
rect 9460 3841 9467 3861
rect 9486 3841 9544 3861
rect 9563 3841 9571 3861
rect 9460 3819 9571 3841
rect 8827 3767 8862 3768
rect 8259 3599 8750 3628
rect 8259 3533 8296 3599
rect 8717 3598 8750 3599
rect 8806 3760 8862 3767
rect 8806 3740 8835 3760
rect 8855 3740 8862 3760
rect 8806 3735 8862 3740
rect 9036 3765 9080 3769
rect 9036 3745 9047 3765
rect 9070 3745 9080 3765
rect 9036 3738 9080 3745
rect 9253 3763 9285 3770
rect 9253 3743 9259 3763
rect 9280 3743 9285 3763
rect 9036 3736 9079 3738
rect 8254 3524 8296 3533
rect 8254 3502 8263 3524
rect 8289 3502 8296 3524
rect 8521 3551 8632 3568
rect 8521 3531 8528 3551
rect 8547 3531 8605 3551
rect 8624 3531 8632 3551
rect 8521 3509 8632 3531
rect 8806 3529 8840 3735
rect 9253 3715 9285 3743
rect 8873 3707 9285 3715
rect 8873 3681 8879 3707
rect 8905 3681 9285 3707
rect 8873 3679 9285 3681
rect 8875 3678 8915 3679
rect 9253 3614 9285 3679
rect 9253 3594 9257 3614
rect 9278 3594 9285 3614
rect 9253 3587 9285 3594
rect 8806 3521 8841 3529
rect 8254 3492 8296 3502
rect 8806 3501 8814 3521
rect 8834 3501 8841 3521
rect 8806 3496 8841 3501
rect 9460 3516 9570 3531
rect 9460 3513 9537 3516
rect 8254 3491 8295 3492
rect 8098 3432 8106 3449
rect 8126 3432 8136 3449
rect 7867 3219 7901 3425
rect 8098 3422 8136 3432
rect 8314 3453 8346 3460
rect 8314 3433 8320 3453
rect 8341 3433 8346 3453
rect 8806 3444 8840 3496
rect 9460 3486 9463 3513
rect 9492 3489 9537 3513
rect 9566 3489 9570 3516
rect 9492 3486 9570 3489
rect 9460 3472 9570 3486
rect 9756 3516 9798 3526
rect 9756 3497 9764 3516
rect 9789 3497 9798 3516
rect 9756 3444 9798 3497
rect 8314 3405 8346 3433
rect 8804 3418 9800 3444
rect 7934 3397 8346 3405
rect 7934 3371 7940 3397
rect 7966 3371 8346 3397
rect 7934 3369 8346 3371
rect 7936 3368 7976 3369
rect 8314 3304 8346 3369
rect 8314 3284 8318 3304
rect 8339 3284 8346 3304
rect 8314 3277 8346 3284
rect 8732 3311 8790 3312
rect 8732 3292 9069 3311
rect 9459 3307 9570 3324
rect 8732 3279 9070 3292
rect 7867 3211 7902 3219
rect 7867 3191 7875 3211
rect 7895 3191 7902 3211
rect 7867 3186 7902 3191
rect 8521 3206 8631 3221
rect 8521 3203 8598 3206
rect 7867 3143 7901 3186
rect 8521 3176 8524 3203
rect 8553 3179 8598 3203
rect 8627 3179 8631 3206
rect 8553 3176 8631 3179
rect 8521 3162 8631 3176
rect 8732 3143 8769 3279
rect 9038 3262 9070 3279
rect 9459 3287 9466 3307
rect 9485 3287 9543 3307
rect 9562 3287 9570 3307
rect 9459 3265 9570 3287
rect 9038 3216 9069 3262
rect 8826 3213 8861 3214
rect 8805 3206 8861 3213
rect 8805 3186 8834 3206
rect 8854 3186 8861 3206
rect 8805 3181 8861 3186
rect 9038 3209 9077 3216
rect 9038 3189 9044 3209
rect 9069 3189 9077 3209
rect 9038 3183 9077 3189
rect 9252 3209 9284 3216
rect 9252 3189 9258 3209
rect 9279 3189 9284 3209
rect 7813 3119 7818 3140
rect 7750 3108 7818 3119
rect 7866 3108 8770 3143
rect 7867 3107 7901 3108
rect 7615 3012 8030 3046
rect 7615 3010 7665 3012
rect 7248 2948 7298 2955
rect 7248 2934 7262 2948
rect 7254 2930 7262 2934
rect 7282 2934 7298 2948
rect 7282 2930 7292 2934
rect 7778 2933 7813 2934
rect 7254 2923 7292 2930
rect 7757 2926 7813 2933
rect 7255 2922 7290 2923
rect 7020 2813 7025 2845
rect 7052 2813 7055 2845
rect 7020 2795 7055 2813
rect 7181 2772 7221 2773
rect 6811 2770 7223 2772
rect 6209 2753 6244 2755
rect 5245 2750 6244 2753
rect 3148 2719 3152 2739
rect 3173 2719 3180 2739
rect 3722 2735 4024 2737
rect 3148 2712 3180 2719
rect 3661 2706 4024 2735
rect 3661 2704 3722 2706
rect 2701 2653 2736 2654
rect 2178 2643 2234 2650
rect 2699 2646 2737 2653
rect 2178 2642 2213 2643
rect 455 2614 532 2617
rect 422 2599 532 2614
rect 1151 2629 1188 2634
rect 1151 2609 1158 2629
rect 1178 2609 1188 2629
rect 2699 2626 2709 2646
rect 2729 2626 2737 2646
rect 1151 2602 1188 2609
rect 2173 2604 2243 2614
rect 1151 2601 1186 2602
rect 188 2501 196 2530
rect 225 2501 236 2530
rect 188 2496 236 2501
rect 707 2536 739 2543
rect 707 2516 714 2536
rect 735 2516 739 2536
rect 707 2451 739 2516
rect 1077 2451 1117 2452
rect 707 2449 1119 2451
rect 707 2423 1087 2449
rect 1113 2423 1119 2449
rect 707 2415 1119 2423
rect 707 2387 739 2415
rect 1152 2395 1186 2601
rect 2171 2597 2243 2604
rect 1469 2569 1580 2591
rect 1469 2549 1477 2569
rect 1496 2549 1554 2569
rect 1573 2549 1580 2569
rect 1469 2532 1580 2549
rect 2171 2568 2178 2597
rect 2226 2568 2243 2597
rect 2171 2559 2243 2568
rect 2090 2468 2124 2469
rect 1221 2433 2125 2468
rect 707 2367 712 2387
rect 733 2367 739 2387
rect 707 2360 739 2367
rect 914 2387 953 2393
rect 914 2367 922 2387
rect 947 2367 953 2387
rect 914 2360 953 2367
rect 1130 2390 1186 2395
rect 1130 2370 1137 2390
rect 1157 2370 1186 2390
rect 1130 2363 1186 2370
rect 1130 2362 1165 2363
rect 922 2314 953 2360
rect 421 2289 532 2311
rect 421 2269 429 2289
rect 448 2269 506 2289
rect 525 2269 532 2289
rect 921 2297 953 2314
rect 1222 2297 1259 2433
rect 1360 2400 1470 2414
rect 1360 2397 1438 2400
rect 1360 2370 1364 2397
rect 1393 2373 1438 2397
rect 1467 2373 1470 2400
rect 2090 2390 2124 2433
rect 1393 2370 1470 2373
rect 1360 2355 1470 2370
rect 2089 2385 2124 2390
rect 2089 2365 2096 2385
rect 2116 2365 2124 2385
rect 2089 2357 2124 2365
rect 921 2284 1259 2297
rect 421 2252 532 2269
rect 922 2265 1259 2284
rect 1201 2264 1259 2265
rect 1645 2292 1677 2299
rect 1645 2272 1652 2292
rect 1673 2272 1677 2292
rect 1645 2207 1677 2272
rect 2015 2207 2055 2208
rect 1645 2205 2057 2207
rect 1645 2179 2025 2205
rect 2051 2179 2057 2205
rect 1645 2171 2057 2179
rect 191 2132 1187 2158
rect 1645 2143 1677 2171
rect 193 2079 235 2132
rect 193 2060 202 2079
rect 227 2060 235 2079
rect 193 2050 235 2060
rect 421 2090 531 2104
rect 421 2087 499 2090
rect 421 2060 425 2087
rect 454 2063 499 2087
rect 528 2063 531 2090
rect 1151 2080 1185 2132
rect 1645 2123 1650 2143
rect 1671 2123 1677 2143
rect 1645 2116 1677 2123
rect 1855 2144 1893 2154
rect 2090 2151 2124 2357
rect 1855 2127 1865 2144
rect 1885 2127 1893 2144
rect 1696 2084 1737 2085
rect 454 2060 531 2063
rect 421 2045 531 2060
rect 1150 2075 1185 2080
rect 1150 2055 1157 2075
rect 1177 2055 1185 2075
rect 1695 2074 1737 2084
rect 1150 2047 1185 2055
rect 706 1982 738 1989
rect 706 1962 713 1982
rect 734 1962 738 1982
rect 706 1897 738 1962
rect 1076 1897 1116 1898
rect 706 1895 1118 1897
rect 706 1869 1086 1895
rect 1112 1869 1118 1895
rect 706 1861 1118 1869
rect 706 1833 738 1861
rect 1151 1841 1185 2047
rect 1359 2045 1470 2067
rect 1359 2025 1367 2045
rect 1386 2025 1444 2045
rect 1463 2025 1470 2045
rect 1359 2008 1470 2025
rect 1695 2052 1702 2074
rect 1728 2052 1737 2074
rect 1695 2043 1737 2052
rect 912 1838 955 1840
rect 706 1813 711 1833
rect 732 1813 738 1833
rect 706 1806 738 1813
rect 911 1831 955 1838
rect 911 1811 921 1831
rect 944 1811 955 1831
rect 911 1807 955 1811
rect 1129 1836 1185 1841
rect 1129 1816 1136 1836
rect 1156 1816 1185 1836
rect 1129 1809 1185 1816
rect 1241 1977 1274 1978
rect 1695 1977 1732 2043
rect 1241 1948 1732 1977
rect 1129 1808 1164 1809
rect 420 1735 531 1757
rect 420 1715 428 1735
rect 447 1715 505 1735
rect 524 1715 531 1735
rect 420 1698 531 1715
rect 911 1726 953 1807
rect 1241 1728 1274 1948
rect 1695 1946 1732 1948
rect 1501 1808 1611 1822
rect 1501 1805 1579 1808
rect 1501 1778 1505 1805
rect 1534 1781 1579 1805
rect 1608 1781 1611 1808
rect 1534 1778 1611 1781
rect 1501 1763 1611 1778
rect 1855 1789 1893 2127
rect 2068 2146 2124 2151
rect 2068 2126 2075 2146
rect 2095 2126 2124 2146
rect 2068 2119 2124 2126
rect 2068 2118 2103 2119
rect 1990 2018 2034 2022
rect 2171 2018 2221 2559
rect 1990 1985 2221 2018
rect 2699 2013 2737 2626
rect 3355 2641 3465 2656
rect 3355 2638 3432 2641
rect 3355 2611 3358 2638
rect 3387 2614 3432 2638
rect 3461 2614 3465 2641
rect 3387 2611 3465 2614
rect 3355 2597 3465 2611
rect 3203 2484 3240 2486
rect 3661 2484 3694 2704
rect 3982 2625 4024 2706
rect 4404 2717 4515 2733
rect 4404 2697 4411 2717
rect 4430 2697 4488 2717
rect 4507 2697 4515 2717
rect 4404 2675 4515 2697
rect 5244 2726 6244 2750
rect 3771 2623 3806 2624
rect 3203 2455 3694 2484
rect 3203 2389 3240 2455
rect 3661 2454 3694 2455
rect 3750 2616 3806 2623
rect 3750 2596 3779 2616
rect 3799 2596 3806 2616
rect 3750 2591 3806 2596
rect 3980 2621 4024 2625
rect 3980 2601 3991 2621
rect 4014 2601 4024 2621
rect 3980 2594 4024 2601
rect 4197 2619 4229 2626
rect 4197 2599 4203 2619
rect 4224 2599 4229 2619
rect 3980 2592 4023 2594
rect 3198 2380 3240 2389
rect 3198 2358 3207 2380
rect 3233 2358 3240 2380
rect 3465 2407 3576 2424
rect 3465 2387 3472 2407
rect 3491 2387 3549 2407
rect 3568 2387 3576 2407
rect 3465 2365 3576 2387
rect 3750 2385 3784 2591
rect 4197 2571 4229 2599
rect 3817 2563 4229 2571
rect 3817 2537 3823 2563
rect 3849 2537 4229 2563
rect 5244 2571 5292 2726
rect 5478 2685 5588 2699
rect 5478 2682 5556 2685
rect 5478 2655 5482 2682
rect 5511 2658 5556 2682
rect 5585 2658 5588 2685
rect 6209 2675 6244 2726
rect 6811 2744 7191 2770
rect 7217 2744 7223 2770
rect 6811 2736 7223 2744
rect 6811 2708 6843 2736
rect 7256 2716 7290 2922
rect 6811 2688 6816 2708
rect 6837 2688 6843 2708
rect 6811 2681 6843 2688
rect 7234 2711 7290 2716
rect 7234 2691 7241 2711
rect 7261 2691 7290 2711
rect 7757 2906 7786 2926
rect 7806 2906 7813 2926
rect 7757 2901 7813 2906
rect 7985 2929 8030 3012
rect 8411 3027 8522 3044
rect 8411 3007 8418 3027
rect 8437 3007 8495 3027
rect 8514 3007 8522 3027
rect 8411 2985 8522 3007
rect 8805 2975 8839 3181
rect 9252 3161 9284 3189
rect 8872 3153 9284 3161
rect 8872 3127 8878 3153
rect 8904 3127 9284 3153
rect 8872 3125 9284 3127
rect 8874 3124 8914 3125
rect 9252 3060 9284 3125
rect 9252 3040 9256 3060
rect 9277 3040 9284 3060
rect 9252 3033 9284 3040
rect 9755 3075 9803 3080
rect 9755 3046 9766 3075
rect 9795 3046 9803 3075
rect 8805 2974 8840 2975
rect 8803 2967 8840 2974
rect 8803 2947 8813 2967
rect 8833 2947 8840 2967
rect 8803 2942 8840 2947
rect 9459 2962 9569 2977
rect 9459 2959 9536 2962
rect 7985 2910 7994 2929
rect 8023 2910 8030 2929
rect 7757 2695 7791 2901
rect 7985 2898 8030 2910
rect 8204 2929 8236 2936
rect 8204 2909 8210 2929
rect 8231 2909 8236 2929
rect 8204 2881 8236 2909
rect 7824 2873 8236 2881
rect 7824 2847 7830 2873
rect 7856 2847 8236 2873
rect 8803 2891 8838 2942
rect 9459 2932 9462 2959
rect 9491 2935 9536 2959
rect 9565 2935 9569 2962
rect 9491 2932 9569 2935
rect 9459 2918 9569 2932
rect 9755 2891 9803 3046
rect 8803 2867 9803 2891
rect 8803 2864 9802 2867
rect 8803 2862 8838 2864
rect 7824 2845 8236 2847
rect 7826 2844 7866 2845
rect 8204 2780 8236 2845
rect 8204 2760 8208 2780
rect 8229 2760 8236 2780
rect 8778 2776 9080 2778
rect 8204 2753 8236 2760
rect 8717 2747 9080 2776
rect 8717 2745 8778 2747
rect 7757 2694 7792 2695
rect 7234 2684 7290 2691
rect 7755 2687 7793 2694
rect 7234 2683 7269 2684
rect 5511 2655 5588 2658
rect 5478 2640 5588 2655
rect 6207 2670 6244 2675
rect 6207 2650 6214 2670
rect 6234 2650 6244 2670
rect 7755 2667 7765 2687
rect 7785 2667 7793 2687
rect 6207 2643 6244 2650
rect 7229 2645 7299 2655
rect 6207 2642 6242 2643
rect 5244 2542 5252 2571
rect 5281 2542 5292 2571
rect 5244 2537 5292 2542
rect 5763 2577 5795 2584
rect 5763 2557 5770 2577
rect 5791 2557 5795 2577
rect 3817 2535 4229 2537
rect 3819 2534 3859 2535
rect 4197 2470 4229 2535
rect 4197 2450 4201 2470
rect 4222 2450 4229 2470
rect 4197 2443 4229 2450
rect 5763 2492 5795 2557
rect 6133 2492 6173 2493
rect 5763 2490 6175 2492
rect 5763 2464 6143 2490
rect 6169 2464 6175 2490
rect 5763 2456 6175 2464
rect 5763 2428 5795 2456
rect 6208 2436 6242 2642
rect 7227 2638 7299 2645
rect 6525 2610 6636 2632
rect 6525 2590 6533 2610
rect 6552 2590 6610 2610
rect 6629 2590 6636 2610
rect 6525 2573 6636 2590
rect 7227 2609 7234 2638
rect 7282 2609 7299 2638
rect 7227 2600 7299 2609
rect 7146 2509 7180 2510
rect 6277 2474 7181 2509
rect 5763 2408 5768 2428
rect 5789 2408 5795 2428
rect 5763 2401 5795 2408
rect 5970 2428 6009 2434
rect 5970 2408 5978 2428
rect 6003 2408 6009 2428
rect 5970 2401 6009 2408
rect 6186 2431 6242 2436
rect 6186 2411 6193 2431
rect 6213 2411 6242 2431
rect 6186 2404 6242 2411
rect 6186 2403 6221 2404
rect 3750 2377 3785 2385
rect 3198 2348 3240 2358
rect 3750 2357 3758 2377
rect 3778 2357 3785 2377
rect 3750 2352 3785 2357
rect 4404 2372 4514 2387
rect 4404 2369 4481 2372
rect 3198 2347 3239 2348
rect 2832 2313 2867 2314
rect 2811 2306 2867 2313
rect 2811 2286 2840 2306
rect 2860 2286 2867 2306
rect 2811 2281 2867 2286
rect 3258 2309 3290 2316
rect 3258 2289 3264 2309
rect 3285 2289 3290 2309
rect 3750 2300 3784 2352
rect 4404 2342 4407 2369
rect 4436 2345 4481 2369
rect 4510 2345 4514 2372
rect 4436 2342 4514 2345
rect 4404 2328 4514 2342
rect 4700 2372 4742 2382
rect 4700 2353 4708 2372
rect 4733 2353 4742 2372
rect 5978 2355 6009 2401
rect 4700 2300 4742 2353
rect 5477 2330 5588 2352
rect 5477 2310 5485 2330
rect 5504 2310 5562 2330
rect 5581 2310 5588 2330
rect 5977 2338 6009 2355
rect 6278 2338 6315 2474
rect 6416 2441 6526 2455
rect 6416 2438 6494 2441
rect 6416 2411 6420 2438
rect 6449 2414 6494 2438
rect 6523 2414 6526 2441
rect 7146 2431 7180 2474
rect 6449 2411 6526 2414
rect 6416 2396 6526 2411
rect 7145 2426 7180 2431
rect 7145 2406 7152 2426
rect 7172 2406 7180 2426
rect 7145 2398 7180 2406
rect 5977 2325 6315 2338
rect 2811 2075 2845 2281
rect 3258 2261 3290 2289
rect 3748 2274 4744 2300
rect 5477 2293 5588 2310
rect 5978 2306 6315 2325
rect 6257 2305 6315 2306
rect 6701 2333 6733 2340
rect 6701 2313 6708 2333
rect 6729 2313 6733 2333
rect 2878 2253 3290 2261
rect 2878 2227 2884 2253
rect 2910 2227 3290 2253
rect 2878 2225 3290 2227
rect 2880 2224 2920 2225
rect 3040 2189 3079 2204
rect 3040 2148 3051 2189
rect 3072 2148 3079 2189
rect 2810 2067 2846 2075
rect 2810 2047 2819 2067
rect 2839 2047 2846 2067
rect 2810 2046 2846 2047
rect 2810 2035 2844 2046
rect 2700 2005 2737 2013
rect 1990 1983 2197 1985
rect 1990 1829 2034 1983
rect 2700 1971 2944 2005
rect 1855 1772 1863 1789
rect 1883 1772 1893 1789
rect 1855 1766 1893 1772
rect 1213 1726 1274 1728
rect 911 1697 1274 1726
rect 1786 1700 1818 1707
rect 911 1695 1213 1697
rect 1786 1680 1793 1700
rect 1814 1680 1818 1700
rect 1786 1615 1818 1680
rect 1996 1693 2034 1829
rect 2692 1802 2727 1803
rect 2233 1798 2264 1799
rect 2230 1793 2264 1798
rect 2230 1773 2237 1793
rect 2257 1773 2264 1793
rect 2230 1765 2264 1773
rect 1996 1655 2002 1693
rect 2025 1655 2034 1693
rect 1996 1645 2034 1655
rect 2231 1707 2264 1765
rect 2671 1795 2727 1802
rect 2671 1775 2700 1795
rect 2720 1775 2727 1795
rect 2671 1770 2727 1775
rect 2902 1800 2944 1971
rect 3040 1875 3079 2148
rect 3258 2160 3290 2225
rect 6701 2248 6733 2313
rect 7071 2248 7111 2249
rect 6701 2246 7113 2248
rect 6701 2220 7081 2246
rect 7107 2220 7113 2246
rect 6701 2212 7113 2220
rect 3258 2140 3262 2160
rect 3283 2140 3290 2160
rect 3258 2133 3290 2140
rect 3676 2167 3734 2168
rect 3676 2148 4013 2167
rect 4403 2163 4514 2180
rect 5247 2173 6243 2199
rect 6701 2184 6733 2212
rect 3676 2135 4014 2148
rect 3180 2071 3233 2074
rect 3180 2054 3192 2071
rect 3224 2054 3233 2071
rect 3180 2046 3233 2054
rect 3179 1999 3233 2046
rect 3465 2062 3575 2077
rect 3465 2059 3542 2062
rect 3465 2032 3468 2059
rect 3497 2035 3542 2059
rect 3571 2035 3575 2062
rect 3497 2032 3575 2035
rect 3465 2018 3575 2032
rect 3676 1999 3713 2135
rect 3982 2118 4014 2135
rect 4403 2143 4410 2163
rect 4429 2143 4487 2163
rect 4506 2143 4514 2163
rect 4403 2121 4514 2143
rect 5249 2120 5291 2173
rect 3982 2072 4013 2118
rect 5249 2101 5258 2120
rect 5283 2101 5291 2120
rect 5249 2091 5291 2101
rect 5477 2131 5587 2145
rect 5477 2128 5555 2131
rect 5477 2101 5481 2128
rect 5510 2104 5555 2128
rect 5584 2104 5587 2131
rect 6207 2121 6241 2173
rect 6701 2164 6706 2184
rect 6727 2164 6733 2184
rect 6701 2157 6733 2164
rect 6911 2185 6949 2195
rect 7146 2192 7180 2398
rect 6911 2168 6921 2185
rect 6941 2168 6949 2185
rect 6752 2125 6793 2126
rect 5510 2101 5587 2104
rect 5477 2086 5587 2101
rect 6206 2116 6241 2121
rect 6206 2096 6213 2116
rect 6233 2096 6241 2116
rect 6751 2115 6793 2125
rect 6206 2088 6241 2096
rect 3770 2069 3805 2070
rect 3749 2062 3805 2069
rect 3749 2042 3778 2062
rect 3798 2042 3805 2062
rect 3749 2037 3805 2042
rect 3982 2065 4021 2072
rect 3982 2045 3988 2065
rect 4013 2045 4021 2065
rect 3982 2039 4021 2045
rect 4196 2065 4228 2072
rect 4196 2045 4202 2065
rect 4223 2045 4228 2065
rect 3179 1964 3714 1999
rect 3179 1960 3232 1964
rect 3040 1848 3044 1875
rect 3075 1848 3079 1875
rect 3325 1896 3436 1913
rect 3325 1876 3332 1896
rect 3351 1876 3409 1896
rect 3428 1876 3436 1896
rect 3325 1854 3436 1876
rect 3040 1841 3079 1848
rect 3749 1831 3783 2037
rect 4196 2017 4228 2045
rect 3816 2009 4228 2017
rect 3816 1983 3822 2009
rect 3848 1983 4228 2009
rect 3816 1981 4228 1983
rect 3818 1980 3858 1981
rect 4196 1916 4228 1981
rect 5762 2023 5794 2030
rect 5762 2003 5769 2023
rect 5790 2003 5794 2023
rect 5762 1938 5794 2003
rect 6132 1938 6172 1939
rect 5762 1936 6174 1938
rect 4196 1896 4200 1916
rect 4221 1896 4228 1916
rect 4196 1889 4228 1896
rect 4699 1931 4747 1936
rect 4699 1902 4710 1931
rect 4739 1902 4747 1931
rect 3749 1830 3784 1831
rect 3747 1823 3784 1830
rect 2902 1779 2910 1800
rect 2937 1779 2944 1800
rect 2156 1615 2196 1616
rect 1786 1613 2198 1615
rect 1154 1609 1189 1611
rect 190 1606 1189 1609
rect 189 1582 1189 1606
rect 189 1427 237 1582
rect 423 1541 533 1555
rect 423 1538 501 1541
rect 423 1511 427 1538
rect 456 1514 501 1538
rect 530 1514 533 1541
rect 1154 1531 1189 1582
rect 456 1511 533 1514
rect 423 1496 533 1511
rect 1152 1526 1189 1531
rect 1152 1506 1159 1526
rect 1179 1506 1189 1526
rect 1786 1587 2166 1613
rect 2192 1587 2198 1613
rect 1786 1579 2198 1587
rect 1786 1551 1818 1579
rect 2231 1559 2267 1707
rect 1786 1531 1791 1551
rect 1812 1531 1818 1551
rect 1786 1524 1818 1531
rect 2209 1554 2267 1559
rect 2209 1534 2216 1554
rect 2236 1534 2267 1554
rect 2209 1527 2267 1534
rect 2671 1564 2705 1770
rect 2902 1768 2944 1779
rect 3118 1798 3150 1805
rect 3118 1778 3124 1798
rect 3145 1778 3150 1798
rect 3118 1750 3150 1778
rect 2738 1742 3150 1750
rect 2738 1716 2744 1742
rect 2770 1716 3150 1742
rect 3747 1803 3757 1823
rect 3777 1803 3784 1823
rect 3747 1798 3784 1803
rect 4403 1818 4513 1833
rect 4403 1815 4480 1818
rect 3747 1747 3782 1798
rect 4403 1788 4406 1815
rect 4435 1791 4480 1815
rect 4509 1791 4513 1818
rect 4435 1788 4513 1791
rect 4403 1774 4513 1788
rect 4699 1747 4747 1902
rect 5762 1910 6142 1936
rect 6168 1910 6174 1936
rect 5762 1902 6174 1910
rect 5762 1874 5794 1902
rect 6207 1882 6241 2088
rect 6415 2086 6526 2108
rect 6415 2066 6423 2086
rect 6442 2066 6500 2086
rect 6519 2066 6526 2086
rect 6415 2049 6526 2066
rect 6751 2093 6758 2115
rect 6784 2093 6793 2115
rect 6751 2084 6793 2093
rect 5968 1879 6011 1881
rect 5762 1854 5767 1874
rect 5788 1854 5794 1874
rect 5762 1847 5794 1854
rect 5967 1872 6011 1879
rect 5967 1852 5977 1872
rect 6000 1852 6011 1872
rect 5967 1848 6011 1852
rect 6185 1877 6241 1882
rect 6185 1857 6192 1877
rect 6212 1857 6241 1877
rect 6185 1850 6241 1857
rect 6297 2018 6330 2019
rect 6751 2018 6788 2084
rect 6297 1989 6788 2018
rect 6185 1849 6220 1850
rect 3747 1723 4747 1747
rect 5476 1776 5587 1798
rect 5476 1756 5484 1776
rect 5503 1756 5561 1776
rect 5580 1756 5587 1776
rect 5476 1739 5587 1756
rect 5967 1767 6009 1848
rect 6297 1769 6330 1989
rect 6751 1987 6788 1989
rect 6557 1849 6667 1863
rect 6557 1846 6635 1849
rect 6557 1819 6561 1846
rect 6590 1822 6635 1846
rect 6664 1822 6667 1849
rect 6590 1819 6667 1822
rect 6557 1804 6667 1819
rect 6911 1830 6949 2168
rect 7124 2187 7180 2192
rect 7124 2167 7131 2187
rect 7151 2167 7180 2187
rect 7124 2160 7180 2167
rect 7124 2159 7159 2160
rect 7046 2059 7090 2063
rect 7227 2059 7277 2600
rect 7046 2026 7277 2059
rect 7755 2054 7793 2667
rect 8411 2682 8521 2697
rect 8411 2679 8488 2682
rect 8411 2652 8414 2679
rect 8443 2655 8488 2679
rect 8517 2655 8521 2682
rect 8443 2652 8521 2655
rect 8411 2638 8521 2652
rect 8259 2525 8296 2527
rect 8717 2525 8750 2745
rect 9038 2666 9080 2747
rect 9460 2758 9571 2774
rect 9460 2738 9467 2758
rect 9486 2738 9544 2758
rect 9563 2738 9571 2758
rect 9460 2716 9571 2738
rect 8827 2664 8862 2665
rect 8259 2496 8750 2525
rect 8259 2430 8296 2496
rect 8717 2495 8750 2496
rect 8806 2657 8862 2664
rect 8806 2637 8835 2657
rect 8855 2637 8862 2657
rect 8806 2632 8862 2637
rect 9036 2662 9080 2666
rect 9036 2642 9047 2662
rect 9070 2642 9080 2662
rect 9036 2635 9080 2642
rect 9253 2660 9285 2667
rect 9253 2640 9259 2660
rect 9280 2640 9285 2660
rect 9036 2633 9079 2635
rect 8254 2421 8296 2430
rect 8254 2399 8263 2421
rect 8289 2399 8296 2421
rect 8521 2448 8632 2465
rect 8521 2428 8528 2448
rect 8547 2428 8605 2448
rect 8624 2428 8632 2448
rect 8521 2406 8632 2428
rect 8806 2426 8840 2632
rect 9253 2612 9285 2640
rect 8873 2604 9285 2612
rect 8873 2578 8879 2604
rect 8905 2578 9285 2604
rect 8873 2576 9285 2578
rect 8875 2575 8915 2576
rect 9253 2511 9285 2576
rect 9253 2491 9257 2511
rect 9278 2491 9285 2511
rect 9253 2484 9285 2491
rect 8806 2418 8841 2426
rect 8254 2389 8296 2399
rect 8806 2398 8814 2418
rect 8834 2398 8841 2418
rect 8806 2393 8841 2398
rect 9460 2413 9570 2428
rect 9460 2410 9537 2413
rect 8254 2388 8295 2389
rect 7888 2354 7923 2355
rect 7867 2347 7923 2354
rect 7867 2327 7896 2347
rect 7916 2327 7923 2347
rect 7867 2322 7923 2327
rect 8314 2350 8346 2357
rect 8314 2330 8320 2350
rect 8341 2330 8346 2350
rect 8806 2341 8840 2393
rect 9460 2383 9463 2410
rect 9492 2386 9537 2410
rect 9566 2386 9570 2413
rect 9492 2383 9570 2386
rect 9460 2369 9570 2383
rect 9756 2413 9798 2423
rect 9756 2394 9764 2413
rect 9789 2394 9798 2413
rect 9756 2341 9798 2394
rect 7867 2116 7901 2322
rect 8314 2302 8346 2330
rect 8804 2315 9800 2341
rect 7934 2294 8346 2302
rect 7934 2268 7940 2294
rect 7966 2268 8346 2294
rect 7934 2266 8346 2268
rect 7936 2265 7976 2266
rect 8096 2230 8135 2245
rect 8096 2189 8107 2230
rect 8128 2189 8135 2230
rect 7866 2108 7902 2116
rect 7866 2088 7875 2108
rect 7895 2088 7902 2108
rect 7866 2087 7902 2088
rect 7866 2076 7900 2087
rect 7756 2046 7793 2054
rect 7046 2024 7253 2026
rect 7046 1870 7090 2024
rect 7756 2012 8000 2046
rect 6911 1813 6919 1830
rect 6939 1813 6949 1830
rect 6911 1807 6949 1813
rect 6269 1767 6330 1769
rect 5967 1738 6330 1767
rect 6842 1741 6874 1748
rect 5967 1736 6269 1738
rect 3747 1720 4746 1723
rect 6842 1721 6849 1741
rect 6870 1721 6874 1741
rect 3747 1718 3782 1720
rect 2738 1714 3150 1716
rect 2740 1713 2780 1714
rect 3118 1649 3150 1714
rect 6842 1656 6874 1721
rect 7052 1734 7090 1870
rect 7748 1843 7783 1844
rect 7289 1839 7320 1840
rect 7286 1834 7320 1839
rect 7286 1814 7293 1834
rect 7313 1814 7320 1834
rect 7286 1806 7320 1814
rect 7052 1696 7058 1734
rect 7081 1696 7090 1734
rect 7052 1686 7090 1696
rect 7287 1748 7320 1806
rect 7727 1836 7783 1843
rect 7727 1816 7756 1836
rect 7776 1816 7783 1836
rect 7727 1811 7783 1816
rect 7958 1841 8000 2012
rect 8096 1916 8135 2189
rect 8314 2201 8346 2266
rect 8314 2181 8318 2201
rect 8339 2181 8346 2201
rect 8314 2174 8346 2181
rect 8732 2208 8790 2209
rect 8732 2189 9069 2208
rect 9459 2204 9570 2221
rect 8732 2176 9070 2189
rect 8236 2112 8289 2115
rect 8236 2095 8248 2112
rect 8280 2095 8289 2112
rect 8236 2087 8289 2095
rect 8235 2040 8289 2087
rect 8521 2103 8631 2118
rect 8521 2100 8598 2103
rect 8521 2073 8524 2100
rect 8553 2076 8598 2100
rect 8627 2076 8631 2103
rect 8553 2073 8631 2076
rect 8521 2059 8631 2073
rect 8732 2040 8769 2176
rect 9038 2159 9070 2176
rect 9459 2184 9466 2204
rect 9485 2184 9543 2204
rect 9562 2184 9570 2204
rect 9459 2162 9570 2184
rect 9038 2113 9069 2159
rect 8826 2110 8861 2111
rect 8805 2103 8861 2110
rect 8805 2083 8834 2103
rect 8854 2083 8861 2103
rect 8805 2078 8861 2083
rect 9038 2106 9077 2113
rect 9038 2086 9044 2106
rect 9069 2086 9077 2106
rect 9038 2080 9077 2086
rect 9252 2106 9284 2113
rect 9252 2086 9258 2106
rect 9279 2086 9284 2106
rect 8235 2005 8770 2040
rect 8235 2001 8288 2005
rect 8096 1889 8100 1916
rect 8131 1889 8135 1916
rect 8381 1937 8492 1954
rect 8381 1917 8388 1937
rect 8407 1917 8465 1937
rect 8484 1917 8492 1937
rect 8381 1895 8492 1917
rect 8096 1882 8135 1889
rect 8805 1872 8839 2078
rect 9252 2058 9284 2086
rect 8872 2050 9284 2058
rect 8872 2024 8878 2050
rect 8904 2024 9284 2050
rect 8872 2022 9284 2024
rect 8874 2021 8914 2022
rect 9252 1957 9284 2022
rect 9252 1937 9256 1957
rect 9277 1937 9284 1957
rect 9252 1930 9284 1937
rect 9755 1972 9803 1977
rect 9755 1943 9766 1972
rect 9795 1943 9803 1972
rect 8805 1871 8840 1872
rect 8803 1864 8840 1871
rect 7958 1820 7966 1841
rect 7993 1820 8000 1841
rect 7212 1656 7252 1657
rect 6842 1654 7254 1656
rect 6210 1650 6245 1652
rect 3118 1629 3122 1649
rect 3143 1629 3150 1649
rect 5246 1647 6245 1650
rect 3723 1632 4025 1634
rect 3118 1622 3150 1629
rect 3662 1603 4025 1632
rect 3662 1601 3723 1603
rect 2671 1556 2706 1564
rect 2671 1536 2679 1556
rect 2699 1536 2706 1556
rect 2671 1531 2706 1536
rect 3043 1557 3081 1563
rect 3043 1540 3053 1557
rect 3073 1540 3081 1557
rect 2671 1530 2703 1531
rect 2209 1526 2244 1527
rect 1152 1499 1189 1506
rect 1152 1498 1187 1499
rect 189 1398 197 1427
rect 226 1398 237 1427
rect 189 1393 237 1398
rect 708 1433 740 1440
rect 708 1413 715 1433
rect 736 1413 740 1433
rect 708 1348 740 1413
rect 1078 1348 1118 1349
rect 708 1346 1120 1348
rect 708 1320 1088 1346
rect 1114 1320 1120 1346
rect 708 1312 1120 1320
rect 708 1284 740 1312
rect 1153 1292 1187 1498
rect 1857 1481 1896 1488
rect 1500 1453 1611 1475
rect 1500 1433 1508 1453
rect 1527 1433 1585 1453
rect 1604 1433 1611 1453
rect 1500 1416 1611 1433
rect 1857 1454 1861 1481
rect 1892 1454 1896 1481
rect 1704 1365 1757 1369
rect 1222 1330 1757 1365
rect 708 1264 713 1284
rect 734 1264 740 1284
rect 708 1257 740 1264
rect 915 1284 954 1290
rect 915 1264 923 1284
rect 948 1264 954 1284
rect 915 1257 954 1264
rect 1131 1287 1187 1292
rect 1131 1267 1138 1287
rect 1158 1267 1187 1287
rect 1131 1260 1187 1267
rect 1131 1259 1166 1260
rect 923 1211 954 1257
rect 422 1186 533 1208
rect 422 1166 430 1186
rect 449 1166 507 1186
rect 526 1166 533 1186
rect 922 1194 954 1211
rect 1223 1194 1260 1330
rect 1361 1297 1471 1311
rect 1361 1294 1439 1297
rect 1361 1267 1365 1294
rect 1394 1270 1439 1294
rect 1468 1270 1471 1297
rect 1394 1267 1471 1270
rect 1361 1252 1471 1267
rect 1703 1283 1757 1330
rect 1703 1275 1756 1283
rect 1703 1258 1712 1275
rect 1744 1258 1756 1275
rect 1703 1255 1756 1258
rect 922 1181 1260 1194
rect 422 1149 533 1166
rect 923 1162 1260 1181
rect 1202 1161 1260 1162
rect 1646 1189 1678 1196
rect 1646 1169 1653 1189
rect 1674 1169 1678 1189
rect 1646 1104 1678 1169
rect 1857 1181 1896 1454
rect 2092 1283 2126 1294
rect 2090 1282 2126 1283
rect 2090 1262 2097 1282
rect 2117 1262 2126 1282
rect 2090 1254 2126 1262
rect 1857 1140 1864 1181
rect 1885 1140 1896 1181
rect 1857 1125 1896 1140
rect 2016 1104 2056 1105
rect 1646 1102 2058 1104
rect 1646 1076 2026 1102
rect 2052 1076 2058 1102
rect 1646 1068 2058 1076
rect 192 1029 1188 1055
rect 1646 1040 1678 1068
rect 2091 1048 2125 1254
rect 2833 1210 2868 1211
rect 194 976 236 1029
rect 194 957 203 976
rect 228 957 236 976
rect 194 947 236 957
rect 422 987 532 1001
rect 422 984 500 987
rect 422 957 426 984
rect 455 960 500 984
rect 529 960 532 987
rect 1152 977 1186 1029
rect 1646 1020 1651 1040
rect 1672 1020 1678 1040
rect 1646 1013 1678 1020
rect 2069 1043 2125 1048
rect 2069 1023 2076 1043
rect 2096 1023 2125 1043
rect 2069 1016 2125 1023
rect 2812 1203 2868 1210
rect 2812 1183 2841 1203
rect 2861 1183 2868 1203
rect 2812 1178 2868 1183
rect 3043 1202 3081 1540
rect 3325 1551 3435 1566
rect 3325 1548 3402 1551
rect 3325 1521 3328 1548
rect 3357 1524 3402 1548
rect 3431 1524 3435 1551
rect 3357 1521 3435 1524
rect 3325 1507 3435 1521
rect 3204 1381 3241 1383
rect 3662 1381 3695 1601
rect 3983 1522 4025 1603
rect 4405 1614 4516 1631
rect 4405 1594 4412 1614
rect 4431 1594 4489 1614
rect 4508 1594 4516 1614
rect 4405 1572 4516 1594
rect 5245 1623 6245 1647
rect 3772 1520 3807 1521
rect 3204 1352 3695 1381
rect 3204 1286 3241 1352
rect 3662 1351 3695 1352
rect 3751 1513 3807 1520
rect 3751 1493 3780 1513
rect 3800 1493 3807 1513
rect 3751 1488 3807 1493
rect 3981 1518 4025 1522
rect 3981 1498 3992 1518
rect 4015 1498 4025 1518
rect 3981 1491 4025 1498
rect 4198 1516 4230 1523
rect 4198 1496 4204 1516
rect 4225 1496 4230 1516
rect 3981 1489 4024 1491
rect 3199 1277 3241 1286
rect 3199 1255 3208 1277
rect 3234 1255 3241 1277
rect 3466 1304 3577 1321
rect 3466 1284 3473 1304
rect 3492 1284 3550 1304
rect 3569 1284 3577 1304
rect 3466 1262 3577 1284
rect 3751 1282 3785 1488
rect 4198 1468 4230 1496
rect 3818 1460 4230 1468
rect 3818 1434 3824 1460
rect 3850 1434 4230 1460
rect 5245 1468 5293 1623
rect 5479 1582 5589 1596
rect 5479 1579 5557 1582
rect 5479 1552 5483 1579
rect 5512 1555 5557 1579
rect 5586 1555 5589 1582
rect 6210 1572 6245 1623
rect 5512 1552 5589 1555
rect 5479 1537 5589 1552
rect 6208 1567 6245 1572
rect 6208 1547 6215 1567
rect 6235 1547 6245 1567
rect 6842 1628 7222 1654
rect 7248 1628 7254 1654
rect 6842 1620 7254 1628
rect 6842 1592 6874 1620
rect 7287 1600 7323 1748
rect 6842 1572 6847 1592
rect 6868 1572 6874 1592
rect 6842 1565 6874 1572
rect 7265 1595 7323 1600
rect 7265 1575 7272 1595
rect 7292 1575 7323 1595
rect 7265 1568 7323 1575
rect 7727 1605 7761 1811
rect 7958 1809 8000 1820
rect 8174 1839 8206 1846
rect 8174 1819 8180 1839
rect 8201 1819 8206 1839
rect 8174 1791 8206 1819
rect 7794 1783 8206 1791
rect 7794 1757 7800 1783
rect 7826 1757 8206 1783
rect 8803 1844 8813 1864
rect 8833 1844 8840 1864
rect 8803 1839 8840 1844
rect 9459 1859 9569 1874
rect 9459 1856 9536 1859
rect 8803 1788 8838 1839
rect 9459 1829 9462 1856
rect 9491 1832 9536 1856
rect 9565 1832 9569 1859
rect 9491 1829 9569 1832
rect 9459 1815 9569 1829
rect 9755 1788 9803 1943
rect 8803 1764 9803 1788
rect 8803 1761 9802 1764
rect 8803 1759 8838 1761
rect 7794 1755 8206 1757
rect 7796 1754 7836 1755
rect 8174 1690 8206 1755
rect 8174 1670 8178 1690
rect 8199 1670 8206 1690
rect 8779 1673 9081 1675
rect 8174 1663 8206 1670
rect 8718 1644 9081 1673
rect 8718 1642 8779 1644
rect 7727 1597 7762 1605
rect 7727 1577 7735 1597
rect 7755 1577 7762 1597
rect 7727 1572 7762 1577
rect 8099 1598 8137 1604
rect 8099 1581 8109 1598
rect 8129 1581 8137 1598
rect 7727 1571 7759 1572
rect 7265 1567 7300 1568
rect 6208 1540 6245 1547
rect 6208 1539 6243 1540
rect 5245 1439 5253 1468
rect 5282 1439 5293 1468
rect 5245 1434 5293 1439
rect 5764 1474 5796 1481
rect 5764 1454 5771 1474
rect 5792 1454 5796 1474
rect 3818 1432 4230 1434
rect 3820 1431 3860 1432
rect 4198 1367 4230 1432
rect 4198 1347 4202 1367
rect 4223 1347 4230 1367
rect 4198 1340 4230 1347
rect 5764 1389 5796 1454
rect 6134 1389 6174 1390
rect 5764 1387 6176 1389
rect 5764 1361 6144 1387
rect 6170 1361 6176 1387
rect 5764 1353 6176 1361
rect 5764 1325 5796 1353
rect 6209 1333 6243 1539
rect 6913 1522 6952 1529
rect 6556 1494 6667 1516
rect 6556 1474 6564 1494
rect 6583 1474 6641 1494
rect 6660 1474 6667 1494
rect 6556 1457 6667 1474
rect 6913 1495 6917 1522
rect 6948 1495 6952 1522
rect 6760 1406 6813 1410
rect 6278 1371 6813 1406
rect 5764 1305 5769 1325
rect 5790 1305 5796 1325
rect 5764 1298 5796 1305
rect 5971 1325 6010 1331
rect 5971 1305 5979 1325
rect 6004 1305 6010 1325
rect 5971 1298 6010 1305
rect 6187 1328 6243 1333
rect 6187 1308 6194 1328
rect 6214 1308 6243 1328
rect 6187 1301 6243 1308
rect 6187 1300 6222 1301
rect 3751 1274 3786 1282
rect 3199 1245 3241 1255
rect 3751 1254 3759 1274
rect 3779 1254 3786 1274
rect 3751 1249 3786 1254
rect 4405 1269 4515 1284
rect 4405 1266 4482 1269
rect 3199 1244 3240 1245
rect 3043 1185 3051 1202
rect 3071 1185 3081 1202
rect 2069 1015 2104 1016
rect 1697 981 1738 982
rect 455 957 532 960
rect 422 942 532 957
rect 1151 972 1186 977
rect 1151 952 1158 972
rect 1178 952 1186 972
rect 1696 971 1738 981
rect 1151 944 1186 952
rect 707 879 739 886
rect 707 859 714 879
rect 735 859 739 879
rect 707 794 739 859
rect 1077 794 1117 795
rect 707 792 1119 794
rect 707 766 1087 792
rect 1113 766 1119 792
rect 707 758 1119 766
rect 707 730 739 758
rect 1152 738 1186 944
rect 1360 942 1471 964
rect 1360 922 1368 942
rect 1387 922 1445 942
rect 1464 922 1471 942
rect 1360 905 1471 922
rect 1696 949 1703 971
rect 1729 949 1738 971
rect 1696 940 1738 949
rect 2812 972 2846 1178
rect 3043 1175 3081 1185
rect 3259 1206 3291 1213
rect 3259 1186 3265 1206
rect 3286 1186 3291 1206
rect 3751 1197 3785 1249
rect 4405 1239 4408 1266
rect 4437 1242 4482 1266
rect 4511 1242 4515 1269
rect 4437 1239 4515 1242
rect 4405 1225 4515 1239
rect 4701 1269 4743 1279
rect 4701 1250 4709 1269
rect 4734 1250 4743 1269
rect 5979 1252 6010 1298
rect 4701 1197 4743 1250
rect 5478 1227 5589 1249
rect 5478 1207 5486 1227
rect 5505 1207 5563 1227
rect 5582 1207 5589 1227
rect 5978 1235 6010 1252
rect 6279 1235 6316 1371
rect 6417 1338 6527 1352
rect 6417 1335 6495 1338
rect 6417 1308 6421 1335
rect 6450 1311 6495 1335
rect 6524 1311 6527 1338
rect 6450 1308 6527 1311
rect 6417 1293 6527 1308
rect 6759 1324 6813 1371
rect 6759 1316 6812 1324
rect 6759 1299 6768 1316
rect 6800 1299 6812 1316
rect 6759 1296 6812 1299
rect 5978 1222 6316 1235
rect 3259 1158 3291 1186
rect 3749 1171 4745 1197
rect 5478 1190 5589 1207
rect 5979 1203 6316 1222
rect 6258 1202 6316 1203
rect 6702 1230 6734 1237
rect 6702 1210 6709 1230
rect 6730 1210 6734 1230
rect 2879 1150 3291 1158
rect 2879 1124 2885 1150
rect 2911 1124 3291 1150
rect 2879 1122 3291 1124
rect 2881 1121 2921 1122
rect 3259 1057 3291 1122
rect 6702 1145 6734 1210
rect 6913 1222 6952 1495
rect 7148 1324 7182 1335
rect 7146 1323 7182 1324
rect 7146 1303 7153 1323
rect 7173 1303 7182 1323
rect 7146 1295 7182 1303
rect 6913 1181 6920 1222
rect 6941 1181 6952 1222
rect 6913 1166 6952 1181
rect 7072 1145 7112 1146
rect 6702 1143 7114 1145
rect 6702 1117 7082 1143
rect 7108 1117 7114 1143
rect 6702 1109 7114 1117
rect 3259 1037 3263 1057
rect 3284 1037 3291 1057
rect 3259 1030 3291 1037
rect 3677 1064 3735 1065
rect 3677 1045 4014 1064
rect 4404 1060 4515 1077
rect 5248 1070 6244 1096
rect 6702 1081 6734 1109
rect 7147 1089 7181 1295
rect 7889 1251 7924 1252
rect 3677 1032 4015 1045
rect 2812 964 2847 972
rect 2812 944 2820 964
rect 2840 944 2847 964
rect 913 735 956 737
rect 707 710 712 730
rect 733 710 739 730
rect 707 703 739 710
rect 912 728 956 735
rect 912 708 922 728
rect 945 708 956 728
rect 912 704 956 708
rect 1130 733 1186 738
rect 1130 713 1137 733
rect 1157 713 1186 733
rect 1130 706 1186 713
rect 1242 874 1275 875
rect 1696 874 1733 940
rect 2812 939 2847 944
rect 3466 959 3576 974
rect 3466 956 3543 959
rect 2812 896 2846 939
rect 3466 929 3469 956
rect 3498 932 3543 956
rect 3572 932 3576 959
rect 3498 929 3576 932
rect 3466 915 3576 929
rect 3677 896 3714 1032
rect 3983 1015 4015 1032
rect 4404 1040 4411 1060
rect 4430 1040 4488 1060
rect 4507 1040 4515 1060
rect 4404 1018 4515 1040
rect 5250 1017 5292 1070
rect 3983 969 4014 1015
rect 5250 998 5259 1017
rect 5284 998 5292 1017
rect 5250 988 5292 998
rect 5478 1028 5588 1042
rect 5478 1025 5556 1028
rect 5478 998 5482 1025
rect 5511 1001 5556 1025
rect 5585 1001 5588 1028
rect 6208 1018 6242 1070
rect 6702 1061 6707 1081
rect 6728 1061 6734 1081
rect 6702 1054 6734 1061
rect 7125 1084 7181 1089
rect 7125 1064 7132 1084
rect 7152 1064 7181 1084
rect 7125 1057 7181 1064
rect 7868 1244 7924 1251
rect 7868 1224 7897 1244
rect 7917 1224 7924 1244
rect 7868 1219 7924 1224
rect 8099 1243 8137 1581
rect 8381 1592 8491 1607
rect 8381 1589 8458 1592
rect 8381 1562 8384 1589
rect 8413 1565 8458 1589
rect 8487 1565 8491 1592
rect 8413 1562 8491 1565
rect 8381 1548 8491 1562
rect 8260 1422 8297 1424
rect 8718 1422 8751 1642
rect 9039 1563 9081 1644
rect 9461 1655 9572 1672
rect 9461 1635 9468 1655
rect 9487 1635 9545 1655
rect 9564 1635 9572 1655
rect 9461 1613 9572 1635
rect 8828 1561 8863 1562
rect 8260 1393 8751 1422
rect 8260 1327 8297 1393
rect 8718 1392 8751 1393
rect 8807 1554 8863 1561
rect 8807 1534 8836 1554
rect 8856 1534 8863 1554
rect 8807 1529 8863 1534
rect 9037 1559 9081 1563
rect 9037 1539 9048 1559
rect 9071 1539 9081 1559
rect 9037 1532 9081 1539
rect 9254 1557 9286 1564
rect 9254 1537 9260 1557
rect 9281 1537 9286 1557
rect 9037 1530 9080 1532
rect 8255 1318 8297 1327
rect 8255 1296 8264 1318
rect 8290 1296 8297 1318
rect 8522 1345 8633 1362
rect 8522 1325 8529 1345
rect 8548 1325 8606 1345
rect 8625 1325 8633 1345
rect 8522 1303 8633 1325
rect 8807 1323 8841 1529
rect 9254 1509 9286 1537
rect 8874 1501 9286 1509
rect 8874 1475 8880 1501
rect 8906 1475 9286 1501
rect 8874 1473 9286 1475
rect 8876 1472 8916 1473
rect 9254 1408 9286 1473
rect 9254 1388 9258 1408
rect 9279 1388 9286 1408
rect 9254 1381 9286 1388
rect 8807 1315 8842 1323
rect 8255 1286 8297 1296
rect 8807 1295 8815 1315
rect 8835 1295 8842 1315
rect 8807 1290 8842 1295
rect 9461 1310 9571 1325
rect 9461 1307 9538 1310
rect 8255 1285 8296 1286
rect 8099 1226 8107 1243
rect 8127 1226 8137 1243
rect 7125 1056 7160 1057
rect 6753 1022 6794 1023
rect 5511 998 5588 1001
rect 5478 983 5588 998
rect 6207 1013 6242 1018
rect 6207 993 6214 1013
rect 6234 993 6242 1013
rect 6752 1012 6794 1022
rect 6207 985 6242 993
rect 3771 966 3806 967
rect 3750 959 3806 966
rect 3750 939 3779 959
rect 3799 939 3806 959
rect 3750 934 3806 939
rect 3983 962 4022 969
rect 3983 942 3989 962
rect 4014 942 4022 962
rect 3983 936 4022 942
rect 4197 962 4229 969
rect 4197 942 4203 962
rect 4224 942 4229 962
rect 1242 845 1733 874
rect 2811 861 3715 896
rect 2812 860 2846 861
rect 1130 705 1165 706
rect 421 634 532 654
rect 421 632 531 634
rect 421 612 429 632
rect 448 612 506 632
rect 525 612 531 632
rect 421 595 531 612
rect 912 623 954 704
rect 1242 625 1275 845
rect 1696 843 1733 845
rect 3750 728 3784 934
rect 4197 914 4229 942
rect 3817 906 4229 914
rect 3817 880 3823 906
rect 3849 880 4229 906
rect 3817 878 4229 880
rect 3819 877 3859 878
rect 4197 813 4229 878
rect 5763 920 5795 927
rect 5763 900 5770 920
rect 5791 900 5795 920
rect 5763 835 5795 900
rect 6133 835 6173 836
rect 5763 833 6175 835
rect 4197 793 4201 813
rect 4222 793 4229 813
rect 4197 786 4229 793
rect 4700 828 4748 833
rect 4700 799 4711 828
rect 4740 799 4748 828
rect 3750 727 3785 728
rect 1214 623 1275 625
rect 912 594 1275 623
rect 3748 720 3785 727
rect 3748 700 3758 720
rect 3778 700 3785 720
rect 3748 695 3785 700
rect 4404 715 4514 730
rect 4404 712 4481 715
rect 3748 644 3783 695
rect 4404 685 4407 712
rect 4436 688 4481 712
rect 4510 688 4514 715
rect 4436 685 4514 688
rect 4404 671 4514 685
rect 4700 644 4748 799
rect 5763 807 6143 833
rect 6169 807 6175 833
rect 5763 799 6175 807
rect 5763 771 5795 799
rect 6208 779 6242 985
rect 6416 983 6527 1005
rect 6416 963 6424 983
rect 6443 963 6501 983
rect 6520 963 6527 983
rect 6416 946 6527 963
rect 6752 990 6759 1012
rect 6785 990 6794 1012
rect 6752 981 6794 990
rect 7868 1013 7902 1219
rect 8099 1216 8137 1226
rect 8315 1247 8347 1254
rect 8315 1227 8321 1247
rect 8342 1227 8347 1247
rect 8807 1238 8841 1290
rect 9461 1280 9464 1307
rect 9493 1283 9538 1307
rect 9567 1283 9571 1310
rect 9493 1280 9571 1283
rect 9461 1266 9571 1280
rect 9757 1310 9799 1320
rect 9757 1291 9765 1310
rect 9790 1291 9799 1310
rect 9757 1238 9799 1291
rect 8315 1199 8347 1227
rect 8805 1212 9801 1238
rect 7935 1191 8347 1199
rect 7935 1165 7941 1191
rect 7967 1165 8347 1191
rect 7935 1163 8347 1165
rect 7937 1162 7977 1163
rect 8315 1098 8347 1163
rect 8315 1078 8319 1098
rect 8340 1078 8347 1098
rect 8315 1071 8347 1078
rect 8733 1105 8791 1106
rect 8733 1086 9070 1105
rect 9460 1101 9571 1118
rect 8733 1073 9071 1086
rect 7868 1005 7903 1013
rect 7868 985 7876 1005
rect 7896 985 7903 1005
rect 5969 776 6012 778
rect 5763 751 5768 771
rect 5789 751 5795 771
rect 5763 744 5795 751
rect 5968 769 6012 776
rect 5968 749 5978 769
rect 6001 749 6012 769
rect 5968 745 6012 749
rect 6186 774 6242 779
rect 6186 754 6193 774
rect 6213 754 6242 774
rect 6186 747 6242 754
rect 6298 915 6331 916
rect 6752 915 6789 981
rect 7868 980 7903 985
rect 8522 1000 8632 1015
rect 8522 997 8599 1000
rect 7868 937 7902 980
rect 8522 970 8525 997
rect 8554 973 8599 997
rect 8628 973 8632 1000
rect 8554 970 8632 973
rect 8522 956 8632 970
rect 8733 937 8770 1073
rect 9039 1056 9071 1073
rect 9460 1081 9467 1101
rect 9486 1081 9544 1101
rect 9563 1081 9571 1101
rect 9460 1059 9571 1081
rect 9039 1010 9070 1056
rect 8827 1007 8862 1008
rect 8806 1000 8862 1007
rect 8806 980 8835 1000
rect 8855 980 8862 1000
rect 8806 975 8862 980
rect 9039 1003 9078 1010
rect 9039 983 9045 1003
rect 9070 983 9078 1003
rect 9039 977 9078 983
rect 9253 1003 9285 1010
rect 9253 983 9259 1003
rect 9280 983 9285 1003
rect 6298 886 6789 915
rect 7867 902 8771 937
rect 7868 901 7902 902
rect 6186 746 6221 747
rect 3748 620 4748 644
rect 5477 675 5588 695
rect 5477 673 5587 675
rect 5477 653 5485 673
rect 5504 653 5562 673
rect 5581 653 5587 673
rect 5477 636 5587 653
rect 5968 664 6010 745
rect 6298 666 6331 886
rect 6752 884 6789 886
rect 8806 769 8840 975
rect 9253 955 9285 983
rect 8873 947 9285 955
rect 8873 921 8879 947
rect 8905 921 9285 947
rect 8873 919 9285 921
rect 8875 918 8915 919
rect 9253 854 9285 919
rect 9253 834 9257 854
rect 9278 834 9285 854
rect 9253 827 9285 834
rect 9756 869 9804 874
rect 9756 840 9767 869
rect 9796 840 9804 869
rect 8806 768 8841 769
rect 6270 664 6331 666
rect 5968 635 6331 664
rect 8804 761 8841 768
rect 8804 741 8814 761
rect 8834 741 8841 761
rect 8804 736 8841 741
rect 9460 756 9570 771
rect 9460 753 9537 756
rect 8804 685 8839 736
rect 9460 726 9463 753
rect 9492 729 9537 753
rect 9566 729 9570 756
rect 9492 726 9570 729
rect 9460 712 9570 726
rect 9756 685 9804 840
rect 8804 661 9804 685
rect 8804 658 9803 661
rect 8804 656 8839 658
rect 5968 633 6270 635
rect 3748 617 4747 620
rect 3748 615 3783 617
rect 5774 604 5853 608
rect 5774 595 9885 604
rect 912 592 1214 594
rect 5774 591 9848 595
rect 5774 570 5813 591
rect 5842 574 9848 591
rect 9877 574 9885 595
rect 5842 570 9885 574
rect 718 563 797 567
rect 718 554 4829 563
rect 718 550 4792 554
rect 718 529 757 550
rect 786 533 4792 550
rect 4821 533 4829 554
rect 5774 562 9885 570
rect 5774 551 5853 562
rect 786 529 4829 533
rect 718 521 4829 529
rect 718 510 797 521
rect 7440 512 7499 528
rect 2384 471 2443 487
rect 1669 428 1779 442
rect 1669 425 1747 428
rect 1669 398 1673 425
rect 1702 401 1747 425
rect 1776 401 1779 428
rect 1702 398 1779 401
rect 1669 383 1779 398
rect 2384 429 2403 471
rect 2435 429 2443 471
rect 2384 413 2443 429
rect 2384 393 2405 413
rect 2425 393 2443 413
rect 2384 388 2443 393
rect 2472 468 2532 488
rect 5351 477 5389 479
rect 2472 405 2484 468
rect 2515 405 2532 468
rect 4311 443 5391 477
rect 6725 469 6835 483
rect 6725 466 6803 469
rect 2472 390 2532 405
rect 2398 385 2433 388
rect 1954 320 1986 327
rect 1954 300 1961 320
rect 1982 300 1986 320
rect 1954 235 1986 300
rect 2324 235 2364 236
rect 1954 233 2366 235
rect 1954 207 2334 233
rect 2360 207 2366 233
rect 1954 199 2366 207
rect 1954 171 1986 199
rect 2399 179 2433 385
rect 1954 151 1959 171
rect 1980 151 1986 171
rect 1954 144 1986 151
rect 2154 170 2212 177
rect 2154 150 2165 170
rect 2199 150 2212 170
rect 1668 73 1779 95
rect 1668 53 1676 73
rect 1695 53 1753 73
rect 1772 53 1779 73
rect 1668 36 1779 53
rect 2154 77 2212 150
rect 2377 174 2433 179
rect 2377 154 2384 174
rect 2404 154 2433 174
rect 2377 147 2433 154
rect 2377 146 2412 147
rect 2472 113 2527 390
rect 2472 92 2486 113
rect 2513 92 2527 113
rect 2472 82 2527 92
rect 2154 66 2215 77
rect 4315 66 4367 443
rect 4619 408 4729 422
rect 4619 405 4697 408
rect 4619 378 4623 405
rect 4652 381 4697 405
rect 4726 381 4729 408
rect 5351 398 5389 443
rect 6725 439 6729 466
rect 6758 442 6803 466
rect 6832 442 6835 469
rect 6758 439 6835 442
rect 6725 424 6835 439
rect 7440 470 7459 512
rect 7491 470 7499 512
rect 7440 454 7499 470
rect 7440 434 7461 454
rect 7481 434 7499 454
rect 7440 429 7499 434
rect 7528 509 7588 529
rect 7528 446 7540 509
rect 7571 446 7588 509
rect 7528 431 7588 446
rect 7454 426 7489 429
rect 4652 378 4729 381
rect 4619 363 4729 378
rect 5348 393 5389 398
rect 5348 373 5355 393
rect 5375 373 5389 393
rect 5348 371 5389 373
rect 5348 365 5383 371
rect 4904 300 4936 307
rect 4904 280 4911 300
rect 4932 280 4936 300
rect 4904 215 4936 280
rect 5274 215 5314 216
rect 4904 213 5316 215
rect 4904 187 5284 213
rect 5310 187 5316 213
rect 4904 179 5316 187
rect 4904 151 4936 179
rect 5349 159 5383 365
rect 7010 361 7042 368
rect 7010 341 7017 361
rect 7038 341 7042 361
rect 7010 276 7042 341
rect 7380 276 7420 277
rect 7010 274 7422 276
rect 7010 248 7390 274
rect 7416 248 7422 274
rect 7010 240 7422 248
rect 7010 212 7042 240
rect 7455 220 7489 426
rect 7010 192 7015 212
rect 7036 192 7042 212
rect 7010 185 7042 192
rect 7210 211 7268 218
rect 7210 191 7221 211
rect 7255 191 7268 211
rect 4904 131 4909 151
rect 4930 131 4936 151
rect 4904 124 4936 131
rect 5327 154 5383 159
rect 5327 134 5334 154
rect 5354 134 5383 154
rect 5327 127 5383 134
rect 5327 126 5362 127
rect 6724 114 6835 136
rect 5413 94 5486 106
rect 2154 49 4367 66
rect 2155 25 4367 49
rect 4315 21 4367 25
rect 4618 53 4729 75
rect 4618 33 4626 53
rect 4645 33 4703 53
rect 4722 33 4729 53
rect 5413 68 5422 94
rect 5481 68 5486 94
rect 6724 94 6732 114
rect 6751 94 6809 114
rect 6828 94 6835 114
rect 6724 77 6835 94
rect 5413 35 5486 68
rect 7210 59 7268 191
rect 7433 215 7489 220
rect 7433 195 7440 215
rect 7460 195 7489 215
rect 7433 188 7489 195
rect 7433 187 7468 188
rect 7528 154 7583 431
rect 7528 133 7542 154
rect 7569 133 7583 154
rect 7528 123 7583 133
rect 7205 35 7270 59
rect 4618 16 4729 33
rect 5406 -17 7275 35
<< via1 >>
rect 2485 5138 2516 5191
rect 7541 5179 7572 5232
rect 2405 4750 2436 4803
rect 7461 4791 7492 4844
rect 2403 429 2435 471
rect 2484 405 2515 468
rect 7459 470 7491 512
rect 7540 446 7571 509
<< metal2 >>
rect 7529 5232 7577 5251
rect 2473 5191 2521 5210
rect 2473 5138 2485 5191
rect 2516 5138 2521 5191
rect 2394 4803 2442 4818
rect 2394 4750 2405 4803
rect 2436 4750 2442 4803
rect 2394 487 2442 4750
rect 2473 488 2521 5138
rect 7529 5179 7541 5232
rect 7572 5179 7577 5232
rect 7450 4844 7498 4859
rect 7450 4791 7461 4844
rect 7492 4791 7498 4844
rect 7450 528 7498 4791
rect 7529 529 7577 5179
rect 7440 512 7499 528
rect 2384 471 2443 487
rect 2384 429 2403 471
rect 2435 429 2443 471
rect 2384 388 2443 429
rect 2472 468 2532 488
rect 2472 405 2484 468
rect 2515 405 2532 468
rect 7440 470 7459 512
rect 7491 470 7499 512
rect 7440 429 7499 470
rect 7528 509 7588 529
rect 7528 446 7540 509
rect 7571 446 7588 509
rect 7528 431 7588 446
rect 2472 390 2532 405
<< labels >>
rlabel locali 290 9043 312 9058 1 d0
rlabel metal1 459 9266 487 9271 1 vdd
rlabel metal1 456 8873 490 8879 1 gnd
rlabel locali 1227 8795 1255 8816 1 d1
rlabel metal1 1394 8629 1428 8635 1 gnd
rlabel metal1 1397 9022 1425 9027 1 vdd
rlabel locali 289 8489 311 8504 1 d0
rlabel metal1 458 8712 486 8717 1 vdd
rlabel metal1 455 8319 489 8325 1 gnd
rlabel locali 110 9328 138 9336 1 vref
rlabel locali 291 7940 313 7955 1 d0
rlabel metal1 460 8163 488 8168 1 vdd
rlabel metal1 457 7770 491 7776 1 gnd
rlabel locali 1228 7692 1256 7713 1 d1
rlabel metal1 1395 7526 1429 7532 1 gnd
rlabel metal1 1398 7919 1426 7924 1 vdd
rlabel locali 290 7386 312 7401 1 d0
rlabel metal1 459 7609 487 7614 1 vdd
rlabel metal1 456 7216 490 7222 1 gnd
rlabel metal1 1538 8430 1566 8435 1 vdd
rlabel metal1 1535 8037 1569 8043 1 gnd
rlabel locali 1366 8202 1387 8221 1 d2
rlabel locali 291 6837 313 6852 1 d0
rlabel metal1 460 7060 488 7065 1 vdd
rlabel metal1 457 6667 491 6673 1 gnd
rlabel locali 1228 6589 1256 6610 1 d1
rlabel metal1 1395 6423 1429 6429 1 gnd
rlabel metal1 1398 6816 1426 6821 1 vdd
rlabel locali 290 6283 312 6298 1 d0
rlabel metal1 459 6506 487 6511 1 vdd
rlabel metal1 456 6113 490 6119 1 gnd
rlabel locali 292 5734 314 5749 1 d0
rlabel metal1 461 5957 489 5962 1 vdd
rlabel metal1 458 5564 492 5570 1 gnd
rlabel locali 1229 5486 1257 5507 1 d1
rlabel metal1 1396 5320 1430 5326 1 gnd
rlabel metal1 1399 5713 1427 5718 1 vdd
rlabel locali 291 5180 313 5195 1 d0
rlabel metal1 460 5403 488 5408 1 vdd
rlabel metal1 457 5010 491 5016 1 gnd
rlabel metal1 1539 6224 1567 6229 1 vdd
rlabel metal1 1536 5831 1570 5837 1 gnd
rlabel locali 1367 5996 1388 6015 1 d2
rlabel metal1 1508 7340 1536 7345 1 vdd
rlabel metal1 1505 6947 1539 6953 1 gnd
rlabel locali 1338 7116 1364 7133 1 d3
rlabel locali 1340 2704 1366 2721 1 d3
rlabel metal1 1507 2535 1541 2541 1 gnd
rlabel metal1 1510 2928 1538 2933 1 vdd
rlabel locali 1369 1584 1390 1603 1 d2
rlabel metal1 1538 1419 1572 1425 1 gnd
rlabel metal1 1541 1812 1569 1817 1 vdd
rlabel metal1 459 598 493 604 1 gnd
rlabel metal1 462 991 490 996 1 vdd
rlabel locali 293 768 315 783 1 d0
rlabel metal1 1401 1301 1429 1306 1 vdd
rlabel metal1 1398 908 1432 914 1 gnd
rlabel locali 1231 1074 1259 1095 1 d1
rlabel metal1 460 1152 494 1158 1 gnd
rlabel metal1 463 1545 491 1550 1 vdd
rlabel locali 294 1322 316 1337 1 d0
rlabel metal1 458 1701 492 1707 1 gnd
rlabel metal1 461 2094 489 2099 1 vdd
rlabel locali 292 1871 314 1886 1 d0
rlabel metal1 1400 2404 1428 2409 1 vdd
rlabel metal1 1397 2011 1431 2017 1 gnd
rlabel locali 1230 2177 1258 2198 1 d1
rlabel metal1 459 2255 493 2261 1 gnd
rlabel metal1 462 2648 490 2653 1 vdd
rlabel locali 293 2425 315 2440 1 d0
rlabel locali 1368 3790 1389 3809 1 d2
rlabel metal1 1537 3625 1571 3631 1 gnd
rlabel metal1 1540 4018 1568 4023 1 vdd
rlabel metal1 458 2804 492 2810 1 gnd
rlabel metal1 461 3197 489 3202 1 vdd
rlabel locali 292 2974 314 2989 1 d0
rlabel metal1 1400 3507 1428 3512 1 vdd
rlabel metal1 1397 3114 1431 3120 1 gnd
rlabel locali 1230 3280 1258 3301 1 d1
rlabel metal1 459 3358 493 3364 1 gnd
rlabel metal1 462 3751 490 3756 1 vdd
rlabel locali 293 3528 315 3543 1 d0
rlabel metal1 457 3907 491 3913 1 gnd
rlabel metal1 460 4300 488 4305 1 vdd
rlabel locali 291 4077 313 4092 1 d0
rlabel metal1 1399 4610 1427 4615 1 vdd
rlabel metal1 1396 4217 1430 4223 1 gnd
rlabel locali 1229 4383 1257 4404 1 d1
rlabel metal1 458 4461 492 4467 1 gnd
rlabel metal1 461 4854 489 4859 1 vdd
rlabel locali 292 4631 314 4646 1 d0
rlabel metal1 1508 5140 1536 5145 1 vdd
rlabel metal1 1505 4747 1539 4753 1 gnd
rlabel locali 1332 4909 1367 4935 1 d4
rlabel locali 4621 889 4643 904 5 d0
rlabel metal1 4446 676 4474 681 5 vdd
rlabel metal1 4443 1068 4477 1074 5 gnd
rlabel locali 3678 1131 3706 1152 5 d1
rlabel metal1 3505 1312 3539 1318 5 gnd
rlabel metal1 3508 920 3536 925 5 vdd
rlabel locali 4622 1443 4644 1458 5 d0
rlabel metal1 4447 1230 4475 1235 5 vdd
rlabel metal1 4444 1622 4478 1628 5 gnd
rlabel locali 4620 1992 4642 2007 5 d0
rlabel metal1 4445 1779 4473 1784 5 vdd
rlabel metal1 4442 2171 4476 2177 5 gnd
rlabel locali 3677 2234 3705 2255 5 d1
rlabel metal1 3504 2415 3538 2421 5 gnd
rlabel metal1 3507 2023 3535 2028 5 vdd
rlabel locali 4621 2546 4643 2561 5 d0
rlabel metal1 4446 2333 4474 2338 5 vdd
rlabel metal1 4443 2725 4477 2731 5 gnd
rlabel metal1 3367 1512 3395 1517 5 vdd
rlabel metal1 3364 1904 3398 1910 5 gnd
rlabel locali 3546 1726 3567 1745 5 d2
rlabel locali 4620 3095 4642 3110 5 d0
rlabel metal1 4445 2882 4473 2887 5 vdd
rlabel metal1 4442 3274 4476 3280 5 gnd
rlabel locali 3677 3337 3705 3358 5 d1
rlabel metal1 3504 3518 3538 3524 5 gnd
rlabel metal1 3507 3126 3535 3131 5 vdd
rlabel locali 4621 3649 4643 3664 5 d0
rlabel metal1 4446 3436 4474 3441 5 vdd
rlabel metal1 4443 3828 4477 3834 5 gnd
rlabel locali 4619 4198 4641 4213 5 d0
rlabel metal1 4444 3985 4472 3990 5 vdd
rlabel metal1 4441 4377 4475 4383 5 gnd
rlabel locali 3676 4440 3704 4461 5 d1
rlabel metal1 3503 4621 3537 4627 5 gnd
rlabel metal1 3506 4229 3534 4234 5 vdd
rlabel locali 4620 4752 4642 4767 5 d0
rlabel metal1 4445 4539 4473 4544 5 vdd
rlabel metal1 4442 4931 4476 4937 5 gnd
rlabel metal1 3366 3718 3394 3723 5 vdd
rlabel metal1 3363 4110 3397 4116 5 gnd
rlabel locali 3545 3932 3566 3951 5 d2
rlabel metal1 3397 2602 3425 2607 5 vdd
rlabel metal1 3394 2994 3428 3000 5 gnd
rlabel locali 3569 2814 3595 2831 5 d3
rlabel locali 3567 7226 3593 7243 5 d3
rlabel metal1 3392 7406 3426 7412 5 gnd
rlabel metal1 3395 7014 3423 7019 5 vdd
rlabel locali 3543 8344 3564 8363 5 d2
rlabel metal1 3361 8522 3395 8528 5 gnd
rlabel metal1 3364 8130 3392 8135 5 vdd
rlabel metal1 4440 9343 4474 9349 5 gnd
rlabel metal1 4443 8951 4471 8956 5 vdd
rlabel locali 4618 9164 4640 9179 5 d0
rlabel metal1 3504 8641 3532 8646 5 vdd
rlabel metal1 3501 9033 3535 9039 5 gnd
rlabel locali 3674 8852 3702 8873 5 d1
rlabel metal1 4439 8789 4473 8795 5 gnd
rlabel metal1 4442 8397 4470 8402 5 vdd
rlabel locali 4617 8610 4639 8625 5 d0
rlabel metal1 4441 8240 4475 8246 5 gnd
rlabel metal1 4444 7848 4472 7853 5 vdd
rlabel locali 4619 8061 4641 8076 5 d0
rlabel metal1 3505 7538 3533 7543 5 vdd
rlabel metal1 3502 7930 3536 7936 5 gnd
rlabel locali 3675 7749 3703 7770 5 d1
rlabel metal1 4440 7686 4474 7692 5 gnd
rlabel metal1 4443 7294 4471 7299 5 vdd
rlabel locali 4618 7507 4640 7522 5 d0
rlabel locali 3544 6138 3565 6157 5 d2
rlabel metal1 3362 6316 3396 6322 5 gnd
rlabel metal1 3365 5924 3393 5929 5 vdd
rlabel metal1 4441 7137 4475 7143 5 gnd
rlabel metal1 4444 6745 4472 6750 5 vdd
rlabel locali 4619 6958 4641 6973 5 d0
rlabel metal1 3505 6435 3533 6440 5 vdd
rlabel metal1 3502 6827 3536 6833 5 gnd
rlabel locali 3675 6646 3703 6667 5 d1
rlabel metal1 4440 6583 4474 6589 5 gnd
rlabel metal1 4443 6191 4471 6196 5 vdd
rlabel locali 4618 6404 4640 6419 5 d0
rlabel metal1 4442 6034 4476 6040 5 gnd
rlabel metal1 4445 5642 4473 5647 5 vdd
rlabel locali 4620 5855 4642 5870 5 d0
rlabel metal1 3506 5332 3534 5337 5 vdd
rlabel metal1 3503 5724 3537 5730 5 gnd
rlabel locali 3676 5543 3704 5564 5 d1
rlabel metal1 4441 5480 4475 5486 5 gnd
rlabel metal1 4444 5088 4472 5093 5 vdd
rlabel locali 4619 5301 4641 5316 5 d0
rlabel metal1 3397 4802 3425 4807 5 vdd
rlabel metal1 3394 5194 3428 5200 5 gnd
rlabel locali 3566 5012 3601 5038 5 d4
rlabel metal1 1709 432 1737 437 1 vdd
rlabel metal1 1706 39 1740 45 1 gnd
rlabel locali 1535 203 1563 225 1 d5
rlabel locali 5346 9084 5368 9099 1 d0
rlabel metal1 5515 9307 5543 9312 1 vdd
rlabel metal1 5512 8914 5546 8920 1 gnd
rlabel locali 6283 8836 6311 8857 1 d1
rlabel metal1 6450 8670 6484 8676 1 gnd
rlabel metal1 6453 9063 6481 9068 1 vdd
rlabel locali 5345 8530 5367 8545 1 d0
rlabel metal1 5514 8753 5542 8758 1 vdd
rlabel metal1 5511 8360 5545 8366 1 gnd
rlabel locali 5347 7981 5369 7996 1 d0
rlabel metal1 5516 8204 5544 8209 1 vdd
rlabel metal1 5513 7811 5547 7817 1 gnd
rlabel locali 6284 7733 6312 7754 1 d1
rlabel metal1 6451 7567 6485 7573 1 gnd
rlabel metal1 6454 7960 6482 7965 1 vdd
rlabel locali 5346 7427 5368 7442 1 d0
rlabel metal1 5515 7650 5543 7655 1 vdd
rlabel metal1 5512 7257 5546 7263 1 gnd
rlabel metal1 6594 8471 6622 8476 1 vdd
rlabel metal1 6591 8078 6625 8084 1 gnd
rlabel locali 6422 8243 6443 8262 1 d2
rlabel locali 5347 6878 5369 6893 1 d0
rlabel metal1 5516 7101 5544 7106 1 vdd
rlabel metal1 5513 6708 5547 6714 1 gnd
rlabel locali 6284 6630 6312 6651 1 d1
rlabel metal1 6451 6464 6485 6470 1 gnd
rlabel metal1 6454 6857 6482 6862 1 vdd
rlabel locali 5346 6324 5368 6339 1 d0
rlabel metal1 5515 6547 5543 6552 1 vdd
rlabel metal1 5512 6154 5546 6160 1 gnd
rlabel locali 5348 5775 5370 5790 1 d0
rlabel metal1 5517 5998 5545 6003 1 vdd
rlabel metal1 5514 5605 5548 5611 1 gnd
rlabel locali 6285 5527 6313 5548 1 d1
rlabel metal1 6452 5361 6486 5367 1 gnd
rlabel metal1 6455 5754 6483 5759 1 vdd
rlabel locali 5347 5221 5369 5236 1 d0
rlabel metal1 5516 5444 5544 5449 1 vdd
rlabel metal1 5513 5051 5547 5057 1 gnd
rlabel metal1 6595 6265 6623 6270 1 vdd
rlabel metal1 6592 5872 6626 5878 1 gnd
rlabel locali 6423 6037 6444 6056 1 d2
rlabel metal1 6564 7381 6592 7386 1 vdd
rlabel metal1 6561 6988 6595 6994 1 gnd
rlabel locali 6394 7157 6420 7174 1 d3
rlabel locali 6396 2745 6422 2762 1 d3
rlabel metal1 6563 2576 6597 2582 1 gnd
rlabel metal1 6566 2969 6594 2974 1 vdd
rlabel locali 6425 1625 6446 1644 1 d2
rlabel metal1 6594 1460 6628 1466 1 gnd
rlabel metal1 6597 1853 6625 1858 1 vdd
rlabel metal1 5515 639 5549 645 1 gnd
rlabel metal1 5518 1032 5546 1037 1 vdd
rlabel locali 5349 809 5371 824 1 d0
rlabel metal1 6457 1342 6485 1347 1 vdd
rlabel metal1 6454 949 6488 955 1 gnd
rlabel locali 6287 1115 6315 1136 1 d1
rlabel metal1 5516 1193 5550 1199 1 gnd
rlabel metal1 5519 1586 5547 1591 1 vdd
rlabel locali 5350 1363 5372 1378 1 d0
rlabel metal1 5514 1742 5548 1748 1 gnd
rlabel metal1 5517 2135 5545 2140 1 vdd
rlabel locali 5348 1912 5370 1927 1 d0
rlabel metal1 6456 2445 6484 2450 1 vdd
rlabel metal1 6453 2052 6487 2058 1 gnd
rlabel locali 6286 2218 6314 2239 1 d1
rlabel metal1 5515 2296 5549 2302 1 gnd
rlabel metal1 5518 2689 5546 2694 1 vdd
rlabel locali 5349 2466 5371 2481 1 d0
rlabel locali 6424 3831 6445 3850 1 d2
rlabel metal1 6593 3666 6627 3672 1 gnd
rlabel metal1 6596 4059 6624 4064 1 vdd
rlabel metal1 5514 2845 5548 2851 1 gnd
rlabel metal1 5517 3238 5545 3243 1 vdd
rlabel locali 5348 3015 5370 3030 1 d0
rlabel metal1 6456 3548 6484 3553 1 vdd
rlabel metal1 6453 3155 6487 3161 1 gnd
rlabel locali 6286 3321 6314 3342 1 d1
rlabel metal1 5515 3399 5549 3405 1 gnd
rlabel metal1 5518 3792 5546 3797 1 vdd
rlabel locali 5349 3569 5371 3584 1 d0
rlabel metal1 5513 3948 5547 3954 1 gnd
rlabel metal1 5516 4341 5544 4346 1 vdd
rlabel locali 5347 4118 5369 4133 1 d0
rlabel metal1 6455 4651 6483 4656 1 vdd
rlabel metal1 6452 4258 6486 4264 1 gnd
rlabel locali 6285 4424 6313 4445 1 d1
rlabel metal1 5514 4502 5548 4508 1 gnd
rlabel metal1 5517 4895 5545 4900 1 vdd
rlabel locali 5348 4672 5370 4687 1 d0
rlabel metal1 6564 5181 6592 5186 1 vdd
rlabel metal1 6561 4788 6595 4794 1 gnd
rlabel locali 6388 4950 6423 4976 1 d4
rlabel locali 9677 930 9699 945 5 d0
rlabel metal1 9502 717 9530 722 5 vdd
rlabel metal1 9499 1109 9533 1115 5 gnd
rlabel locali 8734 1172 8762 1193 5 d1
rlabel metal1 8561 1353 8595 1359 5 gnd
rlabel metal1 8564 961 8592 966 5 vdd
rlabel locali 9678 1484 9700 1499 5 d0
rlabel metal1 9503 1271 9531 1276 5 vdd
rlabel metal1 9500 1663 9534 1669 5 gnd
rlabel locali 9676 2033 9698 2048 5 d0
rlabel metal1 9501 1820 9529 1825 5 vdd
rlabel metal1 9498 2212 9532 2218 5 gnd
rlabel locali 8733 2275 8761 2296 5 d1
rlabel metal1 8560 2456 8594 2462 5 gnd
rlabel metal1 8563 2064 8591 2069 5 vdd
rlabel locali 9677 2587 9699 2602 5 d0
rlabel metal1 9502 2374 9530 2379 5 vdd
rlabel metal1 9499 2766 9533 2772 5 gnd
rlabel metal1 8423 1553 8451 1558 5 vdd
rlabel metal1 8420 1945 8454 1951 5 gnd
rlabel locali 8602 1767 8623 1786 5 d2
rlabel locali 9676 3136 9698 3151 5 d0
rlabel metal1 9501 2923 9529 2928 5 vdd
rlabel metal1 9498 3315 9532 3321 5 gnd
rlabel locali 8733 3378 8761 3399 5 d1
rlabel metal1 8560 3559 8594 3565 5 gnd
rlabel metal1 8563 3167 8591 3172 5 vdd
rlabel locali 9677 3690 9699 3705 5 d0
rlabel metal1 9502 3477 9530 3482 5 vdd
rlabel metal1 9499 3869 9533 3875 5 gnd
rlabel locali 9675 4239 9697 4254 5 d0
rlabel metal1 9500 4026 9528 4031 5 vdd
rlabel metal1 9497 4418 9531 4424 5 gnd
rlabel locali 8732 4481 8760 4502 5 d1
rlabel metal1 8559 4662 8593 4668 5 gnd
rlabel metal1 8562 4270 8590 4275 5 vdd
rlabel locali 9676 4793 9698 4808 5 d0
rlabel metal1 9501 4580 9529 4585 5 vdd
rlabel metal1 9498 4972 9532 4978 5 gnd
rlabel metal1 8422 3759 8450 3764 5 vdd
rlabel metal1 8419 4151 8453 4157 5 gnd
rlabel locali 8601 3973 8622 3992 5 d2
rlabel metal1 8453 2643 8481 2648 5 vdd
rlabel metal1 8450 3035 8484 3041 5 gnd
rlabel locali 8625 2855 8651 2872 5 d3
rlabel locali 8623 7267 8649 7284 5 d3
rlabel metal1 8448 7447 8482 7453 5 gnd
rlabel metal1 8451 7055 8479 7060 5 vdd
rlabel locali 8599 8385 8620 8404 5 d2
rlabel metal1 8417 8563 8451 8569 5 gnd
rlabel metal1 8420 8171 8448 8176 5 vdd
rlabel metal1 9496 9384 9530 9390 5 gnd
rlabel metal1 9499 8992 9527 8997 5 vdd
rlabel locali 9674 9205 9696 9220 5 d0
rlabel metal1 8560 8682 8588 8687 5 vdd
rlabel metal1 8557 9074 8591 9080 5 gnd
rlabel locali 8730 8893 8758 8914 5 d1
rlabel metal1 9495 8830 9529 8836 5 gnd
rlabel metal1 9498 8438 9526 8443 5 vdd
rlabel locali 9673 8651 9695 8666 5 d0
rlabel metal1 9497 8281 9531 8287 5 gnd
rlabel metal1 9500 7889 9528 7894 5 vdd
rlabel locali 9675 8102 9697 8117 5 d0
rlabel metal1 8561 7579 8589 7584 5 vdd
rlabel metal1 8558 7971 8592 7977 5 gnd
rlabel locali 8731 7790 8759 7811 5 d1
rlabel metal1 9496 7727 9530 7733 5 gnd
rlabel metal1 9499 7335 9527 7340 5 vdd
rlabel locali 9674 7548 9696 7563 5 d0
rlabel locali 8600 6179 8621 6198 5 d2
rlabel metal1 8418 6357 8452 6363 5 gnd
rlabel metal1 8421 5965 8449 5970 5 vdd
rlabel metal1 9497 7178 9531 7184 5 gnd
rlabel metal1 9500 6786 9528 6791 5 vdd
rlabel locali 9675 6999 9697 7014 5 d0
rlabel metal1 8561 6476 8589 6481 5 vdd
rlabel metal1 8558 6868 8592 6874 5 gnd
rlabel locali 8731 6687 8759 6708 5 d1
rlabel metal1 9496 6624 9530 6630 5 gnd
rlabel metal1 9499 6232 9527 6237 5 vdd
rlabel locali 9674 6445 9696 6460 5 d0
rlabel metal1 9498 6075 9532 6081 5 gnd
rlabel metal1 9501 5683 9529 5688 5 vdd
rlabel locali 9676 5896 9698 5911 5 d0
rlabel metal1 8562 5373 8590 5378 5 vdd
rlabel metal1 8559 5765 8593 5771 5 gnd
rlabel locali 8732 5584 8760 5605 5 d1
rlabel metal1 9497 5521 9531 5527 5 gnd
rlabel metal1 9500 5129 9528 5134 5 vdd
rlabel locali 9675 5342 9697 5357 5 d0
rlabel metal1 8453 4843 8481 4848 5 vdd
rlabel metal1 8450 5235 8484 5241 5 gnd
rlabel locali 8622 5053 8657 5079 5 d4
rlabel metal1 6765 473 6793 478 1 vdd
rlabel metal1 6762 80 6796 86 1 gnd
rlabel locali 6591 244 6619 266 1 d5
rlabel locali 5120 224 5142 239 1 vout
rlabel metal1 4659 412 4687 417 1 vdd
rlabel metal1 4656 19 4690 25 1 gnd
rlabel locali 4488 182 4515 208 1 d6
<< end >>
