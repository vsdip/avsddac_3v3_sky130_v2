magic
tech sky130A
timestamp 1633159112
<< nwell >>
rect 755 11541 1566 11765
rect 1803 11537 2614 11761
rect 9041 11286 9852 11510
rect 755 10862 1566 11086
rect 3250 10857 4061 11081
rect 7993 10611 8804 10835
rect 9041 10607 9852 10831
rect 755 10094 1566 10318
rect 1803 10090 2614 10314
rect 6546 9844 7357 10068
rect 9041 9839 9852 10063
rect 755 9415 1566 9639
rect 3293 9412 4104 9636
rect 7993 9164 8804 9388
rect 9041 9160 9852 9384
rect 756 8574 1567 8798
rect 1804 8570 2615 8794
rect 6504 8322 7315 8546
rect 9042 8319 9853 8543
rect 756 7895 1567 8119
rect 3251 7890 4062 8114
rect 7994 7644 8805 7868
rect 9042 7640 9853 7864
rect 756 7127 1567 7351
rect 1804 7123 2615 7347
rect 6547 6877 7358 7101
rect 9042 6872 9853 7096
rect 756 6448 1567 6672
rect 4359 6439 5170 6663
rect 7994 6197 8805 6421
rect 9042 6193 9853 6417
rect 753 5533 1564 5757
rect 1801 5529 2612 5753
rect 5436 5287 6247 5511
rect 9039 5278 9850 5502
rect 753 4854 1564 5078
rect 3248 4849 4059 5073
rect 7991 4603 8802 4827
rect 9039 4599 9850 4823
rect 753 4086 1564 4310
rect 1801 4082 2612 4306
rect 6544 3836 7355 4060
rect 9039 3831 9850 4055
rect 753 3407 1564 3631
rect 3291 3404 4102 3628
rect 7991 3156 8802 3380
rect 9039 3152 9850 3376
rect 754 2566 1565 2790
rect 1802 2562 2613 2786
rect 4704 2568 5515 2792
rect 6502 2314 7313 2538
rect 9040 2311 9851 2535
rect 754 1887 1565 2111
rect 3249 1882 4060 2106
rect 7992 1636 8803 1860
rect 9040 1632 9851 1856
rect 754 1119 1565 1343
rect 1802 1115 2613 1339
rect 6545 869 7356 1093
rect 9040 864 9851 1088
rect 754 440 1565 664
rect 7992 189 8803 413
rect 9040 185 9851 409
<< nmos >>
rect 9109 11569 9159 11611
rect 9317 11569 9367 11611
rect 9525 11569 9575 11611
rect 9738 11569 9788 11611
rect 819 11440 869 11482
rect 1032 11440 1082 11482
rect 1240 11440 1290 11482
rect 1448 11440 1498 11482
rect 1867 11436 1917 11478
rect 2080 11436 2130 11478
rect 2288 11436 2338 11478
rect 2496 11436 2546 11478
rect 8061 10894 8111 10936
rect 8269 10894 8319 10936
rect 8477 10894 8527 10936
rect 8690 10894 8740 10936
rect 819 10761 869 10803
rect 1032 10761 1082 10803
rect 1240 10761 1290 10803
rect 1448 10761 1498 10803
rect 9109 10890 9159 10932
rect 9317 10890 9367 10932
rect 9525 10890 9575 10932
rect 9738 10890 9788 10932
rect 3314 10756 3364 10798
rect 3527 10756 3577 10798
rect 3735 10756 3785 10798
rect 3943 10756 3993 10798
rect 6614 10127 6664 10169
rect 6822 10127 6872 10169
rect 7030 10127 7080 10169
rect 7243 10127 7293 10169
rect 819 9993 869 10035
rect 1032 9993 1082 10035
rect 1240 9993 1290 10035
rect 1448 9993 1498 10035
rect 9109 10122 9159 10164
rect 9317 10122 9367 10164
rect 9525 10122 9575 10164
rect 9738 10122 9788 10164
rect 1867 9989 1917 10031
rect 2080 9989 2130 10031
rect 2288 9989 2338 10031
rect 2496 9989 2546 10031
rect 8061 9447 8111 9489
rect 8269 9447 8319 9489
rect 8477 9447 8527 9489
rect 8690 9447 8740 9489
rect 819 9314 869 9356
rect 1032 9314 1082 9356
rect 1240 9314 1290 9356
rect 1448 9314 1498 9356
rect 9109 9443 9159 9485
rect 9317 9443 9367 9485
rect 9525 9443 9575 9485
rect 9738 9443 9788 9485
rect 3357 9311 3407 9353
rect 3570 9311 3620 9353
rect 3778 9311 3828 9353
rect 3986 9311 4036 9353
rect 6572 8605 6622 8647
rect 6780 8605 6830 8647
rect 6988 8605 7038 8647
rect 7201 8605 7251 8647
rect 820 8473 870 8515
rect 1033 8473 1083 8515
rect 1241 8473 1291 8515
rect 1449 8473 1499 8515
rect 9110 8602 9160 8644
rect 9318 8602 9368 8644
rect 9526 8602 9576 8644
rect 9739 8602 9789 8644
rect 1868 8469 1918 8511
rect 2081 8469 2131 8511
rect 2289 8469 2339 8511
rect 2497 8469 2547 8511
rect 8062 7927 8112 7969
rect 8270 7927 8320 7969
rect 8478 7927 8528 7969
rect 8691 7927 8741 7969
rect 820 7794 870 7836
rect 1033 7794 1083 7836
rect 1241 7794 1291 7836
rect 1449 7794 1499 7836
rect 9110 7923 9160 7965
rect 9318 7923 9368 7965
rect 9526 7923 9576 7965
rect 9739 7923 9789 7965
rect 3315 7789 3365 7831
rect 3528 7789 3578 7831
rect 3736 7789 3786 7831
rect 3944 7789 3994 7831
rect 6615 7160 6665 7202
rect 6823 7160 6873 7202
rect 7031 7160 7081 7202
rect 7244 7160 7294 7202
rect 820 7026 870 7068
rect 1033 7026 1083 7068
rect 1241 7026 1291 7068
rect 1449 7026 1499 7068
rect 9110 7155 9160 7197
rect 9318 7155 9368 7197
rect 9526 7155 9576 7197
rect 9739 7155 9789 7197
rect 1868 7022 1918 7064
rect 2081 7022 2131 7064
rect 2289 7022 2339 7064
rect 2497 7022 2547 7064
rect 8062 6480 8112 6522
rect 8270 6480 8320 6522
rect 8478 6480 8528 6522
rect 8691 6480 8741 6522
rect 820 6347 870 6389
rect 1033 6347 1083 6389
rect 1241 6347 1291 6389
rect 1449 6347 1499 6389
rect 9110 6476 9160 6518
rect 9318 6476 9368 6518
rect 9526 6476 9576 6518
rect 9739 6476 9789 6518
rect 4423 6338 4473 6380
rect 4636 6338 4686 6380
rect 4844 6338 4894 6380
rect 5052 6338 5102 6380
rect 5504 5570 5554 5612
rect 5712 5570 5762 5612
rect 5920 5570 5970 5612
rect 6133 5570 6183 5612
rect 817 5432 867 5474
rect 1030 5432 1080 5474
rect 1238 5432 1288 5474
rect 1446 5432 1496 5474
rect 9107 5561 9157 5603
rect 9315 5561 9365 5603
rect 9523 5561 9573 5603
rect 9736 5561 9786 5603
rect 1865 5428 1915 5470
rect 2078 5428 2128 5470
rect 2286 5428 2336 5470
rect 2494 5428 2544 5470
rect 8059 4886 8109 4928
rect 8267 4886 8317 4928
rect 8475 4886 8525 4928
rect 8688 4886 8738 4928
rect 817 4753 867 4795
rect 1030 4753 1080 4795
rect 1238 4753 1288 4795
rect 1446 4753 1496 4795
rect 9107 4882 9157 4924
rect 9315 4882 9365 4924
rect 9523 4882 9573 4924
rect 9736 4882 9786 4924
rect 3312 4748 3362 4790
rect 3525 4748 3575 4790
rect 3733 4748 3783 4790
rect 3941 4748 3991 4790
rect 6612 4119 6662 4161
rect 6820 4119 6870 4161
rect 7028 4119 7078 4161
rect 7241 4119 7291 4161
rect 817 3985 867 4027
rect 1030 3985 1080 4027
rect 1238 3985 1288 4027
rect 1446 3985 1496 4027
rect 9107 4114 9157 4156
rect 9315 4114 9365 4156
rect 9523 4114 9573 4156
rect 9736 4114 9786 4156
rect 1865 3981 1915 4023
rect 2078 3981 2128 4023
rect 2286 3981 2336 4023
rect 2494 3981 2544 4023
rect 8059 3439 8109 3481
rect 8267 3439 8317 3481
rect 8475 3439 8525 3481
rect 8688 3439 8738 3481
rect 817 3306 867 3348
rect 1030 3306 1080 3348
rect 1238 3306 1288 3348
rect 1446 3306 1496 3348
rect 9107 3435 9157 3477
rect 9315 3435 9365 3477
rect 9523 3435 9573 3477
rect 9736 3435 9786 3477
rect 3355 3303 3405 3345
rect 3568 3303 3618 3345
rect 3776 3303 3826 3345
rect 3984 3303 4034 3345
rect 6570 2597 6620 2639
rect 6778 2597 6828 2639
rect 6986 2597 7036 2639
rect 7199 2597 7249 2639
rect 818 2465 868 2507
rect 1031 2465 1081 2507
rect 1239 2465 1289 2507
rect 1447 2465 1497 2507
rect 9108 2594 9158 2636
rect 9316 2594 9366 2636
rect 9524 2594 9574 2636
rect 9737 2594 9787 2636
rect 1866 2461 1916 2503
rect 2079 2461 2129 2503
rect 2287 2461 2337 2503
rect 2495 2461 2545 2503
rect 4768 2467 4818 2509
rect 4981 2467 5031 2509
rect 5189 2467 5239 2509
rect 5397 2467 5447 2509
rect 8060 1919 8110 1961
rect 8268 1919 8318 1961
rect 8476 1919 8526 1961
rect 8689 1919 8739 1961
rect 818 1786 868 1828
rect 1031 1786 1081 1828
rect 1239 1786 1289 1828
rect 1447 1786 1497 1828
rect 9108 1915 9158 1957
rect 9316 1915 9366 1957
rect 9524 1915 9574 1957
rect 9737 1915 9787 1957
rect 3313 1781 3363 1823
rect 3526 1781 3576 1823
rect 3734 1781 3784 1823
rect 3942 1781 3992 1823
rect 6613 1152 6663 1194
rect 6821 1152 6871 1194
rect 7029 1152 7079 1194
rect 7242 1152 7292 1194
rect 818 1018 868 1060
rect 1031 1018 1081 1060
rect 1239 1018 1289 1060
rect 1447 1018 1497 1060
rect 9108 1147 9158 1189
rect 9316 1147 9366 1189
rect 9524 1147 9574 1189
rect 9737 1147 9787 1189
rect 1866 1014 1916 1056
rect 2079 1014 2129 1056
rect 2287 1014 2337 1056
rect 2495 1014 2545 1056
rect 8060 472 8110 514
rect 8268 472 8318 514
rect 8476 472 8526 514
rect 8689 472 8739 514
rect 9108 468 9158 510
rect 9316 468 9366 510
rect 9524 468 9574 510
rect 9737 468 9787 510
rect 818 339 868 381
rect 1031 339 1081 381
rect 1239 339 1289 381
rect 1447 339 1497 381
<< pmos >>
rect 819 11559 869 11659
rect 1032 11559 1082 11659
rect 1240 11559 1290 11659
rect 1448 11559 1498 11659
rect 1867 11555 1917 11655
rect 2080 11555 2130 11655
rect 2288 11555 2338 11655
rect 2496 11555 2546 11655
rect 9109 11392 9159 11492
rect 9317 11392 9367 11492
rect 9525 11392 9575 11492
rect 9738 11392 9788 11492
rect 819 10880 869 10980
rect 1032 10880 1082 10980
rect 1240 10880 1290 10980
rect 1448 10880 1498 10980
rect 3314 10875 3364 10975
rect 3527 10875 3577 10975
rect 3735 10875 3785 10975
rect 3943 10875 3993 10975
rect 8061 10717 8111 10817
rect 8269 10717 8319 10817
rect 8477 10717 8527 10817
rect 8690 10717 8740 10817
rect 9109 10713 9159 10813
rect 9317 10713 9367 10813
rect 9525 10713 9575 10813
rect 9738 10713 9788 10813
rect 819 10112 869 10212
rect 1032 10112 1082 10212
rect 1240 10112 1290 10212
rect 1448 10112 1498 10212
rect 1867 10108 1917 10208
rect 2080 10108 2130 10208
rect 2288 10108 2338 10208
rect 2496 10108 2546 10208
rect 6614 9950 6664 10050
rect 6822 9950 6872 10050
rect 7030 9950 7080 10050
rect 7243 9950 7293 10050
rect 9109 9945 9159 10045
rect 9317 9945 9367 10045
rect 9525 9945 9575 10045
rect 9738 9945 9788 10045
rect 819 9433 869 9533
rect 1032 9433 1082 9533
rect 1240 9433 1290 9533
rect 1448 9433 1498 9533
rect 3357 9430 3407 9530
rect 3570 9430 3620 9530
rect 3778 9430 3828 9530
rect 3986 9430 4036 9530
rect 8061 9270 8111 9370
rect 8269 9270 8319 9370
rect 8477 9270 8527 9370
rect 8690 9270 8740 9370
rect 9109 9266 9159 9366
rect 9317 9266 9367 9366
rect 9525 9266 9575 9366
rect 9738 9266 9788 9366
rect 820 8592 870 8692
rect 1033 8592 1083 8692
rect 1241 8592 1291 8692
rect 1449 8592 1499 8692
rect 1868 8588 1918 8688
rect 2081 8588 2131 8688
rect 2289 8588 2339 8688
rect 2497 8588 2547 8688
rect 6572 8428 6622 8528
rect 6780 8428 6830 8528
rect 6988 8428 7038 8528
rect 7201 8428 7251 8528
rect 9110 8425 9160 8525
rect 9318 8425 9368 8525
rect 9526 8425 9576 8525
rect 9739 8425 9789 8525
rect 820 7913 870 8013
rect 1033 7913 1083 8013
rect 1241 7913 1291 8013
rect 1449 7913 1499 8013
rect 3315 7908 3365 8008
rect 3528 7908 3578 8008
rect 3736 7908 3786 8008
rect 3944 7908 3994 8008
rect 8062 7750 8112 7850
rect 8270 7750 8320 7850
rect 8478 7750 8528 7850
rect 8691 7750 8741 7850
rect 9110 7746 9160 7846
rect 9318 7746 9368 7846
rect 9526 7746 9576 7846
rect 9739 7746 9789 7846
rect 820 7145 870 7245
rect 1033 7145 1083 7245
rect 1241 7145 1291 7245
rect 1449 7145 1499 7245
rect 1868 7141 1918 7241
rect 2081 7141 2131 7241
rect 2289 7141 2339 7241
rect 2497 7141 2547 7241
rect 6615 6983 6665 7083
rect 6823 6983 6873 7083
rect 7031 6983 7081 7083
rect 7244 6983 7294 7083
rect 9110 6978 9160 7078
rect 9318 6978 9368 7078
rect 9526 6978 9576 7078
rect 9739 6978 9789 7078
rect 820 6466 870 6566
rect 1033 6466 1083 6566
rect 1241 6466 1291 6566
rect 1449 6466 1499 6566
rect 4423 6457 4473 6557
rect 4636 6457 4686 6557
rect 4844 6457 4894 6557
rect 5052 6457 5102 6557
rect 8062 6303 8112 6403
rect 8270 6303 8320 6403
rect 8478 6303 8528 6403
rect 8691 6303 8741 6403
rect 9110 6299 9160 6399
rect 9318 6299 9368 6399
rect 9526 6299 9576 6399
rect 9739 6299 9789 6399
rect 817 5551 867 5651
rect 1030 5551 1080 5651
rect 1238 5551 1288 5651
rect 1446 5551 1496 5651
rect 1865 5547 1915 5647
rect 2078 5547 2128 5647
rect 2286 5547 2336 5647
rect 2494 5547 2544 5647
rect 5504 5393 5554 5493
rect 5712 5393 5762 5493
rect 5920 5393 5970 5493
rect 6133 5393 6183 5493
rect 9107 5384 9157 5484
rect 9315 5384 9365 5484
rect 9523 5384 9573 5484
rect 9736 5384 9786 5484
rect 817 4872 867 4972
rect 1030 4872 1080 4972
rect 1238 4872 1288 4972
rect 1446 4872 1496 4972
rect 3312 4867 3362 4967
rect 3525 4867 3575 4967
rect 3733 4867 3783 4967
rect 3941 4867 3991 4967
rect 8059 4709 8109 4809
rect 8267 4709 8317 4809
rect 8475 4709 8525 4809
rect 8688 4709 8738 4809
rect 9107 4705 9157 4805
rect 9315 4705 9365 4805
rect 9523 4705 9573 4805
rect 9736 4705 9786 4805
rect 817 4104 867 4204
rect 1030 4104 1080 4204
rect 1238 4104 1288 4204
rect 1446 4104 1496 4204
rect 1865 4100 1915 4200
rect 2078 4100 2128 4200
rect 2286 4100 2336 4200
rect 2494 4100 2544 4200
rect 6612 3942 6662 4042
rect 6820 3942 6870 4042
rect 7028 3942 7078 4042
rect 7241 3942 7291 4042
rect 9107 3937 9157 4037
rect 9315 3937 9365 4037
rect 9523 3937 9573 4037
rect 9736 3937 9786 4037
rect 817 3425 867 3525
rect 1030 3425 1080 3525
rect 1238 3425 1288 3525
rect 1446 3425 1496 3525
rect 3355 3422 3405 3522
rect 3568 3422 3618 3522
rect 3776 3422 3826 3522
rect 3984 3422 4034 3522
rect 8059 3262 8109 3362
rect 8267 3262 8317 3362
rect 8475 3262 8525 3362
rect 8688 3262 8738 3362
rect 9107 3258 9157 3358
rect 9315 3258 9365 3358
rect 9523 3258 9573 3358
rect 9736 3258 9786 3358
rect 818 2584 868 2684
rect 1031 2584 1081 2684
rect 1239 2584 1289 2684
rect 1447 2584 1497 2684
rect 1866 2580 1916 2680
rect 2079 2580 2129 2680
rect 2287 2580 2337 2680
rect 2495 2580 2545 2680
rect 4768 2586 4818 2686
rect 4981 2586 5031 2686
rect 5189 2586 5239 2686
rect 5397 2586 5447 2686
rect 6570 2420 6620 2520
rect 6778 2420 6828 2520
rect 6986 2420 7036 2520
rect 7199 2420 7249 2520
rect 9108 2417 9158 2517
rect 9316 2417 9366 2517
rect 9524 2417 9574 2517
rect 9737 2417 9787 2517
rect 818 1905 868 2005
rect 1031 1905 1081 2005
rect 1239 1905 1289 2005
rect 1447 1905 1497 2005
rect 3313 1900 3363 2000
rect 3526 1900 3576 2000
rect 3734 1900 3784 2000
rect 3942 1900 3992 2000
rect 8060 1742 8110 1842
rect 8268 1742 8318 1842
rect 8476 1742 8526 1842
rect 8689 1742 8739 1842
rect 9108 1738 9158 1838
rect 9316 1738 9366 1838
rect 9524 1738 9574 1838
rect 9737 1738 9787 1838
rect 818 1137 868 1237
rect 1031 1137 1081 1237
rect 1239 1137 1289 1237
rect 1447 1137 1497 1237
rect 1866 1133 1916 1233
rect 2079 1133 2129 1233
rect 2287 1133 2337 1233
rect 2495 1133 2545 1233
rect 6613 975 6663 1075
rect 6821 975 6871 1075
rect 7029 975 7079 1075
rect 7242 975 7292 1075
rect 9108 970 9158 1070
rect 9316 970 9366 1070
rect 9524 970 9574 1070
rect 9737 970 9787 1070
rect 818 458 868 558
rect 1031 458 1081 558
rect 1239 458 1289 558
rect 1447 458 1497 558
rect 8060 295 8110 395
rect 8268 295 8318 395
rect 8476 295 8526 395
rect 8689 295 8739 395
rect 9108 291 9158 391
rect 9316 291 9366 391
rect 9524 291 9574 391
rect 9737 291 9787 391
<< ndiff >>
rect 9060 11599 9109 11611
rect 9060 11579 9071 11599
rect 9091 11579 9109 11599
rect 9060 11569 9109 11579
rect 9159 11595 9203 11611
rect 9159 11575 9174 11595
rect 9194 11575 9203 11595
rect 9159 11569 9203 11575
rect 9273 11595 9317 11611
rect 9273 11575 9282 11595
rect 9302 11575 9317 11595
rect 9273 11569 9317 11575
rect 9367 11599 9416 11611
rect 9367 11579 9385 11599
rect 9405 11579 9416 11599
rect 9367 11569 9416 11579
rect 9481 11595 9525 11611
rect 9481 11575 9490 11595
rect 9510 11575 9525 11595
rect 9481 11569 9525 11575
rect 9575 11599 9624 11611
rect 9575 11579 9593 11599
rect 9613 11579 9624 11599
rect 9575 11569 9624 11579
rect 9694 11595 9738 11611
rect 9694 11575 9703 11595
rect 9723 11575 9738 11595
rect 9694 11569 9738 11575
rect 9788 11599 9837 11611
rect 9788 11579 9806 11599
rect 9826 11579 9837 11599
rect 9788 11569 9837 11579
rect 770 11472 819 11482
rect 770 11452 781 11472
rect 801 11452 819 11472
rect 770 11440 819 11452
rect 869 11476 913 11482
rect 869 11456 884 11476
rect 904 11456 913 11476
rect 869 11440 913 11456
rect 983 11472 1032 11482
rect 983 11452 994 11472
rect 1014 11452 1032 11472
rect 983 11440 1032 11452
rect 1082 11476 1126 11482
rect 1082 11456 1097 11476
rect 1117 11456 1126 11476
rect 1082 11440 1126 11456
rect 1191 11472 1240 11482
rect 1191 11452 1202 11472
rect 1222 11452 1240 11472
rect 1191 11440 1240 11452
rect 1290 11476 1334 11482
rect 1290 11456 1305 11476
rect 1325 11456 1334 11476
rect 1290 11440 1334 11456
rect 1404 11476 1448 11482
rect 1404 11456 1413 11476
rect 1433 11456 1448 11476
rect 1404 11440 1448 11456
rect 1498 11472 1547 11482
rect 1498 11452 1516 11472
rect 1536 11452 1547 11472
rect 1498 11440 1547 11452
rect 1818 11468 1867 11478
rect 1818 11448 1829 11468
rect 1849 11448 1867 11468
rect 1818 11436 1867 11448
rect 1917 11472 1961 11478
rect 1917 11452 1932 11472
rect 1952 11452 1961 11472
rect 1917 11436 1961 11452
rect 2031 11468 2080 11478
rect 2031 11448 2042 11468
rect 2062 11448 2080 11468
rect 2031 11436 2080 11448
rect 2130 11472 2174 11478
rect 2130 11452 2145 11472
rect 2165 11452 2174 11472
rect 2130 11436 2174 11452
rect 2239 11468 2288 11478
rect 2239 11448 2250 11468
rect 2270 11448 2288 11468
rect 2239 11436 2288 11448
rect 2338 11472 2382 11478
rect 2338 11452 2353 11472
rect 2373 11452 2382 11472
rect 2338 11436 2382 11452
rect 2452 11472 2496 11478
rect 2452 11452 2461 11472
rect 2481 11452 2496 11472
rect 2452 11436 2496 11452
rect 2546 11468 2595 11478
rect 2546 11448 2564 11468
rect 2584 11448 2595 11468
rect 2546 11436 2595 11448
rect 8012 10924 8061 10936
rect 8012 10904 8023 10924
rect 8043 10904 8061 10924
rect 8012 10894 8061 10904
rect 8111 10920 8155 10936
rect 8111 10900 8126 10920
rect 8146 10900 8155 10920
rect 8111 10894 8155 10900
rect 8225 10920 8269 10936
rect 8225 10900 8234 10920
rect 8254 10900 8269 10920
rect 8225 10894 8269 10900
rect 8319 10924 8368 10936
rect 8319 10904 8337 10924
rect 8357 10904 8368 10924
rect 8319 10894 8368 10904
rect 8433 10920 8477 10936
rect 8433 10900 8442 10920
rect 8462 10900 8477 10920
rect 8433 10894 8477 10900
rect 8527 10924 8576 10936
rect 8527 10904 8545 10924
rect 8565 10904 8576 10924
rect 8527 10894 8576 10904
rect 8646 10920 8690 10936
rect 8646 10900 8655 10920
rect 8675 10900 8690 10920
rect 8646 10894 8690 10900
rect 8740 10924 8789 10936
rect 8740 10904 8758 10924
rect 8778 10904 8789 10924
rect 8740 10894 8789 10904
rect 9060 10920 9109 10932
rect 9060 10900 9071 10920
rect 9091 10900 9109 10920
rect 770 10793 819 10803
rect 770 10773 781 10793
rect 801 10773 819 10793
rect 770 10761 819 10773
rect 869 10797 913 10803
rect 869 10777 884 10797
rect 904 10777 913 10797
rect 869 10761 913 10777
rect 983 10793 1032 10803
rect 983 10773 994 10793
rect 1014 10773 1032 10793
rect 983 10761 1032 10773
rect 1082 10797 1126 10803
rect 1082 10777 1097 10797
rect 1117 10777 1126 10797
rect 1082 10761 1126 10777
rect 1191 10793 1240 10803
rect 1191 10773 1202 10793
rect 1222 10773 1240 10793
rect 1191 10761 1240 10773
rect 1290 10797 1334 10803
rect 1290 10777 1305 10797
rect 1325 10777 1334 10797
rect 1290 10761 1334 10777
rect 1404 10797 1448 10803
rect 1404 10777 1413 10797
rect 1433 10777 1448 10797
rect 1404 10761 1448 10777
rect 1498 10793 1547 10803
rect 9060 10890 9109 10900
rect 9159 10916 9203 10932
rect 9159 10896 9174 10916
rect 9194 10896 9203 10916
rect 9159 10890 9203 10896
rect 9273 10916 9317 10932
rect 9273 10896 9282 10916
rect 9302 10896 9317 10916
rect 9273 10890 9317 10896
rect 9367 10920 9416 10932
rect 9367 10900 9385 10920
rect 9405 10900 9416 10920
rect 9367 10890 9416 10900
rect 9481 10916 9525 10932
rect 9481 10896 9490 10916
rect 9510 10896 9525 10916
rect 9481 10890 9525 10896
rect 9575 10920 9624 10932
rect 9575 10900 9593 10920
rect 9613 10900 9624 10920
rect 9575 10890 9624 10900
rect 9694 10916 9738 10932
rect 9694 10896 9703 10916
rect 9723 10896 9738 10916
rect 9694 10890 9738 10896
rect 9788 10920 9837 10932
rect 9788 10900 9806 10920
rect 9826 10900 9837 10920
rect 9788 10890 9837 10900
rect 1498 10773 1516 10793
rect 1536 10773 1547 10793
rect 1498 10761 1547 10773
rect 3265 10788 3314 10798
rect 3265 10768 3276 10788
rect 3296 10768 3314 10788
rect 3265 10756 3314 10768
rect 3364 10792 3408 10798
rect 3364 10772 3379 10792
rect 3399 10772 3408 10792
rect 3364 10756 3408 10772
rect 3478 10788 3527 10798
rect 3478 10768 3489 10788
rect 3509 10768 3527 10788
rect 3478 10756 3527 10768
rect 3577 10792 3621 10798
rect 3577 10772 3592 10792
rect 3612 10772 3621 10792
rect 3577 10756 3621 10772
rect 3686 10788 3735 10798
rect 3686 10768 3697 10788
rect 3717 10768 3735 10788
rect 3686 10756 3735 10768
rect 3785 10792 3829 10798
rect 3785 10772 3800 10792
rect 3820 10772 3829 10792
rect 3785 10756 3829 10772
rect 3899 10792 3943 10798
rect 3899 10772 3908 10792
rect 3928 10772 3943 10792
rect 3899 10756 3943 10772
rect 3993 10788 4042 10798
rect 3993 10768 4011 10788
rect 4031 10768 4042 10788
rect 3993 10756 4042 10768
rect 6565 10157 6614 10169
rect 6565 10137 6576 10157
rect 6596 10137 6614 10157
rect 6565 10127 6614 10137
rect 6664 10153 6708 10169
rect 6664 10133 6679 10153
rect 6699 10133 6708 10153
rect 6664 10127 6708 10133
rect 6778 10153 6822 10169
rect 6778 10133 6787 10153
rect 6807 10133 6822 10153
rect 6778 10127 6822 10133
rect 6872 10157 6921 10169
rect 6872 10137 6890 10157
rect 6910 10137 6921 10157
rect 6872 10127 6921 10137
rect 6986 10153 7030 10169
rect 6986 10133 6995 10153
rect 7015 10133 7030 10153
rect 6986 10127 7030 10133
rect 7080 10157 7129 10169
rect 7080 10137 7098 10157
rect 7118 10137 7129 10157
rect 7080 10127 7129 10137
rect 7199 10153 7243 10169
rect 7199 10133 7208 10153
rect 7228 10133 7243 10153
rect 7199 10127 7243 10133
rect 7293 10157 7342 10169
rect 7293 10137 7311 10157
rect 7331 10137 7342 10157
rect 7293 10127 7342 10137
rect 9060 10152 9109 10164
rect 9060 10132 9071 10152
rect 9091 10132 9109 10152
rect 770 10025 819 10035
rect 770 10005 781 10025
rect 801 10005 819 10025
rect 770 9993 819 10005
rect 869 10029 913 10035
rect 869 10009 884 10029
rect 904 10009 913 10029
rect 869 9993 913 10009
rect 983 10025 1032 10035
rect 983 10005 994 10025
rect 1014 10005 1032 10025
rect 983 9993 1032 10005
rect 1082 10029 1126 10035
rect 1082 10009 1097 10029
rect 1117 10009 1126 10029
rect 1082 9993 1126 10009
rect 1191 10025 1240 10035
rect 1191 10005 1202 10025
rect 1222 10005 1240 10025
rect 1191 9993 1240 10005
rect 1290 10029 1334 10035
rect 1290 10009 1305 10029
rect 1325 10009 1334 10029
rect 1290 9993 1334 10009
rect 1404 10029 1448 10035
rect 1404 10009 1413 10029
rect 1433 10009 1448 10029
rect 1404 9993 1448 10009
rect 1498 10025 1547 10035
rect 9060 10122 9109 10132
rect 9159 10148 9203 10164
rect 9159 10128 9174 10148
rect 9194 10128 9203 10148
rect 9159 10122 9203 10128
rect 9273 10148 9317 10164
rect 9273 10128 9282 10148
rect 9302 10128 9317 10148
rect 9273 10122 9317 10128
rect 9367 10152 9416 10164
rect 9367 10132 9385 10152
rect 9405 10132 9416 10152
rect 9367 10122 9416 10132
rect 9481 10148 9525 10164
rect 9481 10128 9490 10148
rect 9510 10128 9525 10148
rect 9481 10122 9525 10128
rect 9575 10152 9624 10164
rect 9575 10132 9593 10152
rect 9613 10132 9624 10152
rect 9575 10122 9624 10132
rect 9694 10148 9738 10164
rect 9694 10128 9703 10148
rect 9723 10128 9738 10148
rect 9694 10122 9738 10128
rect 9788 10152 9837 10164
rect 9788 10132 9806 10152
rect 9826 10132 9837 10152
rect 9788 10122 9837 10132
rect 1498 10005 1516 10025
rect 1536 10005 1547 10025
rect 1498 9993 1547 10005
rect 1818 10021 1867 10031
rect 1818 10001 1829 10021
rect 1849 10001 1867 10021
rect 1818 9989 1867 10001
rect 1917 10025 1961 10031
rect 1917 10005 1932 10025
rect 1952 10005 1961 10025
rect 1917 9989 1961 10005
rect 2031 10021 2080 10031
rect 2031 10001 2042 10021
rect 2062 10001 2080 10021
rect 2031 9989 2080 10001
rect 2130 10025 2174 10031
rect 2130 10005 2145 10025
rect 2165 10005 2174 10025
rect 2130 9989 2174 10005
rect 2239 10021 2288 10031
rect 2239 10001 2250 10021
rect 2270 10001 2288 10021
rect 2239 9989 2288 10001
rect 2338 10025 2382 10031
rect 2338 10005 2353 10025
rect 2373 10005 2382 10025
rect 2338 9989 2382 10005
rect 2452 10025 2496 10031
rect 2452 10005 2461 10025
rect 2481 10005 2496 10025
rect 2452 9989 2496 10005
rect 2546 10021 2595 10031
rect 2546 10001 2564 10021
rect 2584 10001 2595 10021
rect 2546 9989 2595 10001
rect 8012 9477 8061 9489
rect 8012 9457 8023 9477
rect 8043 9457 8061 9477
rect 8012 9447 8061 9457
rect 8111 9473 8155 9489
rect 8111 9453 8126 9473
rect 8146 9453 8155 9473
rect 8111 9447 8155 9453
rect 8225 9473 8269 9489
rect 8225 9453 8234 9473
rect 8254 9453 8269 9473
rect 8225 9447 8269 9453
rect 8319 9477 8368 9489
rect 8319 9457 8337 9477
rect 8357 9457 8368 9477
rect 8319 9447 8368 9457
rect 8433 9473 8477 9489
rect 8433 9453 8442 9473
rect 8462 9453 8477 9473
rect 8433 9447 8477 9453
rect 8527 9477 8576 9489
rect 8527 9457 8545 9477
rect 8565 9457 8576 9477
rect 8527 9447 8576 9457
rect 8646 9473 8690 9489
rect 8646 9453 8655 9473
rect 8675 9453 8690 9473
rect 8646 9447 8690 9453
rect 8740 9477 8789 9489
rect 8740 9457 8758 9477
rect 8778 9457 8789 9477
rect 8740 9447 8789 9457
rect 9060 9473 9109 9485
rect 9060 9453 9071 9473
rect 9091 9453 9109 9473
rect 770 9346 819 9356
rect 770 9326 781 9346
rect 801 9326 819 9346
rect 770 9314 819 9326
rect 869 9350 913 9356
rect 869 9330 884 9350
rect 904 9330 913 9350
rect 869 9314 913 9330
rect 983 9346 1032 9356
rect 983 9326 994 9346
rect 1014 9326 1032 9346
rect 983 9314 1032 9326
rect 1082 9350 1126 9356
rect 1082 9330 1097 9350
rect 1117 9330 1126 9350
rect 1082 9314 1126 9330
rect 1191 9346 1240 9356
rect 1191 9326 1202 9346
rect 1222 9326 1240 9346
rect 1191 9314 1240 9326
rect 1290 9350 1334 9356
rect 1290 9330 1305 9350
rect 1325 9330 1334 9350
rect 1290 9314 1334 9330
rect 1404 9350 1448 9356
rect 1404 9330 1413 9350
rect 1433 9330 1448 9350
rect 1404 9314 1448 9330
rect 1498 9346 1547 9356
rect 9060 9443 9109 9453
rect 9159 9469 9203 9485
rect 9159 9449 9174 9469
rect 9194 9449 9203 9469
rect 9159 9443 9203 9449
rect 9273 9469 9317 9485
rect 9273 9449 9282 9469
rect 9302 9449 9317 9469
rect 9273 9443 9317 9449
rect 9367 9473 9416 9485
rect 9367 9453 9385 9473
rect 9405 9453 9416 9473
rect 9367 9443 9416 9453
rect 9481 9469 9525 9485
rect 9481 9449 9490 9469
rect 9510 9449 9525 9469
rect 9481 9443 9525 9449
rect 9575 9473 9624 9485
rect 9575 9453 9593 9473
rect 9613 9453 9624 9473
rect 9575 9443 9624 9453
rect 9694 9469 9738 9485
rect 9694 9449 9703 9469
rect 9723 9449 9738 9469
rect 9694 9443 9738 9449
rect 9788 9473 9837 9485
rect 9788 9453 9806 9473
rect 9826 9453 9837 9473
rect 9788 9443 9837 9453
rect 1498 9326 1516 9346
rect 1536 9326 1547 9346
rect 1498 9314 1547 9326
rect 3308 9343 3357 9353
rect 3308 9323 3319 9343
rect 3339 9323 3357 9343
rect 3308 9311 3357 9323
rect 3407 9347 3451 9353
rect 3407 9327 3422 9347
rect 3442 9327 3451 9347
rect 3407 9311 3451 9327
rect 3521 9343 3570 9353
rect 3521 9323 3532 9343
rect 3552 9323 3570 9343
rect 3521 9311 3570 9323
rect 3620 9347 3664 9353
rect 3620 9327 3635 9347
rect 3655 9327 3664 9347
rect 3620 9311 3664 9327
rect 3729 9343 3778 9353
rect 3729 9323 3740 9343
rect 3760 9323 3778 9343
rect 3729 9311 3778 9323
rect 3828 9347 3872 9353
rect 3828 9327 3843 9347
rect 3863 9327 3872 9347
rect 3828 9311 3872 9327
rect 3942 9347 3986 9353
rect 3942 9327 3951 9347
rect 3971 9327 3986 9347
rect 3942 9311 3986 9327
rect 4036 9343 4085 9353
rect 4036 9323 4054 9343
rect 4074 9323 4085 9343
rect 4036 9311 4085 9323
rect 6523 8635 6572 8647
rect 6523 8615 6534 8635
rect 6554 8615 6572 8635
rect 6523 8605 6572 8615
rect 6622 8631 6666 8647
rect 6622 8611 6637 8631
rect 6657 8611 6666 8631
rect 6622 8605 6666 8611
rect 6736 8631 6780 8647
rect 6736 8611 6745 8631
rect 6765 8611 6780 8631
rect 6736 8605 6780 8611
rect 6830 8635 6879 8647
rect 6830 8615 6848 8635
rect 6868 8615 6879 8635
rect 6830 8605 6879 8615
rect 6944 8631 6988 8647
rect 6944 8611 6953 8631
rect 6973 8611 6988 8631
rect 6944 8605 6988 8611
rect 7038 8635 7087 8647
rect 7038 8615 7056 8635
rect 7076 8615 7087 8635
rect 7038 8605 7087 8615
rect 7157 8631 7201 8647
rect 7157 8611 7166 8631
rect 7186 8611 7201 8631
rect 7157 8605 7201 8611
rect 7251 8635 7300 8647
rect 7251 8615 7269 8635
rect 7289 8615 7300 8635
rect 7251 8605 7300 8615
rect 9061 8632 9110 8644
rect 9061 8612 9072 8632
rect 9092 8612 9110 8632
rect 771 8505 820 8515
rect 771 8485 782 8505
rect 802 8485 820 8505
rect 771 8473 820 8485
rect 870 8509 914 8515
rect 870 8489 885 8509
rect 905 8489 914 8509
rect 870 8473 914 8489
rect 984 8505 1033 8515
rect 984 8485 995 8505
rect 1015 8485 1033 8505
rect 984 8473 1033 8485
rect 1083 8509 1127 8515
rect 1083 8489 1098 8509
rect 1118 8489 1127 8509
rect 1083 8473 1127 8489
rect 1192 8505 1241 8515
rect 1192 8485 1203 8505
rect 1223 8485 1241 8505
rect 1192 8473 1241 8485
rect 1291 8509 1335 8515
rect 1291 8489 1306 8509
rect 1326 8489 1335 8509
rect 1291 8473 1335 8489
rect 1405 8509 1449 8515
rect 1405 8489 1414 8509
rect 1434 8489 1449 8509
rect 1405 8473 1449 8489
rect 1499 8505 1548 8515
rect 9061 8602 9110 8612
rect 9160 8628 9204 8644
rect 9160 8608 9175 8628
rect 9195 8608 9204 8628
rect 9160 8602 9204 8608
rect 9274 8628 9318 8644
rect 9274 8608 9283 8628
rect 9303 8608 9318 8628
rect 9274 8602 9318 8608
rect 9368 8632 9417 8644
rect 9368 8612 9386 8632
rect 9406 8612 9417 8632
rect 9368 8602 9417 8612
rect 9482 8628 9526 8644
rect 9482 8608 9491 8628
rect 9511 8608 9526 8628
rect 9482 8602 9526 8608
rect 9576 8632 9625 8644
rect 9576 8612 9594 8632
rect 9614 8612 9625 8632
rect 9576 8602 9625 8612
rect 9695 8628 9739 8644
rect 9695 8608 9704 8628
rect 9724 8608 9739 8628
rect 9695 8602 9739 8608
rect 9789 8632 9838 8644
rect 9789 8612 9807 8632
rect 9827 8612 9838 8632
rect 9789 8602 9838 8612
rect 1499 8485 1517 8505
rect 1537 8485 1548 8505
rect 1499 8473 1548 8485
rect 1819 8501 1868 8511
rect 1819 8481 1830 8501
rect 1850 8481 1868 8501
rect 1819 8469 1868 8481
rect 1918 8505 1962 8511
rect 1918 8485 1933 8505
rect 1953 8485 1962 8505
rect 1918 8469 1962 8485
rect 2032 8501 2081 8511
rect 2032 8481 2043 8501
rect 2063 8481 2081 8501
rect 2032 8469 2081 8481
rect 2131 8505 2175 8511
rect 2131 8485 2146 8505
rect 2166 8485 2175 8505
rect 2131 8469 2175 8485
rect 2240 8501 2289 8511
rect 2240 8481 2251 8501
rect 2271 8481 2289 8501
rect 2240 8469 2289 8481
rect 2339 8505 2383 8511
rect 2339 8485 2354 8505
rect 2374 8485 2383 8505
rect 2339 8469 2383 8485
rect 2453 8505 2497 8511
rect 2453 8485 2462 8505
rect 2482 8485 2497 8505
rect 2453 8469 2497 8485
rect 2547 8501 2596 8511
rect 2547 8481 2565 8501
rect 2585 8481 2596 8501
rect 2547 8469 2596 8481
rect 8013 7957 8062 7969
rect 8013 7937 8024 7957
rect 8044 7937 8062 7957
rect 8013 7927 8062 7937
rect 8112 7953 8156 7969
rect 8112 7933 8127 7953
rect 8147 7933 8156 7953
rect 8112 7927 8156 7933
rect 8226 7953 8270 7969
rect 8226 7933 8235 7953
rect 8255 7933 8270 7953
rect 8226 7927 8270 7933
rect 8320 7957 8369 7969
rect 8320 7937 8338 7957
rect 8358 7937 8369 7957
rect 8320 7927 8369 7937
rect 8434 7953 8478 7969
rect 8434 7933 8443 7953
rect 8463 7933 8478 7953
rect 8434 7927 8478 7933
rect 8528 7957 8577 7969
rect 8528 7937 8546 7957
rect 8566 7937 8577 7957
rect 8528 7927 8577 7937
rect 8647 7953 8691 7969
rect 8647 7933 8656 7953
rect 8676 7933 8691 7953
rect 8647 7927 8691 7933
rect 8741 7957 8790 7969
rect 8741 7937 8759 7957
rect 8779 7937 8790 7957
rect 8741 7927 8790 7937
rect 9061 7953 9110 7965
rect 9061 7933 9072 7953
rect 9092 7933 9110 7953
rect 771 7826 820 7836
rect 771 7806 782 7826
rect 802 7806 820 7826
rect 771 7794 820 7806
rect 870 7830 914 7836
rect 870 7810 885 7830
rect 905 7810 914 7830
rect 870 7794 914 7810
rect 984 7826 1033 7836
rect 984 7806 995 7826
rect 1015 7806 1033 7826
rect 984 7794 1033 7806
rect 1083 7830 1127 7836
rect 1083 7810 1098 7830
rect 1118 7810 1127 7830
rect 1083 7794 1127 7810
rect 1192 7826 1241 7836
rect 1192 7806 1203 7826
rect 1223 7806 1241 7826
rect 1192 7794 1241 7806
rect 1291 7830 1335 7836
rect 1291 7810 1306 7830
rect 1326 7810 1335 7830
rect 1291 7794 1335 7810
rect 1405 7830 1449 7836
rect 1405 7810 1414 7830
rect 1434 7810 1449 7830
rect 1405 7794 1449 7810
rect 1499 7826 1548 7836
rect 9061 7923 9110 7933
rect 9160 7949 9204 7965
rect 9160 7929 9175 7949
rect 9195 7929 9204 7949
rect 9160 7923 9204 7929
rect 9274 7949 9318 7965
rect 9274 7929 9283 7949
rect 9303 7929 9318 7949
rect 9274 7923 9318 7929
rect 9368 7953 9417 7965
rect 9368 7933 9386 7953
rect 9406 7933 9417 7953
rect 9368 7923 9417 7933
rect 9482 7949 9526 7965
rect 9482 7929 9491 7949
rect 9511 7929 9526 7949
rect 9482 7923 9526 7929
rect 9576 7953 9625 7965
rect 9576 7933 9594 7953
rect 9614 7933 9625 7953
rect 9576 7923 9625 7933
rect 9695 7949 9739 7965
rect 9695 7929 9704 7949
rect 9724 7929 9739 7949
rect 9695 7923 9739 7929
rect 9789 7953 9838 7965
rect 9789 7933 9807 7953
rect 9827 7933 9838 7953
rect 9789 7923 9838 7933
rect 1499 7806 1517 7826
rect 1537 7806 1548 7826
rect 1499 7794 1548 7806
rect 3266 7821 3315 7831
rect 3266 7801 3277 7821
rect 3297 7801 3315 7821
rect 3266 7789 3315 7801
rect 3365 7825 3409 7831
rect 3365 7805 3380 7825
rect 3400 7805 3409 7825
rect 3365 7789 3409 7805
rect 3479 7821 3528 7831
rect 3479 7801 3490 7821
rect 3510 7801 3528 7821
rect 3479 7789 3528 7801
rect 3578 7825 3622 7831
rect 3578 7805 3593 7825
rect 3613 7805 3622 7825
rect 3578 7789 3622 7805
rect 3687 7821 3736 7831
rect 3687 7801 3698 7821
rect 3718 7801 3736 7821
rect 3687 7789 3736 7801
rect 3786 7825 3830 7831
rect 3786 7805 3801 7825
rect 3821 7805 3830 7825
rect 3786 7789 3830 7805
rect 3900 7825 3944 7831
rect 3900 7805 3909 7825
rect 3929 7805 3944 7825
rect 3900 7789 3944 7805
rect 3994 7821 4043 7831
rect 3994 7801 4012 7821
rect 4032 7801 4043 7821
rect 3994 7789 4043 7801
rect 6566 7190 6615 7202
rect 6566 7170 6577 7190
rect 6597 7170 6615 7190
rect 6566 7160 6615 7170
rect 6665 7186 6709 7202
rect 6665 7166 6680 7186
rect 6700 7166 6709 7186
rect 6665 7160 6709 7166
rect 6779 7186 6823 7202
rect 6779 7166 6788 7186
rect 6808 7166 6823 7186
rect 6779 7160 6823 7166
rect 6873 7190 6922 7202
rect 6873 7170 6891 7190
rect 6911 7170 6922 7190
rect 6873 7160 6922 7170
rect 6987 7186 7031 7202
rect 6987 7166 6996 7186
rect 7016 7166 7031 7186
rect 6987 7160 7031 7166
rect 7081 7190 7130 7202
rect 7081 7170 7099 7190
rect 7119 7170 7130 7190
rect 7081 7160 7130 7170
rect 7200 7186 7244 7202
rect 7200 7166 7209 7186
rect 7229 7166 7244 7186
rect 7200 7160 7244 7166
rect 7294 7190 7343 7202
rect 7294 7170 7312 7190
rect 7332 7170 7343 7190
rect 7294 7160 7343 7170
rect 9061 7185 9110 7197
rect 9061 7165 9072 7185
rect 9092 7165 9110 7185
rect 771 7058 820 7068
rect 771 7038 782 7058
rect 802 7038 820 7058
rect 771 7026 820 7038
rect 870 7062 914 7068
rect 870 7042 885 7062
rect 905 7042 914 7062
rect 870 7026 914 7042
rect 984 7058 1033 7068
rect 984 7038 995 7058
rect 1015 7038 1033 7058
rect 984 7026 1033 7038
rect 1083 7062 1127 7068
rect 1083 7042 1098 7062
rect 1118 7042 1127 7062
rect 1083 7026 1127 7042
rect 1192 7058 1241 7068
rect 1192 7038 1203 7058
rect 1223 7038 1241 7058
rect 1192 7026 1241 7038
rect 1291 7062 1335 7068
rect 1291 7042 1306 7062
rect 1326 7042 1335 7062
rect 1291 7026 1335 7042
rect 1405 7062 1449 7068
rect 1405 7042 1414 7062
rect 1434 7042 1449 7062
rect 1405 7026 1449 7042
rect 1499 7058 1548 7068
rect 9061 7155 9110 7165
rect 9160 7181 9204 7197
rect 9160 7161 9175 7181
rect 9195 7161 9204 7181
rect 9160 7155 9204 7161
rect 9274 7181 9318 7197
rect 9274 7161 9283 7181
rect 9303 7161 9318 7181
rect 9274 7155 9318 7161
rect 9368 7185 9417 7197
rect 9368 7165 9386 7185
rect 9406 7165 9417 7185
rect 9368 7155 9417 7165
rect 9482 7181 9526 7197
rect 9482 7161 9491 7181
rect 9511 7161 9526 7181
rect 9482 7155 9526 7161
rect 9576 7185 9625 7197
rect 9576 7165 9594 7185
rect 9614 7165 9625 7185
rect 9576 7155 9625 7165
rect 9695 7181 9739 7197
rect 9695 7161 9704 7181
rect 9724 7161 9739 7181
rect 9695 7155 9739 7161
rect 9789 7185 9838 7197
rect 9789 7165 9807 7185
rect 9827 7165 9838 7185
rect 9789 7155 9838 7165
rect 1499 7038 1517 7058
rect 1537 7038 1548 7058
rect 1499 7026 1548 7038
rect 1819 7054 1868 7064
rect 1819 7034 1830 7054
rect 1850 7034 1868 7054
rect 1819 7022 1868 7034
rect 1918 7058 1962 7064
rect 1918 7038 1933 7058
rect 1953 7038 1962 7058
rect 1918 7022 1962 7038
rect 2032 7054 2081 7064
rect 2032 7034 2043 7054
rect 2063 7034 2081 7054
rect 2032 7022 2081 7034
rect 2131 7058 2175 7064
rect 2131 7038 2146 7058
rect 2166 7038 2175 7058
rect 2131 7022 2175 7038
rect 2240 7054 2289 7064
rect 2240 7034 2251 7054
rect 2271 7034 2289 7054
rect 2240 7022 2289 7034
rect 2339 7058 2383 7064
rect 2339 7038 2354 7058
rect 2374 7038 2383 7058
rect 2339 7022 2383 7038
rect 2453 7058 2497 7064
rect 2453 7038 2462 7058
rect 2482 7038 2497 7058
rect 2453 7022 2497 7038
rect 2547 7054 2596 7064
rect 2547 7034 2565 7054
rect 2585 7034 2596 7054
rect 2547 7022 2596 7034
rect 8013 6510 8062 6522
rect 8013 6490 8024 6510
rect 8044 6490 8062 6510
rect 8013 6480 8062 6490
rect 8112 6506 8156 6522
rect 8112 6486 8127 6506
rect 8147 6486 8156 6506
rect 8112 6480 8156 6486
rect 8226 6506 8270 6522
rect 8226 6486 8235 6506
rect 8255 6486 8270 6506
rect 8226 6480 8270 6486
rect 8320 6510 8369 6522
rect 8320 6490 8338 6510
rect 8358 6490 8369 6510
rect 8320 6480 8369 6490
rect 8434 6506 8478 6522
rect 8434 6486 8443 6506
rect 8463 6486 8478 6506
rect 8434 6480 8478 6486
rect 8528 6510 8577 6522
rect 8528 6490 8546 6510
rect 8566 6490 8577 6510
rect 8528 6480 8577 6490
rect 8647 6506 8691 6522
rect 8647 6486 8656 6506
rect 8676 6486 8691 6506
rect 8647 6480 8691 6486
rect 8741 6510 8790 6522
rect 8741 6490 8759 6510
rect 8779 6490 8790 6510
rect 8741 6480 8790 6490
rect 9061 6506 9110 6518
rect 9061 6486 9072 6506
rect 9092 6486 9110 6506
rect 771 6379 820 6389
rect 771 6359 782 6379
rect 802 6359 820 6379
rect 771 6347 820 6359
rect 870 6383 914 6389
rect 870 6363 885 6383
rect 905 6363 914 6383
rect 870 6347 914 6363
rect 984 6379 1033 6389
rect 984 6359 995 6379
rect 1015 6359 1033 6379
rect 984 6347 1033 6359
rect 1083 6383 1127 6389
rect 1083 6363 1098 6383
rect 1118 6363 1127 6383
rect 1083 6347 1127 6363
rect 1192 6379 1241 6389
rect 1192 6359 1203 6379
rect 1223 6359 1241 6379
rect 1192 6347 1241 6359
rect 1291 6383 1335 6389
rect 1291 6363 1306 6383
rect 1326 6363 1335 6383
rect 1291 6347 1335 6363
rect 1405 6383 1449 6389
rect 1405 6363 1414 6383
rect 1434 6363 1449 6383
rect 1405 6347 1449 6363
rect 1499 6379 1548 6389
rect 9061 6476 9110 6486
rect 9160 6502 9204 6518
rect 9160 6482 9175 6502
rect 9195 6482 9204 6502
rect 9160 6476 9204 6482
rect 9274 6502 9318 6518
rect 9274 6482 9283 6502
rect 9303 6482 9318 6502
rect 9274 6476 9318 6482
rect 9368 6506 9417 6518
rect 9368 6486 9386 6506
rect 9406 6486 9417 6506
rect 9368 6476 9417 6486
rect 9482 6502 9526 6518
rect 9482 6482 9491 6502
rect 9511 6482 9526 6502
rect 9482 6476 9526 6482
rect 9576 6506 9625 6518
rect 9576 6486 9594 6506
rect 9614 6486 9625 6506
rect 9576 6476 9625 6486
rect 9695 6502 9739 6518
rect 9695 6482 9704 6502
rect 9724 6482 9739 6502
rect 9695 6476 9739 6482
rect 9789 6506 9838 6518
rect 9789 6486 9807 6506
rect 9827 6486 9838 6506
rect 9789 6476 9838 6486
rect 1499 6359 1517 6379
rect 1537 6359 1548 6379
rect 1499 6347 1548 6359
rect 4374 6370 4423 6380
rect 4374 6350 4385 6370
rect 4405 6350 4423 6370
rect 4374 6338 4423 6350
rect 4473 6374 4517 6380
rect 4473 6354 4488 6374
rect 4508 6354 4517 6374
rect 4473 6338 4517 6354
rect 4587 6370 4636 6380
rect 4587 6350 4598 6370
rect 4618 6350 4636 6370
rect 4587 6338 4636 6350
rect 4686 6374 4730 6380
rect 4686 6354 4701 6374
rect 4721 6354 4730 6374
rect 4686 6338 4730 6354
rect 4795 6370 4844 6380
rect 4795 6350 4806 6370
rect 4826 6350 4844 6370
rect 4795 6338 4844 6350
rect 4894 6374 4938 6380
rect 4894 6354 4909 6374
rect 4929 6354 4938 6374
rect 4894 6338 4938 6354
rect 5008 6374 5052 6380
rect 5008 6354 5017 6374
rect 5037 6354 5052 6374
rect 5008 6338 5052 6354
rect 5102 6370 5151 6380
rect 5102 6350 5120 6370
rect 5140 6350 5151 6370
rect 5102 6338 5151 6350
rect 5455 5600 5504 5612
rect 5455 5580 5466 5600
rect 5486 5580 5504 5600
rect 5455 5570 5504 5580
rect 5554 5596 5598 5612
rect 5554 5576 5569 5596
rect 5589 5576 5598 5596
rect 5554 5570 5598 5576
rect 5668 5596 5712 5612
rect 5668 5576 5677 5596
rect 5697 5576 5712 5596
rect 5668 5570 5712 5576
rect 5762 5600 5811 5612
rect 5762 5580 5780 5600
rect 5800 5580 5811 5600
rect 5762 5570 5811 5580
rect 5876 5596 5920 5612
rect 5876 5576 5885 5596
rect 5905 5576 5920 5596
rect 5876 5570 5920 5576
rect 5970 5600 6019 5612
rect 5970 5580 5988 5600
rect 6008 5580 6019 5600
rect 5970 5570 6019 5580
rect 6089 5596 6133 5612
rect 6089 5576 6098 5596
rect 6118 5576 6133 5596
rect 6089 5570 6133 5576
rect 6183 5600 6232 5612
rect 6183 5580 6201 5600
rect 6221 5580 6232 5600
rect 6183 5570 6232 5580
rect 9058 5591 9107 5603
rect 9058 5571 9069 5591
rect 9089 5571 9107 5591
rect 768 5464 817 5474
rect 768 5444 779 5464
rect 799 5444 817 5464
rect 768 5432 817 5444
rect 867 5468 911 5474
rect 867 5448 882 5468
rect 902 5448 911 5468
rect 867 5432 911 5448
rect 981 5464 1030 5474
rect 981 5444 992 5464
rect 1012 5444 1030 5464
rect 981 5432 1030 5444
rect 1080 5468 1124 5474
rect 1080 5448 1095 5468
rect 1115 5448 1124 5468
rect 1080 5432 1124 5448
rect 1189 5464 1238 5474
rect 1189 5444 1200 5464
rect 1220 5444 1238 5464
rect 1189 5432 1238 5444
rect 1288 5468 1332 5474
rect 1288 5448 1303 5468
rect 1323 5448 1332 5468
rect 1288 5432 1332 5448
rect 1402 5468 1446 5474
rect 1402 5448 1411 5468
rect 1431 5448 1446 5468
rect 1402 5432 1446 5448
rect 1496 5464 1545 5474
rect 9058 5561 9107 5571
rect 9157 5587 9201 5603
rect 9157 5567 9172 5587
rect 9192 5567 9201 5587
rect 9157 5561 9201 5567
rect 9271 5587 9315 5603
rect 9271 5567 9280 5587
rect 9300 5567 9315 5587
rect 9271 5561 9315 5567
rect 9365 5591 9414 5603
rect 9365 5571 9383 5591
rect 9403 5571 9414 5591
rect 9365 5561 9414 5571
rect 9479 5587 9523 5603
rect 9479 5567 9488 5587
rect 9508 5567 9523 5587
rect 9479 5561 9523 5567
rect 9573 5591 9622 5603
rect 9573 5571 9591 5591
rect 9611 5571 9622 5591
rect 9573 5561 9622 5571
rect 9692 5587 9736 5603
rect 9692 5567 9701 5587
rect 9721 5567 9736 5587
rect 9692 5561 9736 5567
rect 9786 5591 9835 5603
rect 9786 5571 9804 5591
rect 9824 5571 9835 5591
rect 9786 5561 9835 5571
rect 1496 5444 1514 5464
rect 1534 5444 1545 5464
rect 1496 5432 1545 5444
rect 1816 5460 1865 5470
rect 1816 5440 1827 5460
rect 1847 5440 1865 5460
rect 1816 5428 1865 5440
rect 1915 5464 1959 5470
rect 1915 5444 1930 5464
rect 1950 5444 1959 5464
rect 1915 5428 1959 5444
rect 2029 5460 2078 5470
rect 2029 5440 2040 5460
rect 2060 5440 2078 5460
rect 2029 5428 2078 5440
rect 2128 5464 2172 5470
rect 2128 5444 2143 5464
rect 2163 5444 2172 5464
rect 2128 5428 2172 5444
rect 2237 5460 2286 5470
rect 2237 5440 2248 5460
rect 2268 5440 2286 5460
rect 2237 5428 2286 5440
rect 2336 5464 2380 5470
rect 2336 5444 2351 5464
rect 2371 5444 2380 5464
rect 2336 5428 2380 5444
rect 2450 5464 2494 5470
rect 2450 5444 2459 5464
rect 2479 5444 2494 5464
rect 2450 5428 2494 5444
rect 2544 5460 2593 5470
rect 2544 5440 2562 5460
rect 2582 5440 2593 5460
rect 2544 5428 2593 5440
rect 8010 4916 8059 4928
rect 8010 4896 8021 4916
rect 8041 4896 8059 4916
rect 8010 4886 8059 4896
rect 8109 4912 8153 4928
rect 8109 4892 8124 4912
rect 8144 4892 8153 4912
rect 8109 4886 8153 4892
rect 8223 4912 8267 4928
rect 8223 4892 8232 4912
rect 8252 4892 8267 4912
rect 8223 4886 8267 4892
rect 8317 4916 8366 4928
rect 8317 4896 8335 4916
rect 8355 4896 8366 4916
rect 8317 4886 8366 4896
rect 8431 4912 8475 4928
rect 8431 4892 8440 4912
rect 8460 4892 8475 4912
rect 8431 4886 8475 4892
rect 8525 4916 8574 4928
rect 8525 4896 8543 4916
rect 8563 4896 8574 4916
rect 8525 4886 8574 4896
rect 8644 4912 8688 4928
rect 8644 4892 8653 4912
rect 8673 4892 8688 4912
rect 8644 4886 8688 4892
rect 8738 4916 8787 4928
rect 8738 4896 8756 4916
rect 8776 4896 8787 4916
rect 8738 4886 8787 4896
rect 9058 4912 9107 4924
rect 9058 4892 9069 4912
rect 9089 4892 9107 4912
rect 768 4785 817 4795
rect 768 4765 779 4785
rect 799 4765 817 4785
rect 768 4753 817 4765
rect 867 4789 911 4795
rect 867 4769 882 4789
rect 902 4769 911 4789
rect 867 4753 911 4769
rect 981 4785 1030 4795
rect 981 4765 992 4785
rect 1012 4765 1030 4785
rect 981 4753 1030 4765
rect 1080 4789 1124 4795
rect 1080 4769 1095 4789
rect 1115 4769 1124 4789
rect 1080 4753 1124 4769
rect 1189 4785 1238 4795
rect 1189 4765 1200 4785
rect 1220 4765 1238 4785
rect 1189 4753 1238 4765
rect 1288 4789 1332 4795
rect 1288 4769 1303 4789
rect 1323 4769 1332 4789
rect 1288 4753 1332 4769
rect 1402 4789 1446 4795
rect 1402 4769 1411 4789
rect 1431 4769 1446 4789
rect 1402 4753 1446 4769
rect 1496 4785 1545 4795
rect 9058 4882 9107 4892
rect 9157 4908 9201 4924
rect 9157 4888 9172 4908
rect 9192 4888 9201 4908
rect 9157 4882 9201 4888
rect 9271 4908 9315 4924
rect 9271 4888 9280 4908
rect 9300 4888 9315 4908
rect 9271 4882 9315 4888
rect 9365 4912 9414 4924
rect 9365 4892 9383 4912
rect 9403 4892 9414 4912
rect 9365 4882 9414 4892
rect 9479 4908 9523 4924
rect 9479 4888 9488 4908
rect 9508 4888 9523 4908
rect 9479 4882 9523 4888
rect 9573 4912 9622 4924
rect 9573 4892 9591 4912
rect 9611 4892 9622 4912
rect 9573 4882 9622 4892
rect 9692 4908 9736 4924
rect 9692 4888 9701 4908
rect 9721 4888 9736 4908
rect 9692 4882 9736 4888
rect 9786 4912 9835 4924
rect 9786 4892 9804 4912
rect 9824 4892 9835 4912
rect 9786 4882 9835 4892
rect 1496 4765 1514 4785
rect 1534 4765 1545 4785
rect 1496 4753 1545 4765
rect 3263 4780 3312 4790
rect 3263 4760 3274 4780
rect 3294 4760 3312 4780
rect 3263 4748 3312 4760
rect 3362 4784 3406 4790
rect 3362 4764 3377 4784
rect 3397 4764 3406 4784
rect 3362 4748 3406 4764
rect 3476 4780 3525 4790
rect 3476 4760 3487 4780
rect 3507 4760 3525 4780
rect 3476 4748 3525 4760
rect 3575 4784 3619 4790
rect 3575 4764 3590 4784
rect 3610 4764 3619 4784
rect 3575 4748 3619 4764
rect 3684 4780 3733 4790
rect 3684 4760 3695 4780
rect 3715 4760 3733 4780
rect 3684 4748 3733 4760
rect 3783 4784 3827 4790
rect 3783 4764 3798 4784
rect 3818 4764 3827 4784
rect 3783 4748 3827 4764
rect 3897 4784 3941 4790
rect 3897 4764 3906 4784
rect 3926 4764 3941 4784
rect 3897 4748 3941 4764
rect 3991 4780 4040 4790
rect 3991 4760 4009 4780
rect 4029 4760 4040 4780
rect 3991 4748 4040 4760
rect 6563 4149 6612 4161
rect 6563 4129 6574 4149
rect 6594 4129 6612 4149
rect 6563 4119 6612 4129
rect 6662 4145 6706 4161
rect 6662 4125 6677 4145
rect 6697 4125 6706 4145
rect 6662 4119 6706 4125
rect 6776 4145 6820 4161
rect 6776 4125 6785 4145
rect 6805 4125 6820 4145
rect 6776 4119 6820 4125
rect 6870 4149 6919 4161
rect 6870 4129 6888 4149
rect 6908 4129 6919 4149
rect 6870 4119 6919 4129
rect 6984 4145 7028 4161
rect 6984 4125 6993 4145
rect 7013 4125 7028 4145
rect 6984 4119 7028 4125
rect 7078 4149 7127 4161
rect 7078 4129 7096 4149
rect 7116 4129 7127 4149
rect 7078 4119 7127 4129
rect 7197 4145 7241 4161
rect 7197 4125 7206 4145
rect 7226 4125 7241 4145
rect 7197 4119 7241 4125
rect 7291 4149 7340 4161
rect 7291 4129 7309 4149
rect 7329 4129 7340 4149
rect 7291 4119 7340 4129
rect 9058 4144 9107 4156
rect 9058 4124 9069 4144
rect 9089 4124 9107 4144
rect 768 4017 817 4027
rect 768 3997 779 4017
rect 799 3997 817 4017
rect 768 3985 817 3997
rect 867 4021 911 4027
rect 867 4001 882 4021
rect 902 4001 911 4021
rect 867 3985 911 4001
rect 981 4017 1030 4027
rect 981 3997 992 4017
rect 1012 3997 1030 4017
rect 981 3985 1030 3997
rect 1080 4021 1124 4027
rect 1080 4001 1095 4021
rect 1115 4001 1124 4021
rect 1080 3985 1124 4001
rect 1189 4017 1238 4027
rect 1189 3997 1200 4017
rect 1220 3997 1238 4017
rect 1189 3985 1238 3997
rect 1288 4021 1332 4027
rect 1288 4001 1303 4021
rect 1323 4001 1332 4021
rect 1288 3985 1332 4001
rect 1402 4021 1446 4027
rect 1402 4001 1411 4021
rect 1431 4001 1446 4021
rect 1402 3985 1446 4001
rect 1496 4017 1545 4027
rect 9058 4114 9107 4124
rect 9157 4140 9201 4156
rect 9157 4120 9172 4140
rect 9192 4120 9201 4140
rect 9157 4114 9201 4120
rect 9271 4140 9315 4156
rect 9271 4120 9280 4140
rect 9300 4120 9315 4140
rect 9271 4114 9315 4120
rect 9365 4144 9414 4156
rect 9365 4124 9383 4144
rect 9403 4124 9414 4144
rect 9365 4114 9414 4124
rect 9479 4140 9523 4156
rect 9479 4120 9488 4140
rect 9508 4120 9523 4140
rect 9479 4114 9523 4120
rect 9573 4144 9622 4156
rect 9573 4124 9591 4144
rect 9611 4124 9622 4144
rect 9573 4114 9622 4124
rect 9692 4140 9736 4156
rect 9692 4120 9701 4140
rect 9721 4120 9736 4140
rect 9692 4114 9736 4120
rect 9786 4144 9835 4156
rect 9786 4124 9804 4144
rect 9824 4124 9835 4144
rect 9786 4114 9835 4124
rect 1496 3997 1514 4017
rect 1534 3997 1545 4017
rect 1496 3985 1545 3997
rect 1816 4013 1865 4023
rect 1816 3993 1827 4013
rect 1847 3993 1865 4013
rect 1816 3981 1865 3993
rect 1915 4017 1959 4023
rect 1915 3997 1930 4017
rect 1950 3997 1959 4017
rect 1915 3981 1959 3997
rect 2029 4013 2078 4023
rect 2029 3993 2040 4013
rect 2060 3993 2078 4013
rect 2029 3981 2078 3993
rect 2128 4017 2172 4023
rect 2128 3997 2143 4017
rect 2163 3997 2172 4017
rect 2128 3981 2172 3997
rect 2237 4013 2286 4023
rect 2237 3993 2248 4013
rect 2268 3993 2286 4013
rect 2237 3981 2286 3993
rect 2336 4017 2380 4023
rect 2336 3997 2351 4017
rect 2371 3997 2380 4017
rect 2336 3981 2380 3997
rect 2450 4017 2494 4023
rect 2450 3997 2459 4017
rect 2479 3997 2494 4017
rect 2450 3981 2494 3997
rect 2544 4013 2593 4023
rect 2544 3993 2562 4013
rect 2582 3993 2593 4013
rect 2544 3981 2593 3993
rect 8010 3469 8059 3481
rect 8010 3449 8021 3469
rect 8041 3449 8059 3469
rect 8010 3439 8059 3449
rect 8109 3465 8153 3481
rect 8109 3445 8124 3465
rect 8144 3445 8153 3465
rect 8109 3439 8153 3445
rect 8223 3465 8267 3481
rect 8223 3445 8232 3465
rect 8252 3445 8267 3465
rect 8223 3439 8267 3445
rect 8317 3469 8366 3481
rect 8317 3449 8335 3469
rect 8355 3449 8366 3469
rect 8317 3439 8366 3449
rect 8431 3465 8475 3481
rect 8431 3445 8440 3465
rect 8460 3445 8475 3465
rect 8431 3439 8475 3445
rect 8525 3469 8574 3481
rect 8525 3449 8543 3469
rect 8563 3449 8574 3469
rect 8525 3439 8574 3449
rect 8644 3465 8688 3481
rect 8644 3445 8653 3465
rect 8673 3445 8688 3465
rect 8644 3439 8688 3445
rect 8738 3469 8787 3481
rect 8738 3449 8756 3469
rect 8776 3449 8787 3469
rect 8738 3439 8787 3449
rect 9058 3465 9107 3477
rect 9058 3445 9069 3465
rect 9089 3445 9107 3465
rect 768 3338 817 3348
rect 768 3318 779 3338
rect 799 3318 817 3338
rect 768 3306 817 3318
rect 867 3342 911 3348
rect 867 3322 882 3342
rect 902 3322 911 3342
rect 867 3306 911 3322
rect 981 3338 1030 3348
rect 981 3318 992 3338
rect 1012 3318 1030 3338
rect 981 3306 1030 3318
rect 1080 3342 1124 3348
rect 1080 3322 1095 3342
rect 1115 3322 1124 3342
rect 1080 3306 1124 3322
rect 1189 3338 1238 3348
rect 1189 3318 1200 3338
rect 1220 3318 1238 3338
rect 1189 3306 1238 3318
rect 1288 3342 1332 3348
rect 1288 3322 1303 3342
rect 1323 3322 1332 3342
rect 1288 3306 1332 3322
rect 1402 3342 1446 3348
rect 1402 3322 1411 3342
rect 1431 3322 1446 3342
rect 1402 3306 1446 3322
rect 1496 3338 1545 3348
rect 9058 3435 9107 3445
rect 9157 3461 9201 3477
rect 9157 3441 9172 3461
rect 9192 3441 9201 3461
rect 9157 3435 9201 3441
rect 9271 3461 9315 3477
rect 9271 3441 9280 3461
rect 9300 3441 9315 3461
rect 9271 3435 9315 3441
rect 9365 3465 9414 3477
rect 9365 3445 9383 3465
rect 9403 3445 9414 3465
rect 9365 3435 9414 3445
rect 9479 3461 9523 3477
rect 9479 3441 9488 3461
rect 9508 3441 9523 3461
rect 9479 3435 9523 3441
rect 9573 3465 9622 3477
rect 9573 3445 9591 3465
rect 9611 3445 9622 3465
rect 9573 3435 9622 3445
rect 9692 3461 9736 3477
rect 9692 3441 9701 3461
rect 9721 3441 9736 3461
rect 9692 3435 9736 3441
rect 9786 3465 9835 3477
rect 9786 3445 9804 3465
rect 9824 3445 9835 3465
rect 9786 3435 9835 3445
rect 1496 3318 1514 3338
rect 1534 3318 1545 3338
rect 1496 3306 1545 3318
rect 3306 3335 3355 3345
rect 3306 3315 3317 3335
rect 3337 3315 3355 3335
rect 3306 3303 3355 3315
rect 3405 3339 3449 3345
rect 3405 3319 3420 3339
rect 3440 3319 3449 3339
rect 3405 3303 3449 3319
rect 3519 3335 3568 3345
rect 3519 3315 3530 3335
rect 3550 3315 3568 3335
rect 3519 3303 3568 3315
rect 3618 3339 3662 3345
rect 3618 3319 3633 3339
rect 3653 3319 3662 3339
rect 3618 3303 3662 3319
rect 3727 3335 3776 3345
rect 3727 3315 3738 3335
rect 3758 3315 3776 3335
rect 3727 3303 3776 3315
rect 3826 3339 3870 3345
rect 3826 3319 3841 3339
rect 3861 3319 3870 3339
rect 3826 3303 3870 3319
rect 3940 3339 3984 3345
rect 3940 3319 3949 3339
rect 3969 3319 3984 3339
rect 3940 3303 3984 3319
rect 4034 3335 4083 3345
rect 4034 3315 4052 3335
rect 4072 3315 4083 3335
rect 4034 3303 4083 3315
rect 6521 2627 6570 2639
rect 6521 2607 6532 2627
rect 6552 2607 6570 2627
rect 6521 2597 6570 2607
rect 6620 2623 6664 2639
rect 6620 2603 6635 2623
rect 6655 2603 6664 2623
rect 6620 2597 6664 2603
rect 6734 2623 6778 2639
rect 6734 2603 6743 2623
rect 6763 2603 6778 2623
rect 6734 2597 6778 2603
rect 6828 2627 6877 2639
rect 6828 2607 6846 2627
rect 6866 2607 6877 2627
rect 6828 2597 6877 2607
rect 6942 2623 6986 2639
rect 6942 2603 6951 2623
rect 6971 2603 6986 2623
rect 6942 2597 6986 2603
rect 7036 2627 7085 2639
rect 7036 2607 7054 2627
rect 7074 2607 7085 2627
rect 7036 2597 7085 2607
rect 7155 2623 7199 2639
rect 7155 2603 7164 2623
rect 7184 2603 7199 2623
rect 7155 2597 7199 2603
rect 7249 2627 7298 2639
rect 7249 2607 7267 2627
rect 7287 2607 7298 2627
rect 7249 2597 7298 2607
rect 9059 2624 9108 2636
rect 9059 2604 9070 2624
rect 9090 2604 9108 2624
rect 769 2497 818 2507
rect 769 2477 780 2497
rect 800 2477 818 2497
rect 769 2465 818 2477
rect 868 2501 912 2507
rect 868 2481 883 2501
rect 903 2481 912 2501
rect 868 2465 912 2481
rect 982 2497 1031 2507
rect 982 2477 993 2497
rect 1013 2477 1031 2497
rect 982 2465 1031 2477
rect 1081 2501 1125 2507
rect 1081 2481 1096 2501
rect 1116 2481 1125 2501
rect 1081 2465 1125 2481
rect 1190 2497 1239 2507
rect 1190 2477 1201 2497
rect 1221 2477 1239 2497
rect 1190 2465 1239 2477
rect 1289 2501 1333 2507
rect 1289 2481 1304 2501
rect 1324 2481 1333 2501
rect 1289 2465 1333 2481
rect 1403 2501 1447 2507
rect 1403 2481 1412 2501
rect 1432 2481 1447 2501
rect 1403 2465 1447 2481
rect 1497 2497 1546 2507
rect 9059 2594 9108 2604
rect 9158 2620 9202 2636
rect 9158 2600 9173 2620
rect 9193 2600 9202 2620
rect 9158 2594 9202 2600
rect 9272 2620 9316 2636
rect 9272 2600 9281 2620
rect 9301 2600 9316 2620
rect 9272 2594 9316 2600
rect 9366 2624 9415 2636
rect 9366 2604 9384 2624
rect 9404 2604 9415 2624
rect 9366 2594 9415 2604
rect 9480 2620 9524 2636
rect 9480 2600 9489 2620
rect 9509 2600 9524 2620
rect 9480 2594 9524 2600
rect 9574 2624 9623 2636
rect 9574 2604 9592 2624
rect 9612 2604 9623 2624
rect 9574 2594 9623 2604
rect 9693 2620 9737 2636
rect 9693 2600 9702 2620
rect 9722 2600 9737 2620
rect 9693 2594 9737 2600
rect 9787 2624 9836 2636
rect 9787 2604 9805 2624
rect 9825 2604 9836 2624
rect 9787 2594 9836 2604
rect 1497 2477 1515 2497
rect 1535 2477 1546 2497
rect 1497 2465 1546 2477
rect 1817 2493 1866 2503
rect 1817 2473 1828 2493
rect 1848 2473 1866 2493
rect 1817 2461 1866 2473
rect 1916 2497 1960 2503
rect 1916 2477 1931 2497
rect 1951 2477 1960 2497
rect 1916 2461 1960 2477
rect 2030 2493 2079 2503
rect 2030 2473 2041 2493
rect 2061 2473 2079 2493
rect 2030 2461 2079 2473
rect 2129 2497 2173 2503
rect 2129 2477 2144 2497
rect 2164 2477 2173 2497
rect 2129 2461 2173 2477
rect 2238 2493 2287 2503
rect 2238 2473 2249 2493
rect 2269 2473 2287 2493
rect 2238 2461 2287 2473
rect 2337 2497 2381 2503
rect 2337 2477 2352 2497
rect 2372 2477 2381 2497
rect 2337 2461 2381 2477
rect 2451 2497 2495 2503
rect 2451 2477 2460 2497
rect 2480 2477 2495 2497
rect 2451 2461 2495 2477
rect 2545 2493 2594 2503
rect 2545 2473 2563 2493
rect 2583 2473 2594 2493
rect 2545 2461 2594 2473
rect 4719 2499 4768 2509
rect 4719 2479 4730 2499
rect 4750 2479 4768 2499
rect 4719 2467 4768 2479
rect 4818 2503 4862 2509
rect 4818 2483 4833 2503
rect 4853 2483 4862 2503
rect 4818 2467 4862 2483
rect 4932 2499 4981 2509
rect 4932 2479 4943 2499
rect 4963 2479 4981 2499
rect 4932 2467 4981 2479
rect 5031 2503 5075 2509
rect 5031 2483 5046 2503
rect 5066 2483 5075 2503
rect 5031 2467 5075 2483
rect 5140 2499 5189 2509
rect 5140 2479 5151 2499
rect 5171 2479 5189 2499
rect 5140 2467 5189 2479
rect 5239 2503 5283 2509
rect 5239 2483 5254 2503
rect 5274 2483 5283 2503
rect 5239 2467 5283 2483
rect 5353 2503 5397 2509
rect 5353 2483 5362 2503
rect 5382 2483 5397 2503
rect 5353 2467 5397 2483
rect 5447 2499 5496 2509
rect 5447 2479 5465 2499
rect 5485 2479 5496 2499
rect 5447 2467 5496 2479
rect 8011 1949 8060 1961
rect 8011 1929 8022 1949
rect 8042 1929 8060 1949
rect 8011 1919 8060 1929
rect 8110 1945 8154 1961
rect 8110 1925 8125 1945
rect 8145 1925 8154 1945
rect 8110 1919 8154 1925
rect 8224 1945 8268 1961
rect 8224 1925 8233 1945
rect 8253 1925 8268 1945
rect 8224 1919 8268 1925
rect 8318 1949 8367 1961
rect 8318 1929 8336 1949
rect 8356 1929 8367 1949
rect 8318 1919 8367 1929
rect 8432 1945 8476 1961
rect 8432 1925 8441 1945
rect 8461 1925 8476 1945
rect 8432 1919 8476 1925
rect 8526 1949 8575 1961
rect 8526 1929 8544 1949
rect 8564 1929 8575 1949
rect 8526 1919 8575 1929
rect 8645 1945 8689 1961
rect 8645 1925 8654 1945
rect 8674 1925 8689 1945
rect 8645 1919 8689 1925
rect 8739 1949 8788 1961
rect 8739 1929 8757 1949
rect 8777 1929 8788 1949
rect 8739 1919 8788 1929
rect 9059 1945 9108 1957
rect 9059 1925 9070 1945
rect 9090 1925 9108 1945
rect 769 1818 818 1828
rect 769 1798 780 1818
rect 800 1798 818 1818
rect 769 1786 818 1798
rect 868 1822 912 1828
rect 868 1802 883 1822
rect 903 1802 912 1822
rect 868 1786 912 1802
rect 982 1818 1031 1828
rect 982 1798 993 1818
rect 1013 1798 1031 1818
rect 982 1786 1031 1798
rect 1081 1822 1125 1828
rect 1081 1802 1096 1822
rect 1116 1802 1125 1822
rect 1081 1786 1125 1802
rect 1190 1818 1239 1828
rect 1190 1798 1201 1818
rect 1221 1798 1239 1818
rect 1190 1786 1239 1798
rect 1289 1822 1333 1828
rect 1289 1802 1304 1822
rect 1324 1802 1333 1822
rect 1289 1786 1333 1802
rect 1403 1822 1447 1828
rect 1403 1802 1412 1822
rect 1432 1802 1447 1822
rect 1403 1786 1447 1802
rect 1497 1818 1546 1828
rect 9059 1915 9108 1925
rect 9158 1941 9202 1957
rect 9158 1921 9173 1941
rect 9193 1921 9202 1941
rect 9158 1915 9202 1921
rect 9272 1941 9316 1957
rect 9272 1921 9281 1941
rect 9301 1921 9316 1941
rect 9272 1915 9316 1921
rect 9366 1945 9415 1957
rect 9366 1925 9384 1945
rect 9404 1925 9415 1945
rect 9366 1915 9415 1925
rect 9480 1941 9524 1957
rect 9480 1921 9489 1941
rect 9509 1921 9524 1941
rect 9480 1915 9524 1921
rect 9574 1945 9623 1957
rect 9574 1925 9592 1945
rect 9612 1925 9623 1945
rect 9574 1915 9623 1925
rect 9693 1941 9737 1957
rect 9693 1921 9702 1941
rect 9722 1921 9737 1941
rect 9693 1915 9737 1921
rect 9787 1945 9836 1957
rect 9787 1925 9805 1945
rect 9825 1925 9836 1945
rect 9787 1915 9836 1925
rect 1497 1798 1515 1818
rect 1535 1798 1546 1818
rect 1497 1786 1546 1798
rect 3264 1813 3313 1823
rect 3264 1793 3275 1813
rect 3295 1793 3313 1813
rect 3264 1781 3313 1793
rect 3363 1817 3407 1823
rect 3363 1797 3378 1817
rect 3398 1797 3407 1817
rect 3363 1781 3407 1797
rect 3477 1813 3526 1823
rect 3477 1793 3488 1813
rect 3508 1793 3526 1813
rect 3477 1781 3526 1793
rect 3576 1817 3620 1823
rect 3576 1797 3591 1817
rect 3611 1797 3620 1817
rect 3576 1781 3620 1797
rect 3685 1813 3734 1823
rect 3685 1793 3696 1813
rect 3716 1793 3734 1813
rect 3685 1781 3734 1793
rect 3784 1817 3828 1823
rect 3784 1797 3799 1817
rect 3819 1797 3828 1817
rect 3784 1781 3828 1797
rect 3898 1817 3942 1823
rect 3898 1797 3907 1817
rect 3927 1797 3942 1817
rect 3898 1781 3942 1797
rect 3992 1813 4041 1823
rect 3992 1793 4010 1813
rect 4030 1793 4041 1813
rect 3992 1781 4041 1793
rect 6564 1182 6613 1194
rect 6564 1162 6575 1182
rect 6595 1162 6613 1182
rect 6564 1152 6613 1162
rect 6663 1178 6707 1194
rect 6663 1158 6678 1178
rect 6698 1158 6707 1178
rect 6663 1152 6707 1158
rect 6777 1178 6821 1194
rect 6777 1158 6786 1178
rect 6806 1158 6821 1178
rect 6777 1152 6821 1158
rect 6871 1182 6920 1194
rect 6871 1162 6889 1182
rect 6909 1162 6920 1182
rect 6871 1152 6920 1162
rect 6985 1178 7029 1194
rect 6985 1158 6994 1178
rect 7014 1158 7029 1178
rect 6985 1152 7029 1158
rect 7079 1182 7128 1194
rect 7079 1162 7097 1182
rect 7117 1162 7128 1182
rect 7079 1152 7128 1162
rect 7198 1178 7242 1194
rect 7198 1158 7207 1178
rect 7227 1158 7242 1178
rect 7198 1152 7242 1158
rect 7292 1182 7341 1194
rect 7292 1162 7310 1182
rect 7330 1162 7341 1182
rect 7292 1152 7341 1162
rect 9059 1177 9108 1189
rect 9059 1157 9070 1177
rect 9090 1157 9108 1177
rect 769 1050 818 1060
rect 769 1030 780 1050
rect 800 1030 818 1050
rect 769 1018 818 1030
rect 868 1054 912 1060
rect 868 1034 883 1054
rect 903 1034 912 1054
rect 868 1018 912 1034
rect 982 1050 1031 1060
rect 982 1030 993 1050
rect 1013 1030 1031 1050
rect 982 1018 1031 1030
rect 1081 1054 1125 1060
rect 1081 1034 1096 1054
rect 1116 1034 1125 1054
rect 1081 1018 1125 1034
rect 1190 1050 1239 1060
rect 1190 1030 1201 1050
rect 1221 1030 1239 1050
rect 1190 1018 1239 1030
rect 1289 1054 1333 1060
rect 1289 1034 1304 1054
rect 1324 1034 1333 1054
rect 1289 1018 1333 1034
rect 1403 1054 1447 1060
rect 1403 1034 1412 1054
rect 1432 1034 1447 1054
rect 1403 1018 1447 1034
rect 1497 1050 1546 1060
rect 9059 1147 9108 1157
rect 9158 1173 9202 1189
rect 9158 1153 9173 1173
rect 9193 1153 9202 1173
rect 9158 1147 9202 1153
rect 9272 1173 9316 1189
rect 9272 1153 9281 1173
rect 9301 1153 9316 1173
rect 9272 1147 9316 1153
rect 9366 1177 9415 1189
rect 9366 1157 9384 1177
rect 9404 1157 9415 1177
rect 9366 1147 9415 1157
rect 9480 1173 9524 1189
rect 9480 1153 9489 1173
rect 9509 1153 9524 1173
rect 9480 1147 9524 1153
rect 9574 1177 9623 1189
rect 9574 1157 9592 1177
rect 9612 1157 9623 1177
rect 9574 1147 9623 1157
rect 9693 1173 9737 1189
rect 9693 1153 9702 1173
rect 9722 1153 9737 1173
rect 9693 1147 9737 1153
rect 9787 1177 9836 1189
rect 9787 1157 9805 1177
rect 9825 1157 9836 1177
rect 9787 1147 9836 1157
rect 1497 1030 1515 1050
rect 1535 1030 1546 1050
rect 1497 1018 1546 1030
rect 1817 1046 1866 1056
rect 1817 1026 1828 1046
rect 1848 1026 1866 1046
rect 1817 1014 1866 1026
rect 1916 1050 1960 1056
rect 1916 1030 1931 1050
rect 1951 1030 1960 1050
rect 1916 1014 1960 1030
rect 2030 1046 2079 1056
rect 2030 1026 2041 1046
rect 2061 1026 2079 1046
rect 2030 1014 2079 1026
rect 2129 1050 2173 1056
rect 2129 1030 2144 1050
rect 2164 1030 2173 1050
rect 2129 1014 2173 1030
rect 2238 1046 2287 1056
rect 2238 1026 2249 1046
rect 2269 1026 2287 1046
rect 2238 1014 2287 1026
rect 2337 1050 2381 1056
rect 2337 1030 2352 1050
rect 2372 1030 2381 1050
rect 2337 1014 2381 1030
rect 2451 1050 2495 1056
rect 2451 1030 2460 1050
rect 2480 1030 2495 1050
rect 2451 1014 2495 1030
rect 2545 1046 2594 1056
rect 2545 1026 2563 1046
rect 2583 1026 2594 1046
rect 2545 1014 2594 1026
rect 8011 502 8060 514
rect 8011 482 8022 502
rect 8042 482 8060 502
rect 8011 472 8060 482
rect 8110 498 8154 514
rect 8110 478 8125 498
rect 8145 478 8154 498
rect 8110 472 8154 478
rect 8224 498 8268 514
rect 8224 478 8233 498
rect 8253 478 8268 498
rect 8224 472 8268 478
rect 8318 502 8367 514
rect 8318 482 8336 502
rect 8356 482 8367 502
rect 8318 472 8367 482
rect 8432 498 8476 514
rect 8432 478 8441 498
rect 8461 478 8476 498
rect 8432 472 8476 478
rect 8526 502 8575 514
rect 8526 482 8544 502
rect 8564 482 8575 502
rect 8526 472 8575 482
rect 8645 498 8689 514
rect 8645 478 8654 498
rect 8674 478 8689 498
rect 8645 472 8689 478
rect 8739 502 8788 514
rect 8739 482 8757 502
rect 8777 482 8788 502
rect 8739 472 8788 482
rect 9059 498 9108 510
rect 9059 478 9070 498
rect 9090 478 9108 498
rect 9059 468 9108 478
rect 9158 494 9202 510
rect 9158 474 9173 494
rect 9193 474 9202 494
rect 9158 468 9202 474
rect 9272 494 9316 510
rect 9272 474 9281 494
rect 9301 474 9316 494
rect 9272 468 9316 474
rect 9366 498 9415 510
rect 9366 478 9384 498
rect 9404 478 9415 498
rect 9366 468 9415 478
rect 9480 494 9524 510
rect 9480 474 9489 494
rect 9509 474 9524 494
rect 9480 468 9524 474
rect 9574 498 9623 510
rect 9574 478 9592 498
rect 9612 478 9623 498
rect 9574 468 9623 478
rect 9693 494 9737 510
rect 9693 474 9702 494
rect 9722 474 9737 494
rect 9693 468 9737 474
rect 9787 498 9836 510
rect 9787 478 9805 498
rect 9825 478 9836 498
rect 9787 468 9836 478
rect 769 371 818 381
rect 769 351 780 371
rect 800 351 818 371
rect 769 339 818 351
rect 868 375 912 381
rect 868 355 883 375
rect 903 355 912 375
rect 868 339 912 355
rect 982 371 1031 381
rect 982 351 993 371
rect 1013 351 1031 371
rect 982 339 1031 351
rect 1081 375 1125 381
rect 1081 355 1096 375
rect 1116 355 1125 375
rect 1081 339 1125 355
rect 1190 371 1239 381
rect 1190 351 1201 371
rect 1221 351 1239 371
rect 1190 339 1239 351
rect 1289 375 1333 381
rect 1289 355 1304 375
rect 1324 355 1333 375
rect 1289 339 1333 355
rect 1403 375 1447 381
rect 1403 355 1412 375
rect 1432 355 1447 375
rect 1403 339 1447 355
rect 1497 371 1546 381
rect 1497 351 1515 371
rect 1535 351 1546 371
rect 1497 339 1546 351
<< pdiff >>
rect 775 11621 819 11659
rect 775 11601 787 11621
rect 807 11601 819 11621
rect 775 11559 819 11601
rect 869 11621 911 11659
rect 869 11601 883 11621
rect 903 11601 911 11621
rect 869 11559 911 11601
rect 988 11621 1032 11659
rect 988 11601 1000 11621
rect 1020 11601 1032 11621
rect 988 11559 1032 11601
rect 1082 11621 1124 11659
rect 1082 11601 1096 11621
rect 1116 11601 1124 11621
rect 1082 11559 1124 11601
rect 1196 11621 1240 11659
rect 1196 11601 1208 11621
rect 1228 11601 1240 11621
rect 1196 11559 1240 11601
rect 1290 11621 1332 11659
rect 1290 11601 1304 11621
rect 1324 11601 1332 11621
rect 1290 11559 1332 11601
rect 1406 11621 1448 11659
rect 1406 11601 1414 11621
rect 1434 11601 1448 11621
rect 1406 11559 1448 11601
rect 1498 11628 1543 11659
rect 1498 11621 1542 11628
rect 1498 11601 1510 11621
rect 1530 11601 1542 11621
rect 1498 11559 1542 11601
rect 1823 11617 1867 11655
rect 1823 11597 1835 11617
rect 1855 11597 1867 11617
rect 1823 11555 1867 11597
rect 1917 11617 1959 11655
rect 1917 11597 1931 11617
rect 1951 11597 1959 11617
rect 1917 11555 1959 11597
rect 2036 11617 2080 11655
rect 2036 11597 2048 11617
rect 2068 11597 2080 11617
rect 2036 11555 2080 11597
rect 2130 11617 2172 11655
rect 2130 11597 2144 11617
rect 2164 11597 2172 11617
rect 2130 11555 2172 11597
rect 2244 11617 2288 11655
rect 2244 11597 2256 11617
rect 2276 11597 2288 11617
rect 2244 11555 2288 11597
rect 2338 11617 2380 11655
rect 2338 11597 2352 11617
rect 2372 11597 2380 11617
rect 2338 11555 2380 11597
rect 2454 11617 2496 11655
rect 2454 11597 2462 11617
rect 2482 11597 2496 11617
rect 2454 11555 2496 11597
rect 2546 11624 2591 11655
rect 2546 11617 2590 11624
rect 2546 11597 2558 11617
rect 2578 11597 2590 11617
rect 2546 11555 2590 11597
rect 9065 11450 9109 11492
rect 9065 11430 9077 11450
rect 9097 11430 9109 11450
rect 9065 11423 9109 11430
rect 9064 11392 9109 11423
rect 9159 11450 9201 11492
rect 9159 11430 9173 11450
rect 9193 11430 9201 11450
rect 9159 11392 9201 11430
rect 9275 11450 9317 11492
rect 9275 11430 9283 11450
rect 9303 11430 9317 11450
rect 9275 11392 9317 11430
rect 9367 11450 9411 11492
rect 9367 11430 9379 11450
rect 9399 11430 9411 11450
rect 9367 11392 9411 11430
rect 9483 11450 9525 11492
rect 9483 11430 9491 11450
rect 9511 11430 9525 11450
rect 9483 11392 9525 11430
rect 9575 11450 9619 11492
rect 9575 11430 9587 11450
rect 9607 11430 9619 11450
rect 9575 11392 9619 11430
rect 9696 11450 9738 11492
rect 9696 11430 9704 11450
rect 9724 11430 9738 11450
rect 9696 11392 9738 11430
rect 9788 11450 9832 11492
rect 9788 11430 9800 11450
rect 9820 11430 9832 11450
rect 9788 11392 9832 11430
rect 775 10942 819 10980
rect 775 10922 787 10942
rect 807 10922 819 10942
rect 775 10880 819 10922
rect 869 10942 911 10980
rect 869 10922 883 10942
rect 903 10922 911 10942
rect 869 10880 911 10922
rect 988 10942 1032 10980
rect 988 10922 1000 10942
rect 1020 10922 1032 10942
rect 988 10880 1032 10922
rect 1082 10942 1124 10980
rect 1082 10922 1096 10942
rect 1116 10922 1124 10942
rect 1082 10880 1124 10922
rect 1196 10942 1240 10980
rect 1196 10922 1208 10942
rect 1228 10922 1240 10942
rect 1196 10880 1240 10922
rect 1290 10942 1332 10980
rect 1290 10922 1304 10942
rect 1324 10922 1332 10942
rect 1290 10880 1332 10922
rect 1406 10942 1448 10980
rect 1406 10922 1414 10942
rect 1434 10922 1448 10942
rect 1406 10880 1448 10922
rect 1498 10949 1543 10980
rect 1498 10942 1542 10949
rect 1498 10922 1510 10942
rect 1530 10922 1542 10942
rect 1498 10880 1542 10922
rect 3270 10937 3314 10975
rect 3270 10917 3282 10937
rect 3302 10917 3314 10937
rect 3270 10875 3314 10917
rect 3364 10937 3406 10975
rect 3364 10917 3378 10937
rect 3398 10917 3406 10937
rect 3364 10875 3406 10917
rect 3483 10937 3527 10975
rect 3483 10917 3495 10937
rect 3515 10917 3527 10937
rect 3483 10875 3527 10917
rect 3577 10937 3619 10975
rect 3577 10917 3591 10937
rect 3611 10917 3619 10937
rect 3577 10875 3619 10917
rect 3691 10937 3735 10975
rect 3691 10917 3703 10937
rect 3723 10917 3735 10937
rect 3691 10875 3735 10917
rect 3785 10937 3827 10975
rect 3785 10917 3799 10937
rect 3819 10917 3827 10937
rect 3785 10875 3827 10917
rect 3901 10937 3943 10975
rect 3901 10917 3909 10937
rect 3929 10917 3943 10937
rect 3901 10875 3943 10917
rect 3993 10944 4038 10975
rect 3993 10937 4037 10944
rect 3993 10917 4005 10937
rect 4025 10917 4037 10937
rect 3993 10875 4037 10917
rect 8017 10775 8061 10817
rect 8017 10755 8029 10775
rect 8049 10755 8061 10775
rect 8017 10748 8061 10755
rect 8016 10717 8061 10748
rect 8111 10775 8153 10817
rect 8111 10755 8125 10775
rect 8145 10755 8153 10775
rect 8111 10717 8153 10755
rect 8227 10775 8269 10817
rect 8227 10755 8235 10775
rect 8255 10755 8269 10775
rect 8227 10717 8269 10755
rect 8319 10775 8363 10817
rect 8319 10755 8331 10775
rect 8351 10755 8363 10775
rect 8319 10717 8363 10755
rect 8435 10775 8477 10817
rect 8435 10755 8443 10775
rect 8463 10755 8477 10775
rect 8435 10717 8477 10755
rect 8527 10775 8571 10817
rect 8527 10755 8539 10775
rect 8559 10755 8571 10775
rect 8527 10717 8571 10755
rect 8648 10775 8690 10817
rect 8648 10755 8656 10775
rect 8676 10755 8690 10775
rect 8648 10717 8690 10755
rect 8740 10775 8784 10817
rect 8740 10755 8752 10775
rect 8772 10755 8784 10775
rect 8740 10717 8784 10755
rect 9065 10771 9109 10813
rect 9065 10751 9077 10771
rect 9097 10751 9109 10771
rect 9065 10744 9109 10751
rect 9064 10713 9109 10744
rect 9159 10771 9201 10813
rect 9159 10751 9173 10771
rect 9193 10751 9201 10771
rect 9159 10713 9201 10751
rect 9275 10771 9317 10813
rect 9275 10751 9283 10771
rect 9303 10751 9317 10771
rect 9275 10713 9317 10751
rect 9367 10771 9411 10813
rect 9367 10751 9379 10771
rect 9399 10751 9411 10771
rect 9367 10713 9411 10751
rect 9483 10771 9525 10813
rect 9483 10751 9491 10771
rect 9511 10751 9525 10771
rect 9483 10713 9525 10751
rect 9575 10771 9619 10813
rect 9575 10751 9587 10771
rect 9607 10751 9619 10771
rect 9575 10713 9619 10751
rect 9696 10771 9738 10813
rect 9696 10751 9704 10771
rect 9724 10751 9738 10771
rect 9696 10713 9738 10751
rect 9788 10771 9832 10813
rect 9788 10751 9800 10771
rect 9820 10751 9832 10771
rect 9788 10713 9832 10751
rect 775 10174 819 10212
rect 775 10154 787 10174
rect 807 10154 819 10174
rect 775 10112 819 10154
rect 869 10174 911 10212
rect 869 10154 883 10174
rect 903 10154 911 10174
rect 869 10112 911 10154
rect 988 10174 1032 10212
rect 988 10154 1000 10174
rect 1020 10154 1032 10174
rect 988 10112 1032 10154
rect 1082 10174 1124 10212
rect 1082 10154 1096 10174
rect 1116 10154 1124 10174
rect 1082 10112 1124 10154
rect 1196 10174 1240 10212
rect 1196 10154 1208 10174
rect 1228 10154 1240 10174
rect 1196 10112 1240 10154
rect 1290 10174 1332 10212
rect 1290 10154 1304 10174
rect 1324 10154 1332 10174
rect 1290 10112 1332 10154
rect 1406 10174 1448 10212
rect 1406 10154 1414 10174
rect 1434 10154 1448 10174
rect 1406 10112 1448 10154
rect 1498 10181 1543 10212
rect 1498 10174 1542 10181
rect 1498 10154 1510 10174
rect 1530 10154 1542 10174
rect 1498 10112 1542 10154
rect 1823 10170 1867 10208
rect 1823 10150 1835 10170
rect 1855 10150 1867 10170
rect 1823 10108 1867 10150
rect 1917 10170 1959 10208
rect 1917 10150 1931 10170
rect 1951 10150 1959 10170
rect 1917 10108 1959 10150
rect 2036 10170 2080 10208
rect 2036 10150 2048 10170
rect 2068 10150 2080 10170
rect 2036 10108 2080 10150
rect 2130 10170 2172 10208
rect 2130 10150 2144 10170
rect 2164 10150 2172 10170
rect 2130 10108 2172 10150
rect 2244 10170 2288 10208
rect 2244 10150 2256 10170
rect 2276 10150 2288 10170
rect 2244 10108 2288 10150
rect 2338 10170 2380 10208
rect 2338 10150 2352 10170
rect 2372 10150 2380 10170
rect 2338 10108 2380 10150
rect 2454 10170 2496 10208
rect 2454 10150 2462 10170
rect 2482 10150 2496 10170
rect 2454 10108 2496 10150
rect 2546 10177 2591 10208
rect 2546 10170 2590 10177
rect 2546 10150 2558 10170
rect 2578 10150 2590 10170
rect 2546 10108 2590 10150
rect 6570 10008 6614 10050
rect 6570 9988 6582 10008
rect 6602 9988 6614 10008
rect 6570 9981 6614 9988
rect 6569 9950 6614 9981
rect 6664 10008 6706 10050
rect 6664 9988 6678 10008
rect 6698 9988 6706 10008
rect 6664 9950 6706 9988
rect 6780 10008 6822 10050
rect 6780 9988 6788 10008
rect 6808 9988 6822 10008
rect 6780 9950 6822 9988
rect 6872 10008 6916 10050
rect 6872 9988 6884 10008
rect 6904 9988 6916 10008
rect 6872 9950 6916 9988
rect 6988 10008 7030 10050
rect 6988 9988 6996 10008
rect 7016 9988 7030 10008
rect 6988 9950 7030 9988
rect 7080 10008 7124 10050
rect 7080 9988 7092 10008
rect 7112 9988 7124 10008
rect 7080 9950 7124 9988
rect 7201 10008 7243 10050
rect 7201 9988 7209 10008
rect 7229 9988 7243 10008
rect 7201 9950 7243 9988
rect 7293 10008 7337 10050
rect 7293 9988 7305 10008
rect 7325 9988 7337 10008
rect 7293 9950 7337 9988
rect 9065 10003 9109 10045
rect 9065 9983 9077 10003
rect 9097 9983 9109 10003
rect 9065 9976 9109 9983
rect 9064 9945 9109 9976
rect 9159 10003 9201 10045
rect 9159 9983 9173 10003
rect 9193 9983 9201 10003
rect 9159 9945 9201 9983
rect 9275 10003 9317 10045
rect 9275 9983 9283 10003
rect 9303 9983 9317 10003
rect 9275 9945 9317 9983
rect 9367 10003 9411 10045
rect 9367 9983 9379 10003
rect 9399 9983 9411 10003
rect 9367 9945 9411 9983
rect 9483 10003 9525 10045
rect 9483 9983 9491 10003
rect 9511 9983 9525 10003
rect 9483 9945 9525 9983
rect 9575 10003 9619 10045
rect 9575 9983 9587 10003
rect 9607 9983 9619 10003
rect 9575 9945 9619 9983
rect 9696 10003 9738 10045
rect 9696 9983 9704 10003
rect 9724 9983 9738 10003
rect 9696 9945 9738 9983
rect 9788 10003 9832 10045
rect 9788 9983 9800 10003
rect 9820 9983 9832 10003
rect 9788 9945 9832 9983
rect 775 9495 819 9533
rect 775 9475 787 9495
rect 807 9475 819 9495
rect 775 9433 819 9475
rect 869 9495 911 9533
rect 869 9475 883 9495
rect 903 9475 911 9495
rect 869 9433 911 9475
rect 988 9495 1032 9533
rect 988 9475 1000 9495
rect 1020 9475 1032 9495
rect 988 9433 1032 9475
rect 1082 9495 1124 9533
rect 1082 9475 1096 9495
rect 1116 9475 1124 9495
rect 1082 9433 1124 9475
rect 1196 9495 1240 9533
rect 1196 9475 1208 9495
rect 1228 9475 1240 9495
rect 1196 9433 1240 9475
rect 1290 9495 1332 9533
rect 1290 9475 1304 9495
rect 1324 9475 1332 9495
rect 1290 9433 1332 9475
rect 1406 9495 1448 9533
rect 1406 9475 1414 9495
rect 1434 9475 1448 9495
rect 1406 9433 1448 9475
rect 1498 9502 1543 9533
rect 1498 9495 1542 9502
rect 1498 9475 1510 9495
rect 1530 9475 1542 9495
rect 1498 9433 1542 9475
rect 3313 9492 3357 9530
rect 3313 9472 3325 9492
rect 3345 9472 3357 9492
rect 3313 9430 3357 9472
rect 3407 9492 3449 9530
rect 3407 9472 3421 9492
rect 3441 9472 3449 9492
rect 3407 9430 3449 9472
rect 3526 9492 3570 9530
rect 3526 9472 3538 9492
rect 3558 9472 3570 9492
rect 3526 9430 3570 9472
rect 3620 9492 3662 9530
rect 3620 9472 3634 9492
rect 3654 9472 3662 9492
rect 3620 9430 3662 9472
rect 3734 9492 3778 9530
rect 3734 9472 3746 9492
rect 3766 9472 3778 9492
rect 3734 9430 3778 9472
rect 3828 9492 3870 9530
rect 3828 9472 3842 9492
rect 3862 9472 3870 9492
rect 3828 9430 3870 9472
rect 3944 9492 3986 9530
rect 3944 9472 3952 9492
rect 3972 9472 3986 9492
rect 3944 9430 3986 9472
rect 4036 9499 4081 9530
rect 4036 9492 4080 9499
rect 4036 9472 4048 9492
rect 4068 9472 4080 9492
rect 4036 9430 4080 9472
rect 8017 9328 8061 9370
rect 8017 9308 8029 9328
rect 8049 9308 8061 9328
rect 8017 9301 8061 9308
rect 8016 9270 8061 9301
rect 8111 9328 8153 9370
rect 8111 9308 8125 9328
rect 8145 9308 8153 9328
rect 8111 9270 8153 9308
rect 8227 9328 8269 9370
rect 8227 9308 8235 9328
rect 8255 9308 8269 9328
rect 8227 9270 8269 9308
rect 8319 9328 8363 9370
rect 8319 9308 8331 9328
rect 8351 9308 8363 9328
rect 8319 9270 8363 9308
rect 8435 9328 8477 9370
rect 8435 9308 8443 9328
rect 8463 9308 8477 9328
rect 8435 9270 8477 9308
rect 8527 9328 8571 9370
rect 8527 9308 8539 9328
rect 8559 9308 8571 9328
rect 8527 9270 8571 9308
rect 8648 9328 8690 9370
rect 8648 9308 8656 9328
rect 8676 9308 8690 9328
rect 8648 9270 8690 9308
rect 8740 9328 8784 9370
rect 8740 9308 8752 9328
rect 8772 9308 8784 9328
rect 8740 9270 8784 9308
rect 9065 9324 9109 9366
rect 9065 9304 9077 9324
rect 9097 9304 9109 9324
rect 9065 9297 9109 9304
rect 9064 9266 9109 9297
rect 9159 9324 9201 9366
rect 9159 9304 9173 9324
rect 9193 9304 9201 9324
rect 9159 9266 9201 9304
rect 9275 9324 9317 9366
rect 9275 9304 9283 9324
rect 9303 9304 9317 9324
rect 9275 9266 9317 9304
rect 9367 9324 9411 9366
rect 9367 9304 9379 9324
rect 9399 9304 9411 9324
rect 9367 9266 9411 9304
rect 9483 9324 9525 9366
rect 9483 9304 9491 9324
rect 9511 9304 9525 9324
rect 9483 9266 9525 9304
rect 9575 9324 9619 9366
rect 9575 9304 9587 9324
rect 9607 9304 9619 9324
rect 9575 9266 9619 9304
rect 9696 9324 9738 9366
rect 9696 9304 9704 9324
rect 9724 9304 9738 9324
rect 9696 9266 9738 9304
rect 9788 9324 9832 9366
rect 9788 9304 9800 9324
rect 9820 9304 9832 9324
rect 9788 9266 9832 9304
rect 776 8654 820 8692
rect 776 8634 788 8654
rect 808 8634 820 8654
rect 776 8592 820 8634
rect 870 8654 912 8692
rect 870 8634 884 8654
rect 904 8634 912 8654
rect 870 8592 912 8634
rect 989 8654 1033 8692
rect 989 8634 1001 8654
rect 1021 8634 1033 8654
rect 989 8592 1033 8634
rect 1083 8654 1125 8692
rect 1083 8634 1097 8654
rect 1117 8634 1125 8654
rect 1083 8592 1125 8634
rect 1197 8654 1241 8692
rect 1197 8634 1209 8654
rect 1229 8634 1241 8654
rect 1197 8592 1241 8634
rect 1291 8654 1333 8692
rect 1291 8634 1305 8654
rect 1325 8634 1333 8654
rect 1291 8592 1333 8634
rect 1407 8654 1449 8692
rect 1407 8634 1415 8654
rect 1435 8634 1449 8654
rect 1407 8592 1449 8634
rect 1499 8661 1544 8692
rect 1499 8654 1543 8661
rect 1499 8634 1511 8654
rect 1531 8634 1543 8654
rect 1499 8592 1543 8634
rect 1824 8650 1868 8688
rect 1824 8630 1836 8650
rect 1856 8630 1868 8650
rect 1824 8588 1868 8630
rect 1918 8650 1960 8688
rect 1918 8630 1932 8650
rect 1952 8630 1960 8650
rect 1918 8588 1960 8630
rect 2037 8650 2081 8688
rect 2037 8630 2049 8650
rect 2069 8630 2081 8650
rect 2037 8588 2081 8630
rect 2131 8650 2173 8688
rect 2131 8630 2145 8650
rect 2165 8630 2173 8650
rect 2131 8588 2173 8630
rect 2245 8650 2289 8688
rect 2245 8630 2257 8650
rect 2277 8630 2289 8650
rect 2245 8588 2289 8630
rect 2339 8650 2381 8688
rect 2339 8630 2353 8650
rect 2373 8630 2381 8650
rect 2339 8588 2381 8630
rect 2455 8650 2497 8688
rect 2455 8630 2463 8650
rect 2483 8630 2497 8650
rect 2455 8588 2497 8630
rect 2547 8657 2592 8688
rect 2547 8650 2591 8657
rect 2547 8630 2559 8650
rect 2579 8630 2591 8650
rect 2547 8588 2591 8630
rect 6528 8486 6572 8528
rect 6528 8466 6540 8486
rect 6560 8466 6572 8486
rect 6528 8459 6572 8466
rect 6527 8428 6572 8459
rect 6622 8486 6664 8528
rect 6622 8466 6636 8486
rect 6656 8466 6664 8486
rect 6622 8428 6664 8466
rect 6738 8486 6780 8528
rect 6738 8466 6746 8486
rect 6766 8466 6780 8486
rect 6738 8428 6780 8466
rect 6830 8486 6874 8528
rect 6830 8466 6842 8486
rect 6862 8466 6874 8486
rect 6830 8428 6874 8466
rect 6946 8486 6988 8528
rect 6946 8466 6954 8486
rect 6974 8466 6988 8486
rect 6946 8428 6988 8466
rect 7038 8486 7082 8528
rect 7038 8466 7050 8486
rect 7070 8466 7082 8486
rect 7038 8428 7082 8466
rect 7159 8486 7201 8528
rect 7159 8466 7167 8486
rect 7187 8466 7201 8486
rect 7159 8428 7201 8466
rect 7251 8486 7295 8528
rect 7251 8466 7263 8486
rect 7283 8466 7295 8486
rect 7251 8428 7295 8466
rect 9066 8483 9110 8525
rect 9066 8463 9078 8483
rect 9098 8463 9110 8483
rect 9066 8456 9110 8463
rect 9065 8425 9110 8456
rect 9160 8483 9202 8525
rect 9160 8463 9174 8483
rect 9194 8463 9202 8483
rect 9160 8425 9202 8463
rect 9276 8483 9318 8525
rect 9276 8463 9284 8483
rect 9304 8463 9318 8483
rect 9276 8425 9318 8463
rect 9368 8483 9412 8525
rect 9368 8463 9380 8483
rect 9400 8463 9412 8483
rect 9368 8425 9412 8463
rect 9484 8483 9526 8525
rect 9484 8463 9492 8483
rect 9512 8463 9526 8483
rect 9484 8425 9526 8463
rect 9576 8483 9620 8525
rect 9576 8463 9588 8483
rect 9608 8463 9620 8483
rect 9576 8425 9620 8463
rect 9697 8483 9739 8525
rect 9697 8463 9705 8483
rect 9725 8463 9739 8483
rect 9697 8425 9739 8463
rect 9789 8483 9833 8525
rect 9789 8463 9801 8483
rect 9821 8463 9833 8483
rect 9789 8425 9833 8463
rect 776 7975 820 8013
rect 776 7955 788 7975
rect 808 7955 820 7975
rect 776 7913 820 7955
rect 870 7975 912 8013
rect 870 7955 884 7975
rect 904 7955 912 7975
rect 870 7913 912 7955
rect 989 7975 1033 8013
rect 989 7955 1001 7975
rect 1021 7955 1033 7975
rect 989 7913 1033 7955
rect 1083 7975 1125 8013
rect 1083 7955 1097 7975
rect 1117 7955 1125 7975
rect 1083 7913 1125 7955
rect 1197 7975 1241 8013
rect 1197 7955 1209 7975
rect 1229 7955 1241 7975
rect 1197 7913 1241 7955
rect 1291 7975 1333 8013
rect 1291 7955 1305 7975
rect 1325 7955 1333 7975
rect 1291 7913 1333 7955
rect 1407 7975 1449 8013
rect 1407 7955 1415 7975
rect 1435 7955 1449 7975
rect 1407 7913 1449 7955
rect 1499 7982 1544 8013
rect 1499 7975 1543 7982
rect 1499 7955 1511 7975
rect 1531 7955 1543 7975
rect 1499 7913 1543 7955
rect 3271 7970 3315 8008
rect 3271 7950 3283 7970
rect 3303 7950 3315 7970
rect 3271 7908 3315 7950
rect 3365 7970 3407 8008
rect 3365 7950 3379 7970
rect 3399 7950 3407 7970
rect 3365 7908 3407 7950
rect 3484 7970 3528 8008
rect 3484 7950 3496 7970
rect 3516 7950 3528 7970
rect 3484 7908 3528 7950
rect 3578 7970 3620 8008
rect 3578 7950 3592 7970
rect 3612 7950 3620 7970
rect 3578 7908 3620 7950
rect 3692 7970 3736 8008
rect 3692 7950 3704 7970
rect 3724 7950 3736 7970
rect 3692 7908 3736 7950
rect 3786 7970 3828 8008
rect 3786 7950 3800 7970
rect 3820 7950 3828 7970
rect 3786 7908 3828 7950
rect 3902 7970 3944 8008
rect 3902 7950 3910 7970
rect 3930 7950 3944 7970
rect 3902 7908 3944 7950
rect 3994 7977 4039 8008
rect 3994 7970 4038 7977
rect 3994 7950 4006 7970
rect 4026 7950 4038 7970
rect 3994 7908 4038 7950
rect 8018 7808 8062 7850
rect 8018 7788 8030 7808
rect 8050 7788 8062 7808
rect 8018 7781 8062 7788
rect 8017 7750 8062 7781
rect 8112 7808 8154 7850
rect 8112 7788 8126 7808
rect 8146 7788 8154 7808
rect 8112 7750 8154 7788
rect 8228 7808 8270 7850
rect 8228 7788 8236 7808
rect 8256 7788 8270 7808
rect 8228 7750 8270 7788
rect 8320 7808 8364 7850
rect 8320 7788 8332 7808
rect 8352 7788 8364 7808
rect 8320 7750 8364 7788
rect 8436 7808 8478 7850
rect 8436 7788 8444 7808
rect 8464 7788 8478 7808
rect 8436 7750 8478 7788
rect 8528 7808 8572 7850
rect 8528 7788 8540 7808
rect 8560 7788 8572 7808
rect 8528 7750 8572 7788
rect 8649 7808 8691 7850
rect 8649 7788 8657 7808
rect 8677 7788 8691 7808
rect 8649 7750 8691 7788
rect 8741 7808 8785 7850
rect 8741 7788 8753 7808
rect 8773 7788 8785 7808
rect 8741 7750 8785 7788
rect 9066 7804 9110 7846
rect 9066 7784 9078 7804
rect 9098 7784 9110 7804
rect 9066 7777 9110 7784
rect 9065 7746 9110 7777
rect 9160 7804 9202 7846
rect 9160 7784 9174 7804
rect 9194 7784 9202 7804
rect 9160 7746 9202 7784
rect 9276 7804 9318 7846
rect 9276 7784 9284 7804
rect 9304 7784 9318 7804
rect 9276 7746 9318 7784
rect 9368 7804 9412 7846
rect 9368 7784 9380 7804
rect 9400 7784 9412 7804
rect 9368 7746 9412 7784
rect 9484 7804 9526 7846
rect 9484 7784 9492 7804
rect 9512 7784 9526 7804
rect 9484 7746 9526 7784
rect 9576 7804 9620 7846
rect 9576 7784 9588 7804
rect 9608 7784 9620 7804
rect 9576 7746 9620 7784
rect 9697 7804 9739 7846
rect 9697 7784 9705 7804
rect 9725 7784 9739 7804
rect 9697 7746 9739 7784
rect 9789 7804 9833 7846
rect 9789 7784 9801 7804
rect 9821 7784 9833 7804
rect 9789 7746 9833 7784
rect 776 7207 820 7245
rect 776 7187 788 7207
rect 808 7187 820 7207
rect 776 7145 820 7187
rect 870 7207 912 7245
rect 870 7187 884 7207
rect 904 7187 912 7207
rect 870 7145 912 7187
rect 989 7207 1033 7245
rect 989 7187 1001 7207
rect 1021 7187 1033 7207
rect 989 7145 1033 7187
rect 1083 7207 1125 7245
rect 1083 7187 1097 7207
rect 1117 7187 1125 7207
rect 1083 7145 1125 7187
rect 1197 7207 1241 7245
rect 1197 7187 1209 7207
rect 1229 7187 1241 7207
rect 1197 7145 1241 7187
rect 1291 7207 1333 7245
rect 1291 7187 1305 7207
rect 1325 7187 1333 7207
rect 1291 7145 1333 7187
rect 1407 7207 1449 7245
rect 1407 7187 1415 7207
rect 1435 7187 1449 7207
rect 1407 7145 1449 7187
rect 1499 7214 1544 7245
rect 1499 7207 1543 7214
rect 1499 7187 1511 7207
rect 1531 7187 1543 7207
rect 1499 7145 1543 7187
rect 1824 7203 1868 7241
rect 1824 7183 1836 7203
rect 1856 7183 1868 7203
rect 1824 7141 1868 7183
rect 1918 7203 1960 7241
rect 1918 7183 1932 7203
rect 1952 7183 1960 7203
rect 1918 7141 1960 7183
rect 2037 7203 2081 7241
rect 2037 7183 2049 7203
rect 2069 7183 2081 7203
rect 2037 7141 2081 7183
rect 2131 7203 2173 7241
rect 2131 7183 2145 7203
rect 2165 7183 2173 7203
rect 2131 7141 2173 7183
rect 2245 7203 2289 7241
rect 2245 7183 2257 7203
rect 2277 7183 2289 7203
rect 2245 7141 2289 7183
rect 2339 7203 2381 7241
rect 2339 7183 2353 7203
rect 2373 7183 2381 7203
rect 2339 7141 2381 7183
rect 2455 7203 2497 7241
rect 2455 7183 2463 7203
rect 2483 7183 2497 7203
rect 2455 7141 2497 7183
rect 2547 7210 2592 7241
rect 2547 7203 2591 7210
rect 2547 7183 2559 7203
rect 2579 7183 2591 7203
rect 2547 7141 2591 7183
rect 6571 7041 6615 7083
rect 6571 7021 6583 7041
rect 6603 7021 6615 7041
rect 6571 7014 6615 7021
rect 6570 6983 6615 7014
rect 6665 7041 6707 7083
rect 6665 7021 6679 7041
rect 6699 7021 6707 7041
rect 6665 6983 6707 7021
rect 6781 7041 6823 7083
rect 6781 7021 6789 7041
rect 6809 7021 6823 7041
rect 6781 6983 6823 7021
rect 6873 7041 6917 7083
rect 6873 7021 6885 7041
rect 6905 7021 6917 7041
rect 6873 6983 6917 7021
rect 6989 7041 7031 7083
rect 6989 7021 6997 7041
rect 7017 7021 7031 7041
rect 6989 6983 7031 7021
rect 7081 7041 7125 7083
rect 7081 7021 7093 7041
rect 7113 7021 7125 7041
rect 7081 6983 7125 7021
rect 7202 7041 7244 7083
rect 7202 7021 7210 7041
rect 7230 7021 7244 7041
rect 7202 6983 7244 7021
rect 7294 7041 7338 7083
rect 7294 7021 7306 7041
rect 7326 7021 7338 7041
rect 7294 6983 7338 7021
rect 9066 7036 9110 7078
rect 9066 7016 9078 7036
rect 9098 7016 9110 7036
rect 9066 7009 9110 7016
rect 9065 6978 9110 7009
rect 9160 7036 9202 7078
rect 9160 7016 9174 7036
rect 9194 7016 9202 7036
rect 9160 6978 9202 7016
rect 9276 7036 9318 7078
rect 9276 7016 9284 7036
rect 9304 7016 9318 7036
rect 9276 6978 9318 7016
rect 9368 7036 9412 7078
rect 9368 7016 9380 7036
rect 9400 7016 9412 7036
rect 9368 6978 9412 7016
rect 9484 7036 9526 7078
rect 9484 7016 9492 7036
rect 9512 7016 9526 7036
rect 9484 6978 9526 7016
rect 9576 7036 9620 7078
rect 9576 7016 9588 7036
rect 9608 7016 9620 7036
rect 9576 6978 9620 7016
rect 9697 7036 9739 7078
rect 9697 7016 9705 7036
rect 9725 7016 9739 7036
rect 9697 6978 9739 7016
rect 9789 7036 9833 7078
rect 9789 7016 9801 7036
rect 9821 7016 9833 7036
rect 9789 6978 9833 7016
rect 776 6528 820 6566
rect 776 6508 788 6528
rect 808 6508 820 6528
rect 776 6466 820 6508
rect 870 6528 912 6566
rect 870 6508 884 6528
rect 904 6508 912 6528
rect 870 6466 912 6508
rect 989 6528 1033 6566
rect 989 6508 1001 6528
rect 1021 6508 1033 6528
rect 989 6466 1033 6508
rect 1083 6528 1125 6566
rect 1083 6508 1097 6528
rect 1117 6508 1125 6528
rect 1083 6466 1125 6508
rect 1197 6528 1241 6566
rect 1197 6508 1209 6528
rect 1229 6508 1241 6528
rect 1197 6466 1241 6508
rect 1291 6528 1333 6566
rect 1291 6508 1305 6528
rect 1325 6508 1333 6528
rect 1291 6466 1333 6508
rect 1407 6528 1449 6566
rect 1407 6508 1415 6528
rect 1435 6508 1449 6528
rect 1407 6466 1449 6508
rect 1499 6535 1544 6566
rect 1499 6528 1543 6535
rect 1499 6508 1511 6528
rect 1531 6508 1543 6528
rect 1499 6466 1543 6508
rect 4379 6519 4423 6557
rect 4379 6499 4391 6519
rect 4411 6499 4423 6519
rect 4379 6457 4423 6499
rect 4473 6519 4515 6557
rect 4473 6499 4487 6519
rect 4507 6499 4515 6519
rect 4473 6457 4515 6499
rect 4592 6519 4636 6557
rect 4592 6499 4604 6519
rect 4624 6499 4636 6519
rect 4592 6457 4636 6499
rect 4686 6519 4728 6557
rect 4686 6499 4700 6519
rect 4720 6499 4728 6519
rect 4686 6457 4728 6499
rect 4800 6519 4844 6557
rect 4800 6499 4812 6519
rect 4832 6499 4844 6519
rect 4800 6457 4844 6499
rect 4894 6519 4936 6557
rect 4894 6499 4908 6519
rect 4928 6499 4936 6519
rect 4894 6457 4936 6499
rect 5010 6519 5052 6557
rect 5010 6499 5018 6519
rect 5038 6499 5052 6519
rect 5010 6457 5052 6499
rect 5102 6526 5147 6557
rect 5102 6519 5146 6526
rect 5102 6499 5114 6519
rect 5134 6499 5146 6519
rect 5102 6457 5146 6499
rect 8018 6361 8062 6403
rect 8018 6341 8030 6361
rect 8050 6341 8062 6361
rect 8018 6334 8062 6341
rect 8017 6303 8062 6334
rect 8112 6361 8154 6403
rect 8112 6341 8126 6361
rect 8146 6341 8154 6361
rect 8112 6303 8154 6341
rect 8228 6361 8270 6403
rect 8228 6341 8236 6361
rect 8256 6341 8270 6361
rect 8228 6303 8270 6341
rect 8320 6361 8364 6403
rect 8320 6341 8332 6361
rect 8352 6341 8364 6361
rect 8320 6303 8364 6341
rect 8436 6361 8478 6403
rect 8436 6341 8444 6361
rect 8464 6341 8478 6361
rect 8436 6303 8478 6341
rect 8528 6361 8572 6403
rect 8528 6341 8540 6361
rect 8560 6341 8572 6361
rect 8528 6303 8572 6341
rect 8649 6361 8691 6403
rect 8649 6341 8657 6361
rect 8677 6341 8691 6361
rect 8649 6303 8691 6341
rect 8741 6361 8785 6403
rect 8741 6341 8753 6361
rect 8773 6341 8785 6361
rect 8741 6303 8785 6341
rect 9066 6357 9110 6399
rect 9066 6337 9078 6357
rect 9098 6337 9110 6357
rect 9066 6330 9110 6337
rect 9065 6299 9110 6330
rect 9160 6357 9202 6399
rect 9160 6337 9174 6357
rect 9194 6337 9202 6357
rect 9160 6299 9202 6337
rect 9276 6357 9318 6399
rect 9276 6337 9284 6357
rect 9304 6337 9318 6357
rect 9276 6299 9318 6337
rect 9368 6357 9412 6399
rect 9368 6337 9380 6357
rect 9400 6337 9412 6357
rect 9368 6299 9412 6337
rect 9484 6357 9526 6399
rect 9484 6337 9492 6357
rect 9512 6337 9526 6357
rect 9484 6299 9526 6337
rect 9576 6357 9620 6399
rect 9576 6337 9588 6357
rect 9608 6337 9620 6357
rect 9576 6299 9620 6337
rect 9697 6357 9739 6399
rect 9697 6337 9705 6357
rect 9725 6337 9739 6357
rect 9697 6299 9739 6337
rect 9789 6357 9833 6399
rect 9789 6337 9801 6357
rect 9821 6337 9833 6357
rect 9789 6299 9833 6337
rect 773 5613 817 5651
rect 773 5593 785 5613
rect 805 5593 817 5613
rect 773 5551 817 5593
rect 867 5613 909 5651
rect 867 5593 881 5613
rect 901 5593 909 5613
rect 867 5551 909 5593
rect 986 5613 1030 5651
rect 986 5593 998 5613
rect 1018 5593 1030 5613
rect 986 5551 1030 5593
rect 1080 5613 1122 5651
rect 1080 5593 1094 5613
rect 1114 5593 1122 5613
rect 1080 5551 1122 5593
rect 1194 5613 1238 5651
rect 1194 5593 1206 5613
rect 1226 5593 1238 5613
rect 1194 5551 1238 5593
rect 1288 5613 1330 5651
rect 1288 5593 1302 5613
rect 1322 5593 1330 5613
rect 1288 5551 1330 5593
rect 1404 5613 1446 5651
rect 1404 5593 1412 5613
rect 1432 5593 1446 5613
rect 1404 5551 1446 5593
rect 1496 5620 1541 5651
rect 1496 5613 1540 5620
rect 1496 5593 1508 5613
rect 1528 5593 1540 5613
rect 1496 5551 1540 5593
rect 1821 5609 1865 5647
rect 1821 5589 1833 5609
rect 1853 5589 1865 5609
rect 1821 5547 1865 5589
rect 1915 5609 1957 5647
rect 1915 5589 1929 5609
rect 1949 5589 1957 5609
rect 1915 5547 1957 5589
rect 2034 5609 2078 5647
rect 2034 5589 2046 5609
rect 2066 5589 2078 5609
rect 2034 5547 2078 5589
rect 2128 5609 2170 5647
rect 2128 5589 2142 5609
rect 2162 5589 2170 5609
rect 2128 5547 2170 5589
rect 2242 5609 2286 5647
rect 2242 5589 2254 5609
rect 2274 5589 2286 5609
rect 2242 5547 2286 5589
rect 2336 5609 2378 5647
rect 2336 5589 2350 5609
rect 2370 5589 2378 5609
rect 2336 5547 2378 5589
rect 2452 5609 2494 5647
rect 2452 5589 2460 5609
rect 2480 5589 2494 5609
rect 2452 5547 2494 5589
rect 2544 5616 2589 5647
rect 2544 5609 2588 5616
rect 2544 5589 2556 5609
rect 2576 5589 2588 5609
rect 2544 5547 2588 5589
rect 5460 5451 5504 5493
rect 5460 5431 5472 5451
rect 5492 5431 5504 5451
rect 5460 5424 5504 5431
rect 5459 5393 5504 5424
rect 5554 5451 5596 5493
rect 5554 5431 5568 5451
rect 5588 5431 5596 5451
rect 5554 5393 5596 5431
rect 5670 5451 5712 5493
rect 5670 5431 5678 5451
rect 5698 5431 5712 5451
rect 5670 5393 5712 5431
rect 5762 5451 5806 5493
rect 5762 5431 5774 5451
rect 5794 5431 5806 5451
rect 5762 5393 5806 5431
rect 5878 5451 5920 5493
rect 5878 5431 5886 5451
rect 5906 5431 5920 5451
rect 5878 5393 5920 5431
rect 5970 5451 6014 5493
rect 5970 5431 5982 5451
rect 6002 5431 6014 5451
rect 5970 5393 6014 5431
rect 6091 5451 6133 5493
rect 6091 5431 6099 5451
rect 6119 5431 6133 5451
rect 6091 5393 6133 5431
rect 6183 5451 6227 5493
rect 6183 5431 6195 5451
rect 6215 5431 6227 5451
rect 6183 5393 6227 5431
rect 9063 5442 9107 5484
rect 9063 5422 9075 5442
rect 9095 5422 9107 5442
rect 9063 5415 9107 5422
rect 9062 5384 9107 5415
rect 9157 5442 9199 5484
rect 9157 5422 9171 5442
rect 9191 5422 9199 5442
rect 9157 5384 9199 5422
rect 9273 5442 9315 5484
rect 9273 5422 9281 5442
rect 9301 5422 9315 5442
rect 9273 5384 9315 5422
rect 9365 5442 9409 5484
rect 9365 5422 9377 5442
rect 9397 5422 9409 5442
rect 9365 5384 9409 5422
rect 9481 5442 9523 5484
rect 9481 5422 9489 5442
rect 9509 5422 9523 5442
rect 9481 5384 9523 5422
rect 9573 5442 9617 5484
rect 9573 5422 9585 5442
rect 9605 5422 9617 5442
rect 9573 5384 9617 5422
rect 9694 5442 9736 5484
rect 9694 5422 9702 5442
rect 9722 5422 9736 5442
rect 9694 5384 9736 5422
rect 9786 5442 9830 5484
rect 9786 5422 9798 5442
rect 9818 5422 9830 5442
rect 9786 5384 9830 5422
rect 773 4934 817 4972
rect 773 4914 785 4934
rect 805 4914 817 4934
rect 773 4872 817 4914
rect 867 4934 909 4972
rect 867 4914 881 4934
rect 901 4914 909 4934
rect 867 4872 909 4914
rect 986 4934 1030 4972
rect 986 4914 998 4934
rect 1018 4914 1030 4934
rect 986 4872 1030 4914
rect 1080 4934 1122 4972
rect 1080 4914 1094 4934
rect 1114 4914 1122 4934
rect 1080 4872 1122 4914
rect 1194 4934 1238 4972
rect 1194 4914 1206 4934
rect 1226 4914 1238 4934
rect 1194 4872 1238 4914
rect 1288 4934 1330 4972
rect 1288 4914 1302 4934
rect 1322 4914 1330 4934
rect 1288 4872 1330 4914
rect 1404 4934 1446 4972
rect 1404 4914 1412 4934
rect 1432 4914 1446 4934
rect 1404 4872 1446 4914
rect 1496 4941 1541 4972
rect 1496 4934 1540 4941
rect 1496 4914 1508 4934
rect 1528 4914 1540 4934
rect 1496 4872 1540 4914
rect 3268 4929 3312 4967
rect 3268 4909 3280 4929
rect 3300 4909 3312 4929
rect 3268 4867 3312 4909
rect 3362 4929 3404 4967
rect 3362 4909 3376 4929
rect 3396 4909 3404 4929
rect 3362 4867 3404 4909
rect 3481 4929 3525 4967
rect 3481 4909 3493 4929
rect 3513 4909 3525 4929
rect 3481 4867 3525 4909
rect 3575 4929 3617 4967
rect 3575 4909 3589 4929
rect 3609 4909 3617 4929
rect 3575 4867 3617 4909
rect 3689 4929 3733 4967
rect 3689 4909 3701 4929
rect 3721 4909 3733 4929
rect 3689 4867 3733 4909
rect 3783 4929 3825 4967
rect 3783 4909 3797 4929
rect 3817 4909 3825 4929
rect 3783 4867 3825 4909
rect 3899 4929 3941 4967
rect 3899 4909 3907 4929
rect 3927 4909 3941 4929
rect 3899 4867 3941 4909
rect 3991 4936 4036 4967
rect 3991 4929 4035 4936
rect 3991 4909 4003 4929
rect 4023 4909 4035 4929
rect 3991 4867 4035 4909
rect 8015 4767 8059 4809
rect 8015 4747 8027 4767
rect 8047 4747 8059 4767
rect 8015 4740 8059 4747
rect 8014 4709 8059 4740
rect 8109 4767 8151 4809
rect 8109 4747 8123 4767
rect 8143 4747 8151 4767
rect 8109 4709 8151 4747
rect 8225 4767 8267 4809
rect 8225 4747 8233 4767
rect 8253 4747 8267 4767
rect 8225 4709 8267 4747
rect 8317 4767 8361 4809
rect 8317 4747 8329 4767
rect 8349 4747 8361 4767
rect 8317 4709 8361 4747
rect 8433 4767 8475 4809
rect 8433 4747 8441 4767
rect 8461 4747 8475 4767
rect 8433 4709 8475 4747
rect 8525 4767 8569 4809
rect 8525 4747 8537 4767
rect 8557 4747 8569 4767
rect 8525 4709 8569 4747
rect 8646 4767 8688 4809
rect 8646 4747 8654 4767
rect 8674 4747 8688 4767
rect 8646 4709 8688 4747
rect 8738 4767 8782 4809
rect 8738 4747 8750 4767
rect 8770 4747 8782 4767
rect 8738 4709 8782 4747
rect 9063 4763 9107 4805
rect 9063 4743 9075 4763
rect 9095 4743 9107 4763
rect 9063 4736 9107 4743
rect 9062 4705 9107 4736
rect 9157 4763 9199 4805
rect 9157 4743 9171 4763
rect 9191 4743 9199 4763
rect 9157 4705 9199 4743
rect 9273 4763 9315 4805
rect 9273 4743 9281 4763
rect 9301 4743 9315 4763
rect 9273 4705 9315 4743
rect 9365 4763 9409 4805
rect 9365 4743 9377 4763
rect 9397 4743 9409 4763
rect 9365 4705 9409 4743
rect 9481 4763 9523 4805
rect 9481 4743 9489 4763
rect 9509 4743 9523 4763
rect 9481 4705 9523 4743
rect 9573 4763 9617 4805
rect 9573 4743 9585 4763
rect 9605 4743 9617 4763
rect 9573 4705 9617 4743
rect 9694 4763 9736 4805
rect 9694 4743 9702 4763
rect 9722 4743 9736 4763
rect 9694 4705 9736 4743
rect 9786 4763 9830 4805
rect 9786 4743 9798 4763
rect 9818 4743 9830 4763
rect 9786 4705 9830 4743
rect 773 4166 817 4204
rect 773 4146 785 4166
rect 805 4146 817 4166
rect 773 4104 817 4146
rect 867 4166 909 4204
rect 867 4146 881 4166
rect 901 4146 909 4166
rect 867 4104 909 4146
rect 986 4166 1030 4204
rect 986 4146 998 4166
rect 1018 4146 1030 4166
rect 986 4104 1030 4146
rect 1080 4166 1122 4204
rect 1080 4146 1094 4166
rect 1114 4146 1122 4166
rect 1080 4104 1122 4146
rect 1194 4166 1238 4204
rect 1194 4146 1206 4166
rect 1226 4146 1238 4166
rect 1194 4104 1238 4146
rect 1288 4166 1330 4204
rect 1288 4146 1302 4166
rect 1322 4146 1330 4166
rect 1288 4104 1330 4146
rect 1404 4166 1446 4204
rect 1404 4146 1412 4166
rect 1432 4146 1446 4166
rect 1404 4104 1446 4146
rect 1496 4173 1541 4204
rect 1496 4166 1540 4173
rect 1496 4146 1508 4166
rect 1528 4146 1540 4166
rect 1496 4104 1540 4146
rect 1821 4162 1865 4200
rect 1821 4142 1833 4162
rect 1853 4142 1865 4162
rect 1821 4100 1865 4142
rect 1915 4162 1957 4200
rect 1915 4142 1929 4162
rect 1949 4142 1957 4162
rect 1915 4100 1957 4142
rect 2034 4162 2078 4200
rect 2034 4142 2046 4162
rect 2066 4142 2078 4162
rect 2034 4100 2078 4142
rect 2128 4162 2170 4200
rect 2128 4142 2142 4162
rect 2162 4142 2170 4162
rect 2128 4100 2170 4142
rect 2242 4162 2286 4200
rect 2242 4142 2254 4162
rect 2274 4142 2286 4162
rect 2242 4100 2286 4142
rect 2336 4162 2378 4200
rect 2336 4142 2350 4162
rect 2370 4142 2378 4162
rect 2336 4100 2378 4142
rect 2452 4162 2494 4200
rect 2452 4142 2460 4162
rect 2480 4142 2494 4162
rect 2452 4100 2494 4142
rect 2544 4169 2589 4200
rect 2544 4162 2588 4169
rect 2544 4142 2556 4162
rect 2576 4142 2588 4162
rect 2544 4100 2588 4142
rect 6568 4000 6612 4042
rect 6568 3980 6580 4000
rect 6600 3980 6612 4000
rect 6568 3973 6612 3980
rect 6567 3942 6612 3973
rect 6662 4000 6704 4042
rect 6662 3980 6676 4000
rect 6696 3980 6704 4000
rect 6662 3942 6704 3980
rect 6778 4000 6820 4042
rect 6778 3980 6786 4000
rect 6806 3980 6820 4000
rect 6778 3942 6820 3980
rect 6870 4000 6914 4042
rect 6870 3980 6882 4000
rect 6902 3980 6914 4000
rect 6870 3942 6914 3980
rect 6986 4000 7028 4042
rect 6986 3980 6994 4000
rect 7014 3980 7028 4000
rect 6986 3942 7028 3980
rect 7078 4000 7122 4042
rect 7078 3980 7090 4000
rect 7110 3980 7122 4000
rect 7078 3942 7122 3980
rect 7199 4000 7241 4042
rect 7199 3980 7207 4000
rect 7227 3980 7241 4000
rect 7199 3942 7241 3980
rect 7291 4000 7335 4042
rect 7291 3980 7303 4000
rect 7323 3980 7335 4000
rect 7291 3942 7335 3980
rect 9063 3995 9107 4037
rect 9063 3975 9075 3995
rect 9095 3975 9107 3995
rect 9063 3968 9107 3975
rect 9062 3937 9107 3968
rect 9157 3995 9199 4037
rect 9157 3975 9171 3995
rect 9191 3975 9199 3995
rect 9157 3937 9199 3975
rect 9273 3995 9315 4037
rect 9273 3975 9281 3995
rect 9301 3975 9315 3995
rect 9273 3937 9315 3975
rect 9365 3995 9409 4037
rect 9365 3975 9377 3995
rect 9397 3975 9409 3995
rect 9365 3937 9409 3975
rect 9481 3995 9523 4037
rect 9481 3975 9489 3995
rect 9509 3975 9523 3995
rect 9481 3937 9523 3975
rect 9573 3995 9617 4037
rect 9573 3975 9585 3995
rect 9605 3975 9617 3995
rect 9573 3937 9617 3975
rect 9694 3995 9736 4037
rect 9694 3975 9702 3995
rect 9722 3975 9736 3995
rect 9694 3937 9736 3975
rect 9786 3995 9830 4037
rect 9786 3975 9798 3995
rect 9818 3975 9830 3995
rect 9786 3937 9830 3975
rect 773 3487 817 3525
rect 773 3467 785 3487
rect 805 3467 817 3487
rect 773 3425 817 3467
rect 867 3487 909 3525
rect 867 3467 881 3487
rect 901 3467 909 3487
rect 867 3425 909 3467
rect 986 3487 1030 3525
rect 986 3467 998 3487
rect 1018 3467 1030 3487
rect 986 3425 1030 3467
rect 1080 3487 1122 3525
rect 1080 3467 1094 3487
rect 1114 3467 1122 3487
rect 1080 3425 1122 3467
rect 1194 3487 1238 3525
rect 1194 3467 1206 3487
rect 1226 3467 1238 3487
rect 1194 3425 1238 3467
rect 1288 3487 1330 3525
rect 1288 3467 1302 3487
rect 1322 3467 1330 3487
rect 1288 3425 1330 3467
rect 1404 3487 1446 3525
rect 1404 3467 1412 3487
rect 1432 3467 1446 3487
rect 1404 3425 1446 3467
rect 1496 3494 1541 3525
rect 1496 3487 1540 3494
rect 1496 3467 1508 3487
rect 1528 3467 1540 3487
rect 1496 3425 1540 3467
rect 3311 3484 3355 3522
rect 3311 3464 3323 3484
rect 3343 3464 3355 3484
rect 3311 3422 3355 3464
rect 3405 3484 3447 3522
rect 3405 3464 3419 3484
rect 3439 3464 3447 3484
rect 3405 3422 3447 3464
rect 3524 3484 3568 3522
rect 3524 3464 3536 3484
rect 3556 3464 3568 3484
rect 3524 3422 3568 3464
rect 3618 3484 3660 3522
rect 3618 3464 3632 3484
rect 3652 3464 3660 3484
rect 3618 3422 3660 3464
rect 3732 3484 3776 3522
rect 3732 3464 3744 3484
rect 3764 3464 3776 3484
rect 3732 3422 3776 3464
rect 3826 3484 3868 3522
rect 3826 3464 3840 3484
rect 3860 3464 3868 3484
rect 3826 3422 3868 3464
rect 3942 3484 3984 3522
rect 3942 3464 3950 3484
rect 3970 3464 3984 3484
rect 3942 3422 3984 3464
rect 4034 3491 4079 3522
rect 4034 3484 4078 3491
rect 4034 3464 4046 3484
rect 4066 3464 4078 3484
rect 4034 3422 4078 3464
rect 8015 3320 8059 3362
rect 8015 3300 8027 3320
rect 8047 3300 8059 3320
rect 8015 3293 8059 3300
rect 8014 3262 8059 3293
rect 8109 3320 8151 3362
rect 8109 3300 8123 3320
rect 8143 3300 8151 3320
rect 8109 3262 8151 3300
rect 8225 3320 8267 3362
rect 8225 3300 8233 3320
rect 8253 3300 8267 3320
rect 8225 3262 8267 3300
rect 8317 3320 8361 3362
rect 8317 3300 8329 3320
rect 8349 3300 8361 3320
rect 8317 3262 8361 3300
rect 8433 3320 8475 3362
rect 8433 3300 8441 3320
rect 8461 3300 8475 3320
rect 8433 3262 8475 3300
rect 8525 3320 8569 3362
rect 8525 3300 8537 3320
rect 8557 3300 8569 3320
rect 8525 3262 8569 3300
rect 8646 3320 8688 3362
rect 8646 3300 8654 3320
rect 8674 3300 8688 3320
rect 8646 3262 8688 3300
rect 8738 3320 8782 3362
rect 8738 3300 8750 3320
rect 8770 3300 8782 3320
rect 8738 3262 8782 3300
rect 9063 3316 9107 3358
rect 9063 3296 9075 3316
rect 9095 3296 9107 3316
rect 9063 3289 9107 3296
rect 9062 3258 9107 3289
rect 9157 3316 9199 3358
rect 9157 3296 9171 3316
rect 9191 3296 9199 3316
rect 9157 3258 9199 3296
rect 9273 3316 9315 3358
rect 9273 3296 9281 3316
rect 9301 3296 9315 3316
rect 9273 3258 9315 3296
rect 9365 3316 9409 3358
rect 9365 3296 9377 3316
rect 9397 3296 9409 3316
rect 9365 3258 9409 3296
rect 9481 3316 9523 3358
rect 9481 3296 9489 3316
rect 9509 3296 9523 3316
rect 9481 3258 9523 3296
rect 9573 3316 9617 3358
rect 9573 3296 9585 3316
rect 9605 3296 9617 3316
rect 9573 3258 9617 3296
rect 9694 3316 9736 3358
rect 9694 3296 9702 3316
rect 9722 3296 9736 3316
rect 9694 3258 9736 3296
rect 9786 3316 9830 3358
rect 9786 3296 9798 3316
rect 9818 3296 9830 3316
rect 9786 3258 9830 3296
rect 774 2646 818 2684
rect 774 2626 786 2646
rect 806 2626 818 2646
rect 774 2584 818 2626
rect 868 2646 910 2684
rect 868 2626 882 2646
rect 902 2626 910 2646
rect 868 2584 910 2626
rect 987 2646 1031 2684
rect 987 2626 999 2646
rect 1019 2626 1031 2646
rect 987 2584 1031 2626
rect 1081 2646 1123 2684
rect 1081 2626 1095 2646
rect 1115 2626 1123 2646
rect 1081 2584 1123 2626
rect 1195 2646 1239 2684
rect 1195 2626 1207 2646
rect 1227 2626 1239 2646
rect 1195 2584 1239 2626
rect 1289 2646 1331 2684
rect 1289 2626 1303 2646
rect 1323 2626 1331 2646
rect 1289 2584 1331 2626
rect 1405 2646 1447 2684
rect 1405 2626 1413 2646
rect 1433 2626 1447 2646
rect 1405 2584 1447 2626
rect 1497 2653 1542 2684
rect 1497 2646 1541 2653
rect 1497 2626 1509 2646
rect 1529 2626 1541 2646
rect 1497 2584 1541 2626
rect 1822 2642 1866 2680
rect 1822 2622 1834 2642
rect 1854 2622 1866 2642
rect 1822 2580 1866 2622
rect 1916 2642 1958 2680
rect 1916 2622 1930 2642
rect 1950 2622 1958 2642
rect 1916 2580 1958 2622
rect 2035 2642 2079 2680
rect 2035 2622 2047 2642
rect 2067 2622 2079 2642
rect 2035 2580 2079 2622
rect 2129 2642 2171 2680
rect 2129 2622 2143 2642
rect 2163 2622 2171 2642
rect 2129 2580 2171 2622
rect 2243 2642 2287 2680
rect 2243 2622 2255 2642
rect 2275 2622 2287 2642
rect 2243 2580 2287 2622
rect 2337 2642 2379 2680
rect 2337 2622 2351 2642
rect 2371 2622 2379 2642
rect 2337 2580 2379 2622
rect 2453 2642 2495 2680
rect 2453 2622 2461 2642
rect 2481 2622 2495 2642
rect 2453 2580 2495 2622
rect 2545 2649 2590 2680
rect 2545 2642 2589 2649
rect 2545 2622 2557 2642
rect 2577 2622 2589 2642
rect 2545 2580 2589 2622
rect 4724 2648 4768 2686
rect 4724 2628 4736 2648
rect 4756 2628 4768 2648
rect 4724 2586 4768 2628
rect 4818 2648 4860 2686
rect 4818 2628 4832 2648
rect 4852 2628 4860 2648
rect 4818 2586 4860 2628
rect 4937 2648 4981 2686
rect 4937 2628 4949 2648
rect 4969 2628 4981 2648
rect 4937 2586 4981 2628
rect 5031 2648 5073 2686
rect 5031 2628 5045 2648
rect 5065 2628 5073 2648
rect 5031 2586 5073 2628
rect 5145 2648 5189 2686
rect 5145 2628 5157 2648
rect 5177 2628 5189 2648
rect 5145 2586 5189 2628
rect 5239 2648 5281 2686
rect 5239 2628 5253 2648
rect 5273 2628 5281 2648
rect 5239 2586 5281 2628
rect 5355 2648 5397 2686
rect 5355 2628 5363 2648
rect 5383 2628 5397 2648
rect 5355 2586 5397 2628
rect 5447 2655 5492 2686
rect 5447 2648 5491 2655
rect 5447 2628 5459 2648
rect 5479 2628 5491 2648
rect 5447 2586 5491 2628
rect 6526 2478 6570 2520
rect 6526 2458 6538 2478
rect 6558 2458 6570 2478
rect 6526 2451 6570 2458
rect 6525 2420 6570 2451
rect 6620 2478 6662 2520
rect 6620 2458 6634 2478
rect 6654 2458 6662 2478
rect 6620 2420 6662 2458
rect 6736 2478 6778 2520
rect 6736 2458 6744 2478
rect 6764 2458 6778 2478
rect 6736 2420 6778 2458
rect 6828 2478 6872 2520
rect 6828 2458 6840 2478
rect 6860 2458 6872 2478
rect 6828 2420 6872 2458
rect 6944 2478 6986 2520
rect 6944 2458 6952 2478
rect 6972 2458 6986 2478
rect 6944 2420 6986 2458
rect 7036 2478 7080 2520
rect 7036 2458 7048 2478
rect 7068 2458 7080 2478
rect 7036 2420 7080 2458
rect 7157 2478 7199 2520
rect 7157 2458 7165 2478
rect 7185 2458 7199 2478
rect 7157 2420 7199 2458
rect 7249 2478 7293 2520
rect 7249 2458 7261 2478
rect 7281 2458 7293 2478
rect 7249 2420 7293 2458
rect 9064 2475 9108 2517
rect 9064 2455 9076 2475
rect 9096 2455 9108 2475
rect 9064 2448 9108 2455
rect 9063 2417 9108 2448
rect 9158 2475 9200 2517
rect 9158 2455 9172 2475
rect 9192 2455 9200 2475
rect 9158 2417 9200 2455
rect 9274 2475 9316 2517
rect 9274 2455 9282 2475
rect 9302 2455 9316 2475
rect 9274 2417 9316 2455
rect 9366 2475 9410 2517
rect 9366 2455 9378 2475
rect 9398 2455 9410 2475
rect 9366 2417 9410 2455
rect 9482 2475 9524 2517
rect 9482 2455 9490 2475
rect 9510 2455 9524 2475
rect 9482 2417 9524 2455
rect 9574 2475 9618 2517
rect 9574 2455 9586 2475
rect 9606 2455 9618 2475
rect 9574 2417 9618 2455
rect 9695 2475 9737 2517
rect 9695 2455 9703 2475
rect 9723 2455 9737 2475
rect 9695 2417 9737 2455
rect 9787 2475 9831 2517
rect 9787 2455 9799 2475
rect 9819 2455 9831 2475
rect 9787 2417 9831 2455
rect 774 1967 818 2005
rect 774 1947 786 1967
rect 806 1947 818 1967
rect 774 1905 818 1947
rect 868 1967 910 2005
rect 868 1947 882 1967
rect 902 1947 910 1967
rect 868 1905 910 1947
rect 987 1967 1031 2005
rect 987 1947 999 1967
rect 1019 1947 1031 1967
rect 987 1905 1031 1947
rect 1081 1967 1123 2005
rect 1081 1947 1095 1967
rect 1115 1947 1123 1967
rect 1081 1905 1123 1947
rect 1195 1967 1239 2005
rect 1195 1947 1207 1967
rect 1227 1947 1239 1967
rect 1195 1905 1239 1947
rect 1289 1967 1331 2005
rect 1289 1947 1303 1967
rect 1323 1947 1331 1967
rect 1289 1905 1331 1947
rect 1405 1967 1447 2005
rect 1405 1947 1413 1967
rect 1433 1947 1447 1967
rect 1405 1905 1447 1947
rect 1497 1974 1542 2005
rect 1497 1967 1541 1974
rect 1497 1947 1509 1967
rect 1529 1947 1541 1967
rect 1497 1905 1541 1947
rect 3269 1962 3313 2000
rect 3269 1942 3281 1962
rect 3301 1942 3313 1962
rect 3269 1900 3313 1942
rect 3363 1962 3405 2000
rect 3363 1942 3377 1962
rect 3397 1942 3405 1962
rect 3363 1900 3405 1942
rect 3482 1962 3526 2000
rect 3482 1942 3494 1962
rect 3514 1942 3526 1962
rect 3482 1900 3526 1942
rect 3576 1962 3618 2000
rect 3576 1942 3590 1962
rect 3610 1942 3618 1962
rect 3576 1900 3618 1942
rect 3690 1962 3734 2000
rect 3690 1942 3702 1962
rect 3722 1942 3734 1962
rect 3690 1900 3734 1942
rect 3784 1962 3826 2000
rect 3784 1942 3798 1962
rect 3818 1942 3826 1962
rect 3784 1900 3826 1942
rect 3900 1962 3942 2000
rect 3900 1942 3908 1962
rect 3928 1942 3942 1962
rect 3900 1900 3942 1942
rect 3992 1969 4037 2000
rect 3992 1962 4036 1969
rect 3992 1942 4004 1962
rect 4024 1942 4036 1962
rect 3992 1900 4036 1942
rect 8016 1800 8060 1842
rect 8016 1780 8028 1800
rect 8048 1780 8060 1800
rect 8016 1773 8060 1780
rect 8015 1742 8060 1773
rect 8110 1800 8152 1842
rect 8110 1780 8124 1800
rect 8144 1780 8152 1800
rect 8110 1742 8152 1780
rect 8226 1800 8268 1842
rect 8226 1780 8234 1800
rect 8254 1780 8268 1800
rect 8226 1742 8268 1780
rect 8318 1800 8362 1842
rect 8318 1780 8330 1800
rect 8350 1780 8362 1800
rect 8318 1742 8362 1780
rect 8434 1800 8476 1842
rect 8434 1780 8442 1800
rect 8462 1780 8476 1800
rect 8434 1742 8476 1780
rect 8526 1800 8570 1842
rect 8526 1780 8538 1800
rect 8558 1780 8570 1800
rect 8526 1742 8570 1780
rect 8647 1800 8689 1842
rect 8647 1780 8655 1800
rect 8675 1780 8689 1800
rect 8647 1742 8689 1780
rect 8739 1800 8783 1842
rect 8739 1780 8751 1800
rect 8771 1780 8783 1800
rect 8739 1742 8783 1780
rect 9064 1796 9108 1838
rect 9064 1776 9076 1796
rect 9096 1776 9108 1796
rect 9064 1769 9108 1776
rect 9063 1738 9108 1769
rect 9158 1796 9200 1838
rect 9158 1776 9172 1796
rect 9192 1776 9200 1796
rect 9158 1738 9200 1776
rect 9274 1796 9316 1838
rect 9274 1776 9282 1796
rect 9302 1776 9316 1796
rect 9274 1738 9316 1776
rect 9366 1796 9410 1838
rect 9366 1776 9378 1796
rect 9398 1776 9410 1796
rect 9366 1738 9410 1776
rect 9482 1796 9524 1838
rect 9482 1776 9490 1796
rect 9510 1776 9524 1796
rect 9482 1738 9524 1776
rect 9574 1796 9618 1838
rect 9574 1776 9586 1796
rect 9606 1776 9618 1796
rect 9574 1738 9618 1776
rect 9695 1796 9737 1838
rect 9695 1776 9703 1796
rect 9723 1776 9737 1796
rect 9695 1738 9737 1776
rect 9787 1796 9831 1838
rect 9787 1776 9799 1796
rect 9819 1776 9831 1796
rect 9787 1738 9831 1776
rect 774 1199 818 1237
rect 774 1179 786 1199
rect 806 1179 818 1199
rect 774 1137 818 1179
rect 868 1199 910 1237
rect 868 1179 882 1199
rect 902 1179 910 1199
rect 868 1137 910 1179
rect 987 1199 1031 1237
rect 987 1179 999 1199
rect 1019 1179 1031 1199
rect 987 1137 1031 1179
rect 1081 1199 1123 1237
rect 1081 1179 1095 1199
rect 1115 1179 1123 1199
rect 1081 1137 1123 1179
rect 1195 1199 1239 1237
rect 1195 1179 1207 1199
rect 1227 1179 1239 1199
rect 1195 1137 1239 1179
rect 1289 1199 1331 1237
rect 1289 1179 1303 1199
rect 1323 1179 1331 1199
rect 1289 1137 1331 1179
rect 1405 1199 1447 1237
rect 1405 1179 1413 1199
rect 1433 1179 1447 1199
rect 1405 1137 1447 1179
rect 1497 1206 1542 1237
rect 1497 1199 1541 1206
rect 1497 1179 1509 1199
rect 1529 1179 1541 1199
rect 1497 1137 1541 1179
rect 1822 1195 1866 1233
rect 1822 1175 1834 1195
rect 1854 1175 1866 1195
rect 1822 1133 1866 1175
rect 1916 1195 1958 1233
rect 1916 1175 1930 1195
rect 1950 1175 1958 1195
rect 1916 1133 1958 1175
rect 2035 1195 2079 1233
rect 2035 1175 2047 1195
rect 2067 1175 2079 1195
rect 2035 1133 2079 1175
rect 2129 1195 2171 1233
rect 2129 1175 2143 1195
rect 2163 1175 2171 1195
rect 2129 1133 2171 1175
rect 2243 1195 2287 1233
rect 2243 1175 2255 1195
rect 2275 1175 2287 1195
rect 2243 1133 2287 1175
rect 2337 1195 2379 1233
rect 2337 1175 2351 1195
rect 2371 1175 2379 1195
rect 2337 1133 2379 1175
rect 2453 1195 2495 1233
rect 2453 1175 2461 1195
rect 2481 1175 2495 1195
rect 2453 1133 2495 1175
rect 2545 1202 2590 1233
rect 2545 1195 2589 1202
rect 2545 1175 2557 1195
rect 2577 1175 2589 1195
rect 2545 1133 2589 1175
rect 6569 1033 6613 1075
rect 6569 1013 6581 1033
rect 6601 1013 6613 1033
rect 6569 1006 6613 1013
rect 6568 975 6613 1006
rect 6663 1033 6705 1075
rect 6663 1013 6677 1033
rect 6697 1013 6705 1033
rect 6663 975 6705 1013
rect 6779 1033 6821 1075
rect 6779 1013 6787 1033
rect 6807 1013 6821 1033
rect 6779 975 6821 1013
rect 6871 1033 6915 1075
rect 6871 1013 6883 1033
rect 6903 1013 6915 1033
rect 6871 975 6915 1013
rect 6987 1033 7029 1075
rect 6987 1013 6995 1033
rect 7015 1013 7029 1033
rect 6987 975 7029 1013
rect 7079 1033 7123 1075
rect 7079 1013 7091 1033
rect 7111 1013 7123 1033
rect 7079 975 7123 1013
rect 7200 1033 7242 1075
rect 7200 1013 7208 1033
rect 7228 1013 7242 1033
rect 7200 975 7242 1013
rect 7292 1033 7336 1075
rect 7292 1013 7304 1033
rect 7324 1013 7336 1033
rect 7292 975 7336 1013
rect 9064 1028 9108 1070
rect 9064 1008 9076 1028
rect 9096 1008 9108 1028
rect 9064 1001 9108 1008
rect 9063 970 9108 1001
rect 9158 1028 9200 1070
rect 9158 1008 9172 1028
rect 9192 1008 9200 1028
rect 9158 970 9200 1008
rect 9274 1028 9316 1070
rect 9274 1008 9282 1028
rect 9302 1008 9316 1028
rect 9274 970 9316 1008
rect 9366 1028 9410 1070
rect 9366 1008 9378 1028
rect 9398 1008 9410 1028
rect 9366 970 9410 1008
rect 9482 1028 9524 1070
rect 9482 1008 9490 1028
rect 9510 1008 9524 1028
rect 9482 970 9524 1008
rect 9574 1028 9618 1070
rect 9574 1008 9586 1028
rect 9606 1008 9618 1028
rect 9574 970 9618 1008
rect 9695 1028 9737 1070
rect 9695 1008 9703 1028
rect 9723 1008 9737 1028
rect 9695 970 9737 1008
rect 9787 1028 9831 1070
rect 9787 1008 9799 1028
rect 9819 1008 9831 1028
rect 9787 970 9831 1008
rect 774 520 818 558
rect 774 500 786 520
rect 806 500 818 520
rect 774 458 818 500
rect 868 520 910 558
rect 868 500 882 520
rect 902 500 910 520
rect 868 458 910 500
rect 987 520 1031 558
rect 987 500 999 520
rect 1019 500 1031 520
rect 987 458 1031 500
rect 1081 520 1123 558
rect 1081 500 1095 520
rect 1115 500 1123 520
rect 1081 458 1123 500
rect 1195 520 1239 558
rect 1195 500 1207 520
rect 1227 500 1239 520
rect 1195 458 1239 500
rect 1289 520 1331 558
rect 1289 500 1303 520
rect 1323 500 1331 520
rect 1289 458 1331 500
rect 1405 520 1447 558
rect 1405 500 1413 520
rect 1433 500 1447 520
rect 1405 458 1447 500
rect 1497 527 1542 558
rect 1497 520 1541 527
rect 1497 500 1509 520
rect 1529 500 1541 520
rect 1497 458 1541 500
rect 8016 353 8060 395
rect 8016 333 8028 353
rect 8048 333 8060 353
rect 8016 326 8060 333
rect 8015 295 8060 326
rect 8110 353 8152 395
rect 8110 333 8124 353
rect 8144 333 8152 353
rect 8110 295 8152 333
rect 8226 353 8268 395
rect 8226 333 8234 353
rect 8254 333 8268 353
rect 8226 295 8268 333
rect 8318 353 8362 395
rect 8318 333 8330 353
rect 8350 333 8362 353
rect 8318 295 8362 333
rect 8434 353 8476 395
rect 8434 333 8442 353
rect 8462 333 8476 353
rect 8434 295 8476 333
rect 8526 353 8570 395
rect 8526 333 8538 353
rect 8558 333 8570 353
rect 8526 295 8570 333
rect 8647 353 8689 395
rect 8647 333 8655 353
rect 8675 333 8689 353
rect 8647 295 8689 333
rect 8739 353 8783 395
rect 8739 333 8751 353
rect 8771 333 8783 353
rect 8739 295 8783 333
rect 9064 349 9108 391
rect 9064 329 9076 349
rect 9096 329 9108 349
rect 9064 322 9108 329
rect 9063 291 9108 322
rect 9158 349 9200 391
rect 9158 329 9172 349
rect 9192 329 9200 349
rect 9158 291 9200 329
rect 9274 349 9316 391
rect 9274 329 9282 349
rect 9302 329 9316 349
rect 9274 291 9316 329
rect 9366 349 9410 391
rect 9366 329 9378 349
rect 9398 329 9410 349
rect 9366 291 9410 329
rect 9482 349 9524 391
rect 9482 329 9490 349
rect 9510 329 9524 349
rect 9482 291 9524 329
rect 9574 349 9618 391
rect 9574 329 9586 349
rect 9606 329 9618 349
rect 9574 291 9618 329
rect 9695 349 9737 391
rect 9695 329 9703 349
rect 9723 329 9737 349
rect 9695 291 9737 329
rect 9787 349 9831 391
rect 9787 329 9799 349
rect 9819 329 9831 349
rect 9787 291 9831 329
<< ndiffc >>
rect 461 11775 479 11793
rect 463 11676 481 11694
rect 461 11519 479 11537
rect 9071 11579 9091 11599
rect 9174 11575 9194 11595
rect 9282 11575 9302 11595
rect 9385 11579 9405 11599
rect 9490 11575 9510 11595
rect 9593 11579 9613 11599
rect 9703 11575 9723 11595
rect 9806 11579 9826 11599
rect 10126 11584 10144 11602
rect 781 11452 801 11472
rect 884 11456 904 11476
rect 994 11452 1014 11472
rect 1097 11456 1117 11476
rect 1202 11452 1222 11472
rect 1305 11456 1325 11476
rect 1413 11456 1433 11476
rect 1516 11452 1536 11472
rect 1829 11448 1849 11468
rect 463 11420 481 11438
rect 1932 11452 1952 11472
rect 2042 11448 2062 11468
rect 2145 11452 2165 11472
rect 2250 11448 2270 11468
rect 2353 11452 2373 11472
rect 2461 11452 2481 11472
rect 2564 11448 2584 11468
rect 10128 11485 10146 11503
rect 10126 11329 10144 11347
rect 10128 11230 10146 11248
rect 461 11124 479 11142
rect 463 11025 481 11043
rect 461 10869 479 10887
rect 8023 10904 8043 10924
rect 8126 10900 8146 10920
rect 8234 10900 8254 10920
rect 8337 10904 8357 10924
rect 8442 10900 8462 10920
rect 8545 10904 8565 10924
rect 8655 10900 8675 10920
rect 10126 10934 10144 10952
rect 8758 10904 8778 10924
rect 9071 10900 9091 10920
rect 463 10770 481 10788
rect 781 10773 801 10793
rect 884 10777 904 10797
rect 994 10773 1014 10793
rect 1097 10777 1117 10797
rect 1202 10773 1222 10793
rect 1305 10777 1325 10797
rect 1413 10777 1433 10797
rect 9174 10896 9194 10916
rect 9282 10896 9302 10916
rect 9385 10900 9405 10920
rect 9490 10896 9510 10916
rect 9593 10900 9613 10920
rect 9703 10896 9723 10916
rect 9806 10900 9826 10920
rect 1516 10773 1536 10793
rect 3276 10768 3296 10788
rect 3379 10772 3399 10792
rect 3489 10768 3509 10788
rect 3592 10772 3612 10792
rect 3697 10768 3717 10788
rect 3800 10772 3820 10792
rect 3908 10772 3928 10792
rect 4011 10768 4031 10788
rect 10128 10835 10146 10853
rect 10126 10678 10144 10696
rect 10128 10579 10146 10597
rect 461 10328 479 10346
rect 463 10229 481 10247
rect 461 10072 479 10090
rect 6576 10137 6596 10157
rect 6679 10133 6699 10153
rect 6787 10133 6807 10153
rect 6890 10137 6910 10157
rect 6995 10133 7015 10153
rect 7098 10137 7118 10157
rect 7208 10133 7228 10153
rect 7311 10137 7331 10157
rect 9071 10132 9091 10152
rect 781 10005 801 10025
rect 884 10009 904 10029
rect 994 10005 1014 10025
rect 1097 10009 1117 10029
rect 1202 10005 1222 10025
rect 1305 10009 1325 10029
rect 1413 10009 1433 10029
rect 9174 10128 9194 10148
rect 9282 10128 9302 10148
rect 9385 10132 9405 10152
rect 9490 10128 9510 10148
rect 9593 10132 9613 10152
rect 9703 10128 9723 10148
rect 9806 10132 9826 10152
rect 10126 10137 10144 10155
rect 1516 10005 1536 10025
rect 1829 10001 1849 10021
rect 463 9973 481 9991
rect 1932 10005 1952 10025
rect 2042 10001 2062 10021
rect 2145 10005 2165 10025
rect 2250 10001 2270 10021
rect 2353 10005 2373 10025
rect 2461 10005 2481 10025
rect 2564 10001 2584 10021
rect 10128 10038 10146 10056
rect 10126 9882 10144 9900
rect 10128 9783 10146 9801
rect 461 9677 479 9695
rect 463 9578 481 9596
rect 461 9422 479 9440
rect 8023 9457 8043 9477
rect 8126 9453 8146 9473
rect 8234 9453 8254 9473
rect 8337 9457 8357 9477
rect 8442 9453 8462 9473
rect 8545 9457 8565 9477
rect 8655 9453 8675 9473
rect 10126 9487 10144 9505
rect 8758 9457 8778 9477
rect 9071 9453 9091 9473
rect 463 9323 481 9341
rect 781 9326 801 9346
rect 884 9330 904 9350
rect 994 9326 1014 9346
rect 1097 9330 1117 9350
rect 1202 9326 1222 9346
rect 1305 9330 1325 9350
rect 1413 9330 1433 9350
rect 9174 9449 9194 9469
rect 9282 9449 9302 9469
rect 9385 9453 9405 9473
rect 9490 9449 9510 9469
rect 9593 9453 9613 9473
rect 9703 9449 9723 9469
rect 9806 9453 9826 9473
rect 1516 9326 1536 9346
rect 3319 9323 3339 9343
rect 3422 9327 3442 9347
rect 3532 9323 3552 9343
rect 3635 9327 3655 9347
rect 3740 9323 3760 9343
rect 3843 9327 3863 9347
rect 3951 9327 3971 9347
rect 4054 9323 4074 9343
rect 10128 9388 10146 9406
rect 10126 9231 10144 9249
rect 10128 9132 10146 9150
rect 462 8808 480 8826
rect 464 8709 482 8727
rect 462 8552 480 8570
rect 6534 8615 6554 8635
rect 6637 8611 6657 8631
rect 6745 8611 6765 8631
rect 6848 8615 6868 8635
rect 6953 8611 6973 8631
rect 7056 8615 7076 8635
rect 7166 8611 7186 8631
rect 7269 8615 7289 8635
rect 9072 8612 9092 8632
rect 782 8485 802 8505
rect 885 8489 905 8509
rect 995 8485 1015 8505
rect 1098 8489 1118 8509
rect 1203 8485 1223 8505
rect 1306 8489 1326 8509
rect 1414 8489 1434 8509
rect 9175 8608 9195 8628
rect 9283 8608 9303 8628
rect 9386 8612 9406 8632
rect 9491 8608 9511 8628
rect 9594 8612 9614 8632
rect 9704 8608 9724 8628
rect 9807 8612 9827 8632
rect 10127 8617 10145 8635
rect 1517 8485 1537 8505
rect 1830 8481 1850 8501
rect 464 8453 482 8471
rect 1933 8485 1953 8505
rect 2043 8481 2063 8501
rect 2146 8485 2166 8505
rect 2251 8481 2271 8501
rect 2354 8485 2374 8505
rect 2462 8485 2482 8505
rect 2565 8481 2585 8501
rect 10129 8518 10147 8536
rect 10127 8362 10145 8380
rect 10129 8263 10147 8281
rect 462 8157 480 8175
rect 464 8058 482 8076
rect 462 7902 480 7920
rect 8024 7937 8044 7957
rect 8127 7933 8147 7953
rect 8235 7933 8255 7953
rect 8338 7937 8358 7957
rect 8443 7933 8463 7953
rect 8546 7937 8566 7957
rect 8656 7933 8676 7953
rect 10127 7967 10145 7985
rect 8759 7937 8779 7957
rect 9072 7933 9092 7953
rect 464 7803 482 7821
rect 782 7806 802 7826
rect 885 7810 905 7830
rect 995 7806 1015 7826
rect 1098 7810 1118 7830
rect 1203 7806 1223 7826
rect 1306 7810 1326 7830
rect 1414 7810 1434 7830
rect 9175 7929 9195 7949
rect 9283 7929 9303 7949
rect 9386 7933 9406 7953
rect 9491 7929 9511 7949
rect 9594 7933 9614 7953
rect 9704 7929 9724 7949
rect 9807 7933 9827 7953
rect 1517 7806 1537 7826
rect 3277 7801 3297 7821
rect 3380 7805 3400 7825
rect 3490 7801 3510 7821
rect 3593 7805 3613 7825
rect 3698 7801 3718 7821
rect 3801 7805 3821 7825
rect 3909 7805 3929 7825
rect 4012 7801 4032 7821
rect 10129 7868 10147 7886
rect 10127 7711 10145 7729
rect 10129 7612 10147 7630
rect 462 7361 480 7379
rect 464 7262 482 7280
rect 462 7105 480 7123
rect 6577 7170 6597 7190
rect 6680 7166 6700 7186
rect 6788 7166 6808 7186
rect 6891 7170 6911 7190
rect 6996 7166 7016 7186
rect 7099 7170 7119 7190
rect 7209 7166 7229 7186
rect 7312 7170 7332 7190
rect 9072 7165 9092 7185
rect 782 7038 802 7058
rect 885 7042 905 7062
rect 995 7038 1015 7058
rect 1098 7042 1118 7062
rect 1203 7038 1223 7058
rect 1306 7042 1326 7062
rect 1414 7042 1434 7062
rect 9175 7161 9195 7181
rect 9283 7161 9303 7181
rect 9386 7165 9406 7185
rect 9491 7161 9511 7181
rect 9594 7165 9614 7185
rect 9704 7161 9724 7181
rect 9807 7165 9827 7185
rect 10127 7170 10145 7188
rect 1517 7038 1537 7058
rect 1830 7034 1850 7054
rect 464 7006 482 7024
rect 1933 7038 1953 7058
rect 2043 7034 2063 7054
rect 2146 7038 2166 7058
rect 2251 7034 2271 7054
rect 2354 7038 2374 7058
rect 2462 7038 2482 7058
rect 2565 7034 2585 7054
rect 10129 7071 10147 7089
rect 10127 6915 10145 6933
rect 10129 6816 10147 6834
rect 462 6710 480 6728
rect 464 6611 482 6629
rect 462 6455 480 6473
rect 8024 6490 8044 6510
rect 8127 6486 8147 6506
rect 8235 6486 8255 6506
rect 8338 6490 8358 6510
rect 8443 6486 8463 6506
rect 8546 6490 8566 6510
rect 8656 6486 8676 6506
rect 10127 6520 10145 6538
rect 8759 6490 8779 6510
rect 9072 6486 9092 6506
rect 464 6356 482 6374
rect 782 6359 802 6379
rect 885 6363 905 6383
rect 995 6359 1015 6379
rect 1098 6363 1118 6383
rect 1203 6359 1223 6379
rect 1306 6363 1326 6383
rect 1414 6363 1434 6383
rect 9175 6482 9195 6502
rect 9283 6482 9303 6502
rect 9386 6486 9406 6506
rect 9491 6482 9511 6502
rect 9594 6486 9614 6506
rect 9704 6482 9724 6502
rect 9807 6486 9827 6506
rect 1517 6359 1537 6379
rect 4385 6350 4405 6370
rect 4488 6354 4508 6374
rect 4598 6350 4618 6370
rect 4701 6354 4721 6374
rect 4806 6350 4826 6370
rect 4909 6354 4929 6374
rect 5017 6354 5037 6374
rect 5120 6350 5140 6370
rect 10129 6421 10147 6439
rect 10127 6264 10145 6282
rect 10129 6165 10147 6183
rect 459 5767 477 5785
rect 461 5668 479 5686
rect 459 5511 477 5529
rect 5466 5580 5486 5600
rect 5569 5576 5589 5596
rect 5677 5576 5697 5596
rect 5780 5580 5800 5600
rect 5885 5576 5905 5596
rect 5988 5580 6008 5600
rect 6098 5576 6118 5596
rect 6201 5580 6221 5600
rect 9069 5571 9089 5591
rect 779 5444 799 5464
rect 882 5448 902 5468
rect 992 5444 1012 5464
rect 1095 5448 1115 5468
rect 1200 5444 1220 5464
rect 1303 5448 1323 5468
rect 1411 5448 1431 5468
rect 9172 5567 9192 5587
rect 9280 5567 9300 5587
rect 9383 5571 9403 5591
rect 9488 5567 9508 5587
rect 9591 5571 9611 5591
rect 9701 5567 9721 5587
rect 9804 5571 9824 5591
rect 10124 5576 10142 5594
rect 1514 5444 1534 5464
rect 1827 5440 1847 5460
rect 461 5412 479 5430
rect 1930 5444 1950 5464
rect 2040 5440 2060 5460
rect 2143 5444 2163 5464
rect 2248 5440 2268 5460
rect 2351 5444 2371 5464
rect 2459 5444 2479 5464
rect 2562 5440 2582 5460
rect 10126 5477 10144 5495
rect 10124 5321 10142 5339
rect 10126 5222 10144 5240
rect 459 5116 477 5134
rect 461 5017 479 5035
rect 459 4861 477 4879
rect 8021 4896 8041 4916
rect 8124 4892 8144 4912
rect 8232 4892 8252 4912
rect 8335 4896 8355 4916
rect 8440 4892 8460 4912
rect 8543 4896 8563 4916
rect 8653 4892 8673 4912
rect 10124 4926 10142 4944
rect 8756 4896 8776 4916
rect 9069 4892 9089 4912
rect 461 4762 479 4780
rect 779 4765 799 4785
rect 882 4769 902 4789
rect 992 4765 1012 4785
rect 1095 4769 1115 4789
rect 1200 4765 1220 4785
rect 1303 4769 1323 4789
rect 1411 4769 1431 4789
rect 9172 4888 9192 4908
rect 9280 4888 9300 4908
rect 9383 4892 9403 4912
rect 9488 4888 9508 4908
rect 9591 4892 9611 4912
rect 9701 4888 9721 4908
rect 9804 4892 9824 4912
rect 1514 4765 1534 4785
rect 3274 4760 3294 4780
rect 3377 4764 3397 4784
rect 3487 4760 3507 4780
rect 3590 4764 3610 4784
rect 3695 4760 3715 4780
rect 3798 4764 3818 4784
rect 3906 4764 3926 4784
rect 4009 4760 4029 4780
rect 10126 4827 10144 4845
rect 10124 4670 10142 4688
rect 10126 4571 10144 4589
rect 459 4320 477 4338
rect 461 4221 479 4239
rect 459 4064 477 4082
rect 6574 4129 6594 4149
rect 6677 4125 6697 4145
rect 6785 4125 6805 4145
rect 6888 4129 6908 4149
rect 6993 4125 7013 4145
rect 7096 4129 7116 4149
rect 7206 4125 7226 4145
rect 7309 4129 7329 4149
rect 9069 4124 9089 4144
rect 779 3997 799 4017
rect 882 4001 902 4021
rect 992 3997 1012 4017
rect 1095 4001 1115 4021
rect 1200 3997 1220 4017
rect 1303 4001 1323 4021
rect 1411 4001 1431 4021
rect 9172 4120 9192 4140
rect 9280 4120 9300 4140
rect 9383 4124 9403 4144
rect 9488 4120 9508 4140
rect 9591 4124 9611 4144
rect 9701 4120 9721 4140
rect 9804 4124 9824 4144
rect 10124 4129 10142 4147
rect 1514 3997 1534 4017
rect 1827 3993 1847 4013
rect 461 3965 479 3983
rect 1930 3997 1950 4017
rect 2040 3993 2060 4013
rect 2143 3997 2163 4017
rect 2248 3993 2268 4013
rect 2351 3997 2371 4017
rect 2459 3997 2479 4017
rect 2562 3993 2582 4013
rect 10126 4030 10144 4048
rect 10124 3874 10142 3892
rect 10126 3775 10144 3793
rect 459 3669 477 3687
rect 461 3570 479 3588
rect 459 3414 477 3432
rect 8021 3449 8041 3469
rect 8124 3445 8144 3465
rect 8232 3445 8252 3465
rect 8335 3449 8355 3469
rect 8440 3445 8460 3465
rect 8543 3449 8563 3469
rect 8653 3445 8673 3465
rect 10124 3479 10142 3497
rect 8756 3449 8776 3469
rect 9069 3445 9089 3465
rect 461 3315 479 3333
rect 779 3318 799 3338
rect 882 3322 902 3342
rect 992 3318 1012 3338
rect 1095 3322 1115 3342
rect 1200 3318 1220 3338
rect 1303 3322 1323 3342
rect 1411 3322 1431 3342
rect 9172 3441 9192 3461
rect 9280 3441 9300 3461
rect 9383 3445 9403 3465
rect 9488 3441 9508 3461
rect 9591 3445 9611 3465
rect 9701 3441 9721 3461
rect 9804 3445 9824 3465
rect 1514 3318 1534 3338
rect 3317 3315 3337 3335
rect 3420 3319 3440 3339
rect 3530 3315 3550 3335
rect 3633 3319 3653 3339
rect 3738 3315 3758 3335
rect 3841 3319 3861 3339
rect 3949 3319 3969 3339
rect 4052 3315 4072 3335
rect 10126 3380 10144 3398
rect 10124 3223 10142 3241
rect 10126 3124 10144 3142
rect 460 2800 478 2818
rect 462 2701 480 2719
rect 460 2544 478 2562
rect 6532 2607 6552 2627
rect 6635 2603 6655 2623
rect 6743 2603 6763 2623
rect 6846 2607 6866 2627
rect 6951 2603 6971 2623
rect 7054 2607 7074 2627
rect 7164 2603 7184 2623
rect 7267 2607 7287 2627
rect 9070 2604 9090 2624
rect 780 2477 800 2497
rect 883 2481 903 2501
rect 993 2477 1013 2497
rect 1096 2481 1116 2501
rect 1201 2477 1221 2497
rect 1304 2481 1324 2501
rect 1412 2481 1432 2501
rect 9173 2600 9193 2620
rect 9281 2600 9301 2620
rect 9384 2604 9404 2624
rect 9489 2600 9509 2620
rect 9592 2604 9612 2624
rect 9702 2600 9722 2620
rect 9805 2604 9825 2624
rect 10125 2609 10143 2627
rect 1515 2477 1535 2497
rect 1828 2473 1848 2493
rect 462 2445 480 2463
rect 1931 2477 1951 2497
rect 2041 2473 2061 2493
rect 2144 2477 2164 2497
rect 2249 2473 2269 2493
rect 2352 2477 2372 2497
rect 2460 2477 2480 2497
rect 2563 2473 2583 2493
rect 4730 2479 4750 2499
rect 4833 2483 4853 2503
rect 4943 2479 4963 2499
rect 5046 2483 5066 2503
rect 5151 2479 5171 2499
rect 5254 2483 5274 2503
rect 5362 2483 5382 2503
rect 5465 2479 5485 2499
rect 10127 2510 10145 2528
rect 10125 2354 10143 2372
rect 10127 2255 10145 2273
rect 460 2149 478 2167
rect 462 2050 480 2068
rect 460 1894 478 1912
rect 8022 1929 8042 1949
rect 8125 1925 8145 1945
rect 8233 1925 8253 1945
rect 8336 1929 8356 1949
rect 8441 1925 8461 1945
rect 8544 1929 8564 1949
rect 8654 1925 8674 1945
rect 10125 1959 10143 1977
rect 8757 1929 8777 1949
rect 9070 1925 9090 1945
rect 462 1795 480 1813
rect 780 1798 800 1818
rect 883 1802 903 1822
rect 993 1798 1013 1818
rect 1096 1802 1116 1822
rect 1201 1798 1221 1818
rect 1304 1802 1324 1822
rect 1412 1802 1432 1822
rect 9173 1921 9193 1941
rect 9281 1921 9301 1941
rect 9384 1925 9404 1945
rect 9489 1921 9509 1941
rect 9592 1925 9612 1945
rect 9702 1921 9722 1941
rect 9805 1925 9825 1945
rect 1515 1798 1535 1818
rect 3275 1793 3295 1813
rect 3378 1797 3398 1817
rect 3488 1793 3508 1813
rect 3591 1797 3611 1817
rect 3696 1793 3716 1813
rect 3799 1797 3819 1817
rect 3907 1797 3927 1817
rect 4010 1793 4030 1813
rect 10127 1860 10145 1878
rect 10125 1703 10143 1721
rect 10127 1604 10145 1622
rect 460 1353 478 1371
rect 462 1254 480 1272
rect 460 1097 478 1115
rect 6575 1162 6595 1182
rect 6678 1158 6698 1178
rect 6786 1158 6806 1178
rect 6889 1162 6909 1182
rect 6994 1158 7014 1178
rect 7097 1162 7117 1182
rect 7207 1158 7227 1178
rect 7310 1162 7330 1182
rect 9070 1157 9090 1177
rect 780 1030 800 1050
rect 883 1034 903 1054
rect 993 1030 1013 1050
rect 1096 1034 1116 1054
rect 1201 1030 1221 1050
rect 1304 1034 1324 1054
rect 1412 1034 1432 1054
rect 9173 1153 9193 1173
rect 9281 1153 9301 1173
rect 9384 1157 9404 1177
rect 9489 1153 9509 1173
rect 9592 1157 9612 1177
rect 9702 1153 9722 1173
rect 9805 1157 9825 1177
rect 10125 1162 10143 1180
rect 1515 1030 1535 1050
rect 1828 1026 1848 1046
rect 462 998 480 1016
rect 1931 1030 1951 1050
rect 2041 1026 2061 1046
rect 2144 1030 2164 1050
rect 2249 1026 2269 1046
rect 2352 1030 2372 1050
rect 2460 1030 2480 1050
rect 2563 1026 2583 1046
rect 10127 1063 10145 1081
rect 10125 907 10143 925
rect 10127 808 10145 826
rect 460 702 478 720
rect 462 603 480 621
rect 460 447 478 465
rect 8022 482 8042 502
rect 8125 478 8145 498
rect 8233 478 8253 498
rect 8336 482 8356 502
rect 8441 478 8461 498
rect 8544 482 8564 502
rect 8654 478 8674 498
rect 10125 512 10143 530
rect 8757 482 8777 502
rect 9070 478 9090 498
rect 9173 474 9193 494
rect 9281 474 9301 494
rect 9384 478 9404 498
rect 9489 474 9509 494
rect 9592 478 9612 498
rect 9702 474 9722 494
rect 9805 478 9825 498
rect 462 348 480 366
rect 780 351 800 371
rect 883 355 903 375
rect 993 351 1013 371
rect 1096 355 1116 375
rect 1201 351 1221 371
rect 1304 355 1324 375
rect 1412 355 1432 375
rect 1515 351 1535 371
rect 10127 413 10145 431
rect 10125 256 10143 274
rect 10127 157 10145 175
<< pdiffc >>
rect 787 11601 807 11621
rect 883 11601 903 11621
rect 1000 11601 1020 11621
rect 1096 11601 1116 11621
rect 1208 11601 1228 11621
rect 1304 11601 1324 11621
rect 1414 11601 1434 11621
rect 1510 11601 1530 11621
rect 1835 11597 1855 11617
rect 1931 11597 1951 11617
rect 2048 11597 2068 11617
rect 2144 11597 2164 11617
rect 2256 11597 2276 11617
rect 2352 11597 2372 11617
rect 2462 11597 2482 11617
rect 2558 11597 2578 11617
rect 9077 11430 9097 11450
rect 9173 11430 9193 11450
rect 9283 11430 9303 11450
rect 9379 11430 9399 11450
rect 9491 11430 9511 11450
rect 9587 11430 9607 11450
rect 9704 11430 9724 11450
rect 9800 11430 9820 11450
rect 787 10922 807 10942
rect 883 10922 903 10942
rect 1000 10922 1020 10942
rect 1096 10922 1116 10942
rect 1208 10922 1228 10942
rect 1304 10922 1324 10942
rect 1414 10922 1434 10942
rect 1510 10922 1530 10942
rect 3282 10917 3302 10937
rect 3378 10917 3398 10937
rect 3495 10917 3515 10937
rect 3591 10917 3611 10937
rect 3703 10917 3723 10937
rect 3799 10917 3819 10937
rect 3909 10917 3929 10937
rect 4005 10917 4025 10937
rect 8029 10755 8049 10775
rect 8125 10755 8145 10775
rect 8235 10755 8255 10775
rect 8331 10755 8351 10775
rect 8443 10755 8463 10775
rect 8539 10755 8559 10775
rect 8656 10755 8676 10775
rect 8752 10755 8772 10775
rect 9077 10751 9097 10771
rect 9173 10751 9193 10771
rect 9283 10751 9303 10771
rect 9379 10751 9399 10771
rect 9491 10751 9511 10771
rect 9587 10751 9607 10771
rect 9704 10751 9724 10771
rect 9800 10751 9820 10771
rect 787 10154 807 10174
rect 883 10154 903 10174
rect 1000 10154 1020 10174
rect 1096 10154 1116 10174
rect 1208 10154 1228 10174
rect 1304 10154 1324 10174
rect 1414 10154 1434 10174
rect 1510 10154 1530 10174
rect 1835 10150 1855 10170
rect 1931 10150 1951 10170
rect 2048 10150 2068 10170
rect 2144 10150 2164 10170
rect 2256 10150 2276 10170
rect 2352 10150 2372 10170
rect 2462 10150 2482 10170
rect 2558 10150 2578 10170
rect 6582 9988 6602 10008
rect 6678 9988 6698 10008
rect 6788 9988 6808 10008
rect 6884 9988 6904 10008
rect 6996 9988 7016 10008
rect 7092 9988 7112 10008
rect 7209 9988 7229 10008
rect 7305 9988 7325 10008
rect 9077 9983 9097 10003
rect 9173 9983 9193 10003
rect 9283 9983 9303 10003
rect 9379 9983 9399 10003
rect 9491 9983 9511 10003
rect 9587 9983 9607 10003
rect 9704 9983 9724 10003
rect 9800 9983 9820 10003
rect 787 9475 807 9495
rect 883 9475 903 9495
rect 1000 9475 1020 9495
rect 1096 9475 1116 9495
rect 1208 9475 1228 9495
rect 1304 9475 1324 9495
rect 1414 9475 1434 9495
rect 1510 9475 1530 9495
rect 3325 9472 3345 9492
rect 3421 9472 3441 9492
rect 3538 9472 3558 9492
rect 3634 9472 3654 9492
rect 3746 9472 3766 9492
rect 3842 9472 3862 9492
rect 3952 9472 3972 9492
rect 4048 9472 4068 9492
rect 8029 9308 8049 9328
rect 8125 9308 8145 9328
rect 8235 9308 8255 9328
rect 8331 9308 8351 9328
rect 8443 9308 8463 9328
rect 8539 9308 8559 9328
rect 8656 9308 8676 9328
rect 8752 9308 8772 9328
rect 9077 9304 9097 9324
rect 9173 9304 9193 9324
rect 9283 9304 9303 9324
rect 9379 9304 9399 9324
rect 9491 9304 9511 9324
rect 9587 9304 9607 9324
rect 9704 9304 9724 9324
rect 9800 9304 9820 9324
rect 788 8634 808 8654
rect 884 8634 904 8654
rect 1001 8634 1021 8654
rect 1097 8634 1117 8654
rect 1209 8634 1229 8654
rect 1305 8634 1325 8654
rect 1415 8634 1435 8654
rect 1511 8634 1531 8654
rect 1836 8630 1856 8650
rect 1932 8630 1952 8650
rect 2049 8630 2069 8650
rect 2145 8630 2165 8650
rect 2257 8630 2277 8650
rect 2353 8630 2373 8650
rect 2463 8630 2483 8650
rect 2559 8630 2579 8650
rect 6540 8466 6560 8486
rect 6636 8466 6656 8486
rect 6746 8466 6766 8486
rect 6842 8466 6862 8486
rect 6954 8466 6974 8486
rect 7050 8466 7070 8486
rect 7167 8466 7187 8486
rect 7263 8466 7283 8486
rect 9078 8463 9098 8483
rect 9174 8463 9194 8483
rect 9284 8463 9304 8483
rect 9380 8463 9400 8483
rect 9492 8463 9512 8483
rect 9588 8463 9608 8483
rect 9705 8463 9725 8483
rect 9801 8463 9821 8483
rect 788 7955 808 7975
rect 884 7955 904 7975
rect 1001 7955 1021 7975
rect 1097 7955 1117 7975
rect 1209 7955 1229 7975
rect 1305 7955 1325 7975
rect 1415 7955 1435 7975
rect 1511 7955 1531 7975
rect 3283 7950 3303 7970
rect 3379 7950 3399 7970
rect 3496 7950 3516 7970
rect 3592 7950 3612 7970
rect 3704 7950 3724 7970
rect 3800 7950 3820 7970
rect 3910 7950 3930 7970
rect 4006 7950 4026 7970
rect 8030 7788 8050 7808
rect 8126 7788 8146 7808
rect 8236 7788 8256 7808
rect 8332 7788 8352 7808
rect 8444 7788 8464 7808
rect 8540 7788 8560 7808
rect 8657 7788 8677 7808
rect 8753 7788 8773 7808
rect 9078 7784 9098 7804
rect 9174 7784 9194 7804
rect 9284 7784 9304 7804
rect 9380 7784 9400 7804
rect 9492 7784 9512 7804
rect 9588 7784 9608 7804
rect 9705 7784 9725 7804
rect 9801 7784 9821 7804
rect 788 7187 808 7207
rect 884 7187 904 7207
rect 1001 7187 1021 7207
rect 1097 7187 1117 7207
rect 1209 7187 1229 7207
rect 1305 7187 1325 7207
rect 1415 7187 1435 7207
rect 1511 7187 1531 7207
rect 1836 7183 1856 7203
rect 1932 7183 1952 7203
rect 2049 7183 2069 7203
rect 2145 7183 2165 7203
rect 2257 7183 2277 7203
rect 2353 7183 2373 7203
rect 2463 7183 2483 7203
rect 2559 7183 2579 7203
rect 6583 7021 6603 7041
rect 6679 7021 6699 7041
rect 6789 7021 6809 7041
rect 6885 7021 6905 7041
rect 6997 7021 7017 7041
rect 7093 7021 7113 7041
rect 7210 7021 7230 7041
rect 7306 7021 7326 7041
rect 9078 7016 9098 7036
rect 9174 7016 9194 7036
rect 9284 7016 9304 7036
rect 9380 7016 9400 7036
rect 9492 7016 9512 7036
rect 9588 7016 9608 7036
rect 9705 7016 9725 7036
rect 9801 7016 9821 7036
rect 788 6508 808 6528
rect 884 6508 904 6528
rect 1001 6508 1021 6528
rect 1097 6508 1117 6528
rect 1209 6508 1229 6528
rect 1305 6508 1325 6528
rect 1415 6508 1435 6528
rect 1511 6508 1531 6528
rect 4391 6499 4411 6519
rect 4487 6499 4507 6519
rect 4604 6499 4624 6519
rect 4700 6499 4720 6519
rect 4812 6499 4832 6519
rect 4908 6499 4928 6519
rect 5018 6499 5038 6519
rect 5114 6499 5134 6519
rect 8030 6341 8050 6361
rect 8126 6341 8146 6361
rect 8236 6341 8256 6361
rect 8332 6341 8352 6361
rect 8444 6341 8464 6361
rect 8540 6341 8560 6361
rect 8657 6341 8677 6361
rect 8753 6341 8773 6361
rect 9078 6337 9098 6357
rect 9174 6337 9194 6357
rect 9284 6337 9304 6357
rect 9380 6337 9400 6357
rect 9492 6337 9512 6357
rect 9588 6337 9608 6357
rect 9705 6337 9725 6357
rect 9801 6337 9821 6357
rect 785 5593 805 5613
rect 881 5593 901 5613
rect 998 5593 1018 5613
rect 1094 5593 1114 5613
rect 1206 5593 1226 5613
rect 1302 5593 1322 5613
rect 1412 5593 1432 5613
rect 1508 5593 1528 5613
rect 1833 5589 1853 5609
rect 1929 5589 1949 5609
rect 2046 5589 2066 5609
rect 2142 5589 2162 5609
rect 2254 5589 2274 5609
rect 2350 5589 2370 5609
rect 2460 5589 2480 5609
rect 2556 5589 2576 5609
rect 5472 5431 5492 5451
rect 5568 5431 5588 5451
rect 5678 5431 5698 5451
rect 5774 5431 5794 5451
rect 5886 5431 5906 5451
rect 5982 5431 6002 5451
rect 6099 5431 6119 5451
rect 6195 5431 6215 5451
rect 9075 5422 9095 5442
rect 9171 5422 9191 5442
rect 9281 5422 9301 5442
rect 9377 5422 9397 5442
rect 9489 5422 9509 5442
rect 9585 5422 9605 5442
rect 9702 5422 9722 5442
rect 9798 5422 9818 5442
rect 785 4914 805 4934
rect 881 4914 901 4934
rect 998 4914 1018 4934
rect 1094 4914 1114 4934
rect 1206 4914 1226 4934
rect 1302 4914 1322 4934
rect 1412 4914 1432 4934
rect 1508 4914 1528 4934
rect 3280 4909 3300 4929
rect 3376 4909 3396 4929
rect 3493 4909 3513 4929
rect 3589 4909 3609 4929
rect 3701 4909 3721 4929
rect 3797 4909 3817 4929
rect 3907 4909 3927 4929
rect 4003 4909 4023 4929
rect 8027 4747 8047 4767
rect 8123 4747 8143 4767
rect 8233 4747 8253 4767
rect 8329 4747 8349 4767
rect 8441 4747 8461 4767
rect 8537 4747 8557 4767
rect 8654 4747 8674 4767
rect 8750 4747 8770 4767
rect 9075 4743 9095 4763
rect 9171 4743 9191 4763
rect 9281 4743 9301 4763
rect 9377 4743 9397 4763
rect 9489 4743 9509 4763
rect 9585 4743 9605 4763
rect 9702 4743 9722 4763
rect 9798 4743 9818 4763
rect 785 4146 805 4166
rect 881 4146 901 4166
rect 998 4146 1018 4166
rect 1094 4146 1114 4166
rect 1206 4146 1226 4166
rect 1302 4146 1322 4166
rect 1412 4146 1432 4166
rect 1508 4146 1528 4166
rect 1833 4142 1853 4162
rect 1929 4142 1949 4162
rect 2046 4142 2066 4162
rect 2142 4142 2162 4162
rect 2254 4142 2274 4162
rect 2350 4142 2370 4162
rect 2460 4142 2480 4162
rect 2556 4142 2576 4162
rect 6580 3980 6600 4000
rect 6676 3980 6696 4000
rect 6786 3980 6806 4000
rect 6882 3980 6902 4000
rect 6994 3980 7014 4000
rect 7090 3980 7110 4000
rect 7207 3980 7227 4000
rect 7303 3980 7323 4000
rect 9075 3975 9095 3995
rect 9171 3975 9191 3995
rect 9281 3975 9301 3995
rect 9377 3975 9397 3995
rect 9489 3975 9509 3995
rect 9585 3975 9605 3995
rect 9702 3975 9722 3995
rect 9798 3975 9818 3995
rect 785 3467 805 3487
rect 881 3467 901 3487
rect 998 3467 1018 3487
rect 1094 3467 1114 3487
rect 1206 3467 1226 3487
rect 1302 3467 1322 3487
rect 1412 3467 1432 3487
rect 1508 3467 1528 3487
rect 3323 3464 3343 3484
rect 3419 3464 3439 3484
rect 3536 3464 3556 3484
rect 3632 3464 3652 3484
rect 3744 3464 3764 3484
rect 3840 3464 3860 3484
rect 3950 3464 3970 3484
rect 4046 3464 4066 3484
rect 8027 3300 8047 3320
rect 8123 3300 8143 3320
rect 8233 3300 8253 3320
rect 8329 3300 8349 3320
rect 8441 3300 8461 3320
rect 8537 3300 8557 3320
rect 8654 3300 8674 3320
rect 8750 3300 8770 3320
rect 9075 3296 9095 3316
rect 9171 3296 9191 3316
rect 9281 3296 9301 3316
rect 9377 3296 9397 3316
rect 9489 3296 9509 3316
rect 9585 3296 9605 3316
rect 9702 3296 9722 3316
rect 9798 3296 9818 3316
rect 786 2626 806 2646
rect 882 2626 902 2646
rect 999 2626 1019 2646
rect 1095 2626 1115 2646
rect 1207 2626 1227 2646
rect 1303 2626 1323 2646
rect 1413 2626 1433 2646
rect 1509 2626 1529 2646
rect 1834 2622 1854 2642
rect 1930 2622 1950 2642
rect 2047 2622 2067 2642
rect 2143 2622 2163 2642
rect 2255 2622 2275 2642
rect 2351 2622 2371 2642
rect 2461 2622 2481 2642
rect 2557 2622 2577 2642
rect 4736 2628 4756 2648
rect 4832 2628 4852 2648
rect 4949 2628 4969 2648
rect 5045 2628 5065 2648
rect 5157 2628 5177 2648
rect 5253 2628 5273 2648
rect 5363 2628 5383 2648
rect 5459 2628 5479 2648
rect 6538 2458 6558 2478
rect 6634 2458 6654 2478
rect 6744 2458 6764 2478
rect 6840 2458 6860 2478
rect 6952 2458 6972 2478
rect 7048 2458 7068 2478
rect 7165 2458 7185 2478
rect 7261 2458 7281 2478
rect 9076 2455 9096 2475
rect 9172 2455 9192 2475
rect 9282 2455 9302 2475
rect 9378 2455 9398 2475
rect 9490 2455 9510 2475
rect 9586 2455 9606 2475
rect 9703 2455 9723 2475
rect 9799 2455 9819 2475
rect 786 1947 806 1967
rect 882 1947 902 1967
rect 999 1947 1019 1967
rect 1095 1947 1115 1967
rect 1207 1947 1227 1967
rect 1303 1947 1323 1967
rect 1413 1947 1433 1967
rect 1509 1947 1529 1967
rect 3281 1942 3301 1962
rect 3377 1942 3397 1962
rect 3494 1942 3514 1962
rect 3590 1942 3610 1962
rect 3702 1942 3722 1962
rect 3798 1942 3818 1962
rect 3908 1942 3928 1962
rect 4004 1942 4024 1962
rect 8028 1780 8048 1800
rect 8124 1780 8144 1800
rect 8234 1780 8254 1800
rect 8330 1780 8350 1800
rect 8442 1780 8462 1800
rect 8538 1780 8558 1800
rect 8655 1780 8675 1800
rect 8751 1780 8771 1800
rect 9076 1776 9096 1796
rect 9172 1776 9192 1796
rect 9282 1776 9302 1796
rect 9378 1776 9398 1796
rect 9490 1776 9510 1796
rect 9586 1776 9606 1796
rect 9703 1776 9723 1796
rect 9799 1776 9819 1796
rect 786 1179 806 1199
rect 882 1179 902 1199
rect 999 1179 1019 1199
rect 1095 1179 1115 1199
rect 1207 1179 1227 1199
rect 1303 1179 1323 1199
rect 1413 1179 1433 1199
rect 1509 1179 1529 1199
rect 1834 1175 1854 1195
rect 1930 1175 1950 1195
rect 2047 1175 2067 1195
rect 2143 1175 2163 1195
rect 2255 1175 2275 1195
rect 2351 1175 2371 1195
rect 2461 1175 2481 1195
rect 2557 1175 2577 1195
rect 6581 1013 6601 1033
rect 6677 1013 6697 1033
rect 6787 1013 6807 1033
rect 6883 1013 6903 1033
rect 6995 1013 7015 1033
rect 7091 1013 7111 1033
rect 7208 1013 7228 1033
rect 7304 1013 7324 1033
rect 9076 1008 9096 1028
rect 9172 1008 9192 1028
rect 9282 1008 9302 1028
rect 9378 1008 9398 1028
rect 9490 1008 9510 1028
rect 9586 1008 9606 1028
rect 9703 1008 9723 1028
rect 9799 1008 9819 1028
rect 786 500 806 520
rect 882 500 902 520
rect 999 500 1019 520
rect 1095 500 1115 520
rect 1207 500 1227 520
rect 1303 500 1323 520
rect 1413 500 1433 520
rect 1509 500 1529 520
rect 8028 333 8048 353
rect 8124 333 8144 353
rect 8234 333 8254 353
rect 8330 333 8350 353
rect 8442 333 8462 353
rect 8538 333 8558 353
rect 8655 333 8675 353
rect 8751 333 8771 353
rect 9076 329 9096 349
rect 9172 329 9192 349
rect 9282 329 9302 349
rect 9378 329 9398 349
rect 9490 329 9510 349
rect 9586 329 9606 349
rect 9703 329 9723 349
rect 9799 329 9819 349
<< psubdiff >>
rect 9641 11696 9752 11711
rect 9641 11666 9683 11696
rect 9711 11666 9752 11696
rect 9641 11652 9752 11666
rect 855 11385 966 11399
rect 855 11355 896 11385
rect 924 11355 966 11385
rect 855 11340 966 11355
rect 1903 11381 2014 11395
rect 1903 11351 1944 11381
rect 1972 11351 2014 11381
rect 1903 11336 2014 11351
rect 8593 11021 8704 11036
rect 8593 10991 8635 11021
rect 8663 10991 8704 11021
rect 8593 10977 8704 10991
rect 9641 11017 9752 11032
rect 9641 10987 9683 11017
rect 9711 10987 9752 11017
rect 9641 10973 9752 10987
rect 855 10706 966 10720
rect 855 10676 896 10706
rect 924 10676 966 10706
rect 855 10663 966 10676
rect 3350 10701 3461 10715
rect 3350 10671 3391 10701
rect 3419 10671 3461 10701
rect 3350 10656 3461 10671
rect 7146 10254 7257 10269
rect 7146 10224 7188 10254
rect 7216 10224 7257 10254
rect 7146 10210 7257 10224
rect 9641 10249 9752 10262
rect 9641 10219 9683 10249
rect 9711 10219 9752 10249
rect 9641 10205 9752 10219
rect 855 9938 966 9952
rect 855 9908 896 9938
rect 924 9908 966 9938
rect 855 9893 966 9908
rect 1903 9934 2014 9948
rect 1903 9904 1944 9934
rect 1972 9904 2014 9934
rect 1903 9889 2014 9904
rect 8593 9574 8704 9589
rect 8593 9544 8635 9574
rect 8663 9544 8704 9574
rect 8593 9530 8704 9544
rect 9641 9570 9752 9585
rect 9641 9540 9683 9570
rect 9711 9540 9752 9570
rect 9641 9526 9752 9540
rect 855 9259 966 9273
rect 855 9229 896 9259
rect 924 9229 966 9259
rect 855 9214 966 9229
rect 3393 9256 3504 9270
rect 3393 9226 3434 9256
rect 3462 9226 3504 9256
rect 3393 9211 3504 9226
rect 7104 8732 7215 8747
rect 7104 8702 7146 8732
rect 7174 8702 7215 8732
rect 7104 8688 7215 8702
rect 9642 8729 9753 8744
rect 9642 8699 9684 8729
rect 9712 8699 9753 8729
rect 9642 8685 9753 8699
rect 856 8418 967 8432
rect 856 8388 897 8418
rect 925 8388 967 8418
rect 856 8373 967 8388
rect 1904 8414 2015 8428
rect 1904 8384 1945 8414
rect 1973 8384 2015 8414
rect 1904 8369 2015 8384
rect 8594 8054 8705 8069
rect 8594 8024 8636 8054
rect 8664 8024 8705 8054
rect 8594 8010 8705 8024
rect 9642 8050 9753 8065
rect 9642 8020 9684 8050
rect 9712 8020 9753 8050
rect 9642 8006 9753 8020
rect 856 7739 967 7753
rect 856 7709 897 7739
rect 925 7709 967 7739
rect 856 7696 967 7709
rect 3351 7734 3462 7748
rect 3351 7704 3392 7734
rect 3420 7704 3462 7734
rect 3351 7689 3462 7704
rect 7147 7287 7258 7302
rect 7147 7257 7189 7287
rect 7217 7257 7258 7287
rect 7147 7243 7258 7257
rect 9642 7282 9753 7295
rect 9642 7252 9684 7282
rect 9712 7252 9753 7282
rect 9642 7238 9753 7252
rect 856 6971 967 6985
rect 856 6941 897 6971
rect 925 6941 967 6971
rect 856 6926 967 6941
rect 1904 6967 2015 6981
rect 1904 6937 1945 6967
rect 1973 6937 2015 6967
rect 1904 6922 2015 6937
rect 8594 6607 8705 6622
rect 8594 6577 8636 6607
rect 8664 6577 8705 6607
rect 8594 6563 8705 6577
rect 9642 6603 9753 6618
rect 9642 6573 9684 6603
rect 9712 6573 9753 6603
rect 9642 6559 9753 6573
rect 856 6292 967 6306
rect 856 6262 897 6292
rect 925 6262 967 6292
rect 856 6247 967 6262
rect 4459 6283 4570 6297
rect 4459 6253 4500 6283
rect 4528 6253 4570 6283
rect 4459 6238 4570 6253
rect 6036 5697 6147 5712
rect 6036 5667 6078 5697
rect 6106 5667 6147 5697
rect 6036 5653 6147 5667
rect 9639 5688 9750 5703
rect 9639 5658 9681 5688
rect 9709 5658 9750 5688
rect 9639 5644 9750 5658
rect 853 5377 964 5391
rect 853 5347 894 5377
rect 922 5347 964 5377
rect 853 5332 964 5347
rect 1901 5373 2012 5387
rect 1901 5343 1942 5373
rect 1970 5343 2012 5373
rect 1901 5328 2012 5343
rect 8591 5013 8702 5028
rect 8591 4983 8633 5013
rect 8661 4983 8702 5013
rect 8591 4969 8702 4983
rect 9639 5009 9750 5024
rect 9639 4979 9681 5009
rect 9709 4979 9750 5009
rect 9639 4965 9750 4979
rect 853 4698 964 4712
rect 853 4668 894 4698
rect 922 4668 964 4698
rect 853 4655 964 4668
rect 3348 4693 3459 4707
rect 3348 4663 3389 4693
rect 3417 4663 3459 4693
rect 3348 4648 3459 4663
rect 7144 4246 7255 4261
rect 7144 4216 7186 4246
rect 7214 4216 7255 4246
rect 7144 4202 7255 4216
rect 9639 4241 9750 4254
rect 9639 4211 9681 4241
rect 9709 4211 9750 4241
rect 9639 4197 9750 4211
rect 853 3930 964 3944
rect 853 3900 894 3930
rect 922 3900 964 3930
rect 853 3885 964 3900
rect 1901 3926 2012 3940
rect 1901 3896 1942 3926
rect 1970 3896 2012 3926
rect 1901 3881 2012 3896
rect 8591 3566 8702 3581
rect 8591 3536 8633 3566
rect 8661 3536 8702 3566
rect 8591 3522 8702 3536
rect 9639 3562 9750 3577
rect 9639 3532 9681 3562
rect 9709 3532 9750 3562
rect 9639 3518 9750 3532
rect 853 3251 964 3265
rect 853 3221 894 3251
rect 922 3221 964 3251
rect 853 3206 964 3221
rect 3391 3248 3502 3262
rect 3391 3218 3432 3248
rect 3460 3218 3502 3248
rect 3391 3203 3502 3218
rect 7102 2724 7213 2739
rect 7102 2694 7144 2724
rect 7172 2694 7213 2724
rect 7102 2680 7213 2694
rect 9640 2721 9751 2736
rect 9640 2691 9682 2721
rect 9710 2691 9751 2721
rect 9640 2677 9751 2691
rect 854 2410 965 2424
rect 854 2380 895 2410
rect 923 2380 965 2410
rect 854 2365 965 2380
rect 1902 2406 2013 2420
rect 1902 2376 1943 2406
rect 1971 2376 2013 2406
rect 1902 2361 2013 2376
rect 4804 2412 4915 2426
rect 4804 2382 4845 2412
rect 4873 2382 4915 2412
rect 4804 2367 4915 2382
rect 8592 2046 8703 2061
rect 8592 2016 8634 2046
rect 8662 2016 8703 2046
rect 8592 2002 8703 2016
rect 9640 2042 9751 2057
rect 9640 2012 9682 2042
rect 9710 2012 9751 2042
rect 9640 1998 9751 2012
rect 854 1731 965 1745
rect 854 1701 895 1731
rect 923 1701 965 1731
rect 854 1688 965 1701
rect 3349 1726 3460 1740
rect 3349 1696 3390 1726
rect 3418 1696 3460 1726
rect 3349 1681 3460 1696
rect 7145 1279 7256 1294
rect 7145 1249 7187 1279
rect 7215 1249 7256 1279
rect 7145 1235 7256 1249
rect 9640 1274 9751 1287
rect 9640 1244 9682 1274
rect 9710 1244 9751 1274
rect 9640 1230 9751 1244
rect 854 963 965 977
rect 854 933 895 963
rect 923 933 965 963
rect 854 918 965 933
rect 1902 959 2013 973
rect 1902 929 1943 959
rect 1971 929 2013 959
rect 1902 914 2013 929
rect 8592 599 8703 614
rect 8592 569 8634 599
rect 8662 569 8703 599
rect 8592 555 8703 569
rect 9640 595 9751 610
rect 9640 565 9682 595
rect 9710 565 9751 595
rect 9640 551 9751 565
rect 854 284 965 298
rect 854 254 895 284
rect 923 254 965 284
rect 854 239 965 254
<< nsubdiff >>
rect 856 11732 966 11746
rect 856 11702 899 11732
rect 927 11702 966 11732
rect 856 11687 966 11702
rect 1904 11728 2014 11742
rect 1904 11698 1947 11728
rect 1975 11698 2014 11728
rect 1904 11683 2014 11698
rect 9641 11349 9751 11364
rect 9641 11319 9680 11349
rect 9708 11319 9751 11349
rect 9641 11305 9751 11319
rect 856 11053 966 11067
rect 856 11023 899 11053
rect 927 11023 966 11053
rect 856 11008 966 11023
rect 3351 11048 3461 11062
rect 3351 11018 3394 11048
rect 3422 11018 3461 11048
rect 3351 11003 3461 11018
rect 8593 10674 8703 10689
rect 8593 10644 8632 10674
rect 8660 10644 8703 10674
rect 8593 10630 8703 10644
rect 9641 10670 9751 10685
rect 9641 10640 9680 10670
rect 9708 10640 9751 10670
rect 9641 10626 9751 10640
rect 856 10285 966 10299
rect 856 10255 899 10285
rect 927 10255 966 10285
rect 856 10240 966 10255
rect 1904 10281 2014 10295
rect 1904 10251 1947 10281
rect 1975 10251 2014 10281
rect 1904 10236 2014 10251
rect 7146 9907 7256 9922
rect 7146 9877 7185 9907
rect 7213 9877 7256 9907
rect 7146 9863 7256 9877
rect 9641 9902 9751 9917
rect 9641 9872 9680 9902
rect 9708 9872 9751 9902
rect 9641 9858 9751 9872
rect 856 9606 966 9620
rect 856 9576 899 9606
rect 927 9576 966 9606
rect 856 9561 966 9576
rect 3394 9603 3504 9617
rect 3394 9573 3437 9603
rect 3465 9573 3504 9603
rect 3394 9558 3504 9573
rect 8593 9227 8703 9242
rect 8593 9197 8632 9227
rect 8660 9197 8703 9227
rect 8593 9183 8703 9197
rect 9641 9223 9751 9238
rect 9641 9193 9680 9223
rect 9708 9193 9751 9223
rect 9641 9179 9751 9193
rect 857 8765 967 8779
rect 857 8735 900 8765
rect 928 8735 967 8765
rect 857 8720 967 8735
rect 1905 8761 2015 8775
rect 1905 8731 1948 8761
rect 1976 8731 2015 8761
rect 1905 8716 2015 8731
rect 7104 8385 7214 8400
rect 7104 8355 7143 8385
rect 7171 8355 7214 8385
rect 7104 8341 7214 8355
rect 9642 8382 9752 8397
rect 9642 8352 9681 8382
rect 9709 8352 9752 8382
rect 9642 8338 9752 8352
rect 857 8086 967 8100
rect 857 8056 900 8086
rect 928 8056 967 8086
rect 857 8041 967 8056
rect 3352 8081 3462 8095
rect 3352 8051 3395 8081
rect 3423 8051 3462 8081
rect 3352 8036 3462 8051
rect 8594 7707 8704 7722
rect 8594 7677 8633 7707
rect 8661 7677 8704 7707
rect 8594 7663 8704 7677
rect 9642 7703 9752 7718
rect 9642 7673 9681 7703
rect 9709 7673 9752 7703
rect 9642 7659 9752 7673
rect 857 7318 967 7332
rect 857 7288 900 7318
rect 928 7288 967 7318
rect 857 7273 967 7288
rect 1905 7314 2015 7328
rect 1905 7284 1948 7314
rect 1976 7284 2015 7314
rect 1905 7269 2015 7284
rect 7147 6940 7257 6955
rect 7147 6910 7186 6940
rect 7214 6910 7257 6940
rect 7147 6896 7257 6910
rect 9642 6935 9752 6950
rect 9642 6905 9681 6935
rect 9709 6905 9752 6935
rect 9642 6891 9752 6905
rect 857 6639 967 6653
rect 857 6609 900 6639
rect 928 6609 967 6639
rect 857 6594 967 6609
rect 4460 6630 4570 6644
rect 4460 6600 4503 6630
rect 4531 6600 4570 6630
rect 4460 6585 4570 6600
rect 8594 6260 8704 6275
rect 8594 6230 8633 6260
rect 8661 6230 8704 6260
rect 8594 6216 8704 6230
rect 9642 6256 9752 6271
rect 9642 6226 9681 6256
rect 9709 6226 9752 6256
rect 9642 6212 9752 6226
rect 854 5724 964 5738
rect 854 5694 897 5724
rect 925 5694 964 5724
rect 854 5679 964 5694
rect 1902 5720 2012 5734
rect 1902 5690 1945 5720
rect 1973 5690 2012 5720
rect 1902 5675 2012 5690
rect 6036 5350 6146 5365
rect 6036 5320 6075 5350
rect 6103 5320 6146 5350
rect 6036 5306 6146 5320
rect 9639 5341 9749 5356
rect 9639 5311 9678 5341
rect 9706 5311 9749 5341
rect 9639 5297 9749 5311
rect 854 5045 964 5059
rect 854 5015 897 5045
rect 925 5015 964 5045
rect 854 5000 964 5015
rect 3349 5040 3459 5054
rect 3349 5010 3392 5040
rect 3420 5010 3459 5040
rect 3349 4995 3459 5010
rect 8591 4666 8701 4681
rect 8591 4636 8630 4666
rect 8658 4636 8701 4666
rect 8591 4622 8701 4636
rect 9639 4662 9749 4677
rect 9639 4632 9678 4662
rect 9706 4632 9749 4662
rect 9639 4618 9749 4632
rect 854 4277 964 4291
rect 854 4247 897 4277
rect 925 4247 964 4277
rect 854 4232 964 4247
rect 1902 4273 2012 4287
rect 1902 4243 1945 4273
rect 1973 4243 2012 4273
rect 1902 4228 2012 4243
rect 7144 3899 7254 3914
rect 7144 3869 7183 3899
rect 7211 3869 7254 3899
rect 7144 3855 7254 3869
rect 9639 3894 9749 3909
rect 9639 3864 9678 3894
rect 9706 3864 9749 3894
rect 9639 3850 9749 3864
rect 854 3598 964 3612
rect 854 3568 897 3598
rect 925 3568 964 3598
rect 854 3553 964 3568
rect 3392 3595 3502 3609
rect 3392 3565 3435 3595
rect 3463 3565 3502 3595
rect 3392 3550 3502 3565
rect 8591 3219 8701 3234
rect 8591 3189 8630 3219
rect 8658 3189 8701 3219
rect 8591 3175 8701 3189
rect 9639 3215 9749 3230
rect 9639 3185 9678 3215
rect 9706 3185 9749 3215
rect 9639 3171 9749 3185
rect 855 2757 965 2771
rect 855 2727 898 2757
rect 926 2727 965 2757
rect 855 2712 965 2727
rect 1903 2753 2013 2767
rect 1903 2723 1946 2753
rect 1974 2723 2013 2753
rect 1903 2708 2013 2723
rect 4805 2759 4915 2773
rect 4805 2729 4848 2759
rect 4876 2729 4915 2759
rect 4805 2714 4915 2729
rect 7102 2377 7212 2392
rect 7102 2347 7141 2377
rect 7169 2347 7212 2377
rect 7102 2333 7212 2347
rect 9640 2374 9750 2389
rect 9640 2344 9679 2374
rect 9707 2344 9750 2374
rect 9640 2330 9750 2344
rect 855 2078 965 2092
rect 855 2048 898 2078
rect 926 2048 965 2078
rect 855 2033 965 2048
rect 3350 2073 3460 2087
rect 3350 2043 3393 2073
rect 3421 2043 3460 2073
rect 3350 2028 3460 2043
rect 8592 1699 8702 1714
rect 8592 1669 8631 1699
rect 8659 1669 8702 1699
rect 8592 1655 8702 1669
rect 9640 1695 9750 1710
rect 9640 1665 9679 1695
rect 9707 1665 9750 1695
rect 9640 1651 9750 1665
rect 855 1310 965 1324
rect 855 1280 898 1310
rect 926 1280 965 1310
rect 855 1265 965 1280
rect 1903 1306 2013 1320
rect 1903 1276 1946 1306
rect 1974 1276 2013 1306
rect 1903 1261 2013 1276
rect 7145 932 7255 947
rect 7145 902 7184 932
rect 7212 902 7255 932
rect 7145 888 7255 902
rect 9640 927 9750 942
rect 9640 897 9679 927
rect 9707 897 9750 927
rect 9640 883 9750 897
rect 855 631 965 645
rect 855 601 898 631
rect 926 601 965 631
rect 855 586 965 601
rect 8592 252 8702 267
rect 8592 222 8631 252
rect 8659 222 8702 252
rect 8592 208 8702 222
rect 9640 248 9750 263
rect 9640 218 9679 248
rect 9707 218 9750 248
rect 9640 204 9750 218
<< psubdiffcont >>
rect 9683 11666 9711 11696
rect 896 11355 924 11385
rect 1944 11351 1972 11381
rect 8635 10991 8663 11021
rect 9683 10987 9711 11017
rect 896 10676 924 10706
rect 3391 10671 3419 10701
rect 7188 10224 7216 10254
rect 9683 10219 9711 10249
rect 896 9908 924 9938
rect 1944 9904 1972 9934
rect 8635 9544 8663 9574
rect 9683 9540 9711 9570
rect 896 9229 924 9259
rect 3434 9226 3462 9256
rect 7146 8702 7174 8732
rect 9684 8699 9712 8729
rect 897 8388 925 8418
rect 1945 8384 1973 8414
rect 8636 8024 8664 8054
rect 9684 8020 9712 8050
rect 897 7709 925 7739
rect 3392 7704 3420 7734
rect 7189 7257 7217 7287
rect 9684 7252 9712 7282
rect 897 6941 925 6971
rect 1945 6937 1973 6967
rect 8636 6577 8664 6607
rect 9684 6573 9712 6603
rect 897 6262 925 6292
rect 4500 6253 4528 6283
rect 6078 5667 6106 5697
rect 9681 5658 9709 5688
rect 894 5347 922 5377
rect 1942 5343 1970 5373
rect 8633 4983 8661 5013
rect 9681 4979 9709 5009
rect 894 4668 922 4698
rect 3389 4663 3417 4693
rect 7186 4216 7214 4246
rect 9681 4211 9709 4241
rect 894 3900 922 3930
rect 1942 3896 1970 3926
rect 8633 3536 8661 3566
rect 9681 3532 9709 3562
rect 894 3221 922 3251
rect 3432 3218 3460 3248
rect 7144 2694 7172 2724
rect 9682 2691 9710 2721
rect 895 2380 923 2410
rect 1943 2376 1971 2406
rect 4845 2382 4873 2412
rect 8634 2016 8662 2046
rect 9682 2012 9710 2042
rect 895 1701 923 1731
rect 3390 1696 3418 1726
rect 7187 1249 7215 1279
rect 9682 1244 9710 1274
rect 895 933 923 963
rect 1943 929 1971 959
rect 8634 569 8662 599
rect 9682 565 9710 595
rect 895 254 923 284
<< nsubdiffcont >>
rect 899 11702 927 11732
rect 1947 11698 1975 11728
rect 9680 11319 9708 11349
rect 899 11023 927 11053
rect 3394 11018 3422 11048
rect 8632 10644 8660 10674
rect 9680 10640 9708 10670
rect 899 10255 927 10285
rect 1947 10251 1975 10281
rect 7185 9877 7213 9907
rect 9680 9872 9708 9902
rect 899 9576 927 9606
rect 3437 9573 3465 9603
rect 8632 9197 8660 9227
rect 9680 9193 9708 9223
rect 900 8735 928 8765
rect 1948 8731 1976 8761
rect 7143 8355 7171 8385
rect 9681 8352 9709 8382
rect 900 8056 928 8086
rect 3395 8051 3423 8081
rect 8633 7677 8661 7707
rect 9681 7673 9709 7703
rect 900 7288 928 7318
rect 1948 7284 1976 7314
rect 7186 6910 7214 6940
rect 9681 6905 9709 6935
rect 900 6609 928 6639
rect 4503 6600 4531 6630
rect 8633 6230 8661 6260
rect 9681 6226 9709 6256
rect 897 5694 925 5724
rect 1945 5690 1973 5720
rect 6075 5320 6103 5350
rect 9678 5311 9706 5341
rect 897 5015 925 5045
rect 3392 5010 3420 5040
rect 8630 4636 8658 4666
rect 9678 4632 9706 4662
rect 897 4247 925 4277
rect 1945 4243 1973 4273
rect 7183 3869 7211 3899
rect 9678 3864 9706 3894
rect 897 3568 925 3598
rect 3435 3565 3463 3595
rect 8630 3189 8658 3219
rect 9678 3185 9706 3215
rect 898 2727 926 2757
rect 1946 2723 1974 2753
rect 4848 2729 4876 2759
rect 7141 2347 7169 2377
rect 9679 2344 9707 2374
rect 898 2048 926 2078
rect 3393 2043 3421 2073
rect 8631 1669 8659 1699
rect 9679 1665 9707 1695
rect 898 1280 926 1310
rect 1946 1276 1974 1306
rect 7184 902 7212 932
rect 9679 897 9707 927
rect 898 601 926 631
rect 8631 222 8659 252
rect 9679 218 9707 248
<< poly >>
rect 819 11659 869 11672
rect 1032 11659 1082 11672
rect 1240 11659 1290 11672
rect 1448 11659 1498 11672
rect 1867 11655 1917 11668
rect 2080 11655 2130 11668
rect 2288 11655 2338 11668
rect 2496 11655 2546 11668
rect 819 11531 869 11559
rect 819 11511 832 11531
rect 852 11511 869 11531
rect 819 11482 869 11511
rect 1032 11530 1082 11559
rect 1032 11506 1043 11530
rect 1067 11506 1082 11530
rect 1032 11482 1082 11506
rect 1240 11535 1290 11559
rect 1240 11511 1252 11535
rect 1276 11511 1290 11535
rect 1240 11482 1290 11511
rect 1448 11533 1498 11559
rect 9109 11611 9159 11627
rect 9317 11611 9367 11627
rect 9525 11611 9575 11627
rect 9738 11611 9788 11627
rect 1448 11507 1466 11533
rect 1492 11507 1498 11533
rect 1448 11482 1498 11507
rect 1867 11527 1917 11555
rect 1867 11507 1880 11527
rect 1900 11507 1917 11527
rect 1867 11478 1917 11507
rect 2080 11526 2130 11555
rect 2080 11502 2091 11526
rect 2115 11502 2130 11526
rect 2080 11478 2130 11502
rect 2288 11531 2338 11555
rect 2288 11507 2300 11531
rect 2324 11507 2338 11531
rect 2288 11478 2338 11507
rect 2496 11529 2546 11555
rect 2496 11503 2514 11529
rect 2540 11503 2546 11529
rect 2496 11478 2546 11503
rect 9109 11544 9159 11569
rect 9109 11518 9115 11544
rect 9141 11518 9159 11544
rect 9109 11492 9159 11518
rect 9317 11540 9367 11569
rect 9317 11516 9331 11540
rect 9355 11516 9367 11540
rect 9317 11492 9367 11516
rect 9525 11545 9575 11569
rect 9525 11521 9540 11545
rect 9564 11521 9575 11545
rect 9525 11492 9575 11521
rect 9738 11540 9788 11569
rect 9738 11520 9755 11540
rect 9775 11520 9788 11540
rect 9738 11492 9788 11520
rect 819 11424 869 11440
rect 1032 11424 1082 11440
rect 1240 11424 1290 11440
rect 1448 11424 1498 11440
rect 1867 11420 1917 11436
rect 2080 11420 2130 11436
rect 2288 11420 2338 11436
rect 2496 11420 2546 11436
rect 9109 11379 9159 11392
rect 9317 11379 9367 11392
rect 9525 11379 9575 11392
rect 9738 11379 9788 11392
rect 819 10980 869 10993
rect 1032 10980 1082 10993
rect 1240 10980 1290 10993
rect 1448 10980 1498 10993
rect 3314 10975 3364 10988
rect 3527 10975 3577 10988
rect 3735 10975 3785 10988
rect 3943 10975 3993 10988
rect 819 10852 869 10880
rect 819 10832 832 10852
rect 852 10832 869 10852
rect 819 10803 869 10832
rect 1032 10851 1082 10880
rect 1032 10827 1043 10851
rect 1067 10827 1082 10851
rect 1032 10803 1082 10827
rect 1240 10856 1290 10880
rect 1240 10832 1252 10856
rect 1276 10832 1290 10856
rect 1240 10803 1290 10832
rect 1448 10854 1498 10880
rect 8061 10936 8111 10952
rect 8269 10936 8319 10952
rect 8477 10936 8527 10952
rect 8690 10936 8740 10952
rect 9109 10932 9159 10948
rect 9317 10932 9367 10948
rect 9525 10932 9575 10948
rect 9738 10932 9788 10948
rect 1448 10828 1466 10854
rect 1492 10828 1498 10854
rect 1448 10803 1498 10828
rect 3314 10847 3364 10875
rect 3314 10827 3327 10847
rect 3347 10827 3364 10847
rect 3314 10798 3364 10827
rect 3527 10846 3577 10875
rect 3527 10822 3538 10846
rect 3562 10822 3577 10846
rect 3527 10798 3577 10822
rect 3735 10851 3785 10875
rect 3735 10827 3747 10851
rect 3771 10827 3785 10851
rect 3735 10798 3785 10827
rect 3943 10849 3993 10875
rect 3943 10823 3961 10849
rect 3987 10823 3993 10849
rect 3943 10798 3993 10823
rect 8061 10869 8111 10894
rect 8061 10843 8067 10869
rect 8093 10843 8111 10869
rect 8061 10817 8111 10843
rect 8269 10865 8319 10894
rect 8269 10841 8283 10865
rect 8307 10841 8319 10865
rect 8269 10817 8319 10841
rect 8477 10870 8527 10894
rect 8477 10846 8492 10870
rect 8516 10846 8527 10870
rect 8477 10817 8527 10846
rect 8690 10865 8740 10894
rect 8690 10845 8707 10865
rect 8727 10845 8740 10865
rect 8690 10817 8740 10845
rect 9109 10865 9159 10890
rect 9109 10839 9115 10865
rect 9141 10839 9159 10865
rect 819 10745 869 10761
rect 1032 10745 1082 10761
rect 1240 10745 1290 10761
rect 1448 10745 1498 10761
rect 3314 10740 3364 10756
rect 3527 10740 3577 10756
rect 3735 10740 3785 10756
rect 3943 10740 3993 10756
rect 9109 10813 9159 10839
rect 9317 10861 9367 10890
rect 9317 10837 9331 10861
rect 9355 10837 9367 10861
rect 9317 10813 9367 10837
rect 9525 10866 9575 10890
rect 9525 10842 9540 10866
rect 9564 10842 9575 10866
rect 9525 10813 9575 10842
rect 9738 10861 9788 10890
rect 9738 10841 9755 10861
rect 9775 10841 9788 10861
rect 9738 10813 9788 10841
rect 8061 10704 8111 10717
rect 8269 10704 8319 10717
rect 8477 10704 8527 10717
rect 8690 10704 8740 10717
rect 9109 10700 9159 10713
rect 9317 10700 9367 10713
rect 9525 10700 9575 10713
rect 9738 10700 9788 10713
rect 819 10212 869 10225
rect 1032 10212 1082 10225
rect 1240 10212 1290 10225
rect 1448 10212 1498 10225
rect 1867 10208 1917 10221
rect 2080 10208 2130 10221
rect 2288 10208 2338 10221
rect 2496 10208 2546 10221
rect 819 10084 869 10112
rect 819 10064 832 10084
rect 852 10064 869 10084
rect 819 10035 869 10064
rect 1032 10083 1082 10112
rect 1032 10059 1043 10083
rect 1067 10059 1082 10083
rect 1032 10035 1082 10059
rect 1240 10088 1290 10112
rect 1240 10064 1252 10088
rect 1276 10064 1290 10088
rect 1240 10035 1290 10064
rect 1448 10086 1498 10112
rect 6614 10169 6664 10185
rect 6822 10169 6872 10185
rect 7030 10169 7080 10185
rect 7243 10169 7293 10185
rect 9109 10164 9159 10180
rect 9317 10164 9367 10180
rect 9525 10164 9575 10180
rect 9738 10164 9788 10180
rect 1448 10060 1466 10086
rect 1492 10060 1498 10086
rect 1448 10035 1498 10060
rect 1867 10080 1917 10108
rect 1867 10060 1880 10080
rect 1900 10060 1917 10080
rect 1867 10031 1917 10060
rect 2080 10079 2130 10108
rect 2080 10055 2091 10079
rect 2115 10055 2130 10079
rect 2080 10031 2130 10055
rect 2288 10084 2338 10108
rect 2288 10060 2300 10084
rect 2324 10060 2338 10084
rect 2288 10031 2338 10060
rect 2496 10082 2546 10108
rect 2496 10056 2514 10082
rect 2540 10056 2546 10082
rect 2496 10031 2546 10056
rect 6614 10102 6664 10127
rect 6614 10076 6620 10102
rect 6646 10076 6664 10102
rect 6614 10050 6664 10076
rect 6822 10098 6872 10127
rect 6822 10074 6836 10098
rect 6860 10074 6872 10098
rect 6822 10050 6872 10074
rect 7030 10103 7080 10127
rect 7030 10079 7045 10103
rect 7069 10079 7080 10103
rect 7030 10050 7080 10079
rect 7243 10098 7293 10127
rect 7243 10078 7260 10098
rect 7280 10078 7293 10098
rect 7243 10050 7293 10078
rect 9109 10097 9159 10122
rect 9109 10071 9115 10097
rect 9141 10071 9159 10097
rect 819 9977 869 9993
rect 1032 9977 1082 9993
rect 1240 9977 1290 9993
rect 1448 9977 1498 9993
rect 1867 9973 1917 9989
rect 2080 9973 2130 9989
rect 2288 9973 2338 9989
rect 2496 9973 2546 9989
rect 9109 10045 9159 10071
rect 9317 10093 9367 10122
rect 9317 10069 9331 10093
rect 9355 10069 9367 10093
rect 9317 10045 9367 10069
rect 9525 10098 9575 10122
rect 9525 10074 9540 10098
rect 9564 10074 9575 10098
rect 9525 10045 9575 10074
rect 9738 10093 9788 10122
rect 9738 10073 9755 10093
rect 9775 10073 9788 10093
rect 9738 10045 9788 10073
rect 6614 9937 6664 9950
rect 6822 9937 6872 9950
rect 7030 9937 7080 9950
rect 7243 9937 7293 9950
rect 9109 9932 9159 9945
rect 9317 9932 9367 9945
rect 9525 9932 9575 9945
rect 9738 9932 9788 9945
rect 819 9533 869 9546
rect 1032 9533 1082 9546
rect 1240 9533 1290 9546
rect 1448 9533 1498 9546
rect 3357 9530 3407 9543
rect 3570 9530 3620 9543
rect 3778 9530 3828 9543
rect 3986 9530 4036 9543
rect 819 9405 869 9433
rect 819 9385 832 9405
rect 852 9385 869 9405
rect 819 9356 869 9385
rect 1032 9404 1082 9433
rect 1032 9380 1043 9404
rect 1067 9380 1082 9404
rect 1032 9356 1082 9380
rect 1240 9409 1290 9433
rect 1240 9385 1252 9409
rect 1276 9385 1290 9409
rect 1240 9356 1290 9385
rect 1448 9407 1498 9433
rect 8061 9489 8111 9505
rect 8269 9489 8319 9505
rect 8477 9489 8527 9505
rect 8690 9489 8740 9505
rect 9109 9485 9159 9501
rect 9317 9485 9367 9501
rect 9525 9485 9575 9501
rect 9738 9485 9788 9501
rect 1448 9381 1466 9407
rect 1492 9381 1498 9407
rect 1448 9356 1498 9381
rect 3357 9402 3407 9430
rect 3357 9382 3370 9402
rect 3390 9382 3407 9402
rect 3357 9353 3407 9382
rect 3570 9401 3620 9430
rect 3570 9377 3581 9401
rect 3605 9377 3620 9401
rect 3570 9353 3620 9377
rect 3778 9406 3828 9430
rect 3778 9382 3790 9406
rect 3814 9382 3828 9406
rect 3778 9353 3828 9382
rect 3986 9404 4036 9430
rect 3986 9378 4004 9404
rect 4030 9378 4036 9404
rect 3986 9353 4036 9378
rect 8061 9422 8111 9447
rect 8061 9396 8067 9422
rect 8093 9396 8111 9422
rect 8061 9370 8111 9396
rect 8269 9418 8319 9447
rect 8269 9394 8283 9418
rect 8307 9394 8319 9418
rect 8269 9370 8319 9394
rect 8477 9423 8527 9447
rect 8477 9399 8492 9423
rect 8516 9399 8527 9423
rect 8477 9370 8527 9399
rect 8690 9418 8740 9447
rect 8690 9398 8707 9418
rect 8727 9398 8740 9418
rect 8690 9370 8740 9398
rect 9109 9418 9159 9443
rect 9109 9392 9115 9418
rect 9141 9392 9159 9418
rect 819 9298 869 9314
rect 1032 9298 1082 9314
rect 1240 9298 1290 9314
rect 1448 9298 1498 9314
rect 3357 9295 3407 9311
rect 3570 9295 3620 9311
rect 3778 9295 3828 9311
rect 3986 9295 4036 9311
rect 9109 9366 9159 9392
rect 9317 9414 9367 9443
rect 9317 9390 9331 9414
rect 9355 9390 9367 9414
rect 9317 9366 9367 9390
rect 9525 9419 9575 9443
rect 9525 9395 9540 9419
rect 9564 9395 9575 9419
rect 9525 9366 9575 9395
rect 9738 9414 9788 9443
rect 9738 9394 9755 9414
rect 9775 9394 9788 9414
rect 9738 9366 9788 9394
rect 8061 9257 8111 9270
rect 8269 9257 8319 9270
rect 8477 9257 8527 9270
rect 8690 9257 8740 9270
rect 9109 9253 9159 9266
rect 9317 9253 9367 9266
rect 9525 9253 9575 9266
rect 9738 9253 9788 9266
rect 820 8692 870 8705
rect 1033 8692 1083 8705
rect 1241 8692 1291 8705
rect 1449 8692 1499 8705
rect 1868 8688 1918 8701
rect 2081 8688 2131 8701
rect 2289 8688 2339 8701
rect 2497 8688 2547 8701
rect 820 8564 870 8592
rect 820 8544 833 8564
rect 853 8544 870 8564
rect 820 8515 870 8544
rect 1033 8563 1083 8592
rect 1033 8539 1044 8563
rect 1068 8539 1083 8563
rect 1033 8515 1083 8539
rect 1241 8568 1291 8592
rect 1241 8544 1253 8568
rect 1277 8544 1291 8568
rect 1241 8515 1291 8544
rect 1449 8566 1499 8592
rect 6572 8647 6622 8663
rect 6780 8647 6830 8663
rect 6988 8647 7038 8663
rect 7201 8647 7251 8663
rect 9110 8644 9160 8660
rect 9318 8644 9368 8660
rect 9526 8644 9576 8660
rect 9739 8644 9789 8660
rect 1449 8540 1467 8566
rect 1493 8540 1499 8566
rect 1449 8515 1499 8540
rect 1868 8560 1918 8588
rect 1868 8540 1881 8560
rect 1901 8540 1918 8560
rect 1868 8511 1918 8540
rect 2081 8559 2131 8588
rect 2081 8535 2092 8559
rect 2116 8535 2131 8559
rect 2081 8511 2131 8535
rect 2289 8564 2339 8588
rect 2289 8540 2301 8564
rect 2325 8540 2339 8564
rect 2289 8511 2339 8540
rect 2497 8562 2547 8588
rect 2497 8536 2515 8562
rect 2541 8536 2547 8562
rect 2497 8511 2547 8536
rect 6572 8580 6622 8605
rect 6572 8554 6578 8580
rect 6604 8554 6622 8580
rect 6572 8528 6622 8554
rect 6780 8576 6830 8605
rect 6780 8552 6794 8576
rect 6818 8552 6830 8576
rect 6780 8528 6830 8552
rect 6988 8581 7038 8605
rect 6988 8557 7003 8581
rect 7027 8557 7038 8581
rect 6988 8528 7038 8557
rect 7201 8576 7251 8605
rect 7201 8556 7218 8576
rect 7238 8556 7251 8576
rect 7201 8528 7251 8556
rect 9110 8577 9160 8602
rect 9110 8551 9116 8577
rect 9142 8551 9160 8577
rect 820 8457 870 8473
rect 1033 8457 1083 8473
rect 1241 8457 1291 8473
rect 1449 8457 1499 8473
rect 1868 8453 1918 8469
rect 2081 8453 2131 8469
rect 2289 8453 2339 8469
rect 2497 8453 2547 8469
rect 9110 8525 9160 8551
rect 9318 8573 9368 8602
rect 9318 8549 9332 8573
rect 9356 8549 9368 8573
rect 9318 8525 9368 8549
rect 9526 8578 9576 8602
rect 9526 8554 9541 8578
rect 9565 8554 9576 8578
rect 9526 8525 9576 8554
rect 9739 8573 9789 8602
rect 9739 8553 9756 8573
rect 9776 8553 9789 8573
rect 9739 8525 9789 8553
rect 6572 8415 6622 8428
rect 6780 8415 6830 8428
rect 6988 8415 7038 8428
rect 7201 8415 7251 8428
rect 9110 8412 9160 8425
rect 9318 8412 9368 8425
rect 9526 8412 9576 8425
rect 9739 8412 9789 8425
rect 820 8013 870 8026
rect 1033 8013 1083 8026
rect 1241 8013 1291 8026
rect 1449 8013 1499 8026
rect 3315 8008 3365 8021
rect 3528 8008 3578 8021
rect 3736 8008 3786 8021
rect 3944 8008 3994 8021
rect 820 7885 870 7913
rect 820 7865 833 7885
rect 853 7865 870 7885
rect 820 7836 870 7865
rect 1033 7884 1083 7913
rect 1033 7860 1044 7884
rect 1068 7860 1083 7884
rect 1033 7836 1083 7860
rect 1241 7889 1291 7913
rect 1241 7865 1253 7889
rect 1277 7865 1291 7889
rect 1241 7836 1291 7865
rect 1449 7887 1499 7913
rect 8062 7969 8112 7985
rect 8270 7969 8320 7985
rect 8478 7969 8528 7985
rect 8691 7969 8741 7985
rect 9110 7965 9160 7981
rect 9318 7965 9368 7981
rect 9526 7965 9576 7981
rect 9739 7965 9789 7981
rect 1449 7861 1467 7887
rect 1493 7861 1499 7887
rect 1449 7836 1499 7861
rect 3315 7880 3365 7908
rect 3315 7860 3328 7880
rect 3348 7860 3365 7880
rect 3315 7831 3365 7860
rect 3528 7879 3578 7908
rect 3528 7855 3539 7879
rect 3563 7855 3578 7879
rect 3528 7831 3578 7855
rect 3736 7884 3786 7908
rect 3736 7860 3748 7884
rect 3772 7860 3786 7884
rect 3736 7831 3786 7860
rect 3944 7882 3994 7908
rect 3944 7856 3962 7882
rect 3988 7856 3994 7882
rect 3944 7831 3994 7856
rect 8062 7902 8112 7927
rect 8062 7876 8068 7902
rect 8094 7876 8112 7902
rect 8062 7850 8112 7876
rect 8270 7898 8320 7927
rect 8270 7874 8284 7898
rect 8308 7874 8320 7898
rect 8270 7850 8320 7874
rect 8478 7903 8528 7927
rect 8478 7879 8493 7903
rect 8517 7879 8528 7903
rect 8478 7850 8528 7879
rect 8691 7898 8741 7927
rect 8691 7878 8708 7898
rect 8728 7878 8741 7898
rect 8691 7850 8741 7878
rect 9110 7898 9160 7923
rect 9110 7872 9116 7898
rect 9142 7872 9160 7898
rect 820 7778 870 7794
rect 1033 7778 1083 7794
rect 1241 7778 1291 7794
rect 1449 7778 1499 7794
rect 3315 7773 3365 7789
rect 3528 7773 3578 7789
rect 3736 7773 3786 7789
rect 3944 7773 3994 7789
rect 9110 7846 9160 7872
rect 9318 7894 9368 7923
rect 9318 7870 9332 7894
rect 9356 7870 9368 7894
rect 9318 7846 9368 7870
rect 9526 7899 9576 7923
rect 9526 7875 9541 7899
rect 9565 7875 9576 7899
rect 9526 7846 9576 7875
rect 9739 7894 9789 7923
rect 9739 7874 9756 7894
rect 9776 7874 9789 7894
rect 9739 7846 9789 7874
rect 8062 7737 8112 7750
rect 8270 7737 8320 7750
rect 8478 7737 8528 7750
rect 8691 7737 8741 7750
rect 9110 7733 9160 7746
rect 9318 7733 9368 7746
rect 9526 7733 9576 7746
rect 9739 7733 9789 7746
rect 820 7245 870 7258
rect 1033 7245 1083 7258
rect 1241 7245 1291 7258
rect 1449 7245 1499 7258
rect 1868 7241 1918 7254
rect 2081 7241 2131 7254
rect 2289 7241 2339 7254
rect 2497 7241 2547 7254
rect 820 7117 870 7145
rect 820 7097 833 7117
rect 853 7097 870 7117
rect 820 7068 870 7097
rect 1033 7116 1083 7145
rect 1033 7092 1044 7116
rect 1068 7092 1083 7116
rect 1033 7068 1083 7092
rect 1241 7121 1291 7145
rect 1241 7097 1253 7121
rect 1277 7097 1291 7121
rect 1241 7068 1291 7097
rect 1449 7119 1499 7145
rect 6615 7202 6665 7218
rect 6823 7202 6873 7218
rect 7031 7202 7081 7218
rect 7244 7202 7294 7218
rect 9110 7197 9160 7213
rect 9318 7197 9368 7213
rect 9526 7197 9576 7213
rect 9739 7197 9789 7213
rect 1449 7093 1467 7119
rect 1493 7093 1499 7119
rect 1449 7068 1499 7093
rect 1868 7113 1918 7141
rect 1868 7093 1881 7113
rect 1901 7093 1918 7113
rect 1868 7064 1918 7093
rect 2081 7112 2131 7141
rect 2081 7088 2092 7112
rect 2116 7088 2131 7112
rect 2081 7064 2131 7088
rect 2289 7117 2339 7141
rect 2289 7093 2301 7117
rect 2325 7093 2339 7117
rect 2289 7064 2339 7093
rect 2497 7115 2547 7141
rect 2497 7089 2515 7115
rect 2541 7089 2547 7115
rect 2497 7064 2547 7089
rect 6615 7135 6665 7160
rect 6615 7109 6621 7135
rect 6647 7109 6665 7135
rect 6615 7083 6665 7109
rect 6823 7131 6873 7160
rect 6823 7107 6837 7131
rect 6861 7107 6873 7131
rect 6823 7083 6873 7107
rect 7031 7136 7081 7160
rect 7031 7112 7046 7136
rect 7070 7112 7081 7136
rect 7031 7083 7081 7112
rect 7244 7131 7294 7160
rect 7244 7111 7261 7131
rect 7281 7111 7294 7131
rect 7244 7083 7294 7111
rect 9110 7130 9160 7155
rect 9110 7104 9116 7130
rect 9142 7104 9160 7130
rect 820 7010 870 7026
rect 1033 7010 1083 7026
rect 1241 7010 1291 7026
rect 1449 7010 1499 7026
rect 1868 7006 1918 7022
rect 2081 7006 2131 7022
rect 2289 7006 2339 7022
rect 2497 7006 2547 7022
rect 9110 7078 9160 7104
rect 9318 7126 9368 7155
rect 9318 7102 9332 7126
rect 9356 7102 9368 7126
rect 9318 7078 9368 7102
rect 9526 7131 9576 7155
rect 9526 7107 9541 7131
rect 9565 7107 9576 7131
rect 9526 7078 9576 7107
rect 9739 7126 9789 7155
rect 9739 7106 9756 7126
rect 9776 7106 9789 7126
rect 9739 7078 9789 7106
rect 6615 6970 6665 6983
rect 6823 6970 6873 6983
rect 7031 6970 7081 6983
rect 7244 6970 7294 6983
rect 9110 6965 9160 6978
rect 9318 6965 9368 6978
rect 9526 6965 9576 6978
rect 9739 6965 9789 6978
rect 820 6566 870 6579
rect 1033 6566 1083 6579
rect 1241 6566 1291 6579
rect 1449 6566 1499 6579
rect 4423 6557 4473 6570
rect 4636 6557 4686 6570
rect 4844 6557 4894 6570
rect 5052 6557 5102 6570
rect 820 6438 870 6466
rect 820 6418 833 6438
rect 853 6418 870 6438
rect 820 6389 870 6418
rect 1033 6437 1083 6466
rect 1033 6413 1044 6437
rect 1068 6413 1083 6437
rect 1033 6389 1083 6413
rect 1241 6442 1291 6466
rect 1241 6418 1253 6442
rect 1277 6418 1291 6442
rect 1241 6389 1291 6418
rect 1449 6440 1499 6466
rect 8062 6522 8112 6538
rect 8270 6522 8320 6538
rect 8478 6522 8528 6538
rect 8691 6522 8741 6538
rect 9110 6518 9160 6534
rect 9318 6518 9368 6534
rect 9526 6518 9576 6534
rect 9739 6518 9789 6534
rect 1449 6414 1467 6440
rect 1493 6414 1499 6440
rect 1449 6389 1499 6414
rect 4423 6429 4473 6457
rect 4423 6409 4436 6429
rect 4456 6409 4473 6429
rect 4423 6380 4473 6409
rect 4636 6428 4686 6457
rect 4636 6404 4647 6428
rect 4671 6404 4686 6428
rect 4636 6380 4686 6404
rect 4844 6433 4894 6457
rect 4844 6409 4856 6433
rect 4880 6409 4894 6433
rect 4844 6380 4894 6409
rect 5052 6431 5102 6457
rect 5052 6405 5070 6431
rect 5096 6405 5102 6431
rect 5052 6380 5102 6405
rect 8062 6455 8112 6480
rect 8062 6429 8068 6455
rect 8094 6429 8112 6455
rect 8062 6403 8112 6429
rect 8270 6451 8320 6480
rect 8270 6427 8284 6451
rect 8308 6427 8320 6451
rect 8270 6403 8320 6427
rect 8478 6456 8528 6480
rect 8478 6432 8493 6456
rect 8517 6432 8528 6456
rect 8478 6403 8528 6432
rect 8691 6451 8741 6480
rect 8691 6431 8708 6451
rect 8728 6431 8741 6451
rect 8691 6403 8741 6431
rect 9110 6451 9160 6476
rect 9110 6425 9116 6451
rect 9142 6425 9160 6451
rect 820 6331 870 6347
rect 1033 6331 1083 6347
rect 1241 6331 1291 6347
rect 1449 6331 1499 6347
rect 4423 6322 4473 6338
rect 4636 6322 4686 6338
rect 4844 6322 4894 6338
rect 5052 6322 5102 6338
rect 9110 6399 9160 6425
rect 9318 6447 9368 6476
rect 9318 6423 9332 6447
rect 9356 6423 9368 6447
rect 9318 6399 9368 6423
rect 9526 6452 9576 6476
rect 9526 6428 9541 6452
rect 9565 6428 9576 6452
rect 9526 6399 9576 6428
rect 9739 6447 9789 6476
rect 9739 6427 9756 6447
rect 9776 6427 9789 6447
rect 9739 6399 9789 6427
rect 8062 6290 8112 6303
rect 8270 6290 8320 6303
rect 8478 6290 8528 6303
rect 8691 6290 8741 6303
rect 9110 6286 9160 6299
rect 9318 6286 9368 6299
rect 9526 6286 9576 6299
rect 9739 6286 9789 6299
rect 817 5651 867 5664
rect 1030 5651 1080 5664
rect 1238 5651 1288 5664
rect 1446 5651 1496 5664
rect 1865 5647 1915 5660
rect 2078 5647 2128 5660
rect 2286 5647 2336 5660
rect 2494 5647 2544 5660
rect 817 5523 867 5551
rect 817 5503 830 5523
rect 850 5503 867 5523
rect 817 5474 867 5503
rect 1030 5522 1080 5551
rect 1030 5498 1041 5522
rect 1065 5498 1080 5522
rect 1030 5474 1080 5498
rect 1238 5527 1288 5551
rect 1238 5503 1250 5527
rect 1274 5503 1288 5527
rect 1238 5474 1288 5503
rect 1446 5525 1496 5551
rect 5504 5612 5554 5628
rect 5712 5612 5762 5628
rect 5920 5612 5970 5628
rect 6133 5612 6183 5628
rect 9107 5603 9157 5619
rect 9315 5603 9365 5619
rect 9523 5603 9573 5619
rect 9736 5603 9786 5619
rect 1446 5499 1464 5525
rect 1490 5499 1496 5525
rect 1446 5474 1496 5499
rect 1865 5519 1915 5547
rect 1865 5499 1878 5519
rect 1898 5499 1915 5519
rect 1865 5470 1915 5499
rect 2078 5518 2128 5547
rect 2078 5494 2089 5518
rect 2113 5494 2128 5518
rect 2078 5470 2128 5494
rect 2286 5523 2336 5547
rect 2286 5499 2298 5523
rect 2322 5499 2336 5523
rect 2286 5470 2336 5499
rect 2494 5521 2544 5547
rect 2494 5495 2512 5521
rect 2538 5495 2544 5521
rect 2494 5470 2544 5495
rect 5504 5545 5554 5570
rect 5504 5519 5510 5545
rect 5536 5519 5554 5545
rect 5504 5493 5554 5519
rect 5712 5541 5762 5570
rect 5712 5517 5726 5541
rect 5750 5517 5762 5541
rect 5712 5493 5762 5517
rect 5920 5546 5970 5570
rect 5920 5522 5935 5546
rect 5959 5522 5970 5546
rect 5920 5493 5970 5522
rect 6133 5541 6183 5570
rect 6133 5521 6150 5541
rect 6170 5521 6183 5541
rect 6133 5493 6183 5521
rect 9107 5536 9157 5561
rect 9107 5510 9113 5536
rect 9139 5510 9157 5536
rect 817 5416 867 5432
rect 1030 5416 1080 5432
rect 1238 5416 1288 5432
rect 1446 5416 1496 5432
rect 1865 5412 1915 5428
rect 2078 5412 2128 5428
rect 2286 5412 2336 5428
rect 2494 5412 2544 5428
rect 9107 5484 9157 5510
rect 9315 5532 9365 5561
rect 9315 5508 9329 5532
rect 9353 5508 9365 5532
rect 9315 5484 9365 5508
rect 9523 5537 9573 5561
rect 9523 5513 9538 5537
rect 9562 5513 9573 5537
rect 9523 5484 9573 5513
rect 9736 5532 9786 5561
rect 9736 5512 9753 5532
rect 9773 5512 9786 5532
rect 9736 5484 9786 5512
rect 5504 5380 5554 5393
rect 5712 5380 5762 5393
rect 5920 5380 5970 5393
rect 6133 5380 6183 5393
rect 9107 5371 9157 5384
rect 9315 5371 9365 5384
rect 9523 5371 9573 5384
rect 9736 5371 9786 5384
rect 817 4972 867 4985
rect 1030 4972 1080 4985
rect 1238 4972 1288 4985
rect 1446 4972 1496 4985
rect 3312 4967 3362 4980
rect 3525 4967 3575 4980
rect 3733 4967 3783 4980
rect 3941 4967 3991 4980
rect 817 4844 867 4872
rect 817 4824 830 4844
rect 850 4824 867 4844
rect 817 4795 867 4824
rect 1030 4843 1080 4872
rect 1030 4819 1041 4843
rect 1065 4819 1080 4843
rect 1030 4795 1080 4819
rect 1238 4848 1288 4872
rect 1238 4824 1250 4848
rect 1274 4824 1288 4848
rect 1238 4795 1288 4824
rect 1446 4846 1496 4872
rect 8059 4928 8109 4944
rect 8267 4928 8317 4944
rect 8475 4928 8525 4944
rect 8688 4928 8738 4944
rect 9107 4924 9157 4940
rect 9315 4924 9365 4940
rect 9523 4924 9573 4940
rect 9736 4924 9786 4940
rect 1446 4820 1464 4846
rect 1490 4820 1496 4846
rect 1446 4795 1496 4820
rect 3312 4839 3362 4867
rect 3312 4819 3325 4839
rect 3345 4819 3362 4839
rect 3312 4790 3362 4819
rect 3525 4838 3575 4867
rect 3525 4814 3536 4838
rect 3560 4814 3575 4838
rect 3525 4790 3575 4814
rect 3733 4843 3783 4867
rect 3733 4819 3745 4843
rect 3769 4819 3783 4843
rect 3733 4790 3783 4819
rect 3941 4841 3991 4867
rect 3941 4815 3959 4841
rect 3985 4815 3991 4841
rect 3941 4790 3991 4815
rect 8059 4861 8109 4886
rect 8059 4835 8065 4861
rect 8091 4835 8109 4861
rect 8059 4809 8109 4835
rect 8267 4857 8317 4886
rect 8267 4833 8281 4857
rect 8305 4833 8317 4857
rect 8267 4809 8317 4833
rect 8475 4862 8525 4886
rect 8475 4838 8490 4862
rect 8514 4838 8525 4862
rect 8475 4809 8525 4838
rect 8688 4857 8738 4886
rect 8688 4837 8705 4857
rect 8725 4837 8738 4857
rect 8688 4809 8738 4837
rect 9107 4857 9157 4882
rect 9107 4831 9113 4857
rect 9139 4831 9157 4857
rect 817 4737 867 4753
rect 1030 4737 1080 4753
rect 1238 4737 1288 4753
rect 1446 4737 1496 4753
rect 3312 4732 3362 4748
rect 3525 4732 3575 4748
rect 3733 4732 3783 4748
rect 3941 4732 3991 4748
rect 9107 4805 9157 4831
rect 9315 4853 9365 4882
rect 9315 4829 9329 4853
rect 9353 4829 9365 4853
rect 9315 4805 9365 4829
rect 9523 4858 9573 4882
rect 9523 4834 9538 4858
rect 9562 4834 9573 4858
rect 9523 4805 9573 4834
rect 9736 4853 9786 4882
rect 9736 4833 9753 4853
rect 9773 4833 9786 4853
rect 9736 4805 9786 4833
rect 8059 4696 8109 4709
rect 8267 4696 8317 4709
rect 8475 4696 8525 4709
rect 8688 4696 8738 4709
rect 9107 4692 9157 4705
rect 9315 4692 9365 4705
rect 9523 4692 9573 4705
rect 9736 4692 9786 4705
rect 817 4204 867 4217
rect 1030 4204 1080 4217
rect 1238 4204 1288 4217
rect 1446 4204 1496 4217
rect 1865 4200 1915 4213
rect 2078 4200 2128 4213
rect 2286 4200 2336 4213
rect 2494 4200 2544 4213
rect 817 4076 867 4104
rect 817 4056 830 4076
rect 850 4056 867 4076
rect 817 4027 867 4056
rect 1030 4075 1080 4104
rect 1030 4051 1041 4075
rect 1065 4051 1080 4075
rect 1030 4027 1080 4051
rect 1238 4080 1288 4104
rect 1238 4056 1250 4080
rect 1274 4056 1288 4080
rect 1238 4027 1288 4056
rect 1446 4078 1496 4104
rect 6612 4161 6662 4177
rect 6820 4161 6870 4177
rect 7028 4161 7078 4177
rect 7241 4161 7291 4177
rect 9107 4156 9157 4172
rect 9315 4156 9365 4172
rect 9523 4156 9573 4172
rect 9736 4156 9786 4172
rect 1446 4052 1464 4078
rect 1490 4052 1496 4078
rect 1446 4027 1496 4052
rect 1865 4072 1915 4100
rect 1865 4052 1878 4072
rect 1898 4052 1915 4072
rect 1865 4023 1915 4052
rect 2078 4071 2128 4100
rect 2078 4047 2089 4071
rect 2113 4047 2128 4071
rect 2078 4023 2128 4047
rect 2286 4076 2336 4100
rect 2286 4052 2298 4076
rect 2322 4052 2336 4076
rect 2286 4023 2336 4052
rect 2494 4074 2544 4100
rect 2494 4048 2512 4074
rect 2538 4048 2544 4074
rect 2494 4023 2544 4048
rect 6612 4094 6662 4119
rect 6612 4068 6618 4094
rect 6644 4068 6662 4094
rect 6612 4042 6662 4068
rect 6820 4090 6870 4119
rect 6820 4066 6834 4090
rect 6858 4066 6870 4090
rect 6820 4042 6870 4066
rect 7028 4095 7078 4119
rect 7028 4071 7043 4095
rect 7067 4071 7078 4095
rect 7028 4042 7078 4071
rect 7241 4090 7291 4119
rect 7241 4070 7258 4090
rect 7278 4070 7291 4090
rect 7241 4042 7291 4070
rect 9107 4089 9157 4114
rect 9107 4063 9113 4089
rect 9139 4063 9157 4089
rect 817 3969 867 3985
rect 1030 3969 1080 3985
rect 1238 3969 1288 3985
rect 1446 3969 1496 3985
rect 1865 3965 1915 3981
rect 2078 3965 2128 3981
rect 2286 3965 2336 3981
rect 2494 3965 2544 3981
rect 9107 4037 9157 4063
rect 9315 4085 9365 4114
rect 9315 4061 9329 4085
rect 9353 4061 9365 4085
rect 9315 4037 9365 4061
rect 9523 4090 9573 4114
rect 9523 4066 9538 4090
rect 9562 4066 9573 4090
rect 9523 4037 9573 4066
rect 9736 4085 9786 4114
rect 9736 4065 9753 4085
rect 9773 4065 9786 4085
rect 9736 4037 9786 4065
rect 6612 3929 6662 3942
rect 6820 3929 6870 3942
rect 7028 3929 7078 3942
rect 7241 3929 7291 3942
rect 9107 3924 9157 3937
rect 9315 3924 9365 3937
rect 9523 3924 9573 3937
rect 9736 3924 9786 3937
rect 817 3525 867 3538
rect 1030 3525 1080 3538
rect 1238 3525 1288 3538
rect 1446 3525 1496 3538
rect 3355 3522 3405 3535
rect 3568 3522 3618 3535
rect 3776 3522 3826 3535
rect 3984 3522 4034 3535
rect 817 3397 867 3425
rect 817 3377 830 3397
rect 850 3377 867 3397
rect 817 3348 867 3377
rect 1030 3396 1080 3425
rect 1030 3372 1041 3396
rect 1065 3372 1080 3396
rect 1030 3348 1080 3372
rect 1238 3401 1288 3425
rect 1238 3377 1250 3401
rect 1274 3377 1288 3401
rect 1238 3348 1288 3377
rect 1446 3399 1496 3425
rect 8059 3481 8109 3497
rect 8267 3481 8317 3497
rect 8475 3481 8525 3497
rect 8688 3481 8738 3497
rect 9107 3477 9157 3493
rect 9315 3477 9365 3493
rect 9523 3477 9573 3493
rect 9736 3477 9786 3493
rect 1446 3373 1464 3399
rect 1490 3373 1496 3399
rect 1446 3348 1496 3373
rect 3355 3394 3405 3422
rect 3355 3374 3368 3394
rect 3388 3374 3405 3394
rect 3355 3345 3405 3374
rect 3568 3393 3618 3422
rect 3568 3369 3579 3393
rect 3603 3369 3618 3393
rect 3568 3345 3618 3369
rect 3776 3398 3826 3422
rect 3776 3374 3788 3398
rect 3812 3374 3826 3398
rect 3776 3345 3826 3374
rect 3984 3396 4034 3422
rect 3984 3370 4002 3396
rect 4028 3370 4034 3396
rect 3984 3345 4034 3370
rect 8059 3414 8109 3439
rect 8059 3388 8065 3414
rect 8091 3388 8109 3414
rect 8059 3362 8109 3388
rect 8267 3410 8317 3439
rect 8267 3386 8281 3410
rect 8305 3386 8317 3410
rect 8267 3362 8317 3386
rect 8475 3415 8525 3439
rect 8475 3391 8490 3415
rect 8514 3391 8525 3415
rect 8475 3362 8525 3391
rect 8688 3410 8738 3439
rect 8688 3390 8705 3410
rect 8725 3390 8738 3410
rect 8688 3362 8738 3390
rect 9107 3410 9157 3435
rect 9107 3384 9113 3410
rect 9139 3384 9157 3410
rect 817 3290 867 3306
rect 1030 3290 1080 3306
rect 1238 3290 1288 3306
rect 1446 3290 1496 3306
rect 3355 3287 3405 3303
rect 3568 3287 3618 3303
rect 3776 3287 3826 3303
rect 3984 3287 4034 3303
rect 9107 3358 9157 3384
rect 9315 3406 9365 3435
rect 9315 3382 9329 3406
rect 9353 3382 9365 3406
rect 9315 3358 9365 3382
rect 9523 3411 9573 3435
rect 9523 3387 9538 3411
rect 9562 3387 9573 3411
rect 9523 3358 9573 3387
rect 9736 3406 9786 3435
rect 9736 3386 9753 3406
rect 9773 3386 9786 3406
rect 9736 3358 9786 3386
rect 8059 3249 8109 3262
rect 8267 3249 8317 3262
rect 8475 3249 8525 3262
rect 8688 3249 8738 3262
rect 9107 3245 9157 3258
rect 9315 3245 9365 3258
rect 9523 3245 9573 3258
rect 9736 3245 9786 3258
rect 818 2684 868 2697
rect 1031 2684 1081 2697
rect 1239 2684 1289 2697
rect 1447 2684 1497 2697
rect 1866 2680 1916 2693
rect 2079 2680 2129 2693
rect 2287 2680 2337 2693
rect 2495 2680 2545 2693
rect 4768 2686 4818 2699
rect 4981 2686 5031 2699
rect 5189 2686 5239 2699
rect 5397 2686 5447 2699
rect 818 2556 868 2584
rect 818 2536 831 2556
rect 851 2536 868 2556
rect 818 2507 868 2536
rect 1031 2555 1081 2584
rect 1031 2531 1042 2555
rect 1066 2531 1081 2555
rect 1031 2507 1081 2531
rect 1239 2560 1289 2584
rect 1239 2536 1251 2560
rect 1275 2536 1289 2560
rect 1239 2507 1289 2536
rect 1447 2558 1497 2584
rect 6570 2639 6620 2655
rect 6778 2639 6828 2655
rect 6986 2639 7036 2655
rect 7199 2639 7249 2655
rect 9108 2636 9158 2652
rect 9316 2636 9366 2652
rect 9524 2636 9574 2652
rect 9737 2636 9787 2652
rect 1447 2532 1465 2558
rect 1491 2532 1497 2558
rect 1447 2507 1497 2532
rect 1866 2552 1916 2580
rect 1866 2532 1879 2552
rect 1899 2532 1916 2552
rect 1866 2503 1916 2532
rect 2079 2551 2129 2580
rect 2079 2527 2090 2551
rect 2114 2527 2129 2551
rect 2079 2503 2129 2527
rect 2287 2556 2337 2580
rect 2287 2532 2299 2556
rect 2323 2532 2337 2556
rect 2287 2503 2337 2532
rect 2495 2554 2545 2580
rect 2495 2528 2513 2554
rect 2539 2528 2545 2554
rect 2495 2503 2545 2528
rect 4768 2558 4818 2586
rect 4768 2538 4781 2558
rect 4801 2538 4818 2558
rect 4768 2509 4818 2538
rect 4981 2557 5031 2586
rect 4981 2533 4992 2557
rect 5016 2533 5031 2557
rect 4981 2509 5031 2533
rect 5189 2562 5239 2586
rect 5189 2538 5201 2562
rect 5225 2538 5239 2562
rect 5189 2509 5239 2538
rect 5397 2560 5447 2586
rect 5397 2534 5415 2560
rect 5441 2534 5447 2560
rect 5397 2509 5447 2534
rect 6570 2572 6620 2597
rect 6570 2546 6576 2572
rect 6602 2546 6620 2572
rect 6570 2520 6620 2546
rect 6778 2568 6828 2597
rect 6778 2544 6792 2568
rect 6816 2544 6828 2568
rect 6778 2520 6828 2544
rect 6986 2573 7036 2597
rect 6986 2549 7001 2573
rect 7025 2549 7036 2573
rect 6986 2520 7036 2549
rect 7199 2568 7249 2597
rect 7199 2548 7216 2568
rect 7236 2548 7249 2568
rect 7199 2520 7249 2548
rect 9108 2569 9158 2594
rect 9108 2543 9114 2569
rect 9140 2543 9158 2569
rect 818 2449 868 2465
rect 1031 2449 1081 2465
rect 1239 2449 1289 2465
rect 1447 2449 1497 2465
rect 1866 2445 1916 2461
rect 2079 2445 2129 2461
rect 2287 2445 2337 2461
rect 2495 2445 2545 2461
rect 4768 2451 4818 2467
rect 4981 2451 5031 2467
rect 5189 2451 5239 2467
rect 5397 2451 5447 2467
rect 9108 2517 9158 2543
rect 9316 2565 9366 2594
rect 9316 2541 9330 2565
rect 9354 2541 9366 2565
rect 9316 2517 9366 2541
rect 9524 2570 9574 2594
rect 9524 2546 9539 2570
rect 9563 2546 9574 2570
rect 9524 2517 9574 2546
rect 9737 2565 9787 2594
rect 9737 2545 9754 2565
rect 9774 2545 9787 2565
rect 9737 2517 9787 2545
rect 6570 2407 6620 2420
rect 6778 2407 6828 2420
rect 6986 2407 7036 2420
rect 7199 2407 7249 2420
rect 9108 2404 9158 2417
rect 9316 2404 9366 2417
rect 9524 2404 9574 2417
rect 9737 2404 9787 2417
rect 818 2005 868 2018
rect 1031 2005 1081 2018
rect 1239 2005 1289 2018
rect 1447 2005 1497 2018
rect 3313 2000 3363 2013
rect 3526 2000 3576 2013
rect 3734 2000 3784 2013
rect 3942 2000 3992 2013
rect 818 1877 868 1905
rect 818 1857 831 1877
rect 851 1857 868 1877
rect 818 1828 868 1857
rect 1031 1876 1081 1905
rect 1031 1852 1042 1876
rect 1066 1852 1081 1876
rect 1031 1828 1081 1852
rect 1239 1881 1289 1905
rect 1239 1857 1251 1881
rect 1275 1857 1289 1881
rect 1239 1828 1289 1857
rect 1447 1879 1497 1905
rect 8060 1961 8110 1977
rect 8268 1961 8318 1977
rect 8476 1961 8526 1977
rect 8689 1961 8739 1977
rect 9108 1957 9158 1973
rect 9316 1957 9366 1973
rect 9524 1957 9574 1973
rect 9737 1957 9787 1973
rect 1447 1853 1465 1879
rect 1491 1853 1497 1879
rect 1447 1828 1497 1853
rect 3313 1872 3363 1900
rect 3313 1852 3326 1872
rect 3346 1852 3363 1872
rect 3313 1823 3363 1852
rect 3526 1871 3576 1900
rect 3526 1847 3537 1871
rect 3561 1847 3576 1871
rect 3526 1823 3576 1847
rect 3734 1876 3784 1900
rect 3734 1852 3746 1876
rect 3770 1852 3784 1876
rect 3734 1823 3784 1852
rect 3942 1874 3992 1900
rect 3942 1848 3960 1874
rect 3986 1848 3992 1874
rect 3942 1823 3992 1848
rect 8060 1894 8110 1919
rect 8060 1868 8066 1894
rect 8092 1868 8110 1894
rect 8060 1842 8110 1868
rect 8268 1890 8318 1919
rect 8268 1866 8282 1890
rect 8306 1866 8318 1890
rect 8268 1842 8318 1866
rect 8476 1895 8526 1919
rect 8476 1871 8491 1895
rect 8515 1871 8526 1895
rect 8476 1842 8526 1871
rect 8689 1890 8739 1919
rect 8689 1870 8706 1890
rect 8726 1870 8739 1890
rect 8689 1842 8739 1870
rect 9108 1890 9158 1915
rect 9108 1864 9114 1890
rect 9140 1864 9158 1890
rect 818 1770 868 1786
rect 1031 1770 1081 1786
rect 1239 1770 1289 1786
rect 1447 1770 1497 1786
rect 3313 1765 3363 1781
rect 3526 1765 3576 1781
rect 3734 1765 3784 1781
rect 3942 1765 3992 1781
rect 9108 1838 9158 1864
rect 9316 1886 9366 1915
rect 9316 1862 9330 1886
rect 9354 1862 9366 1886
rect 9316 1838 9366 1862
rect 9524 1891 9574 1915
rect 9524 1867 9539 1891
rect 9563 1867 9574 1891
rect 9524 1838 9574 1867
rect 9737 1886 9787 1915
rect 9737 1866 9754 1886
rect 9774 1866 9787 1886
rect 9737 1838 9787 1866
rect 8060 1729 8110 1742
rect 8268 1729 8318 1742
rect 8476 1729 8526 1742
rect 8689 1729 8739 1742
rect 9108 1725 9158 1738
rect 9316 1725 9366 1738
rect 9524 1725 9574 1738
rect 9737 1725 9787 1738
rect 818 1237 868 1250
rect 1031 1237 1081 1250
rect 1239 1237 1289 1250
rect 1447 1237 1497 1250
rect 1866 1233 1916 1246
rect 2079 1233 2129 1246
rect 2287 1233 2337 1246
rect 2495 1233 2545 1246
rect 818 1109 868 1137
rect 818 1089 831 1109
rect 851 1089 868 1109
rect 818 1060 868 1089
rect 1031 1108 1081 1137
rect 1031 1084 1042 1108
rect 1066 1084 1081 1108
rect 1031 1060 1081 1084
rect 1239 1113 1289 1137
rect 1239 1089 1251 1113
rect 1275 1089 1289 1113
rect 1239 1060 1289 1089
rect 1447 1111 1497 1137
rect 6613 1194 6663 1210
rect 6821 1194 6871 1210
rect 7029 1194 7079 1210
rect 7242 1194 7292 1210
rect 9108 1189 9158 1205
rect 9316 1189 9366 1205
rect 9524 1189 9574 1205
rect 9737 1189 9787 1205
rect 1447 1085 1465 1111
rect 1491 1085 1497 1111
rect 1447 1060 1497 1085
rect 1866 1105 1916 1133
rect 1866 1085 1879 1105
rect 1899 1085 1916 1105
rect 1866 1056 1916 1085
rect 2079 1104 2129 1133
rect 2079 1080 2090 1104
rect 2114 1080 2129 1104
rect 2079 1056 2129 1080
rect 2287 1109 2337 1133
rect 2287 1085 2299 1109
rect 2323 1085 2337 1109
rect 2287 1056 2337 1085
rect 2495 1107 2545 1133
rect 2495 1081 2513 1107
rect 2539 1081 2545 1107
rect 2495 1056 2545 1081
rect 6613 1127 6663 1152
rect 6613 1101 6619 1127
rect 6645 1101 6663 1127
rect 6613 1075 6663 1101
rect 6821 1123 6871 1152
rect 6821 1099 6835 1123
rect 6859 1099 6871 1123
rect 6821 1075 6871 1099
rect 7029 1128 7079 1152
rect 7029 1104 7044 1128
rect 7068 1104 7079 1128
rect 7029 1075 7079 1104
rect 7242 1123 7292 1152
rect 7242 1103 7259 1123
rect 7279 1103 7292 1123
rect 7242 1075 7292 1103
rect 9108 1122 9158 1147
rect 9108 1096 9114 1122
rect 9140 1096 9158 1122
rect 818 1002 868 1018
rect 1031 1002 1081 1018
rect 1239 1002 1289 1018
rect 1447 1002 1497 1018
rect 1866 998 1916 1014
rect 2079 998 2129 1014
rect 2287 998 2337 1014
rect 2495 998 2545 1014
rect 9108 1070 9158 1096
rect 9316 1118 9366 1147
rect 9316 1094 9330 1118
rect 9354 1094 9366 1118
rect 9316 1070 9366 1094
rect 9524 1123 9574 1147
rect 9524 1099 9539 1123
rect 9563 1099 9574 1123
rect 9524 1070 9574 1099
rect 9737 1118 9787 1147
rect 9737 1098 9754 1118
rect 9774 1098 9787 1118
rect 9737 1070 9787 1098
rect 6613 962 6663 975
rect 6821 962 6871 975
rect 7029 962 7079 975
rect 7242 962 7292 975
rect 9108 957 9158 970
rect 9316 957 9366 970
rect 9524 957 9574 970
rect 9737 957 9787 970
rect 818 558 868 571
rect 1031 558 1081 571
rect 1239 558 1289 571
rect 1447 558 1497 571
rect 8060 514 8110 530
rect 8268 514 8318 530
rect 8476 514 8526 530
rect 8689 514 8739 530
rect 9108 510 9158 526
rect 9316 510 9366 526
rect 9524 510 9574 526
rect 9737 510 9787 526
rect 818 430 868 458
rect 818 410 831 430
rect 851 410 868 430
rect 818 381 868 410
rect 1031 429 1081 458
rect 1031 405 1042 429
rect 1066 405 1081 429
rect 1031 381 1081 405
rect 1239 434 1289 458
rect 1239 410 1251 434
rect 1275 410 1289 434
rect 1239 381 1289 410
rect 1447 432 1497 458
rect 1447 406 1465 432
rect 1491 406 1497 432
rect 1447 381 1497 406
rect 8060 447 8110 472
rect 8060 421 8066 447
rect 8092 421 8110 447
rect 8060 395 8110 421
rect 8268 443 8318 472
rect 8268 419 8282 443
rect 8306 419 8318 443
rect 8268 395 8318 419
rect 8476 448 8526 472
rect 8476 424 8491 448
rect 8515 424 8526 448
rect 8476 395 8526 424
rect 8689 443 8739 472
rect 8689 423 8706 443
rect 8726 423 8739 443
rect 8689 395 8739 423
rect 9108 443 9158 468
rect 9108 417 9114 443
rect 9140 417 9158 443
rect 818 323 868 339
rect 1031 323 1081 339
rect 1239 323 1289 339
rect 1447 323 1497 339
rect 9108 391 9158 417
rect 9316 439 9366 468
rect 9316 415 9330 439
rect 9354 415 9366 439
rect 9316 391 9366 415
rect 9524 444 9574 468
rect 9524 420 9539 444
rect 9563 420 9574 444
rect 9524 391 9574 420
rect 9737 439 9787 468
rect 9737 419 9754 439
rect 9774 419 9787 439
rect 9737 391 9787 419
rect 8060 282 8110 295
rect 8268 282 8318 295
rect 8476 282 8526 295
rect 8689 282 8739 295
rect 9108 278 9158 291
rect 9316 278 9366 291
rect 9524 278 9574 291
rect 9737 278 9787 291
<< polycont >>
rect 832 11511 852 11531
rect 1043 11506 1067 11530
rect 1252 11511 1276 11535
rect 1466 11507 1492 11533
rect 1880 11507 1900 11527
rect 2091 11502 2115 11526
rect 2300 11507 2324 11531
rect 2514 11503 2540 11529
rect 9115 11518 9141 11544
rect 9331 11516 9355 11540
rect 9540 11521 9564 11545
rect 9755 11520 9775 11540
rect 832 10832 852 10852
rect 1043 10827 1067 10851
rect 1252 10832 1276 10856
rect 1466 10828 1492 10854
rect 3327 10827 3347 10847
rect 3538 10822 3562 10846
rect 3747 10827 3771 10851
rect 3961 10823 3987 10849
rect 8067 10843 8093 10869
rect 8283 10841 8307 10865
rect 8492 10846 8516 10870
rect 8707 10845 8727 10865
rect 9115 10839 9141 10865
rect 9331 10837 9355 10861
rect 9540 10842 9564 10866
rect 9755 10841 9775 10861
rect 832 10064 852 10084
rect 1043 10059 1067 10083
rect 1252 10064 1276 10088
rect 1466 10060 1492 10086
rect 1880 10060 1900 10080
rect 2091 10055 2115 10079
rect 2300 10060 2324 10084
rect 2514 10056 2540 10082
rect 6620 10076 6646 10102
rect 6836 10074 6860 10098
rect 7045 10079 7069 10103
rect 7260 10078 7280 10098
rect 9115 10071 9141 10097
rect 9331 10069 9355 10093
rect 9540 10074 9564 10098
rect 9755 10073 9775 10093
rect 832 9385 852 9405
rect 1043 9380 1067 9404
rect 1252 9385 1276 9409
rect 1466 9381 1492 9407
rect 3370 9382 3390 9402
rect 3581 9377 3605 9401
rect 3790 9382 3814 9406
rect 4004 9378 4030 9404
rect 8067 9396 8093 9422
rect 8283 9394 8307 9418
rect 8492 9399 8516 9423
rect 8707 9398 8727 9418
rect 9115 9392 9141 9418
rect 9331 9390 9355 9414
rect 9540 9395 9564 9419
rect 9755 9394 9775 9414
rect 833 8544 853 8564
rect 1044 8539 1068 8563
rect 1253 8544 1277 8568
rect 1467 8540 1493 8566
rect 1881 8540 1901 8560
rect 2092 8535 2116 8559
rect 2301 8540 2325 8564
rect 2515 8536 2541 8562
rect 6578 8554 6604 8580
rect 6794 8552 6818 8576
rect 7003 8557 7027 8581
rect 7218 8556 7238 8576
rect 9116 8551 9142 8577
rect 9332 8549 9356 8573
rect 9541 8554 9565 8578
rect 9756 8553 9776 8573
rect 833 7865 853 7885
rect 1044 7860 1068 7884
rect 1253 7865 1277 7889
rect 1467 7861 1493 7887
rect 3328 7860 3348 7880
rect 3539 7855 3563 7879
rect 3748 7860 3772 7884
rect 3962 7856 3988 7882
rect 8068 7876 8094 7902
rect 8284 7874 8308 7898
rect 8493 7879 8517 7903
rect 8708 7878 8728 7898
rect 9116 7872 9142 7898
rect 9332 7870 9356 7894
rect 9541 7875 9565 7899
rect 9756 7874 9776 7894
rect 833 7097 853 7117
rect 1044 7092 1068 7116
rect 1253 7097 1277 7121
rect 1467 7093 1493 7119
rect 1881 7093 1901 7113
rect 2092 7088 2116 7112
rect 2301 7093 2325 7117
rect 2515 7089 2541 7115
rect 6621 7109 6647 7135
rect 6837 7107 6861 7131
rect 7046 7112 7070 7136
rect 7261 7111 7281 7131
rect 9116 7104 9142 7130
rect 9332 7102 9356 7126
rect 9541 7107 9565 7131
rect 9756 7106 9776 7126
rect 833 6418 853 6438
rect 1044 6413 1068 6437
rect 1253 6418 1277 6442
rect 1467 6414 1493 6440
rect 4436 6409 4456 6429
rect 4647 6404 4671 6428
rect 4856 6409 4880 6433
rect 5070 6405 5096 6431
rect 8068 6429 8094 6455
rect 8284 6427 8308 6451
rect 8493 6432 8517 6456
rect 8708 6431 8728 6451
rect 9116 6425 9142 6451
rect 9332 6423 9356 6447
rect 9541 6428 9565 6452
rect 9756 6427 9776 6447
rect 830 5503 850 5523
rect 1041 5498 1065 5522
rect 1250 5503 1274 5527
rect 1464 5499 1490 5525
rect 1878 5499 1898 5519
rect 2089 5494 2113 5518
rect 2298 5499 2322 5523
rect 2512 5495 2538 5521
rect 5510 5519 5536 5545
rect 5726 5517 5750 5541
rect 5935 5522 5959 5546
rect 6150 5521 6170 5541
rect 9113 5510 9139 5536
rect 9329 5508 9353 5532
rect 9538 5513 9562 5537
rect 9753 5512 9773 5532
rect 830 4824 850 4844
rect 1041 4819 1065 4843
rect 1250 4824 1274 4848
rect 1464 4820 1490 4846
rect 3325 4819 3345 4839
rect 3536 4814 3560 4838
rect 3745 4819 3769 4843
rect 3959 4815 3985 4841
rect 8065 4835 8091 4861
rect 8281 4833 8305 4857
rect 8490 4838 8514 4862
rect 8705 4837 8725 4857
rect 9113 4831 9139 4857
rect 9329 4829 9353 4853
rect 9538 4834 9562 4858
rect 9753 4833 9773 4853
rect 830 4056 850 4076
rect 1041 4051 1065 4075
rect 1250 4056 1274 4080
rect 1464 4052 1490 4078
rect 1878 4052 1898 4072
rect 2089 4047 2113 4071
rect 2298 4052 2322 4076
rect 2512 4048 2538 4074
rect 6618 4068 6644 4094
rect 6834 4066 6858 4090
rect 7043 4071 7067 4095
rect 7258 4070 7278 4090
rect 9113 4063 9139 4089
rect 9329 4061 9353 4085
rect 9538 4066 9562 4090
rect 9753 4065 9773 4085
rect 830 3377 850 3397
rect 1041 3372 1065 3396
rect 1250 3377 1274 3401
rect 1464 3373 1490 3399
rect 3368 3374 3388 3394
rect 3579 3369 3603 3393
rect 3788 3374 3812 3398
rect 4002 3370 4028 3396
rect 8065 3388 8091 3414
rect 8281 3386 8305 3410
rect 8490 3391 8514 3415
rect 8705 3390 8725 3410
rect 9113 3384 9139 3410
rect 9329 3382 9353 3406
rect 9538 3387 9562 3411
rect 9753 3386 9773 3406
rect 831 2536 851 2556
rect 1042 2531 1066 2555
rect 1251 2536 1275 2560
rect 1465 2532 1491 2558
rect 1879 2532 1899 2552
rect 2090 2527 2114 2551
rect 2299 2532 2323 2556
rect 2513 2528 2539 2554
rect 4781 2538 4801 2558
rect 4992 2533 5016 2557
rect 5201 2538 5225 2562
rect 5415 2534 5441 2560
rect 6576 2546 6602 2572
rect 6792 2544 6816 2568
rect 7001 2549 7025 2573
rect 7216 2548 7236 2568
rect 9114 2543 9140 2569
rect 9330 2541 9354 2565
rect 9539 2546 9563 2570
rect 9754 2545 9774 2565
rect 831 1857 851 1877
rect 1042 1852 1066 1876
rect 1251 1857 1275 1881
rect 1465 1853 1491 1879
rect 3326 1852 3346 1872
rect 3537 1847 3561 1871
rect 3746 1852 3770 1876
rect 3960 1848 3986 1874
rect 8066 1868 8092 1894
rect 8282 1866 8306 1890
rect 8491 1871 8515 1895
rect 8706 1870 8726 1890
rect 9114 1864 9140 1890
rect 9330 1862 9354 1886
rect 9539 1867 9563 1891
rect 9754 1866 9774 1886
rect 831 1089 851 1109
rect 1042 1084 1066 1108
rect 1251 1089 1275 1113
rect 1465 1085 1491 1111
rect 1879 1085 1899 1105
rect 2090 1080 2114 1104
rect 2299 1085 2323 1109
rect 2513 1081 2539 1107
rect 6619 1101 6645 1127
rect 6835 1099 6859 1123
rect 7044 1104 7068 1128
rect 7259 1103 7279 1123
rect 9114 1096 9140 1122
rect 9330 1094 9354 1118
rect 9539 1099 9563 1123
rect 9754 1098 9774 1118
rect 831 410 851 430
rect 1042 405 1066 429
rect 1251 410 1275 434
rect 1465 406 1491 432
rect 8066 421 8092 447
rect 8282 419 8306 443
rect 8491 424 8515 448
rect 8706 423 8726 443
rect 9114 417 9140 443
rect 9330 415 9354 439
rect 9539 420 9563 444
rect 9754 419 9774 439
<< ndiffres >>
rect 440 11793 497 11812
rect 440 11790 461 11793
rect 346 11775 461 11790
rect 479 11775 497 11793
rect 346 11752 497 11775
rect 346 11716 388 11752
rect 345 11715 445 11716
rect 345 11694 501 11715
rect 345 11676 463 11694
rect 481 11676 501 11694
rect 345 11672 501 11676
rect 440 11656 501 11672
rect 440 11537 497 11556
rect 440 11534 461 11537
rect 346 11519 461 11534
rect 479 11519 497 11537
rect 346 11496 497 11519
rect 346 11460 388 11496
rect 10106 11606 10167 11622
rect 10106 11602 10262 11606
rect 10106 11584 10126 11602
rect 10144 11584 10262 11602
rect 345 11459 445 11460
rect 345 11438 501 11459
rect 10106 11563 10262 11584
rect 10162 11562 10262 11563
rect 10219 11526 10261 11562
rect 10110 11503 10261 11526
rect 345 11420 463 11438
rect 481 11420 501 11438
rect 345 11416 501 11420
rect 440 11400 501 11416
rect 10110 11485 10128 11503
rect 10146 11488 10261 11503
rect 10146 11485 10167 11488
rect 10110 11466 10167 11485
rect 10106 11351 10167 11367
rect 10106 11347 10262 11351
rect 10106 11329 10126 11347
rect 10144 11329 10262 11347
rect 10106 11308 10262 11329
rect 10162 11307 10262 11308
rect 10219 11271 10261 11307
rect 10110 11248 10261 11271
rect 10110 11230 10128 11248
rect 10146 11233 10261 11248
rect 10146 11230 10167 11233
rect 10110 11211 10167 11230
rect 440 11142 497 11161
rect 440 11139 461 11142
rect 346 11124 461 11139
rect 479 11124 497 11142
rect 346 11101 497 11124
rect 346 11065 388 11101
rect 345 11064 445 11065
rect 345 11043 501 11064
rect 345 11025 463 11043
rect 481 11025 501 11043
rect 345 11021 501 11025
rect 440 11005 501 11021
rect 440 10887 497 10906
rect 440 10884 461 10887
rect 346 10869 461 10884
rect 479 10869 497 10887
rect 346 10846 497 10869
rect 346 10810 388 10846
rect 345 10809 445 10810
rect 345 10788 501 10809
rect 10106 10956 10167 10972
rect 10106 10952 10262 10956
rect 10106 10934 10126 10952
rect 10144 10934 10262 10952
rect 345 10770 463 10788
rect 481 10770 501 10788
rect 345 10766 501 10770
rect 440 10750 501 10766
rect 10106 10913 10262 10934
rect 10162 10912 10262 10913
rect 10219 10876 10261 10912
rect 10110 10853 10261 10876
rect 10110 10835 10128 10853
rect 10146 10838 10261 10853
rect 10146 10835 10167 10838
rect 10110 10816 10167 10835
rect 10106 10700 10167 10716
rect 10106 10696 10262 10700
rect 10106 10678 10126 10696
rect 10144 10678 10262 10696
rect 10106 10657 10262 10678
rect 10162 10656 10262 10657
rect 10219 10620 10261 10656
rect 10110 10597 10261 10620
rect 10110 10579 10128 10597
rect 10146 10582 10261 10597
rect 10146 10579 10167 10582
rect 10110 10560 10167 10579
rect 440 10346 497 10365
rect 440 10343 461 10346
rect 346 10328 461 10343
rect 479 10328 497 10346
rect 346 10305 497 10328
rect 346 10269 388 10305
rect 345 10268 445 10269
rect 345 10247 501 10268
rect 345 10229 463 10247
rect 481 10229 501 10247
rect 345 10225 501 10229
rect 440 10209 501 10225
rect 440 10090 497 10109
rect 440 10087 461 10090
rect 346 10072 461 10087
rect 479 10072 497 10090
rect 346 10049 497 10072
rect 346 10013 388 10049
rect 345 10012 445 10013
rect 345 9991 501 10012
rect 10106 10159 10167 10175
rect 10106 10155 10262 10159
rect 10106 10137 10126 10155
rect 10144 10137 10262 10155
rect 345 9973 463 9991
rect 481 9973 501 9991
rect 345 9969 501 9973
rect 440 9953 501 9969
rect 10106 10116 10262 10137
rect 10162 10115 10262 10116
rect 10219 10079 10261 10115
rect 10110 10056 10261 10079
rect 10110 10038 10128 10056
rect 10146 10041 10261 10056
rect 10146 10038 10167 10041
rect 10110 10019 10167 10038
rect 10106 9904 10167 9920
rect 10106 9900 10262 9904
rect 10106 9882 10126 9900
rect 10144 9882 10262 9900
rect 10106 9861 10262 9882
rect 10162 9860 10262 9861
rect 10219 9824 10261 9860
rect 10110 9801 10261 9824
rect 10110 9783 10128 9801
rect 10146 9786 10261 9801
rect 10146 9783 10167 9786
rect 10110 9764 10167 9783
rect 440 9695 497 9714
rect 440 9692 461 9695
rect 346 9677 461 9692
rect 479 9677 497 9695
rect 346 9654 497 9677
rect 346 9618 388 9654
rect 345 9617 445 9618
rect 345 9596 501 9617
rect 345 9578 463 9596
rect 481 9578 501 9596
rect 345 9574 501 9578
rect 440 9558 501 9574
rect 440 9440 497 9459
rect 440 9437 461 9440
rect 346 9422 461 9437
rect 479 9422 497 9440
rect 346 9399 497 9422
rect 346 9363 388 9399
rect 345 9362 445 9363
rect 345 9341 501 9362
rect 10106 9509 10167 9525
rect 10106 9505 10262 9509
rect 10106 9487 10126 9505
rect 10144 9487 10262 9505
rect 345 9323 463 9341
rect 481 9323 501 9341
rect 345 9319 501 9323
rect 440 9303 501 9319
rect 10106 9466 10262 9487
rect 10162 9465 10262 9466
rect 10219 9429 10261 9465
rect 10110 9406 10261 9429
rect 10110 9388 10128 9406
rect 10146 9391 10261 9406
rect 10146 9388 10167 9391
rect 10110 9369 10167 9388
rect 10106 9253 10167 9269
rect 10106 9249 10262 9253
rect 10106 9231 10126 9249
rect 10144 9231 10262 9249
rect 10106 9210 10262 9231
rect 10162 9209 10262 9210
rect 10219 9173 10261 9209
rect 10110 9150 10261 9173
rect 10110 9132 10128 9150
rect 10146 9135 10261 9150
rect 10146 9132 10167 9135
rect 10110 9113 10167 9132
rect 441 8826 498 8845
rect 441 8823 462 8826
rect 347 8808 462 8823
rect 480 8808 498 8826
rect 347 8785 498 8808
rect 347 8749 389 8785
rect 346 8748 446 8749
rect 346 8727 502 8748
rect 346 8709 464 8727
rect 482 8709 502 8727
rect 346 8705 502 8709
rect 441 8689 502 8705
rect 441 8570 498 8589
rect 441 8567 462 8570
rect 347 8552 462 8567
rect 480 8552 498 8570
rect 347 8529 498 8552
rect 347 8493 389 8529
rect 346 8492 446 8493
rect 346 8471 502 8492
rect 10107 8639 10168 8655
rect 10107 8635 10263 8639
rect 10107 8617 10127 8635
rect 10145 8617 10263 8635
rect 346 8453 464 8471
rect 482 8453 502 8471
rect 346 8449 502 8453
rect 441 8433 502 8449
rect 10107 8596 10263 8617
rect 10163 8595 10263 8596
rect 10220 8559 10262 8595
rect 10111 8536 10262 8559
rect 10111 8518 10129 8536
rect 10147 8521 10262 8536
rect 10147 8518 10168 8521
rect 10111 8499 10168 8518
rect 10107 8384 10168 8400
rect 10107 8380 10263 8384
rect 10107 8362 10127 8380
rect 10145 8362 10263 8380
rect 10107 8341 10263 8362
rect 10163 8340 10263 8341
rect 10220 8304 10262 8340
rect 10111 8281 10262 8304
rect 10111 8263 10129 8281
rect 10147 8266 10262 8281
rect 10147 8263 10168 8266
rect 10111 8244 10168 8263
rect 441 8175 498 8194
rect 441 8172 462 8175
rect 347 8157 462 8172
rect 480 8157 498 8175
rect 347 8134 498 8157
rect 347 8098 389 8134
rect 346 8097 446 8098
rect 346 8076 502 8097
rect 346 8058 464 8076
rect 482 8058 502 8076
rect 346 8054 502 8058
rect 441 8038 502 8054
rect 441 7920 498 7939
rect 441 7917 462 7920
rect 347 7902 462 7917
rect 480 7902 498 7920
rect 347 7879 498 7902
rect 347 7843 389 7879
rect 346 7842 446 7843
rect 346 7821 502 7842
rect 10107 7989 10168 8005
rect 10107 7985 10263 7989
rect 10107 7967 10127 7985
rect 10145 7967 10263 7985
rect 346 7803 464 7821
rect 482 7803 502 7821
rect 346 7799 502 7803
rect 441 7783 502 7799
rect 10107 7946 10263 7967
rect 10163 7945 10263 7946
rect 10220 7909 10262 7945
rect 10111 7886 10262 7909
rect 10111 7868 10129 7886
rect 10147 7871 10262 7886
rect 10147 7868 10168 7871
rect 10111 7849 10168 7868
rect 10107 7733 10168 7749
rect 10107 7729 10263 7733
rect 10107 7711 10127 7729
rect 10145 7711 10263 7729
rect 10107 7690 10263 7711
rect 10163 7689 10263 7690
rect 10220 7653 10262 7689
rect 10111 7630 10262 7653
rect 10111 7612 10129 7630
rect 10147 7615 10262 7630
rect 10147 7612 10168 7615
rect 10111 7593 10168 7612
rect 441 7379 498 7398
rect 441 7376 462 7379
rect 347 7361 462 7376
rect 480 7361 498 7379
rect 347 7338 498 7361
rect 347 7302 389 7338
rect 346 7301 446 7302
rect 346 7280 502 7301
rect 346 7262 464 7280
rect 482 7262 502 7280
rect 346 7258 502 7262
rect 441 7242 502 7258
rect 441 7123 498 7142
rect 441 7120 462 7123
rect 347 7105 462 7120
rect 480 7105 498 7123
rect 347 7082 498 7105
rect 347 7046 389 7082
rect 346 7045 446 7046
rect 346 7024 502 7045
rect 10107 7192 10168 7208
rect 10107 7188 10263 7192
rect 10107 7170 10127 7188
rect 10145 7170 10263 7188
rect 346 7006 464 7024
rect 482 7006 502 7024
rect 346 7002 502 7006
rect 441 6986 502 7002
rect 10107 7149 10263 7170
rect 10163 7148 10263 7149
rect 10220 7112 10262 7148
rect 10111 7089 10262 7112
rect 10111 7071 10129 7089
rect 10147 7074 10262 7089
rect 10147 7071 10168 7074
rect 10111 7052 10168 7071
rect 10107 6937 10168 6953
rect 10107 6933 10263 6937
rect 10107 6915 10127 6933
rect 10145 6915 10263 6933
rect 10107 6894 10263 6915
rect 10163 6893 10263 6894
rect 10220 6857 10262 6893
rect 10111 6834 10262 6857
rect 10111 6816 10129 6834
rect 10147 6819 10262 6834
rect 10147 6816 10168 6819
rect 10111 6797 10168 6816
rect 441 6728 498 6747
rect 441 6725 462 6728
rect 347 6710 462 6725
rect 480 6710 498 6728
rect 347 6687 498 6710
rect 347 6651 389 6687
rect 346 6650 446 6651
rect 346 6629 502 6650
rect 346 6611 464 6629
rect 482 6611 502 6629
rect 346 6607 502 6611
rect 441 6591 502 6607
rect 441 6473 498 6492
rect 441 6470 462 6473
rect 347 6455 462 6470
rect 480 6455 498 6473
rect 347 6432 498 6455
rect 347 6396 389 6432
rect 346 6395 446 6396
rect 346 6374 502 6395
rect 10107 6542 10168 6558
rect 10107 6538 10263 6542
rect 10107 6520 10127 6538
rect 10145 6520 10263 6538
rect 346 6356 464 6374
rect 482 6356 502 6374
rect 346 6352 502 6356
rect 441 6336 502 6352
rect 10107 6499 10263 6520
rect 10163 6498 10263 6499
rect 10220 6462 10262 6498
rect 10111 6439 10262 6462
rect 10111 6421 10129 6439
rect 10147 6424 10262 6439
rect 10147 6421 10168 6424
rect 10111 6402 10168 6421
rect 10107 6286 10168 6302
rect 10107 6282 10263 6286
rect 10107 6264 10127 6282
rect 10145 6264 10263 6282
rect 10107 6243 10263 6264
rect 10163 6242 10263 6243
rect 10220 6206 10262 6242
rect 10111 6183 10262 6206
rect 10111 6165 10129 6183
rect 10147 6168 10262 6183
rect 10147 6165 10168 6168
rect 10111 6146 10168 6165
rect 438 5785 495 5804
rect 438 5782 459 5785
rect 344 5767 459 5782
rect 477 5767 495 5785
rect 344 5744 495 5767
rect 344 5708 386 5744
rect 343 5707 443 5708
rect 343 5686 499 5707
rect 343 5668 461 5686
rect 479 5668 499 5686
rect 343 5664 499 5668
rect 438 5648 499 5664
rect 438 5529 495 5548
rect 438 5526 459 5529
rect 344 5511 459 5526
rect 477 5511 495 5529
rect 344 5488 495 5511
rect 344 5452 386 5488
rect 343 5451 443 5452
rect 343 5430 499 5451
rect 10104 5598 10165 5614
rect 10104 5594 10260 5598
rect 10104 5576 10124 5594
rect 10142 5576 10260 5594
rect 343 5412 461 5430
rect 479 5412 499 5430
rect 343 5408 499 5412
rect 438 5392 499 5408
rect 10104 5555 10260 5576
rect 10160 5554 10260 5555
rect 10217 5518 10259 5554
rect 10108 5495 10259 5518
rect 10108 5477 10126 5495
rect 10144 5480 10259 5495
rect 10144 5477 10165 5480
rect 10108 5458 10165 5477
rect 10104 5343 10165 5359
rect 10104 5339 10260 5343
rect 10104 5321 10124 5339
rect 10142 5321 10260 5339
rect 10104 5300 10260 5321
rect 10160 5299 10260 5300
rect 10217 5263 10259 5299
rect 10108 5240 10259 5263
rect 10108 5222 10126 5240
rect 10144 5225 10259 5240
rect 10144 5222 10165 5225
rect 10108 5203 10165 5222
rect 438 5134 495 5153
rect 438 5131 459 5134
rect 344 5116 459 5131
rect 477 5116 495 5134
rect 344 5093 495 5116
rect 344 5057 386 5093
rect 343 5056 443 5057
rect 343 5035 499 5056
rect 343 5017 461 5035
rect 479 5017 499 5035
rect 343 5013 499 5017
rect 438 4997 499 5013
rect 438 4879 495 4898
rect 438 4876 459 4879
rect 344 4861 459 4876
rect 477 4861 495 4879
rect 344 4838 495 4861
rect 344 4802 386 4838
rect 343 4801 443 4802
rect 343 4780 499 4801
rect 10104 4948 10165 4964
rect 10104 4944 10260 4948
rect 10104 4926 10124 4944
rect 10142 4926 10260 4944
rect 343 4762 461 4780
rect 479 4762 499 4780
rect 343 4758 499 4762
rect 438 4742 499 4758
rect 10104 4905 10260 4926
rect 10160 4904 10260 4905
rect 10217 4868 10259 4904
rect 10108 4845 10259 4868
rect 10108 4827 10126 4845
rect 10144 4830 10259 4845
rect 10144 4827 10165 4830
rect 10108 4808 10165 4827
rect 10104 4692 10165 4708
rect 10104 4688 10260 4692
rect 10104 4670 10124 4688
rect 10142 4670 10260 4688
rect 10104 4649 10260 4670
rect 10160 4648 10260 4649
rect 10217 4612 10259 4648
rect 10108 4589 10259 4612
rect 10108 4571 10126 4589
rect 10144 4574 10259 4589
rect 10144 4571 10165 4574
rect 10108 4552 10165 4571
rect 438 4338 495 4357
rect 438 4335 459 4338
rect 344 4320 459 4335
rect 477 4320 495 4338
rect 344 4297 495 4320
rect 344 4261 386 4297
rect 343 4260 443 4261
rect 343 4239 499 4260
rect 343 4221 461 4239
rect 479 4221 499 4239
rect 343 4217 499 4221
rect 438 4201 499 4217
rect 438 4082 495 4101
rect 438 4079 459 4082
rect 344 4064 459 4079
rect 477 4064 495 4082
rect 344 4041 495 4064
rect 344 4005 386 4041
rect 343 4004 443 4005
rect 343 3983 499 4004
rect 10104 4151 10165 4167
rect 10104 4147 10260 4151
rect 10104 4129 10124 4147
rect 10142 4129 10260 4147
rect 343 3965 461 3983
rect 479 3965 499 3983
rect 343 3961 499 3965
rect 438 3945 499 3961
rect 10104 4108 10260 4129
rect 10160 4107 10260 4108
rect 10217 4071 10259 4107
rect 10108 4048 10259 4071
rect 10108 4030 10126 4048
rect 10144 4033 10259 4048
rect 10144 4030 10165 4033
rect 10108 4011 10165 4030
rect 10104 3896 10165 3912
rect 10104 3892 10260 3896
rect 10104 3874 10124 3892
rect 10142 3874 10260 3892
rect 10104 3853 10260 3874
rect 10160 3852 10260 3853
rect 10217 3816 10259 3852
rect 10108 3793 10259 3816
rect 10108 3775 10126 3793
rect 10144 3778 10259 3793
rect 10144 3775 10165 3778
rect 10108 3756 10165 3775
rect 438 3687 495 3706
rect 438 3684 459 3687
rect 344 3669 459 3684
rect 477 3669 495 3687
rect 344 3646 495 3669
rect 344 3610 386 3646
rect 343 3609 443 3610
rect 343 3588 499 3609
rect 343 3570 461 3588
rect 479 3570 499 3588
rect 343 3566 499 3570
rect 438 3550 499 3566
rect 438 3432 495 3451
rect 438 3429 459 3432
rect 344 3414 459 3429
rect 477 3414 495 3432
rect 344 3391 495 3414
rect 344 3355 386 3391
rect 343 3354 443 3355
rect 343 3333 499 3354
rect 10104 3501 10165 3517
rect 10104 3497 10260 3501
rect 10104 3479 10124 3497
rect 10142 3479 10260 3497
rect 343 3315 461 3333
rect 479 3315 499 3333
rect 343 3311 499 3315
rect 438 3295 499 3311
rect 10104 3458 10260 3479
rect 10160 3457 10260 3458
rect 10217 3421 10259 3457
rect 10108 3398 10259 3421
rect 10108 3380 10126 3398
rect 10144 3383 10259 3398
rect 10144 3380 10165 3383
rect 10108 3361 10165 3380
rect 10104 3245 10165 3261
rect 10104 3241 10260 3245
rect 10104 3223 10124 3241
rect 10142 3223 10260 3241
rect 10104 3202 10260 3223
rect 10160 3201 10260 3202
rect 10217 3165 10259 3201
rect 10108 3142 10259 3165
rect 10108 3124 10126 3142
rect 10144 3127 10259 3142
rect 10144 3124 10165 3127
rect 10108 3105 10165 3124
rect 439 2818 496 2837
rect 439 2815 460 2818
rect 345 2800 460 2815
rect 478 2800 496 2818
rect 345 2777 496 2800
rect 345 2741 387 2777
rect 344 2740 444 2741
rect 344 2719 500 2740
rect 344 2701 462 2719
rect 480 2701 500 2719
rect 344 2697 500 2701
rect 439 2681 500 2697
rect 439 2562 496 2581
rect 439 2559 460 2562
rect 345 2544 460 2559
rect 478 2544 496 2562
rect 345 2521 496 2544
rect 345 2485 387 2521
rect 344 2484 444 2485
rect 344 2463 500 2484
rect 10105 2631 10166 2647
rect 10105 2627 10261 2631
rect 10105 2609 10125 2627
rect 10143 2609 10261 2627
rect 344 2445 462 2463
rect 480 2445 500 2463
rect 344 2441 500 2445
rect 439 2425 500 2441
rect 10105 2588 10261 2609
rect 10161 2587 10261 2588
rect 10218 2551 10260 2587
rect 10109 2528 10260 2551
rect 10109 2510 10127 2528
rect 10145 2513 10260 2528
rect 10145 2510 10166 2513
rect 10109 2491 10166 2510
rect 10105 2376 10166 2392
rect 10105 2372 10261 2376
rect 10105 2354 10125 2372
rect 10143 2354 10261 2372
rect 10105 2333 10261 2354
rect 10161 2332 10261 2333
rect 10218 2296 10260 2332
rect 10109 2273 10260 2296
rect 10109 2255 10127 2273
rect 10145 2258 10260 2273
rect 10145 2255 10166 2258
rect 10109 2236 10166 2255
rect 439 2167 496 2186
rect 439 2164 460 2167
rect 345 2149 460 2164
rect 478 2149 496 2167
rect 345 2126 496 2149
rect 345 2090 387 2126
rect 344 2089 444 2090
rect 344 2068 500 2089
rect 344 2050 462 2068
rect 480 2050 500 2068
rect 344 2046 500 2050
rect 439 2030 500 2046
rect 439 1912 496 1931
rect 439 1909 460 1912
rect 345 1894 460 1909
rect 478 1894 496 1912
rect 345 1871 496 1894
rect 345 1835 387 1871
rect 344 1834 444 1835
rect 344 1813 500 1834
rect 10105 1981 10166 1997
rect 10105 1977 10261 1981
rect 10105 1959 10125 1977
rect 10143 1959 10261 1977
rect 344 1795 462 1813
rect 480 1795 500 1813
rect 344 1791 500 1795
rect 439 1775 500 1791
rect 10105 1938 10261 1959
rect 10161 1937 10261 1938
rect 10218 1901 10260 1937
rect 10109 1878 10260 1901
rect 10109 1860 10127 1878
rect 10145 1863 10260 1878
rect 10145 1860 10166 1863
rect 10109 1841 10166 1860
rect 10105 1725 10166 1741
rect 10105 1721 10261 1725
rect 10105 1703 10125 1721
rect 10143 1703 10261 1721
rect 10105 1682 10261 1703
rect 10161 1681 10261 1682
rect 10218 1645 10260 1681
rect 10109 1622 10260 1645
rect 10109 1604 10127 1622
rect 10145 1607 10260 1622
rect 10145 1604 10166 1607
rect 10109 1585 10166 1604
rect 439 1371 496 1390
rect 439 1368 460 1371
rect 345 1353 460 1368
rect 478 1353 496 1371
rect 345 1330 496 1353
rect 345 1294 387 1330
rect 344 1293 444 1294
rect 344 1272 500 1293
rect 344 1254 462 1272
rect 480 1254 500 1272
rect 344 1250 500 1254
rect 439 1234 500 1250
rect 439 1115 496 1134
rect 439 1112 460 1115
rect 345 1097 460 1112
rect 478 1097 496 1115
rect 345 1074 496 1097
rect 345 1038 387 1074
rect 344 1037 444 1038
rect 344 1016 500 1037
rect 10105 1184 10166 1200
rect 10105 1180 10261 1184
rect 10105 1162 10125 1180
rect 10143 1162 10261 1180
rect 344 998 462 1016
rect 480 998 500 1016
rect 344 994 500 998
rect 439 978 500 994
rect 10105 1141 10261 1162
rect 10161 1140 10261 1141
rect 10218 1104 10260 1140
rect 10109 1081 10260 1104
rect 10109 1063 10127 1081
rect 10145 1066 10260 1081
rect 10145 1063 10166 1066
rect 10109 1044 10166 1063
rect 10105 929 10166 945
rect 10105 925 10261 929
rect 10105 907 10125 925
rect 10143 907 10261 925
rect 10105 886 10261 907
rect 10161 885 10261 886
rect 10218 849 10260 885
rect 10109 826 10260 849
rect 10109 808 10127 826
rect 10145 811 10260 826
rect 10145 808 10166 811
rect 10109 789 10166 808
rect 439 720 496 739
rect 439 717 460 720
rect 345 702 460 717
rect 478 702 496 720
rect 345 679 496 702
rect 345 643 387 679
rect 344 642 444 643
rect 344 621 500 642
rect 344 603 462 621
rect 480 603 500 621
rect 344 599 500 603
rect 439 583 500 599
rect 439 465 496 484
rect 439 462 460 465
rect 345 447 460 462
rect 478 447 496 465
rect 10105 534 10166 550
rect 10105 530 10261 534
rect 10105 512 10125 530
rect 10143 512 10261 530
rect 345 424 496 447
rect 345 388 387 424
rect 344 387 444 388
rect 344 366 500 387
rect 10105 491 10261 512
rect 10161 490 10261 491
rect 344 348 462 366
rect 480 348 500 366
rect 344 344 500 348
rect 439 328 500 344
rect 10218 454 10260 490
rect 10109 431 10260 454
rect 10109 413 10127 431
rect 10145 416 10260 431
rect 10145 413 10166 416
rect 10109 394 10166 413
rect 10105 278 10166 294
rect 10105 274 10261 278
rect 10105 256 10125 274
rect 10143 256 10261 274
rect 10105 235 10261 256
rect 10161 234 10261 235
rect 10218 198 10260 234
rect 10109 175 10260 198
rect 10109 157 10127 175
rect 10145 160 10260 175
rect 10145 157 10166 160
rect 10109 138 10166 157
<< locali >>
rect 439 11793 498 12176
rect 2816 12167 2881 12178
rect 2816 12119 2829 12167
rect 2866 12119 2881 12167
rect 2816 12106 2881 12119
rect 3029 11876 3740 11878
rect 2402 11875 3740 11876
rect 1352 11874 1424 11875
rect 1351 11866 1450 11874
rect 1351 11863 1403 11866
rect 1351 11828 1359 11863
rect 1384 11828 1403 11863
rect 1428 11855 1450 11866
rect 2401 11867 3740 11875
rect 2401 11864 2453 11867
rect 1428 11854 2295 11855
rect 1428 11828 2296 11854
rect 1351 11818 2296 11828
rect 1351 11816 1450 11818
rect 439 11775 461 11793
rect 479 11775 498 11793
rect 439 11753 498 11775
rect 706 11789 1238 11794
rect 706 11769 1592 11789
rect 1612 11769 1615 11789
rect 2251 11785 2296 11818
rect 2401 11829 2409 11864
rect 2434 11829 2453 11864
rect 2478 11829 3740 11867
rect 2401 11820 3740 11829
rect 2401 11817 2490 11820
rect 3029 11818 3740 11820
rect 706 11765 1615 11769
rect 706 11718 749 11765
rect 1199 11764 1615 11765
rect 2247 11765 2640 11785
rect 2660 11765 2663 11785
rect 1199 11763 1540 11764
rect 856 11732 966 11746
rect 856 11729 899 11732
rect 856 11724 860 11729
rect 694 11717 749 11718
rect 438 11694 749 11717
rect 438 11676 463 11694
rect 481 11682 749 11694
rect 778 11702 860 11724
rect 889 11702 899 11729
rect 927 11705 934 11732
rect 963 11724 966 11732
rect 963 11705 1028 11724
rect 927 11702 1028 11705
rect 778 11700 1028 11702
rect 481 11676 503 11682
rect 438 11537 503 11676
rect 778 11621 815 11700
rect 856 11687 966 11700
rect 930 11631 961 11632
rect 778 11601 787 11621
rect 807 11601 815 11621
rect 438 11519 461 11537
rect 479 11519 503 11537
rect 438 11502 503 11519
rect 658 11583 726 11596
rect 778 11591 815 11601
rect 874 11621 961 11631
rect 874 11601 883 11621
rect 903 11601 961 11621
rect 874 11592 961 11601
rect 874 11591 911 11592
rect 658 11541 665 11583
rect 714 11541 726 11583
rect 658 11538 726 11541
rect 930 11539 961 11592
rect 991 11621 1028 11700
rect 1143 11631 1174 11632
rect 991 11601 1000 11621
rect 1020 11601 1028 11621
rect 991 11591 1028 11601
rect 1087 11624 1174 11631
rect 1087 11621 1148 11624
rect 1087 11601 1096 11621
rect 1116 11604 1148 11621
rect 1169 11604 1174 11624
rect 1116 11601 1174 11604
rect 1087 11594 1174 11601
rect 1199 11621 1236 11763
rect 1502 11762 1539 11763
rect 2247 11760 2663 11765
rect 2247 11759 2588 11760
rect 1904 11728 2014 11742
rect 1904 11725 1947 11728
rect 1904 11720 1908 11725
rect 1826 11698 1908 11720
rect 1937 11698 1947 11725
rect 1975 11701 1982 11728
rect 2011 11720 2014 11728
rect 2011 11701 2076 11720
rect 1975 11698 2076 11701
rect 1826 11696 2076 11698
rect 1351 11631 1387 11632
rect 1199 11601 1208 11621
rect 1228 11601 1236 11621
rect 1087 11592 1143 11594
rect 1087 11591 1124 11592
rect 1199 11591 1236 11601
rect 1295 11621 1443 11631
rect 1543 11628 1639 11630
rect 1295 11601 1304 11621
rect 1324 11601 1414 11621
rect 1434 11601 1443 11621
rect 1295 11595 1443 11601
rect 1295 11592 1359 11595
rect 1295 11591 1332 11592
rect 1351 11565 1359 11592
rect 1380 11592 1443 11595
rect 1501 11621 1639 11628
rect 1501 11601 1510 11621
rect 1530 11601 1639 11621
rect 1501 11592 1639 11601
rect 1826 11617 1863 11696
rect 1904 11683 2014 11696
rect 1978 11627 2009 11628
rect 1826 11597 1835 11617
rect 1855 11597 1863 11617
rect 1380 11565 1387 11592
rect 1406 11591 1443 11592
rect 1502 11591 1539 11592
rect 1351 11540 1387 11565
rect 822 11538 863 11539
rect 658 11531 863 11538
rect 658 11520 832 11531
rect 658 11487 666 11520
rect 659 11478 666 11487
rect 715 11511 832 11520
rect 852 11511 863 11531
rect 715 11503 863 11511
rect 930 11535 1289 11539
rect 930 11530 1252 11535
rect 930 11506 1043 11530
rect 1067 11511 1252 11530
rect 1276 11511 1289 11535
rect 1067 11506 1289 11511
rect 930 11503 1289 11506
rect 1351 11503 1386 11540
rect 1454 11537 1554 11540
rect 1454 11533 1521 11537
rect 1454 11507 1466 11533
rect 1492 11511 1521 11533
rect 1547 11511 1554 11537
rect 1492 11507 1554 11511
rect 1454 11503 1554 11507
rect 715 11487 726 11503
rect 715 11478 723 11487
rect 930 11482 961 11503
rect 1351 11482 1387 11503
rect 773 11481 810 11482
rect 438 11438 503 11457
rect 438 11420 463 11438
rect 481 11420 503 11438
rect 438 11219 503 11420
rect 659 11294 723 11478
rect 772 11472 810 11481
rect 772 11452 781 11472
rect 801 11452 810 11472
rect 772 11444 810 11452
rect 876 11476 961 11482
rect 986 11481 1023 11482
rect 876 11456 884 11476
rect 904 11456 961 11476
rect 876 11448 961 11456
rect 985 11472 1023 11481
rect 985 11452 994 11472
rect 1014 11452 1023 11472
rect 876 11447 912 11448
rect 985 11444 1023 11452
rect 1089 11476 1174 11482
rect 1194 11481 1231 11482
rect 1089 11456 1097 11476
rect 1117 11475 1174 11476
rect 1117 11456 1146 11475
rect 1089 11455 1146 11456
rect 1167 11455 1174 11475
rect 1089 11448 1174 11455
rect 1193 11472 1231 11481
rect 1193 11452 1202 11472
rect 1222 11452 1231 11472
rect 1089 11447 1125 11448
rect 1193 11444 1231 11452
rect 1297 11476 1441 11482
rect 1297 11456 1305 11476
rect 1325 11456 1413 11476
rect 1433 11456 1441 11476
rect 1297 11448 1441 11456
rect 1297 11447 1333 11448
rect 1405 11447 1441 11448
rect 1507 11481 1544 11482
rect 1507 11480 1545 11481
rect 1507 11472 1571 11480
rect 1507 11452 1516 11472
rect 1536 11458 1571 11472
rect 1591 11458 1594 11478
rect 1536 11453 1594 11458
rect 1536 11452 1571 11453
rect 773 11415 810 11444
rect 774 11413 810 11415
rect 986 11413 1023 11444
rect 774 11391 1023 11413
rect 855 11385 966 11391
rect 855 11377 896 11385
rect 855 11357 863 11377
rect 882 11357 896 11377
rect 855 11355 896 11357
rect 924 11377 966 11385
rect 924 11357 940 11377
rect 959 11357 966 11377
rect 924 11355 966 11357
rect 855 11340 966 11355
rect 659 11284 727 11294
rect 659 11251 676 11284
rect 716 11251 727 11284
rect 659 11239 727 11251
rect 659 11237 723 11239
rect 1194 11220 1231 11444
rect 1507 11440 1571 11452
rect 1611 11222 1638 11592
rect 1826 11587 1863 11597
rect 1922 11617 2009 11627
rect 1922 11597 1931 11617
rect 1951 11597 2009 11617
rect 1922 11588 2009 11597
rect 1922 11587 1959 11588
rect 1702 11574 1772 11579
rect 1697 11568 1772 11574
rect 1697 11535 1705 11568
rect 1758 11535 1772 11568
rect 1978 11535 2009 11588
rect 2039 11617 2076 11696
rect 2191 11627 2222 11628
rect 2039 11597 2048 11617
rect 2068 11597 2076 11617
rect 2039 11587 2076 11597
rect 2135 11620 2222 11627
rect 2135 11617 2196 11620
rect 2135 11597 2144 11617
rect 2164 11600 2196 11617
rect 2217 11600 2222 11620
rect 2164 11597 2222 11600
rect 2135 11590 2222 11597
rect 2247 11617 2284 11759
rect 2550 11758 2587 11759
rect 2399 11627 2435 11628
rect 2247 11597 2256 11617
rect 2276 11597 2284 11617
rect 2135 11588 2191 11590
rect 2135 11587 2172 11588
rect 2247 11587 2284 11597
rect 2343 11617 2491 11627
rect 2591 11624 2687 11626
rect 2343 11597 2352 11617
rect 2372 11597 2462 11617
rect 2482 11597 2491 11617
rect 2343 11591 2491 11597
rect 2343 11588 2407 11591
rect 2343 11587 2380 11588
rect 2399 11561 2407 11588
rect 2428 11588 2491 11591
rect 2549 11617 2687 11624
rect 2549 11597 2558 11617
rect 2578 11597 2687 11617
rect 2549 11588 2687 11597
rect 2428 11561 2435 11588
rect 2454 11587 2491 11588
rect 2550 11587 2587 11588
rect 2399 11536 2435 11561
rect 1697 11534 1780 11535
rect 1870 11534 1911 11535
rect 1697 11527 1911 11534
rect 1697 11510 1880 11527
rect 1697 11477 1710 11510
rect 1763 11507 1880 11510
rect 1900 11507 1911 11527
rect 1763 11499 1911 11507
rect 1978 11531 2337 11535
rect 1978 11526 2300 11531
rect 1978 11502 2091 11526
rect 2115 11507 2300 11526
rect 2324 11507 2337 11531
rect 2115 11502 2337 11507
rect 1978 11499 2337 11502
rect 2399 11499 2434 11536
rect 2502 11533 2602 11536
rect 2502 11529 2569 11533
rect 2502 11503 2514 11529
rect 2540 11507 2569 11529
rect 2595 11507 2602 11533
rect 2540 11503 2602 11507
rect 2502 11499 2602 11503
rect 1763 11477 1780 11499
rect 1978 11478 2009 11499
rect 2399 11478 2435 11499
rect 1821 11477 1858 11478
rect 1697 11463 1780 11477
rect 1470 11220 1638 11222
rect 1194 11219 1638 11220
rect 438 11189 1638 11219
rect 1708 11253 1780 11463
rect 1820 11468 1858 11477
rect 1820 11448 1829 11468
rect 1849 11448 1858 11468
rect 1820 11440 1858 11448
rect 1924 11472 2009 11478
rect 2034 11477 2071 11478
rect 1924 11452 1932 11472
rect 1952 11452 2009 11472
rect 1924 11444 2009 11452
rect 2033 11468 2071 11477
rect 2033 11448 2042 11468
rect 2062 11448 2071 11468
rect 1924 11443 1960 11444
rect 2033 11440 2071 11448
rect 2137 11472 2222 11478
rect 2242 11477 2279 11478
rect 2137 11452 2145 11472
rect 2165 11471 2222 11472
rect 2165 11452 2194 11471
rect 2137 11451 2194 11452
rect 2215 11451 2222 11471
rect 2137 11444 2222 11451
rect 2241 11468 2279 11477
rect 2241 11448 2250 11468
rect 2270 11448 2279 11468
rect 2137 11443 2173 11444
rect 2241 11440 2279 11448
rect 2345 11472 2489 11478
rect 2345 11452 2353 11472
rect 2373 11452 2461 11472
rect 2481 11452 2489 11472
rect 2345 11444 2489 11452
rect 2345 11443 2381 11444
rect 2453 11443 2489 11444
rect 2555 11477 2592 11478
rect 2555 11476 2593 11477
rect 2555 11468 2619 11476
rect 2555 11448 2564 11468
rect 2584 11454 2619 11468
rect 2639 11454 2642 11474
rect 2584 11449 2642 11454
rect 2584 11448 2619 11449
rect 1821 11411 1858 11440
rect 1822 11409 1858 11411
rect 2034 11409 2071 11440
rect 1822 11387 2071 11409
rect 1903 11381 2014 11387
rect 1903 11373 1944 11381
rect 1903 11353 1911 11373
rect 1930 11353 1944 11373
rect 1903 11351 1944 11353
rect 1972 11373 2014 11381
rect 1972 11353 1988 11373
rect 2007 11353 2014 11373
rect 1972 11351 2014 11353
rect 1903 11336 2014 11351
rect 1708 11214 1727 11253
rect 1772 11214 1780 11253
rect 1708 11197 1780 11214
rect 2242 11241 2279 11440
rect 2555 11436 2619 11448
rect 2242 11235 2283 11241
rect 2659 11237 2686 11588
rect 2981 11575 3076 11601
rect 2817 11553 2881 11572
rect 2817 11514 2830 11553
rect 2864 11514 2881 11553
rect 2817 11495 2881 11514
rect 2518 11235 2686 11237
rect 2242 11209 2686 11235
rect 438 11142 503 11189
rect 438 11124 461 11142
rect 479 11124 503 11142
rect 1351 11169 1386 11171
rect 1351 11167 1455 11169
rect 2244 11167 2283 11209
rect 2518 11208 2686 11209
rect 1351 11160 2285 11167
rect 1351 11159 1402 11160
rect 1351 11139 1354 11159
rect 1379 11140 1402 11159
rect 1434 11140 2285 11160
rect 1379 11139 2285 11140
rect 1351 11132 2285 11139
rect 1624 11131 2285 11132
rect 438 11103 503 11124
rect 715 11114 755 11117
rect 715 11110 1618 11114
rect 715 11090 1592 11110
rect 1612 11090 1618 11110
rect 715 11087 1618 11090
rect 439 11043 504 11063
rect 439 11025 463 11043
rect 481 11025 504 11043
rect 439 10998 504 11025
rect 715 10998 755 11087
rect 1199 11085 1615 11087
rect 1199 11084 1540 11085
rect 856 11053 966 11067
rect 856 11050 899 11053
rect 856 11045 860 11050
rect 438 10963 755 10998
rect 778 11023 860 11045
rect 889 11023 899 11050
rect 927 11026 934 11053
rect 963 11045 966 11053
rect 963 11026 1028 11045
rect 927 11023 1028 11026
rect 778 11021 1028 11023
rect 439 10887 504 10963
rect 778 10942 815 11021
rect 856 11008 966 11021
rect 930 10952 961 10953
rect 778 10922 787 10942
rect 807 10922 815 10942
rect 778 10912 815 10922
rect 874 10942 961 10952
rect 874 10922 883 10942
rect 903 10922 961 10942
rect 874 10913 961 10922
rect 874 10912 911 10913
rect 439 10869 461 10887
rect 479 10869 504 10887
rect 439 10848 504 10869
rect 652 10867 717 10876
rect 652 10830 662 10867
rect 702 10859 717 10867
rect 930 10860 961 10913
rect 991 10942 1028 11021
rect 1143 10952 1174 10953
rect 991 10922 1000 10942
rect 1020 10922 1028 10942
rect 991 10912 1028 10922
rect 1087 10945 1174 10952
rect 1087 10942 1148 10945
rect 1087 10922 1096 10942
rect 1116 10925 1148 10942
rect 1169 10925 1174 10945
rect 1116 10922 1174 10925
rect 1087 10915 1174 10922
rect 1199 10942 1236 11084
rect 1502 11083 1539 11084
rect 2819 11024 2881 11495
rect 2981 11534 3007 11575
rect 3043 11534 3076 11575
rect 2981 11238 3076 11534
rect 2981 11194 2996 11238
rect 3056 11194 3076 11238
rect 2981 11174 3076 11194
rect 3693 11105 3736 11818
rect 5547 11708 5685 11740
rect 5547 11641 5579 11708
rect 5665 11641 5685 11708
rect 8835 11644 8905 11897
rect 9374 11894 9415 11896
rect 9646 11894 9750 11896
rect 8967 11892 10161 11894
rect 8967 11859 10163 11892
rect 8967 11845 8995 11859
rect 8969 11714 8995 11845
rect 9374 11856 10163 11859
rect 5547 11614 5685 11641
rect 3693 11085 4087 11105
rect 4107 11085 4110 11105
rect 3694 11080 4110 11085
rect 3694 11079 4035 11080
rect 3351 11048 3461 11062
rect 3351 11045 3394 11048
rect 3351 11040 3355 11045
rect 2814 10972 2889 11024
rect 3273 11018 3355 11040
rect 3384 11018 3394 11045
rect 3422 11021 3429 11048
rect 3458 11040 3461 11048
rect 3458 11021 3523 11040
rect 3422 11018 3523 11021
rect 3273 11016 3523 11018
rect 3183 10972 3229 10973
rect 1351 10952 1387 10953
rect 1199 10922 1208 10942
rect 1228 10922 1236 10942
rect 1087 10913 1143 10915
rect 1087 10912 1124 10913
rect 1199 10912 1236 10922
rect 1295 10942 1443 10952
rect 1543 10949 1639 10951
rect 1295 10922 1304 10942
rect 1324 10922 1414 10942
rect 1434 10922 1443 10942
rect 1295 10916 1443 10922
rect 1295 10913 1359 10916
rect 1295 10912 1332 10913
rect 1351 10886 1359 10913
rect 1380 10913 1443 10916
rect 1501 10942 1639 10949
rect 1501 10922 1510 10942
rect 1530 10922 1639 10942
rect 1501 10913 1639 10922
rect 2814 10937 3229 10972
rect 1380 10886 1387 10913
rect 1406 10912 1443 10913
rect 1502 10912 1539 10913
rect 1351 10861 1387 10886
rect 822 10859 863 10860
rect 702 10852 863 10859
rect 702 10832 832 10852
rect 852 10832 863 10852
rect 702 10830 863 10832
rect 652 10824 863 10830
rect 930 10856 1289 10860
rect 930 10851 1252 10856
rect 930 10827 1043 10851
rect 1067 10832 1252 10851
rect 1276 10832 1289 10856
rect 1067 10827 1289 10832
rect 930 10824 1289 10827
rect 1351 10824 1386 10861
rect 1454 10858 1554 10861
rect 1454 10854 1521 10858
rect 1454 10828 1466 10854
rect 1492 10832 1521 10854
rect 1547 10832 1554 10858
rect 1492 10828 1554 10832
rect 1454 10824 1554 10828
rect 652 10811 719 10824
rect 444 10788 500 10808
rect 444 10770 463 10788
rect 481 10770 500 10788
rect 444 10657 500 10770
rect 652 10790 666 10811
rect 702 10790 719 10811
rect 930 10803 961 10824
rect 1351 10803 1387 10824
rect 773 10802 810 10803
rect 652 10783 719 10790
rect 772 10793 810 10802
rect 444 10519 499 10657
rect 652 10631 717 10783
rect 772 10773 781 10793
rect 801 10773 810 10793
rect 772 10765 810 10773
rect 876 10797 961 10803
rect 986 10802 1023 10803
rect 876 10777 884 10797
rect 904 10777 961 10797
rect 876 10769 961 10777
rect 985 10793 1023 10802
rect 985 10773 994 10793
rect 1014 10773 1023 10793
rect 876 10768 912 10769
rect 985 10765 1023 10773
rect 1089 10797 1174 10803
rect 1194 10802 1231 10803
rect 1089 10777 1097 10797
rect 1117 10796 1174 10797
rect 1117 10777 1146 10796
rect 1089 10776 1146 10777
rect 1167 10776 1174 10796
rect 1089 10769 1174 10776
rect 1193 10793 1231 10802
rect 1193 10773 1202 10793
rect 1222 10773 1231 10793
rect 1089 10768 1125 10769
rect 1193 10765 1231 10773
rect 1297 10797 1441 10803
rect 1297 10777 1305 10797
rect 1325 10777 1413 10797
rect 1433 10777 1441 10797
rect 1297 10769 1441 10777
rect 1297 10768 1333 10769
rect 1405 10768 1441 10769
rect 1507 10802 1544 10803
rect 1507 10801 1545 10802
rect 1507 10793 1571 10801
rect 1507 10773 1516 10793
rect 1536 10779 1571 10793
rect 1591 10779 1594 10799
rect 1536 10774 1594 10779
rect 1536 10773 1571 10774
rect 773 10736 810 10765
rect 774 10734 810 10736
rect 986 10734 1023 10765
rect 774 10712 1023 10734
rect 855 10706 966 10712
rect 855 10698 896 10706
rect 855 10678 863 10698
rect 882 10678 896 10698
rect 855 10676 896 10678
rect 924 10698 966 10706
rect 924 10678 940 10698
rect 959 10678 966 10698
rect 924 10676 966 10678
rect 855 10663 966 10676
rect 1194 10666 1231 10765
rect 1507 10761 1571 10773
rect 645 10621 766 10631
rect 645 10619 714 10621
rect 645 10578 658 10619
rect 695 10580 714 10619
rect 751 10580 766 10621
rect 695 10578 766 10580
rect 645 10560 766 10578
rect 437 10516 501 10519
rect 857 10516 961 10522
rect 1192 10516 1233 10666
rect 1611 10658 1638 10913
rect 1700 10903 1780 10914
rect 1700 10877 1717 10903
rect 1757 10877 1780 10903
rect 1700 10850 1780 10877
rect 1700 10824 1721 10850
rect 1761 10824 1780 10850
rect 1700 10805 1780 10824
rect 1700 10779 1724 10805
rect 1764 10779 1780 10805
rect 1700 10728 1780 10779
rect 437 10513 1233 10516
rect 1612 10527 1638 10658
rect 1612 10513 1640 10527
rect 437 10478 1640 10513
rect 1702 10520 1772 10728
rect 2814 10653 2889 10937
rect 3183 10854 3229 10937
rect 3273 10937 3310 11016
rect 3351 11003 3461 11016
rect 3425 10947 3456 10948
rect 3273 10917 3282 10937
rect 3302 10917 3310 10937
rect 3273 10907 3310 10917
rect 3369 10937 3456 10947
rect 3369 10917 3378 10937
rect 3398 10917 3456 10937
rect 3369 10908 3456 10917
rect 3369 10907 3406 10908
rect 3425 10855 3456 10908
rect 3486 10937 3523 11016
rect 3638 10947 3669 10948
rect 3486 10917 3495 10937
rect 3515 10917 3523 10937
rect 3486 10907 3523 10917
rect 3582 10940 3669 10947
rect 3582 10937 3643 10940
rect 3582 10917 3591 10937
rect 3611 10920 3643 10937
rect 3664 10920 3669 10940
rect 3611 10917 3669 10920
rect 3582 10910 3669 10917
rect 3694 10937 3731 11079
rect 3997 11078 4034 11079
rect 3846 10947 3882 10948
rect 3694 10917 3703 10937
rect 3723 10917 3731 10937
rect 3582 10908 3638 10910
rect 3582 10907 3619 10908
rect 3694 10907 3731 10917
rect 3790 10937 3938 10947
rect 4038 10944 4134 10946
rect 3790 10917 3799 10937
rect 3819 10917 3909 10937
rect 3929 10917 3938 10937
rect 3790 10911 3938 10917
rect 3790 10908 3854 10911
rect 3790 10907 3827 10908
rect 3846 10881 3854 10908
rect 3875 10908 3938 10911
rect 3996 10937 4134 10944
rect 3996 10917 4005 10937
rect 4025 10917 4134 10937
rect 3996 10908 4134 10917
rect 3875 10881 3882 10908
rect 3901 10907 3938 10908
rect 3997 10907 4034 10908
rect 3846 10856 3882 10881
rect 3317 10854 3358 10855
rect 3183 10847 3358 10854
rect 2981 10821 3067 10840
rect 2981 10780 2996 10821
rect 3050 10780 3067 10821
rect 3183 10827 3327 10847
rect 3347 10827 3358 10847
rect 3183 10819 3358 10827
rect 3425 10851 3784 10855
rect 3425 10846 3747 10851
rect 3425 10822 3538 10846
rect 3562 10827 3747 10846
rect 3771 10827 3784 10851
rect 3562 10822 3784 10827
rect 3425 10819 3784 10822
rect 3846 10819 3881 10856
rect 3949 10853 4049 10856
rect 3949 10849 4016 10853
rect 3949 10823 3961 10849
rect 3987 10827 4016 10849
rect 4042 10827 4049 10853
rect 3987 10823 4049 10827
rect 3949 10819 4049 10823
rect 3183 10815 3229 10819
rect 3425 10798 3456 10819
rect 3846 10798 3882 10819
rect 3268 10797 3305 10798
rect 2981 10744 3067 10780
rect 3267 10788 3305 10797
rect 3267 10768 3276 10788
rect 3296 10768 3305 10788
rect 3267 10760 3305 10768
rect 3371 10792 3456 10798
rect 3481 10797 3518 10798
rect 3371 10772 3379 10792
rect 3399 10772 3456 10792
rect 3371 10764 3456 10772
rect 3480 10788 3518 10797
rect 3480 10768 3489 10788
rect 3509 10768 3518 10788
rect 3371 10763 3407 10764
rect 3480 10760 3518 10768
rect 3584 10792 3669 10798
rect 3689 10797 3726 10798
rect 3584 10772 3592 10792
rect 3612 10791 3669 10792
rect 3612 10772 3641 10791
rect 3584 10771 3641 10772
rect 3662 10771 3669 10791
rect 3584 10764 3669 10771
rect 3688 10788 3726 10797
rect 3688 10768 3697 10788
rect 3717 10768 3726 10788
rect 3584 10763 3620 10764
rect 3688 10760 3726 10768
rect 3792 10792 3936 10798
rect 3792 10772 3800 10792
rect 3820 10772 3908 10792
rect 3928 10772 3936 10792
rect 3792 10764 3936 10772
rect 3792 10763 3828 10764
rect 437 10417 501 10478
rect 857 10476 961 10478
rect 1192 10476 1233 10478
rect 1702 10475 1723 10520
rect 1703 10454 1723 10475
rect 1753 10475 1772 10520
rect 2809 10611 2889 10653
rect 1753 10454 1770 10475
rect 1703 10435 1770 10454
rect 1352 10427 1424 10428
rect 1351 10419 1450 10427
rect 439 10346 498 10417
rect 1351 10416 1403 10419
rect 1351 10381 1359 10416
rect 1384 10381 1403 10416
rect 1428 10408 1450 10419
rect 1428 10407 2295 10408
rect 1428 10381 2296 10407
rect 1351 10371 2296 10381
rect 1351 10369 1450 10371
rect 439 10328 461 10346
rect 479 10328 498 10346
rect 439 10306 498 10328
rect 706 10342 1238 10347
rect 706 10322 1592 10342
rect 1612 10322 1615 10342
rect 2251 10338 2296 10371
rect 706 10318 1615 10322
rect 706 10271 749 10318
rect 1199 10317 1615 10318
rect 2247 10318 2640 10338
rect 2660 10318 2663 10338
rect 1199 10316 1540 10317
rect 856 10285 966 10299
rect 856 10282 899 10285
rect 856 10277 860 10282
rect 694 10270 749 10271
rect 438 10247 749 10270
rect 438 10229 463 10247
rect 481 10235 749 10247
rect 778 10255 860 10277
rect 889 10255 899 10282
rect 927 10258 934 10285
rect 963 10277 966 10285
rect 963 10258 1028 10277
rect 927 10255 1028 10258
rect 778 10253 1028 10255
rect 481 10229 503 10235
rect 438 10090 503 10229
rect 778 10174 815 10253
rect 856 10240 966 10253
rect 930 10184 961 10185
rect 778 10154 787 10174
rect 807 10154 815 10174
rect 438 10072 461 10090
rect 479 10072 503 10090
rect 438 10055 503 10072
rect 658 10136 726 10149
rect 778 10144 815 10154
rect 874 10174 961 10184
rect 874 10154 883 10174
rect 903 10154 961 10174
rect 874 10145 961 10154
rect 874 10144 911 10145
rect 658 10094 665 10136
rect 714 10094 726 10136
rect 658 10091 726 10094
rect 930 10092 961 10145
rect 991 10174 1028 10253
rect 1143 10184 1174 10185
rect 991 10154 1000 10174
rect 1020 10154 1028 10174
rect 991 10144 1028 10154
rect 1087 10177 1174 10184
rect 1087 10174 1148 10177
rect 1087 10154 1096 10174
rect 1116 10157 1148 10174
rect 1169 10157 1174 10177
rect 1116 10154 1174 10157
rect 1087 10147 1174 10154
rect 1199 10174 1236 10316
rect 1502 10315 1539 10316
rect 2247 10313 2663 10318
rect 2247 10312 2588 10313
rect 1904 10281 2014 10295
rect 1904 10278 1947 10281
rect 1904 10273 1908 10278
rect 1826 10251 1908 10273
rect 1937 10251 1947 10278
rect 1975 10254 1982 10281
rect 2011 10273 2014 10281
rect 2011 10254 2076 10273
rect 1975 10251 2076 10254
rect 1826 10249 2076 10251
rect 1351 10184 1387 10185
rect 1199 10154 1208 10174
rect 1228 10154 1236 10174
rect 1087 10145 1143 10147
rect 1087 10144 1124 10145
rect 1199 10144 1236 10154
rect 1295 10174 1443 10184
rect 1543 10181 1639 10183
rect 1295 10154 1304 10174
rect 1324 10154 1414 10174
rect 1434 10154 1443 10174
rect 1295 10148 1443 10154
rect 1295 10145 1359 10148
rect 1295 10144 1332 10145
rect 1351 10118 1359 10145
rect 1380 10145 1443 10148
rect 1501 10174 1639 10181
rect 1501 10154 1510 10174
rect 1530 10154 1639 10174
rect 1501 10145 1639 10154
rect 1826 10170 1863 10249
rect 1904 10236 2014 10249
rect 1978 10180 2009 10181
rect 1826 10150 1835 10170
rect 1855 10150 1863 10170
rect 1380 10118 1387 10145
rect 1406 10144 1443 10145
rect 1502 10144 1539 10145
rect 1351 10093 1387 10118
rect 822 10091 863 10092
rect 658 10084 863 10091
rect 658 10073 832 10084
rect 658 10040 666 10073
rect 659 10031 666 10040
rect 715 10064 832 10073
rect 852 10064 863 10084
rect 715 10056 863 10064
rect 930 10088 1289 10092
rect 930 10083 1252 10088
rect 930 10059 1043 10083
rect 1067 10064 1252 10083
rect 1276 10064 1289 10088
rect 1067 10059 1289 10064
rect 930 10056 1289 10059
rect 1351 10056 1386 10093
rect 1454 10090 1554 10093
rect 1454 10086 1521 10090
rect 1454 10060 1466 10086
rect 1492 10064 1521 10086
rect 1547 10064 1554 10090
rect 1492 10060 1554 10064
rect 1454 10056 1554 10060
rect 715 10040 726 10056
rect 715 10031 723 10040
rect 930 10035 961 10056
rect 1351 10035 1387 10056
rect 773 10034 810 10035
rect 438 9991 503 10010
rect 438 9973 463 9991
rect 481 9973 503 9991
rect 438 9772 503 9973
rect 659 9847 723 10031
rect 772 10025 810 10034
rect 772 10005 781 10025
rect 801 10005 810 10025
rect 772 9997 810 10005
rect 876 10029 961 10035
rect 986 10034 1023 10035
rect 876 10009 884 10029
rect 904 10009 961 10029
rect 876 10001 961 10009
rect 985 10025 1023 10034
rect 985 10005 994 10025
rect 1014 10005 1023 10025
rect 876 10000 912 10001
rect 985 9997 1023 10005
rect 1089 10029 1174 10035
rect 1194 10034 1231 10035
rect 1089 10009 1097 10029
rect 1117 10028 1174 10029
rect 1117 10009 1146 10028
rect 1089 10008 1146 10009
rect 1167 10008 1174 10028
rect 1089 10001 1174 10008
rect 1193 10025 1231 10034
rect 1193 10005 1202 10025
rect 1222 10005 1231 10025
rect 1089 10000 1125 10001
rect 1193 9997 1231 10005
rect 1297 10029 1441 10035
rect 1297 10009 1305 10029
rect 1325 10009 1413 10029
rect 1433 10009 1441 10029
rect 1297 10001 1441 10009
rect 1297 10000 1333 10001
rect 1405 10000 1441 10001
rect 1507 10034 1544 10035
rect 1507 10033 1545 10034
rect 1507 10025 1571 10033
rect 1507 10005 1516 10025
rect 1536 10011 1571 10025
rect 1591 10011 1594 10031
rect 1536 10006 1594 10011
rect 1536 10005 1571 10006
rect 773 9968 810 9997
rect 774 9966 810 9968
rect 986 9966 1023 9997
rect 774 9944 1023 9966
rect 855 9938 966 9944
rect 855 9930 896 9938
rect 855 9910 863 9930
rect 882 9910 896 9930
rect 855 9908 896 9910
rect 924 9930 966 9938
rect 924 9910 940 9930
rect 959 9910 966 9930
rect 924 9908 966 9910
rect 855 9893 966 9908
rect 659 9837 727 9847
rect 659 9804 676 9837
rect 716 9804 727 9837
rect 659 9792 727 9804
rect 659 9790 723 9792
rect 1194 9773 1231 9997
rect 1507 9993 1571 10005
rect 1611 9775 1638 10145
rect 1826 10140 1863 10150
rect 1922 10170 2009 10180
rect 1922 10150 1931 10170
rect 1951 10150 2009 10170
rect 1922 10141 2009 10150
rect 1922 10140 1959 10141
rect 1702 10127 1772 10132
rect 1697 10121 1772 10127
rect 1697 10088 1705 10121
rect 1758 10088 1772 10121
rect 1978 10088 2009 10141
rect 2039 10170 2076 10249
rect 2191 10180 2222 10181
rect 2039 10150 2048 10170
rect 2068 10150 2076 10170
rect 2039 10140 2076 10150
rect 2135 10173 2222 10180
rect 2135 10170 2196 10173
rect 2135 10150 2144 10170
rect 2164 10153 2196 10170
rect 2217 10153 2222 10173
rect 2164 10150 2222 10153
rect 2135 10143 2222 10150
rect 2247 10170 2284 10312
rect 2550 10311 2587 10312
rect 2399 10180 2435 10181
rect 2247 10150 2256 10170
rect 2276 10150 2284 10170
rect 2135 10141 2191 10143
rect 2135 10140 2172 10141
rect 2247 10140 2284 10150
rect 2343 10170 2491 10180
rect 2591 10177 2687 10179
rect 2343 10150 2352 10170
rect 2372 10150 2462 10170
rect 2482 10150 2491 10170
rect 2343 10144 2491 10150
rect 2343 10141 2407 10144
rect 2343 10140 2380 10141
rect 2399 10114 2407 10141
rect 2428 10141 2491 10144
rect 2549 10170 2687 10177
rect 2549 10150 2558 10170
rect 2578 10150 2687 10170
rect 2549 10141 2687 10150
rect 2428 10114 2435 10141
rect 2454 10140 2491 10141
rect 2550 10140 2587 10141
rect 2399 10089 2435 10114
rect 1697 10087 1780 10088
rect 1870 10087 1911 10088
rect 1697 10080 1911 10087
rect 1697 10063 1880 10080
rect 1697 10030 1710 10063
rect 1763 10060 1880 10063
rect 1900 10060 1911 10080
rect 1763 10052 1911 10060
rect 1978 10084 2337 10088
rect 1978 10079 2300 10084
rect 1978 10055 2091 10079
rect 2115 10060 2300 10079
rect 2324 10060 2337 10084
rect 2115 10055 2337 10060
rect 1978 10052 2337 10055
rect 2399 10052 2434 10089
rect 2502 10086 2602 10089
rect 2502 10082 2569 10086
rect 2502 10056 2514 10082
rect 2540 10060 2569 10082
rect 2595 10060 2602 10086
rect 2540 10056 2602 10060
rect 2502 10052 2602 10056
rect 1763 10030 1780 10052
rect 1978 10031 2009 10052
rect 2399 10031 2435 10052
rect 1821 10030 1858 10031
rect 1697 10016 1780 10030
rect 1470 9773 1638 9775
rect 1194 9772 1638 9773
rect 438 9742 1638 9772
rect 1708 9806 1780 10016
rect 1820 10021 1858 10030
rect 1820 10001 1829 10021
rect 1849 10001 1858 10021
rect 1820 9993 1858 10001
rect 1924 10025 2009 10031
rect 2034 10030 2071 10031
rect 1924 10005 1932 10025
rect 1952 10005 2009 10025
rect 1924 9997 2009 10005
rect 2033 10021 2071 10030
rect 2033 10001 2042 10021
rect 2062 10001 2071 10021
rect 1924 9996 1960 9997
rect 2033 9993 2071 10001
rect 2137 10025 2222 10031
rect 2242 10030 2279 10031
rect 2137 10005 2145 10025
rect 2165 10024 2222 10025
rect 2165 10005 2194 10024
rect 2137 10004 2194 10005
rect 2215 10004 2222 10024
rect 2137 9997 2222 10004
rect 2241 10021 2279 10030
rect 2241 10001 2250 10021
rect 2270 10001 2279 10021
rect 2137 9996 2173 9997
rect 2241 9993 2279 10001
rect 2345 10025 2489 10031
rect 2345 10005 2353 10025
rect 2373 10005 2461 10025
rect 2481 10005 2489 10025
rect 2345 9997 2489 10005
rect 2345 9996 2381 9997
rect 2453 9996 2489 9997
rect 2555 10030 2592 10031
rect 2555 10029 2593 10030
rect 2555 10021 2619 10029
rect 2555 10001 2564 10021
rect 2584 10007 2619 10021
rect 2639 10007 2642 10027
rect 2584 10002 2642 10007
rect 2584 10001 2619 10002
rect 1821 9964 1858 9993
rect 1822 9962 1858 9964
rect 2034 9962 2071 9993
rect 1822 9940 2071 9962
rect 1903 9934 2014 9940
rect 1903 9926 1944 9934
rect 1903 9906 1911 9926
rect 1930 9906 1944 9926
rect 1903 9904 1944 9906
rect 1972 9926 2014 9934
rect 1972 9906 1988 9926
rect 2007 9906 2014 9926
rect 1972 9904 2014 9906
rect 1903 9889 2014 9904
rect 1708 9767 1727 9806
rect 1772 9767 1780 9806
rect 1708 9750 1780 9767
rect 2242 9794 2279 9993
rect 2555 9989 2619 10001
rect 2242 9788 2283 9794
rect 2659 9790 2686 10141
rect 2809 10011 2888 10611
rect 2985 10159 3064 10744
rect 3268 10731 3305 10760
rect 3269 10729 3305 10731
rect 3481 10729 3518 10760
rect 3269 10707 3518 10729
rect 3350 10701 3461 10707
rect 3350 10693 3391 10701
rect 3350 10673 3358 10693
rect 3377 10673 3391 10693
rect 3350 10671 3391 10673
rect 3419 10693 3461 10701
rect 3419 10673 3435 10693
rect 3454 10673 3461 10693
rect 3419 10671 3461 10673
rect 3350 10656 3461 10671
rect 3689 10645 3726 10760
rect 3682 10533 3729 10645
rect 3850 10605 3880 10764
rect 3900 10763 3936 10764
rect 4002 10797 4039 10798
rect 4002 10796 4040 10797
rect 4002 10788 4066 10796
rect 4002 10768 4011 10788
rect 4031 10774 4066 10788
rect 4086 10774 4089 10794
rect 4031 10769 4089 10774
rect 4031 10768 4066 10769
rect 4002 10756 4066 10768
rect 3850 10601 3936 10605
rect 3850 10583 3865 10601
rect 3917 10583 3936 10601
rect 3850 10574 3936 10583
rect 4106 10535 4133 10908
rect 3965 10533 4133 10535
rect 3682 10507 4133 10533
rect 3682 10429 3729 10507
rect 3965 10506 4133 10507
rect 3627 10428 3729 10429
rect 3626 10420 3729 10428
rect 3626 10417 3678 10420
rect 3626 10382 3634 10417
rect 3659 10382 3678 10417
rect 3703 10382 3729 10420
rect 3626 10376 3729 10382
rect 3889 10421 3925 10425
rect 3889 10398 3897 10421
rect 3921 10398 3925 10421
rect 3889 10377 3925 10398
rect 3626 10372 3725 10376
rect 3889 10354 3897 10377
rect 3921 10354 3925 10377
rect 2518 9788 2686 9790
rect 2242 9762 2686 9788
rect 438 9695 503 9742
rect 438 9677 461 9695
rect 479 9677 503 9695
rect 1351 9722 1386 9724
rect 1351 9720 1455 9722
rect 2244 9720 2283 9762
rect 2518 9761 2686 9762
rect 1351 9713 2285 9720
rect 1351 9712 1402 9713
rect 1351 9692 1354 9712
rect 1379 9693 1402 9712
rect 1434 9693 2285 9713
rect 1379 9692 2285 9693
rect 1351 9685 2285 9692
rect 1624 9684 2285 9685
rect 438 9656 503 9677
rect 715 9667 755 9670
rect 715 9663 1618 9667
rect 715 9643 1592 9663
rect 1612 9643 1618 9663
rect 715 9640 1618 9643
rect 439 9596 504 9616
rect 439 9578 463 9596
rect 481 9578 504 9596
rect 439 9551 504 9578
rect 715 9551 755 9640
rect 1199 9638 1615 9640
rect 1199 9637 1540 9638
rect 856 9606 966 9620
rect 856 9603 899 9606
rect 856 9598 860 9603
rect 438 9516 755 9551
rect 778 9576 860 9598
rect 889 9576 899 9603
rect 927 9579 934 9606
rect 963 9598 966 9606
rect 963 9579 1028 9598
rect 927 9576 1028 9579
rect 778 9574 1028 9576
rect 439 9440 504 9516
rect 778 9495 815 9574
rect 856 9561 966 9574
rect 930 9505 961 9506
rect 778 9475 787 9495
rect 807 9475 815 9495
rect 778 9465 815 9475
rect 874 9495 961 9505
rect 874 9475 883 9495
rect 903 9475 961 9495
rect 874 9466 961 9475
rect 874 9465 911 9466
rect 439 9422 461 9440
rect 479 9422 504 9440
rect 439 9401 504 9422
rect 652 9420 717 9429
rect 652 9383 662 9420
rect 702 9412 717 9420
rect 930 9413 961 9466
rect 991 9495 1028 9574
rect 1143 9505 1174 9506
rect 991 9475 1000 9495
rect 1020 9475 1028 9495
rect 991 9465 1028 9475
rect 1087 9498 1174 9505
rect 1087 9495 1148 9498
rect 1087 9475 1096 9495
rect 1116 9478 1148 9495
rect 1169 9478 1174 9498
rect 1116 9475 1174 9478
rect 1087 9468 1174 9475
rect 1199 9495 1236 9637
rect 1502 9636 1539 9637
rect 1351 9505 1387 9506
rect 1199 9475 1208 9495
rect 1228 9475 1236 9495
rect 1087 9466 1143 9468
rect 1087 9465 1124 9466
rect 1199 9465 1236 9475
rect 1295 9495 1443 9505
rect 1543 9502 1639 9504
rect 1295 9475 1304 9495
rect 1324 9475 1414 9495
rect 1434 9475 1443 9495
rect 1295 9469 1443 9475
rect 1295 9466 1359 9469
rect 1295 9465 1332 9466
rect 1351 9439 1359 9466
rect 1380 9466 1443 9469
rect 1501 9495 1639 9502
rect 1501 9475 1510 9495
rect 1530 9475 1639 9495
rect 1501 9466 1639 9475
rect 1380 9439 1387 9466
rect 1406 9465 1443 9466
rect 1502 9465 1539 9466
rect 1351 9414 1387 9439
rect 822 9412 863 9413
rect 702 9405 863 9412
rect 702 9385 832 9405
rect 852 9385 863 9405
rect 702 9383 863 9385
rect 652 9377 863 9383
rect 930 9409 1289 9413
rect 930 9404 1252 9409
rect 930 9380 1043 9404
rect 1067 9385 1252 9404
rect 1276 9385 1289 9409
rect 1067 9380 1289 9385
rect 930 9377 1289 9380
rect 1351 9377 1386 9414
rect 1454 9411 1554 9414
rect 1454 9407 1521 9411
rect 1454 9381 1466 9407
rect 1492 9385 1521 9407
rect 1547 9385 1554 9411
rect 1492 9381 1554 9385
rect 1454 9377 1554 9381
rect 652 9364 719 9377
rect 444 9341 500 9361
rect 444 9323 463 9341
rect 481 9323 500 9341
rect 444 9210 500 9323
rect 652 9343 666 9364
rect 702 9343 719 9364
rect 930 9356 961 9377
rect 1351 9356 1387 9377
rect 773 9355 810 9356
rect 652 9336 719 9343
rect 772 9346 810 9355
rect 444 9081 499 9210
rect 652 9184 717 9336
rect 772 9326 781 9346
rect 801 9326 810 9346
rect 772 9318 810 9326
rect 876 9350 961 9356
rect 986 9355 1023 9356
rect 876 9330 884 9350
rect 904 9330 961 9350
rect 876 9322 961 9330
rect 985 9346 1023 9355
rect 985 9326 994 9346
rect 1014 9326 1023 9346
rect 876 9321 912 9322
rect 985 9318 1023 9326
rect 1089 9350 1174 9356
rect 1194 9355 1231 9356
rect 1089 9330 1097 9350
rect 1117 9349 1174 9350
rect 1117 9330 1146 9349
rect 1089 9329 1146 9330
rect 1167 9329 1174 9349
rect 1089 9322 1174 9329
rect 1193 9346 1231 9355
rect 1193 9326 1202 9346
rect 1222 9326 1231 9346
rect 1089 9321 1125 9322
rect 1193 9318 1231 9326
rect 1297 9350 1441 9356
rect 1297 9330 1305 9350
rect 1325 9330 1413 9350
rect 1433 9330 1441 9350
rect 1297 9322 1441 9330
rect 1297 9321 1333 9322
rect 1405 9321 1441 9322
rect 1507 9355 1544 9356
rect 1507 9354 1545 9355
rect 1507 9346 1571 9354
rect 1507 9326 1516 9346
rect 1536 9332 1571 9346
rect 1591 9332 1594 9352
rect 1536 9327 1594 9332
rect 1536 9326 1571 9327
rect 773 9289 810 9318
rect 774 9287 810 9289
rect 986 9287 1023 9318
rect 774 9265 1023 9287
rect 855 9259 966 9265
rect 855 9251 896 9259
rect 855 9231 863 9251
rect 882 9231 896 9251
rect 855 9229 896 9231
rect 924 9251 966 9259
rect 924 9231 940 9251
rect 959 9231 966 9251
rect 924 9229 966 9231
rect 855 9214 966 9229
rect 1194 9219 1231 9318
rect 1507 9314 1571 9326
rect 857 9205 961 9214
rect 645 9174 766 9184
rect 645 9172 714 9174
rect 645 9131 658 9172
rect 695 9133 714 9172
rect 751 9133 766 9174
rect 695 9131 766 9133
rect 645 9113 766 9131
rect 438 9069 499 9081
rect 1192 9069 1233 9219
rect 1611 9211 1638 9466
rect 1700 9456 1780 9467
rect 1700 9430 1717 9456
rect 1757 9430 1780 9456
rect 1700 9403 1780 9430
rect 1700 9377 1721 9403
rect 1761 9377 1780 9403
rect 1700 9358 1780 9377
rect 1700 9332 1724 9358
rect 1764 9332 1780 9358
rect 1700 9281 1780 9332
rect 438 9066 1233 9069
rect 1612 9080 1638 9211
rect 1702 9125 1772 9281
rect 1701 9109 1777 9125
rect 1612 9066 1640 9080
rect 438 9031 1640 9066
rect 1701 9072 1716 9109
rect 1760 9072 1777 9109
rect 1701 9052 1777 9072
rect 2815 9102 2885 10011
rect 2984 9446 3065 10159
rect 3889 10045 3925 10354
rect 3813 10016 3926 10045
rect 3813 9660 3844 10016
rect 3883 9761 4874 9786
rect 3883 9756 3943 9761
rect 3883 9735 3902 9756
rect 3922 9740 3943 9756
rect 3963 9740 4874 9761
rect 3922 9735 4874 9740
rect 3883 9727 4874 9735
rect 3888 9704 3994 9727
rect 3888 9701 3993 9704
rect 3737 9640 4130 9660
rect 4150 9640 4153 9660
rect 3737 9635 4153 9640
rect 3737 9634 4078 9635
rect 3394 9603 3504 9617
rect 3394 9600 3437 9603
rect 3394 9595 3398 9600
rect 3316 9573 3398 9595
rect 3427 9573 3437 9600
rect 3465 9576 3472 9603
rect 3501 9595 3504 9603
rect 3501 9576 3566 9595
rect 3465 9573 3566 9576
rect 3316 9571 3566 9573
rect 3316 9492 3353 9571
rect 3394 9558 3504 9571
rect 3468 9502 3499 9503
rect 3316 9472 3325 9492
rect 3345 9472 3353 9492
rect 3316 9462 3353 9472
rect 3412 9492 3499 9502
rect 3412 9472 3421 9492
rect 3441 9472 3499 9492
rect 3412 9463 3499 9472
rect 3412 9462 3449 9463
rect 2982 9410 3074 9446
rect 3468 9410 3499 9463
rect 3529 9492 3566 9571
rect 3681 9502 3712 9503
rect 3529 9472 3538 9492
rect 3558 9472 3566 9492
rect 3529 9462 3566 9472
rect 3625 9495 3712 9502
rect 3625 9492 3686 9495
rect 3625 9472 3634 9492
rect 3654 9475 3686 9492
rect 3707 9475 3712 9495
rect 3654 9472 3712 9475
rect 3625 9465 3712 9472
rect 3737 9492 3774 9634
rect 4040 9633 4077 9634
rect 3889 9502 3925 9503
rect 3737 9472 3746 9492
rect 3766 9472 3774 9492
rect 3625 9463 3681 9465
rect 3625 9462 3662 9463
rect 3737 9462 3774 9472
rect 3833 9492 3981 9502
rect 4081 9499 4177 9501
rect 3833 9472 3842 9492
rect 3862 9472 3952 9492
rect 3972 9472 3981 9492
rect 3833 9466 3981 9472
rect 3833 9463 3897 9466
rect 3833 9462 3870 9463
rect 3889 9436 3897 9463
rect 3918 9463 3981 9466
rect 4039 9492 4177 9499
rect 4039 9472 4048 9492
rect 4068 9472 4177 9492
rect 4039 9463 4177 9472
rect 3918 9436 3925 9463
rect 3944 9462 3981 9463
rect 4040 9462 4077 9463
rect 3889 9411 3925 9436
rect 2982 9409 3318 9410
rect 3360 9409 3401 9410
rect 2982 9402 3401 9409
rect 2982 9382 3370 9402
rect 3390 9382 3401 9402
rect 2982 9374 3401 9382
rect 3468 9406 3827 9410
rect 3468 9401 3790 9406
rect 3468 9377 3581 9401
rect 3605 9382 3790 9401
rect 3814 9382 3827 9406
rect 3605 9377 3827 9382
rect 3468 9374 3827 9377
rect 3889 9374 3924 9411
rect 3992 9408 4092 9411
rect 3992 9404 4059 9408
rect 3992 9378 4004 9404
rect 4030 9382 4059 9404
rect 4085 9382 4092 9408
rect 4030 9378 4092 9382
rect 3992 9374 4092 9378
rect 2982 9370 3318 9374
rect 2815 9052 2887 9102
rect 438 8956 499 9031
rect 857 9029 961 9031
rect 1192 9029 1233 9031
rect 1701 8986 1711 9052
rect 1765 8986 1777 9052
rect 1701 8962 1777 8986
rect 440 8826 499 8956
rect 1353 8907 1425 8908
rect 1352 8899 1451 8907
rect 1352 8896 1404 8899
rect 1352 8861 1360 8896
rect 1385 8861 1404 8896
rect 1429 8888 1451 8899
rect 1429 8887 2296 8888
rect 1429 8861 2297 8887
rect 1352 8851 2297 8861
rect 1352 8849 1451 8851
rect 440 8808 462 8826
rect 480 8808 499 8826
rect 440 8786 499 8808
rect 707 8822 1239 8827
rect 707 8802 1593 8822
rect 1613 8802 1616 8822
rect 2252 8818 2297 8851
rect 707 8798 1616 8802
rect 707 8751 750 8798
rect 1200 8797 1616 8798
rect 2248 8798 2641 8818
rect 2661 8798 2664 8818
rect 1200 8796 1541 8797
rect 857 8765 967 8779
rect 857 8762 900 8765
rect 857 8757 861 8762
rect 695 8750 750 8751
rect 439 8727 750 8750
rect 439 8709 464 8727
rect 482 8715 750 8727
rect 779 8735 861 8757
rect 890 8735 900 8762
rect 928 8738 935 8765
rect 964 8757 967 8765
rect 964 8738 1029 8757
rect 928 8735 1029 8738
rect 779 8733 1029 8735
rect 482 8709 504 8715
rect 439 8570 504 8709
rect 779 8654 816 8733
rect 857 8720 967 8733
rect 931 8664 962 8665
rect 779 8634 788 8654
rect 808 8634 816 8654
rect 439 8552 462 8570
rect 480 8552 504 8570
rect 439 8535 504 8552
rect 659 8616 727 8629
rect 779 8624 816 8634
rect 875 8654 962 8664
rect 875 8634 884 8654
rect 904 8634 962 8654
rect 875 8625 962 8634
rect 875 8624 912 8625
rect 659 8574 666 8616
rect 715 8574 727 8616
rect 659 8571 727 8574
rect 931 8572 962 8625
rect 992 8654 1029 8733
rect 1144 8664 1175 8665
rect 992 8634 1001 8654
rect 1021 8634 1029 8654
rect 992 8624 1029 8634
rect 1088 8657 1175 8664
rect 1088 8654 1149 8657
rect 1088 8634 1097 8654
rect 1117 8637 1149 8654
rect 1170 8637 1175 8657
rect 1117 8634 1175 8637
rect 1088 8627 1175 8634
rect 1200 8654 1237 8796
rect 1503 8795 1540 8796
rect 2248 8793 2664 8798
rect 2248 8792 2589 8793
rect 1905 8761 2015 8775
rect 1905 8758 1948 8761
rect 1905 8753 1909 8758
rect 1827 8731 1909 8753
rect 1938 8731 1948 8758
rect 1976 8734 1983 8761
rect 2012 8753 2015 8761
rect 2012 8734 2077 8753
rect 1976 8731 2077 8734
rect 1827 8729 2077 8731
rect 1352 8664 1388 8665
rect 1200 8634 1209 8654
rect 1229 8634 1237 8654
rect 1088 8625 1144 8627
rect 1088 8624 1125 8625
rect 1200 8624 1237 8634
rect 1296 8654 1444 8664
rect 1544 8661 1640 8663
rect 1296 8634 1305 8654
rect 1325 8634 1415 8654
rect 1435 8634 1444 8654
rect 1296 8628 1444 8634
rect 1296 8625 1360 8628
rect 1296 8624 1333 8625
rect 1352 8598 1360 8625
rect 1381 8625 1444 8628
rect 1502 8654 1640 8661
rect 1502 8634 1511 8654
rect 1531 8634 1640 8654
rect 1502 8625 1640 8634
rect 1827 8650 1864 8729
rect 1905 8716 2015 8729
rect 1979 8660 2010 8661
rect 1827 8630 1836 8650
rect 1856 8630 1864 8650
rect 1381 8598 1388 8625
rect 1407 8624 1444 8625
rect 1503 8624 1540 8625
rect 1352 8573 1388 8598
rect 823 8571 864 8572
rect 659 8564 864 8571
rect 659 8553 833 8564
rect 659 8520 667 8553
rect 660 8511 667 8520
rect 716 8544 833 8553
rect 853 8544 864 8564
rect 716 8536 864 8544
rect 931 8568 1290 8572
rect 931 8563 1253 8568
rect 931 8539 1044 8563
rect 1068 8544 1253 8563
rect 1277 8544 1290 8568
rect 1068 8539 1290 8544
rect 931 8536 1290 8539
rect 1352 8536 1387 8573
rect 1455 8570 1555 8573
rect 1455 8566 1522 8570
rect 1455 8540 1467 8566
rect 1493 8544 1522 8566
rect 1548 8544 1555 8570
rect 1493 8540 1555 8544
rect 1455 8536 1555 8540
rect 716 8520 727 8536
rect 716 8511 724 8520
rect 931 8515 962 8536
rect 1352 8515 1388 8536
rect 774 8514 811 8515
rect 439 8471 504 8490
rect 439 8453 464 8471
rect 482 8453 504 8471
rect 439 8252 504 8453
rect 660 8327 724 8511
rect 773 8505 811 8514
rect 773 8485 782 8505
rect 802 8485 811 8505
rect 773 8477 811 8485
rect 877 8509 962 8515
rect 987 8514 1024 8515
rect 877 8489 885 8509
rect 905 8489 962 8509
rect 877 8481 962 8489
rect 986 8505 1024 8514
rect 986 8485 995 8505
rect 1015 8485 1024 8505
rect 877 8480 913 8481
rect 986 8477 1024 8485
rect 1090 8509 1175 8515
rect 1195 8514 1232 8515
rect 1090 8489 1098 8509
rect 1118 8508 1175 8509
rect 1118 8489 1147 8508
rect 1090 8488 1147 8489
rect 1168 8488 1175 8508
rect 1090 8481 1175 8488
rect 1194 8505 1232 8514
rect 1194 8485 1203 8505
rect 1223 8485 1232 8505
rect 1090 8480 1126 8481
rect 1194 8477 1232 8485
rect 1298 8509 1442 8515
rect 1298 8489 1306 8509
rect 1326 8489 1414 8509
rect 1434 8489 1442 8509
rect 1298 8481 1442 8489
rect 1298 8480 1334 8481
rect 1406 8480 1442 8481
rect 1508 8514 1545 8515
rect 1508 8513 1546 8514
rect 1508 8505 1572 8513
rect 1508 8485 1517 8505
rect 1537 8491 1572 8505
rect 1592 8491 1595 8511
rect 1537 8486 1595 8491
rect 1537 8485 1572 8486
rect 774 8448 811 8477
rect 775 8446 811 8448
rect 987 8446 1024 8477
rect 775 8424 1024 8446
rect 856 8418 967 8424
rect 856 8410 897 8418
rect 856 8390 864 8410
rect 883 8390 897 8410
rect 856 8388 897 8390
rect 925 8410 967 8418
rect 925 8390 941 8410
rect 960 8390 967 8410
rect 925 8388 967 8390
rect 856 8373 967 8388
rect 660 8317 728 8327
rect 660 8284 677 8317
rect 717 8284 728 8317
rect 660 8272 728 8284
rect 660 8270 724 8272
rect 1195 8253 1232 8477
rect 1508 8473 1572 8485
rect 1612 8255 1639 8625
rect 1827 8620 1864 8630
rect 1923 8650 2010 8660
rect 1923 8630 1932 8650
rect 1952 8630 2010 8650
rect 1923 8621 2010 8630
rect 1923 8620 1960 8621
rect 1703 8607 1773 8612
rect 1698 8601 1773 8607
rect 1698 8568 1706 8601
rect 1759 8568 1773 8601
rect 1979 8568 2010 8621
rect 2040 8650 2077 8729
rect 2192 8660 2223 8661
rect 2040 8630 2049 8650
rect 2069 8630 2077 8650
rect 2040 8620 2077 8630
rect 2136 8653 2223 8660
rect 2136 8650 2197 8653
rect 2136 8630 2145 8650
rect 2165 8633 2197 8650
rect 2218 8633 2223 8653
rect 2165 8630 2223 8633
rect 2136 8623 2223 8630
rect 2248 8650 2285 8792
rect 2551 8791 2588 8792
rect 2400 8660 2436 8661
rect 2248 8630 2257 8650
rect 2277 8630 2285 8650
rect 2136 8621 2192 8623
rect 2136 8620 2173 8621
rect 2248 8620 2285 8630
rect 2344 8650 2492 8660
rect 2592 8657 2688 8659
rect 2344 8630 2353 8650
rect 2373 8630 2463 8650
rect 2483 8630 2492 8650
rect 2344 8624 2492 8630
rect 2344 8621 2408 8624
rect 2344 8620 2381 8621
rect 2400 8594 2408 8621
rect 2429 8621 2492 8624
rect 2550 8650 2688 8657
rect 2550 8630 2559 8650
rect 2579 8630 2688 8650
rect 2550 8621 2688 8630
rect 2429 8594 2436 8621
rect 2455 8620 2492 8621
rect 2551 8620 2588 8621
rect 2400 8569 2436 8594
rect 1698 8567 1781 8568
rect 1871 8567 1912 8568
rect 1698 8560 1912 8567
rect 1698 8543 1881 8560
rect 1698 8510 1711 8543
rect 1764 8540 1881 8543
rect 1901 8540 1912 8560
rect 1764 8532 1912 8540
rect 1979 8564 2338 8568
rect 1979 8559 2301 8564
rect 1979 8535 2092 8559
rect 2116 8540 2301 8559
rect 2325 8540 2338 8564
rect 2116 8535 2338 8540
rect 1979 8532 2338 8535
rect 2400 8532 2435 8569
rect 2503 8566 2603 8569
rect 2503 8562 2570 8566
rect 2503 8536 2515 8562
rect 2541 8540 2570 8562
rect 2596 8540 2603 8566
rect 2541 8536 2603 8540
rect 2503 8532 2603 8536
rect 1764 8510 1781 8532
rect 1979 8511 2010 8532
rect 2400 8511 2436 8532
rect 1822 8510 1859 8511
rect 1698 8496 1781 8510
rect 1471 8253 1639 8255
rect 1195 8252 1639 8253
rect 439 8222 1639 8252
rect 1709 8286 1781 8496
rect 1821 8501 1859 8510
rect 1821 8481 1830 8501
rect 1850 8481 1859 8501
rect 1821 8473 1859 8481
rect 1925 8505 2010 8511
rect 2035 8510 2072 8511
rect 1925 8485 1933 8505
rect 1953 8485 2010 8505
rect 1925 8477 2010 8485
rect 2034 8501 2072 8510
rect 2034 8481 2043 8501
rect 2063 8481 2072 8501
rect 1925 8476 1961 8477
rect 2034 8473 2072 8481
rect 2138 8505 2223 8511
rect 2243 8510 2280 8511
rect 2138 8485 2146 8505
rect 2166 8504 2223 8505
rect 2166 8485 2195 8504
rect 2138 8484 2195 8485
rect 2216 8484 2223 8504
rect 2138 8477 2223 8484
rect 2242 8501 2280 8510
rect 2242 8481 2251 8501
rect 2271 8481 2280 8501
rect 2138 8476 2174 8477
rect 2242 8473 2280 8481
rect 2346 8505 2490 8511
rect 2346 8485 2354 8505
rect 2374 8485 2462 8505
rect 2482 8485 2490 8505
rect 2346 8477 2490 8485
rect 2346 8476 2382 8477
rect 2454 8476 2490 8477
rect 2556 8510 2593 8511
rect 2556 8509 2594 8510
rect 2556 8501 2620 8509
rect 2556 8481 2565 8501
rect 2585 8487 2620 8501
rect 2640 8487 2643 8507
rect 2585 8482 2643 8487
rect 2585 8481 2620 8482
rect 1822 8444 1859 8473
rect 1823 8442 1859 8444
rect 2035 8442 2072 8473
rect 1823 8420 2072 8442
rect 1904 8414 2015 8420
rect 1904 8406 1945 8414
rect 1904 8386 1912 8406
rect 1931 8386 1945 8406
rect 1904 8384 1945 8386
rect 1973 8406 2015 8414
rect 1973 8386 1989 8406
rect 2008 8386 2015 8406
rect 1973 8384 2015 8386
rect 1904 8369 2015 8384
rect 1709 8247 1728 8286
rect 1773 8247 1781 8286
rect 1709 8230 1781 8247
rect 2243 8274 2280 8473
rect 2556 8469 2620 8481
rect 2243 8268 2284 8274
rect 2660 8270 2687 8621
rect 2816 8573 2887 9052
rect 2816 8489 2885 8573
rect 2519 8268 2687 8270
rect 2243 8242 2687 8268
rect 439 8175 504 8222
rect 439 8157 462 8175
rect 480 8157 504 8175
rect 1352 8202 1387 8204
rect 1352 8200 1456 8202
rect 2245 8200 2284 8242
rect 2519 8241 2687 8242
rect 1352 8193 2286 8200
rect 1352 8192 1403 8193
rect 1352 8172 1355 8192
rect 1380 8173 1403 8192
rect 1435 8173 2286 8193
rect 1380 8172 2286 8173
rect 1352 8165 2286 8172
rect 1625 8164 2286 8165
rect 439 8136 504 8157
rect 716 8147 756 8150
rect 716 8143 1619 8147
rect 716 8123 1593 8143
rect 1613 8123 1619 8143
rect 716 8120 1619 8123
rect 440 8076 505 8096
rect 440 8058 464 8076
rect 482 8058 505 8076
rect 440 8031 505 8058
rect 716 8031 756 8120
rect 1200 8118 1616 8120
rect 1200 8117 1541 8118
rect 857 8086 967 8100
rect 857 8083 900 8086
rect 857 8078 861 8083
rect 439 7996 756 8031
rect 779 8056 861 8078
rect 890 8056 900 8083
rect 928 8059 935 8086
rect 964 8078 967 8086
rect 964 8059 1029 8078
rect 928 8056 1029 8059
rect 779 8054 1029 8056
rect 440 7920 505 7996
rect 779 7975 816 8054
rect 857 8041 967 8054
rect 931 7985 962 7986
rect 779 7955 788 7975
rect 808 7955 816 7975
rect 779 7945 816 7955
rect 875 7975 962 7985
rect 875 7955 884 7975
rect 904 7955 962 7975
rect 875 7946 962 7955
rect 875 7945 912 7946
rect 440 7902 462 7920
rect 480 7902 505 7920
rect 440 7881 505 7902
rect 653 7900 718 7909
rect 653 7863 663 7900
rect 703 7892 718 7900
rect 931 7893 962 7946
rect 992 7975 1029 8054
rect 1144 7985 1175 7986
rect 992 7955 1001 7975
rect 1021 7955 1029 7975
rect 992 7945 1029 7955
rect 1088 7978 1175 7985
rect 1088 7975 1149 7978
rect 1088 7955 1097 7975
rect 1117 7958 1149 7975
rect 1170 7958 1175 7978
rect 1117 7955 1175 7958
rect 1088 7948 1175 7955
rect 1200 7975 1237 8117
rect 1503 8116 1540 8117
rect 1352 7985 1388 7986
rect 1200 7955 1209 7975
rect 1229 7955 1237 7975
rect 1088 7946 1144 7948
rect 1088 7945 1125 7946
rect 1200 7945 1237 7955
rect 1296 7975 1444 7985
rect 1544 7982 1640 7984
rect 1296 7955 1305 7975
rect 1325 7955 1415 7975
rect 1435 7955 1444 7975
rect 1296 7949 1444 7955
rect 1296 7946 1360 7949
rect 1296 7945 1333 7946
rect 1352 7919 1360 7946
rect 1381 7946 1444 7949
rect 1502 7975 1640 7982
rect 1502 7955 1511 7975
rect 1531 7955 1640 7975
rect 2820 7973 2882 8489
rect 1502 7946 1640 7955
rect 1381 7919 1388 7946
rect 1407 7945 1444 7946
rect 1503 7945 1540 7946
rect 1352 7894 1388 7919
rect 823 7892 864 7893
rect 703 7885 864 7892
rect 703 7865 833 7885
rect 853 7865 864 7885
rect 703 7863 864 7865
rect 653 7857 864 7863
rect 931 7889 1290 7893
rect 931 7884 1253 7889
rect 931 7860 1044 7884
rect 1068 7865 1253 7884
rect 1277 7865 1290 7889
rect 1068 7860 1290 7865
rect 931 7857 1290 7860
rect 1352 7857 1387 7894
rect 1455 7891 1555 7894
rect 1455 7887 1522 7891
rect 1455 7861 1467 7887
rect 1493 7865 1522 7887
rect 1548 7865 1555 7891
rect 1493 7861 1555 7865
rect 1455 7857 1555 7861
rect 653 7844 720 7857
rect 445 7821 501 7841
rect 445 7803 464 7821
rect 482 7803 501 7821
rect 445 7690 501 7803
rect 653 7823 667 7844
rect 703 7823 720 7844
rect 931 7836 962 7857
rect 1352 7836 1388 7857
rect 774 7835 811 7836
rect 653 7816 720 7823
rect 773 7826 811 7835
rect 445 7552 500 7690
rect 653 7664 718 7816
rect 773 7806 782 7826
rect 802 7806 811 7826
rect 773 7798 811 7806
rect 877 7830 962 7836
rect 987 7835 1024 7836
rect 877 7810 885 7830
rect 905 7810 962 7830
rect 877 7802 962 7810
rect 986 7826 1024 7835
rect 986 7806 995 7826
rect 1015 7806 1024 7826
rect 877 7801 913 7802
rect 986 7798 1024 7806
rect 1090 7830 1175 7836
rect 1195 7835 1232 7836
rect 1090 7810 1098 7830
rect 1118 7829 1175 7830
rect 1118 7810 1147 7829
rect 1090 7809 1147 7810
rect 1168 7809 1175 7829
rect 1090 7802 1175 7809
rect 1194 7826 1232 7835
rect 1194 7806 1203 7826
rect 1223 7806 1232 7826
rect 1090 7801 1126 7802
rect 1194 7798 1232 7806
rect 1298 7830 1442 7836
rect 1298 7810 1306 7830
rect 1326 7810 1414 7830
rect 1434 7810 1442 7830
rect 1298 7802 1442 7810
rect 1298 7801 1334 7802
rect 1406 7801 1442 7802
rect 1508 7835 1545 7836
rect 1508 7834 1546 7835
rect 1508 7826 1572 7834
rect 1508 7806 1517 7826
rect 1537 7812 1572 7826
rect 1592 7812 1595 7832
rect 1537 7807 1595 7812
rect 1537 7806 1572 7807
rect 774 7769 811 7798
rect 775 7767 811 7769
rect 987 7767 1024 7798
rect 775 7745 1024 7767
rect 856 7739 967 7745
rect 856 7731 897 7739
rect 856 7711 864 7731
rect 883 7711 897 7731
rect 856 7709 897 7711
rect 925 7731 967 7739
rect 925 7711 941 7731
rect 960 7711 967 7731
rect 925 7709 967 7711
rect 856 7696 967 7709
rect 1195 7699 1232 7798
rect 1508 7794 1572 7806
rect 646 7654 767 7664
rect 646 7652 715 7654
rect 646 7611 659 7652
rect 696 7613 715 7652
rect 752 7613 767 7654
rect 696 7611 767 7613
rect 646 7593 767 7611
rect 438 7549 502 7552
rect 858 7549 962 7555
rect 1193 7549 1234 7699
rect 1612 7691 1639 7946
rect 1701 7936 1781 7947
rect 1701 7910 1718 7936
rect 1758 7910 1781 7936
rect 1701 7883 1781 7910
rect 1701 7857 1722 7883
rect 1762 7857 1781 7883
rect 1701 7838 1781 7857
rect 1701 7812 1725 7838
rect 1765 7812 1781 7838
rect 1701 7761 1781 7812
rect 2804 7938 2882 7973
rect 2804 7876 2886 7938
rect 2804 7853 2832 7876
rect 2858 7853 2886 7876
rect 2804 7833 2886 7853
rect 438 7546 1234 7549
rect 1613 7560 1639 7691
rect 1613 7546 1641 7560
rect 438 7511 1641 7546
rect 1703 7553 1773 7761
rect 438 7450 502 7511
rect 858 7509 962 7511
rect 1193 7509 1234 7511
rect 1703 7508 1724 7553
rect 1704 7487 1724 7508
rect 1754 7508 1773 7553
rect 1754 7487 1771 7508
rect 1704 7468 1771 7487
rect 1353 7460 1425 7461
rect 1352 7452 1451 7460
rect 440 7379 499 7450
rect 1352 7449 1404 7452
rect 1352 7414 1360 7449
rect 1385 7414 1404 7449
rect 1429 7441 1451 7452
rect 1429 7440 2296 7441
rect 1429 7414 2297 7440
rect 1352 7404 2297 7414
rect 1352 7402 1451 7404
rect 440 7361 462 7379
rect 480 7361 499 7379
rect 440 7339 499 7361
rect 707 7375 1239 7380
rect 707 7355 1593 7375
rect 1613 7355 1616 7375
rect 2252 7371 2297 7404
rect 707 7351 1616 7355
rect 707 7304 750 7351
rect 1200 7350 1616 7351
rect 2248 7351 2641 7371
rect 2661 7351 2664 7371
rect 1200 7349 1541 7350
rect 857 7318 967 7332
rect 857 7315 900 7318
rect 857 7310 861 7315
rect 695 7303 750 7304
rect 439 7280 750 7303
rect 439 7262 464 7280
rect 482 7268 750 7280
rect 779 7288 861 7310
rect 890 7288 900 7315
rect 928 7291 935 7318
rect 964 7310 967 7318
rect 964 7291 1029 7310
rect 928 7288 1029 7291
rect 779 7286 1029 7288
rect 482 7262 504 7268
rect 439 7123 504 7262
rect 779 7207 816 7286
rect 857 7273 967 7286
rect 931 7217 962 7218
rect 779 7187 788 7207
rect 808 7187 816 7207
rect 439 7105 462 7123
rect 480 7105 504 7123
rect 439 7088 504 7105
rect 659 7169 727 7182
rect 779 7177 816 7187
rect 875 7207 962 7217
rect 875 7187 884 7207
rect 904 7187 962 7207
rect 875 7178 962 7187
rect 875 7177 912 7178
rect 659 7127 666 7169
rect 715 7127 727 7169
rect 659 7124 727 7127
rect 931 7125 962 7178
rect 992 7207 1029 7286
rect 1144 7217 1175 7218
rect 992 7187 1001 7207
rect 1021 7187 1029 7207
rect 992 7177 1029 7187
rect 1088 7210 1175 7217
rect 1088 7207 1149 7210
rect 1088 7187 1097 7207
rect 1117 7190 1149 7207
rect 1170 7190 1175 7210
rect 1117 7187 1175 7190
rect 1088 7180 1175 7187
rect 1200 7207 1237 7349
rect 1503 7348 1540 7349
rect 2248 7346 2664 7351
rect 2248 7345 2589 7346
rect 1905 7314 2015 7328
rect 1905 7311 1948 7314
rect 1905 7306 1909 7311
rect 1827 7284 1909 7306
rect 1938 7284 1948 7311
rect 1976 7287 1983 7314
rect 2012 7306 2015 7314
rect 2012 7287 2077 7306
rect 1976 7284 2077 7287
rect 1827 7282 2077 7284
rect 1352 7217 1388 7218
rect 1200 7187 1209 7207
rect 1229 7187 1237 7207
rect 1088 7178 1144 7180
rect 1088 7177 1125 7178
rect 1200 7177 1237 7187
rect 1296 7207 1444 7217
rect 1544 7214 1640 7216
rect 1296 7187 1305 7207
rect 1325 7187 1415 7207
rect 1435 7187 1444 7207
rect 1296 7181 1444 7187
rect 1296 7178 1360 7181
rect 1296 7177 1333 7178
rect 1352 7151 1360 7178
rect 1381 7178 1444 7181
rect 1502 7207 1640 7214
rect 1502 7187 1511 7207
rect 1531 7187 1640 7207
rect 1502 7178 1640 7187
rect 1827 7203 1864 7282
rect 1905 7269 2015 7282
rect 1979 7213 2010 7214
rect 1827 7183 1836 7203
rect 1856 7183 1864 7203
rect 1381 7151 1388 7178
rect 1407 7177 1444 7178
rect 1503 7177 1540 7178
rect 1352 7126 1388 7151
rect 823 7124 864 7125
rect 659 7117 864 7124
rect 659 7106 833 7117
rect 659 7073 667 7106
rect 660 7064 667 7073
rect 716 7097 833 7106
rect 853 7097 864 7117
rect 716 7089 864 7097
rect 931 7121 1290 7125
rect 931 7116 1253 7121
rect 931 7092 1044 7116
rect 1068 7097 1253 7116
rect 1277 7097 1290 7121
rect 1068 7092 1290 7097
rect 931 7089 1290 7092
rect 1352 7089 1387 7126
rect 1455 7123 1555 7126
rect 1455 7119 1522 7123
rect 1455 7093 1467 7119
rect 1493 7097 1522 7119
rect 1548 7097 1555 7123
rect 1493 7093 1555 7097
rect 1455 7089 1555 7093
rect 716 7073 727 7089
rect 716 7064 724 7073
rect 931 7068 962 7089
rect 1352 7068 1388 7089
rect 774 7067 811 7068
rect 439 7024 504 7043
rect 439 7006 464 7024
rect 482 7006 504 7024
rect 439 6805 504 7006
rect 660 6880 724 7064
rect 773 7058 811 7067
rect 773 7038 782 7058
rect 802 7038 811 7058
rect 773 7030 811 7038
rect 877 7062 962 7068
rect 987 7067 1024 7068
rect 877 7042 885 7062
rect 905 7042 962 7062
rect 877 7034 962 7042
rect 986 7058 1024 7067
rect 986 7038 995 7058
rect 1015 7038 1024 7058
rect 877 7033 913 7034
rect 986 7030 1024 7038
rect 1090 7062 1175 7068
rect 1195 7067 1232 7068
rect 1090 7042 1098 7062
rect 1118 7061 1175 7062
rect 1118 7042 1147 7061
rect 1090 7041 1147 7042
rect 1168 7041 1175 7061
rect 1090 7034 1175 7041
rect 1194 7058 1232 7067
rect 1194 7038 1203 7058
rect 1223 7038 1232 7058
rect 1090 7033 1126 7034
rect 1194 7030 1232 7038
rect 1298 7062 1442 7068
rect 1298 7042 1306 7062
rect 1326 7042 1414 7062
rect 1434 7042 1442 7062
rect 1298 7034 1442 7042
rect 1298 7033 1334 7034
rect 1406 7033 1442 7034
rect 1508 7067 1545 7068
rect 1508 7066 1546 7067
rect 1508 7058 1572 7066
rect 1508 7038 1517 7058
rect 1537 7044 1572 7058
rect 1592 7044 1595 7064
rect 1537 7039 1595 7044
rect 1537 7038 1572 7039
rect 774 7001 811 7030
rect 775 6999 811 7001
rect 987 6999 1024 7030
rect 775 6977 1024 6999
rect 856 6971 967 6977
rect 856 6963 897 6971
rect 856 6943 864 6963
rect 883 6943 897 6963
rect 856 6941 897 6943
rect 925 6963 967 6971
rect 925 6943 941 6963
rect 960 6943 967 6963
rect 925 6941 967 6943
rect 856 6926 967 6941
rect 660 6870 728 6880
rect 660 6837 677 6870
rect 717 6837 728 6870
rect 660 6825 728 6837
rect 660 6823 724 6825
rect 1195 6806 1232 7030
rect 1508 7026 1572 7038
rect 1612 6808 1639 7178
rect 1827 7173 1864 7183
rect 1923 7203 2010 7213
rect 1923 7183 1932 7203
rect 1952 7183 2010 7203
rect 1923 7174 2010 7183
rect 1923 7173 1960 7174
rect 1703 7160 1773 7165
rect 1698 7154 1773 7160
rect 1698 7121 1706 7154
rect 1759 7121 1773 7154
rect 1979 7121 2010 7174
rect 2040 7203 2077 7282
rect 2192 7213 2223 7214
rect 2040 7183 2049 7203
rect 2069 7183 2077 7203
rect 2040 7173 2077 7183
rect 2136 7206 2223 7213
rect 2136 7203 2197 7206
rect 2136 7183 2145 7203
rect 2165 7186 2197 7203
rect 2218 7186 2223 7206
rect 2165 7183 2223 7186
rect 2136 7176 2223 7183
rect 2248 7203 2285 7345
rect 2551 7344 2588 7345
rect 2400 7213 2436 7214
rect 2248 7183 2257 7203
rect 2277 7183 2285 7203
rect 2136 7174 2192 7176
rect 2136 7173 2173 7174
rect 2248 7173 2285 7183
rect 2344 7203 2492 7213
rect 2592 7210 2688 7212
rect 2344 7183 2353 7203
rect 2373 7183 2463 7203
rect 2483 7183 2492 7203
rect 2344 7177 2492 7183
rect 2344 7174 2408 7177
rect 2344 7173 2381 7174
rect 2400 7147 2408 7174
rect 2429 7174 2492 7177
rect 2550 7203 2688 7210
rect 2550 7183 2559 7203
rect 2579 7183 2688 7203
rect 2550 7174 2688 7183
rect 2429 7147 2436 7174
rect 2455 7173 2492 7174
rect 2551 7173 2588 7174
rect 2400 7122 2436 7147
rect 1698 7120 1781 7121
rect 1871 7120 1912 7121
rect 1698 7113 1912 7120
rect 1698 7096 1881 7113
rect 1698 7063 1711 7096
rect 1764 7093 1881 7096
rect 1901 7093 1912 7113
rect 1764 7085 1912 7093
rect 1979 7117 2338 7121
rect 1979 7112 2301 7117
rect 1979 7088 2092 7112
rect 2116 7093 2301 7112
rect 2325 7093 2338 7117
rect 2116 7088 2338 7093
rect 1979 7085 2338 7088
rect 2400 7085 2435 7122
rect 2503 7119 2603 7122
rect 2503 7115 2570 7119
rect 2503 7089 2515 7115
rect 2541 7093 2570 7115
rect 2596 7093 2603 7119
rect 2541 7089 2603 7093
rect 2503 7085 2603 7089
rect 1764 7063 1781 7085
rect 1979 7064 2010 7085
rect 2400 7064 2436 7085
rect 1822 7063 1859 7064
rect 1698 7049 1781 7063
rect 1471 6806 1639 6808
rect 1195 6805 1639 6806
rect 439 6775 1639 6805
rect 1709 6839 1781 7049
rect 1821 7054 1859 7063
rect 1821 7034 1830 7054
rect 1850 7034 1859 7054
rect 1821 7026 1859 7034
rect 1925 7058 2010 7064
rect 2035 7063 2072 7064
rect 1925 7038 1933 7058
rect 1953 7038 2010 7058
rect 1925 7030 2010 7038
rect 2034 7054 2072 7063
rect 2034 7034 2043 7054
rect 2063 7034 2072 7054
rect 1925 7029 1961 7030
rect 2034 7026 2072 7034
rect 2138 7058 2223 7064
rect 2243 7063 2280 7064
rect 2138 7038 2146 7058
rect 2166 7057 2223 7058
rect 2166 7038 2195 7057
rect 2138 7037 2195 7038
rect 2216 7037 2223 7057
rect 2138 7030 2223 7037
rect 2242 7054 2280 7063
rect 2242 7034 2251 7054
rect 2271 7034 2280 7054
rect 2138 7029 2174 7030
rect 2242 7026 2280 7034
rect 2346 7058 2490 7064
rect 2346 7038 2354 7058
rect 2374 7038 2462 7058
rect 2482 7038 2490 7058
rect 2346 7030 2490 7038
rect 2346 7029 2382 7030
rect 2454 7029 2490 7030
rect 2556 7063 2593 7064
rect 2556 7062 2594 7063
rect 2556 7054 2620 7062
rect 2556 7034 2565 7054
rect 2585 7040 2620 7054
rect 2640 7040 2643 7060
rect 2585 7035 2643 7040
rect 2585 7034 2620 7035
rect 1822 6997 1859 7026
rect 1823 6995 1859 6997
rect 2035 6995 2072 7026
rect 1823 6973 2072 6995
rect 1904 6967 2015 6973
rect 1904 6959 1945 6967
rect 1904 6939 1912 6959
rect 1931 6939 1945 6959
rect 1904 6937 1945 6939
rect 1973 6959 2015 6967
rect 1973 6939 1989 6959
rect 2008 6939 2015 6959
rect 1973 6937 2015 6939
rect 1904 6922 2015 6937
rect 1709 6800 1728 6839
rect 1773 6800 1781 6839
rect 1709 6783 1781 6800
rect 2243 6827 2280 7026
rect 2556 7022 2620 7034
rect 2243 6821 2284 6827
rect 2660 6823 2687 7174
rect 2519 6821 2687 6823
rect 2243 6795 2687 6821
rect 439 6728 504 6775
rect 439 6710 462 6728
rect 480 6710 504 6728
rect 1352 6755 1387 6757
rect 1352 6753 1456 6755
rect 2245 6753 2284 6795
rect 2519 6794 2687 6795
rect 1352 6746 2286 6753
rect 1352 6745 1403 6746
rect 1352 6725 1355 6745
rect 1380 6726 1403 6745
rect 1435 6726 2286 6746
rect 1380 6725 2286 6726
rect 1352 6718 2286 6725
rect 1625 6717 2286 6718
rect 439 6689 504 6710
rect 716 6700 756 6703
rect 716 6696 1619 6700
rect 716 6676 1593 6696
rect 1613 6676 1619 6696
rect 716 6673 1619 6676
rect 440 6629 505 6649
rect 440 6611 464 6629
rect 482 6611 505 6629
rect 440 6584 505 6611
rect 716 6584 756 6673
rect 1200 6671 1616 6673
rect 1200 6670 1541 6671
rect 857 6639 967 6653
rect 857 6636 900 6639
rect 857 6631 861 6636
rect 439 6549 756 6584
rect 779 6609 861 6631
rect 890 6609 900 6636
rect 928 6612 935 6639
rect 964 6631 967 6639
rect 964 6612 1029 6631
rect 928 6609 1029 6612
rect 779 6607 1029 6609
rect 440 6473 505 6549
rect 779 6528 816 6607
rect 857 6594 967 6607
rect 931 6538 962 6539
rect 779 6508 788 6528
rect 808 6508 816 6528
rect 779 6498 816 6508
rect 875 6528 962 6538
rect 875 6508 884 6528
rect 904 6508 962 6528
rect 875 6499 962 6508
rect 875 6498 912 6499
rect 440 6455 462 6473
rect 480 6455 505 6473
rect 440 6434 505 6455
rect 653 6453 718 6462
rect 653 6416 663 6453
rect 703 6445 718 6453
rect 931 6446 962 6499
rect 992 6528 1029 6607
rect 1144 6538 1175 6539
rect 992 6508 1001 6528
rect 1021 6508 1029 6528
rect 992 6498 1029 6508
rect 1088 6531 1175 6538
rect 1088 6528 1149 6531
rect 1088 6508 1097 6528
rect 1117 6511 1149 6528
rect 1170 6511 1175 6531
rect 1117 6508 1175 6511
rect 1088 6501 1175 6508
rect 1200 6528 1237 6670
rect 1503 6669 1540 6670
rect 1352 6538 1388 6539
rect 1200 6508 1209 6528
rect 1229 6508 1237 6528
rect 1088 6499 1144 6501
rect 1088 6498 1125 6499
rect 1200 6498 1237 6508
rect 1296 6528 1444 6538
rect 1544 6535 1640 6537
rect 1296 6508 1305 6528
rect 1325 6508 1415 6528
rect 1435 6508 1444 6528
rect 1296 6502 1444 6508
rect 1296 6499 1360 6502
rect 1296 6498 1333 6499
rect 1352 6472 1360 6499
rect 1381 6499 1444 6502
rect 1502 6528 1640 6535
rect 1502 6508 1511 6528
rect 1531 6508 1640 6528
rect 1502 6499 1640 6508
rect 1381 6472 1388 6499
rect 1407 6498 1444 6499
rect 1503 6498 1540 6499
rect 1352 6447 1388 6472
rect 823 6445 864 6446
rect 703 6438 864 6445
rect 703 6418 833 6438
rect 853 6418 864 6438
rect 703 6416 864 6418
rect 653 6410 864 6416
rect 931 6442 1290 6446
rect 931 6437 1253 6442
rect 931 6413 1044 6437
rect 1068 6418 1253 6437
rect 1277 6418 1290 6442
rect 1068 6413 1290 6418
rect 931 6410 1290 6413
rect 1352 6410 1387 6447
rect 1455 6444 1555 6447
rect 1455 6440 1522 6444
rect 1455 6414 1467 6440
rect 1493 6418 1522 6440
rect 1548 6418 1555 6444
rect 1493 6414 1555 6418
rect 1455 6410 1555 6414
rect 653 6397 720 6410
rect 445 6374 501 6394
rect 445 6356 464 6374
rect 482 6356 501 6374
rect 445 6243 501 6356
rect 653 6376 667 6397
rect 703 6376 720 6397
rect 931 6389 962 6410
rect 1352 6389 1388 6410
rect 774 6388 811 6389
rect 653 6369 720 6376
rect 773 6379 811 6388
rect 445 6136 500 6243
rect 653 6217 718 6369
rect 773 6359 782 6379
rect 802 6359 811 6379
rect 773 6351 811 6359
rect 877 6383 962 6389
rect 987 6388 1024 6389
rect 877 6363 885 6383
rect 905 6363 962 6383
rect 877 6355 962 6363
rect 986 6379 1024 6388
rect 986 6359 995 6379
rect 1015 6359 1024 6379
rect 877 6354 913 6355
rect 986 6351 1024 6359
rect 1090 6383 1175 6389
rect 1195 6388 1232 6389
rect 1090 6363 1098 6383
rect 1118 6382 1175 6383
rect 1118 6363 1147 6382
rect 1090 6362 1147 6363
rect 1168 6362 1175 6382
rect 1090 6355 1175 6362
rect 1194 6379 1232 6388
rect 1194 6359 1203 6379
rect 1223 6359 1232 6379
rect 1090 6354 1126 6355
rect 1194 6351 1232 6359
rect 1298 6383 1442 6389
rect 1298 6363 1306 6383
rect 1326 6363 1414 6383
rect 1434 6363 1442 6383
rect 1298 6355 1442 6363
rect 1298 6354 1334 6355
rect 1406 6354 1442 6355
rect 1508 6388 1545 6389
rect 1508 6387 1546 6388
rect 1508 6379 1572 6387
rect 1508 6359 1517 6379
rect 1537 6365 1572 6379
rect 1592 6365 1595 6385
rect 1537 6360 1595 6365
rect 1537 6359 1572 6360
rect 774 6322 811 6351
rect 775 6320 811 6322
rect 987 6320 1024 6351
rect 775 6298 1024 6320
rect 856 6292 967 6298
rect 856 6284 897 6292
rect 856 6264 864 6284
rect 883 6264 897 6284
rect 856 6262 897 6264
rect 925 6284 967 6292
rect 925 6264 941 6284
rect 960 6264 967 6284
rect 925 6262 967 6264
rect 856 6247 967 6262
rect 1195 6252 1232 6351
rect 1508 6347 1572 6359
rect 858 6244 962 6247
rect 646 6207 767 6217
rect 646 6205 715 6207
rect 646 6164 659 6205
rect 696 6166 715 6205
rect 752 6166 767 6207
rect 696 6164 767 6166
rect 646 6146 767 6164
rect 438 6102 503 6136
rect 858 6102 962 6104
rect 1193 6102 1234 6252
rect 1612 6244 1639 6499
rect 1701 6489 1781 6500
rect 1701 6463 1718 6489
rect 1758 6463 1781 6489
rect 1701 6436 1781 6463
rect 1701 6410 1722 6436
rect 1762 6410 1781 6436
rect 1701 6391 1781 6410
rect 1701 6365 1725 6391
rect 1765 6365 1781 6391
rect 1701 6314 1781 6365
rect 438 6099 1234 6102
rect 1613 6113 1639 6244
rect 1703 6114 1773 6314
rect 1613 6099 1641 6113
rect 438 6064 1641 6099
rect 1702 6092 1774 6114
rect 438 5907 503 6064
rect 858 6062 962 6064
rect 1193 6062 1234 6064
rect 1702 6044 1716 6092
rect 1762 6044 1774 6092
rect 1702 6027 1774 6044
rect 2804 5994 2876 7833
rect 2982 6066 3074 9370
rect 3468 9353 3499 9374
rect 3889 9353 3925 9374
rect 3311 9352 3348 9353
rect 3310 9343 3348 9352
rect 3310 9323 3319 9343
rect 3339 9323 3348 9343
rect 3310 9315 3348 9323
rect 3414 9347 3499 9353
rect 3524 9352 3561 9353
rect 3414 9327 3422 9347
rect 3442 9327 3499 9347
rect 3414 9319 3499 9327
rect 3523 9343 3561 9352
rect 3523 9323 3532 9343
rect 3552 9323 3561 9343
rect 3414 9318 3450 9319
rect 3523 9315 3561 9323
rect 3627 9347 3712 9353
rect 3732 9352 3769 9353
rect 3627 9327 3635 9347
rect 3655 9346 3712 9347
rect 3655 9327 3684 9346
rect 3627 9326 3684 9327
rect 3705 9326 3712 9346
rect 3627 9319 3712 9326
rect 3731 9343 3769 9352
rect 3731 9323 3740 9343
rect 3760 9323 3769 9343
rect 3627 9318 3663 9319
rect 3731 9315 3769 9323
rect 3835 9347 3979 9353
rect 3835 9327 3843 9347
rect 3863 9327 3951 9347
rect 3971 9327 3979 9347
rect 3835 9319 3979 9327
rect 3835 9318 3871 9319
rect 3943 9318 3979 9319
rect 4045 9352 4082 9353
rect 4045 9351 4083 9352
rect 4045 9343 4109 9351
rect 4045 9323 4054 9343
rect 4074 9329 4109 9343
rect 4129 9329 4132 9349
rect 4074 9324 4132 9329
rect 4074 9323 4109 9324
rect 3311 9286 3348 9315
rect 3312 9284 3348 9286
rect 3524 9284 3561 9315
rect 3312 9262 3561 9284
rect 3393 9256 3504 9262
rect 3393 9248 3434 9256
rect 3393 9228 3401 9248
rect 3420 9228 3434 9248
rect 3393 9226 3434 9228
rect 3462 9248 3504 9256
rect 3462 9228 3478 9248
rect 3497 9228 3504 9248
rect 3462 9226 3504 9228
rect 3393 9211 3504 9226
rect 3732 9194 3769 9315
rect 4045 9311 4109 9323
rect 3850 9194 3879 9198
rect 4149 9196 4176 9463
rect 4008 9194 4176 9196
rect 3732 9168 4176 9194
rect 3691 8900 3736 8909
rect 3691 8862 3701 8900
rect 3726 8862 3736 8900
rect 3691 8851 3736 8862
rect 3694 8843 3736 8851
rect 3694 8138 3737 8843
rect 3850 8229 3879 9168
rect 4008 9167 4176 9168
rect 3848 8208 3885 8229
rect 3848 8171 3859 8208
rect 3876 8171 3885 8208
rect 3848 8161 3885 8171
rect 3694 8118 4088 8138
rect 4108 8118 4111 8138
rect 3695 8113 4111 8118
rect 3695 8112 4036 8113
rect 3352 8081 3462 8095
rect 3352 8078 3395 8081
rect 3352 8073 3356 8078
rect 3274 8051 3356 8073
rect 3385 8051 3395 8078
rect 3423 8054 3430 8081
rect 3459 8073 3462 8081
rect 3459 8054 3524 8073
rect 3423 8051 3524 8054
rect 3274 8049 3524 8051
rect 3274 7970 3311 8049
rect 3352 8036 3462 8049
rect 3426 7980 3457 7981
rect 3274 7950 3283 7970
rect 3303 7950 3311 7970
rect 3274 7940 3311 7950
rect 3370 7970 3457 7980
rect 3370 7950 3379 7970
rect 3399 7950 3457 7970
rect 3370 7941 3457 7950
rect 3370 7940 3407 7941
rect 3426 7888 3457 7941
rect 3487 7970 3524 8049
rect 3639 7980 3670 7981
rect 3487 7950 3496 7970
rect 3516 7950 3524 7970
rect 3487 7940 3524 7950
rect 3583 7973 3670 7980
rect 3583 7970 3644 7973
rect 3583 7950 3592 7970
rect 3612 7953 3644 7970
rect 3665 7953 3670 7973
rect 3612 7950 3670 7953
rect 3583 7943 3670 7950
rect 3695 7970 3732 8112
rect 3998 8111 4035 8112
rect 3847 7980 3883 7981
rect 3695 7950 3704 7970
rect 3724 7950 3732 7970
rect 3583 7941 3639 7943
rect 3583 7940 3620 7941
rect 3695 7940 3732 7950
rect 3791 7970 3939 7980
rect 4039 7977 4135 7979
rect 3791 7950 3800 7970
rect 3820 7950 3910 7970
rect 3930 7950 3939 7970
rect 3791 7944 3939 7950
rect 3791 7941 3855 7944
rect 3791 7940 3828 7941
rect 3847 7914 3855 7941
rect 3876 7941 3939 7944
rect 3997 7970 4135 7977
rect 3997 7950 4006 7970
rect 4026 7950 4135 7970
rect 3997 7941 4135 7950
rect 3876 7914 3883 7941
rect 3902 7940 3939 7941
rect 3998 7940 4035 7941
rect 3847 7889 3883 7914
rect 3318 7887 3359 7888
rect 3238 7882 3359 7887
rect 3189 7880 3359 7882
rect 3189 7869 3328 7880
rect 3189 7846 3212 7869
rect 3238 7860 3328 7869
rect 3348 7860 3359 7880
rect 3238 7852 3359 7860
rect 3426 7884 3785 7888
rect 3426 7879 3748 7884
rect 3426 7855 3539 7879
rect 3563 7860 3748 7879
rect 3772 7860 3785 7884
rect 3563 7855 3785 7860
rect 3426 7852 3785 7855
rect 3847 7852 3882 7889
rect 3950 7886 4050 7889
rect 3950 7882 4017 7886
rect 3950 7856 3962 7882
rect 3988 7860 4017 7882
rect 4043 7860 4050 7886
rect 3988 7856 4050 7860
rect 3950 7852 4050 7856
rect 3238 7846 3246 7852
rect 3189 7838 3246 7846
rect 3426 7831 3457 7852
rect 3847 7831 3883 7852
rect 3269 7830 3306 7831
rect 3268 7821 3306 7830
rect 3268 7801 3277 7821
rect 3297 7801 3306 7821
rect 3268 7793 3306 7801
rect 3372 7825 3457 7831
rect 3482 7830 3519 7831
rect 3372 7805 3380 7825
rect 3400 7805 3457 7825
rect 3372 7797 3457 7805
rect 3481 7821 3519 7830
rect 3481 7801 3490 7821
rect 3510 7801 3519 7821
rect 3372 7796 3408 7797
rect 3481 7793 3519 7801
rect 3585 7825 3670 7831
rect 3690 7830 3727 7831
rect 3585 7805 3593 7825
rect 3613 7824 3670 7825
rect 3613 7805 3642 7824
rect 3585 7804 3642 7805
rect 3663 7804 3670 7824
rect 3585 7797 3670 7804
rect 3689 7821 3727 7830
rect 3689 7801 3698 7821
rect 3718 7801 3727 7821
rect 3585 7796 3621 7797
rect 3689 7793 3727 7801
rect 3793 7825 3937 7831
rect 3793 7805 3801 7825
rect 3821 7805 3909 7825
rect 3929 7805 3937 7825
rect 3793 7797 3937 7805
rect 3793 7796 3829 7797
rect 3901 7796 3937 7797
rect 4003 7830 4040 7831
rect 4003 7829 4041 7830
rect 4003 7821 4067 7829
rect 4003 7801 4012 7821
rect 4032 7807 4067 7821
rect 4087 7807 4090 7827
rect 4032 7802 4090 7807
rect 4032 7801 4067 7802
rect 3269 7764 3306 7793
rect 3270 7762 3306 7764
rect 3482 7762 3519 7793
rect 3270 7740 3519 7762
rect 3351 7734 3462 7740
rect 3351 7726 3392 7734
rect 3351 7706 3359 7726
rect 3378 7706 3392 7726
rect 3351 7704 3392 7706
rect 3420 7726 3462 7734
rect 3420 7706 3436 7726
rect 3455 7706 3462 7726
rect 3420 7704 3462 7706
rect 3351 7689 3462 7704
rect 3690 7678 3727 7793
rect 4003 7789 4067 7801
rect 3683 7672 3730 7678
rect 4107 7674 4134 7941
rect 3966 7672 4134 7674
rect 3683 7646 4134 7672
rect 3683 7511 3730 7646
rect 3966 7645 4134 7646
rect 3681 7462 3740 7511
rect 3681 7434 3699 7462
rect 3727 7434 3740 7462
rect 3681 7424 3740 7434
rect 4796 6687 4874 9727
rect 4796 6667 5196 6687
rect 5216 6667 5219 6687
rect 4796 6665 5219 6667
rect 4803 6662 5219 6665
rect 4803 6661 5144 6662
rect 4460 6630 4570 6644
rect 4460 6627 4503 6630
rect 4460 6622 4464 6627
rect 4382 6600 4464 6622
rect 4493 6600 4503 6627
rect 4531 6603 4538 6630
rect 4567 6622 4570 6630
rect 4567 6603 4632 6622
rect 4531 6600 4632 6603
rect 4382 6598 4632 6600
rect 4382 6519 4419 6598
rect 4460 6585 4570 6598
rect 4534 6529 4565 6530
rect 4382 6499 4391 6519
rect 4411 6499 4419 6519
rect 4382 6489 4419 6499
rect 4478 6519 4565 6529
rect 4478 6499 4487 6519
rect 4507 6499 4565 6519
rect 4478 6490 4565 6499
rect 4478 6489 4515 6490
rect 4252 6436 4363 6439
rect 4534 6437 4565 6490
rect 4595 6519 4632 6598
rect 4747 6529 4778 6530
rect 4595 6499 4604 6519
rect 4624 6499 4632 6519
rect 4595 6489 4632 6499
rect 4691 6522 4778 6529
rect 4691 6519 4752 6522
rect 4691 6499 4700 6519
rect 4720 6502 4752 6519
rect 4773 6502 4778 6522
rect 4720 6499 4778 6502
rect 4691 6492 4778 6499
rect 4803 6519 4840 6661
rect 5106 6660 5143 6661
rect 4955 6529 4991 6530
rect 4803 6499 4812 6519
rect 4832 6499 4840 6519
rect 4691 6490 4747 6492
rect 4691 6489 4728 6490
rect 4803 6489 4840 6499
rect 4899 6519 5047 6529
rect 5147 6526 5243 6528
rect 4899 6499 4908 6519
rect 4928 6499 5018 6519
rect 5038 6499 5047 6519
rect 4899 6493 5047 6499
rect 4899 6490 4963 6493
rect 4899 6489 4936 6490
rect 4955 6463 4963 6490
rect 4984 6490 5047 6493
rect 5105 6519 5243 6526
rect 5105 6499 5114 6519
rect 5134 6499 5243 6519
rect 5105 6490 5243 6499
rect 4984 6463 4991 6490
rect 5010 6489 5047 6490
rect 5106 6489 5143 6490
rect 4955 6438 4991 6463
rect 4426 6436 4467 6437
rect 4252 6429 4467 6436
rect 4252 6428 4317 6429
rect 4252 6404 4260 6428
rect 4284 6405 4317 6428
rect 4341 6409 4436 6429
rect 4456 6409 4467 6429
rect 4341 6405 4467 6409
rect 4284 6404 4467 6405
rect 4252 6401 4467 6404
rect 4534 6433 4893 6437
rect 4534 6428 4856 6433
rect 4534 6404 4647 6428
rect 4671 6409 4856 6428
rect 4880 6409 4893 6433
rect 4671 6404 4893 6409
rect 4534 6401 4893 6404
rect 4955 6401 4990 6438
rect 5058 6435 5158 6438
rect 5058 6431 5125 6435
rect 5058 6405 5070 6431
rect 5096 6409 5125 6431
rect 5151 6409 5158 6435
rect 5096 6405 5158 6409
rect 5058 6401 5158 6405
rect 4252 6397 4363 6401
rect 4534 6380 4565 6401
rect 4955 6380 4991 6401
rect 4377 6379 4414 6380
rect 4376 6370 4414 6379
rect 4376 6350 4385 6370
rect 4405 6350 4414 6370
rect 4376 6342 4414 6350
rect 4480 6374 4565 6380
rect 4590 6379 4627 6380
rect 4480 6354 4488 6374
rect 4508 6354 4565 6374
rect 4480 6346 4565 6354
rect 4589 6370 4627 6379
rect 4589 6350 4598 6370
rect 4618 6350 4627 6370
rect 4480 6345 4516 6346
rect 4589 6342 4627 6350
rect 4693 6374 4778 6380
rect 4798 6379 4835 6380
rect 4693 6354 4701 6374
rect 4721 6373 4778 6374
rect 4721 6354 4750 6373
rect 4693 6353 4750 6354
rect 4771 6353 4778 6373
rect 4693 6346 4778 6353
rect 4797 6370 4835 6379
rect 4797 6350 4806 6370
rect 4826 6350 4835 6370
rect 4693 6345 4729 6346
rect 4797 6342 4835 6350
rect 4901 6374 5045 6380
rect 4901 6354 4909 6374
rect 4929 6373 5017 6374
rect 4929 6354 4963 6373
rect 4901 6351 4963 6354
rect 4987 6354 5017 6373
rect 5037 6354 5045 6374
rect 4987 6351 5045 6354
rect 4901 6346 5045 6351
rect 4901 6345 4937 6346
rect 5009 6345 5045 6346
rect 5111 6379 5148 6380
rect 5111 6378 5149 6379
rect 5111 6370 5175 6378
rect 5111 6350 5120 6370
rect 5140 6356 5175 6370
rect 5195 6356 5198 6376
rect 5140 6351 5198 6356
rect 5140 6350 5175 6351
rect 4377 6313 4414 6342
rect 4378 6311 4414 6313
rect 4590 6311 4627 6342
rect 4378 6289 4627 6311
rect 4459 6283 4570 6289
rect 4459 6275 4500 6283
rect 4459 6255 4467 6275
rect 4486 6255 4500 6275
rect 4459 6253 4500 6255
rect 4528 6275 4570 6283
rect 4528 6255 4544 6275
rect 4563 6255 4570 6275
rect 4528 6253 4570 6255
rect 4459 6238 4570 6253
rect 4798 6227 4835 6342
rect 5111 6338 5175 6350
rect 4794 6221 4849 6227
rect 5215 6223 5242 6490
rect 5074 6221 5242 6223
rect 4794 6196 5242 6221
rect 5555 6281 5661 11614
rect 8827 11593 8907 11644
rect 8827 11567 8843 11593
rect 8883 11567 8907 11593
rect 8827 11548 8907 11567
rect 8827 11522 8846 11548
rect 8886 11522 8907 11548
rect 8827 11495 8907 11522
rect 8827 11469 8850 11495
rect 8890 11469 8907 11495
rect 8827 11458 8907 11469
rect 8969 11459 8996 11714
rect 9374 11706 9415 11856
rect 9646 11711 9750 11856
rect 9841 11794 9962 11812
rect 9841 11792 9912 11794
rect 9841 11751 9856 11792
rect 9893 11753 9912 11792
rect 9949 11753 9962 11794
rect 9893 11751 9962 11753
rect 9841 11741 9962 11751
rect 9036 11599 9100 11611
rect 9376 11607 9413 11706
rect 9641 11696 9752 11711
rect 9641 11694 9683 11696
rect 9641 11674 9648 11694
rect 9667 11674 9683 11694
rect 9641 11666 9683 11674
rect 9711 11694 9752 11696
rect 9711 11674 9725 11694
rect 9744 11674 9752 11694
rect 9711 11666 9752 11674
rect 9641 11660 9752 11666
rect 9584 11638 9833 11660
rect 9584 11607 9621 11638
rect 9797 11636 9833 11638
rect 9797 11607 9834 11636
rect 9036 11598 9071 11599
rect 9013 11593 9071 11598
rect 9013 11573 9016 11593
rect 9036 11579 9071 11593
rect 9091 11579 9100 11599
rect 9036 11571 9100 11579
rect 9062 11570 9100 11571
rect 9063 11569 9100 11570
rect 9166 11603 9202 11604
rect 9274 11603 9310 11604
rect 9166 11595 9310 11603
rect 9166 11575 9174 11595
rect 9194 11575 9282 11595
rect 9302 11575 9310 11595
rect 9166 11569 9310 11575
rect 9376 11599 9414 11607
rect 9482 11603 9518 11604
rect 9376 11579 9385 11599
rect 9405 11579 9414 11599
rect 9376 11570 9414 11579
rect 9433 11596 9518 11603
rect 9433 11576 9440 11596
rect 9461 11595 9518 11596
rect 9461 11576 9490 11595
rect 9433 11575 9490 11576
rect 9510 11575 9518 11595
rect 9376 11569 9413 11570
rect 9433 11569 9518 11575
rect 9584 11599 9622 11607
rect 9695 11603 9731 11604
rect 9584 11579 9593 11599
rect 9613 11579 9622 11599
rect 9584 11570 9622 11579
rect 9646 11595 9731 11603
rect 9646 11575 9703 11595
rect 9723 11575 9731 11595
rect 9584 11569 9621 11570
rect 9646 11569 9731 11575
rect 9797 11599 9835 11607
rect 9797 11579 9806 11599
rect 9826 11579 9835 11599
rect 9890 11589 9955 11741
rect 10108 11715 10163 11856
rect 9797 11570 9835 11579
rect 9888 11582 9955 11589
rect 9797 11569 9834 11570
rect 9220 11548 9256 11569
rect 9646 11548 9677 11569
rect 9888 11561 9905 11582
rect 9941 11561 9955 11582
rect 10107 11602 10163 11715
rect 10107 11584 10126 11602
rect 10144 11584 10163 11602
rect 10107 11564 10163 11584
rect 9888 11548 9955 11561
rect 9053 11544 9153 11548
rect 9053 11540 9115 11544
rect 9053 11514 9060 11540
rect 9086 11518 9115 11540
rect 9141 11518 9153 11544
rect 9086 11514 9153 11518
rect 9053 11511 9153 11514
rect 9221 11511 9256 11548
rect 9318 11545 9677 11548
rect 9318 11540 9540 11545
rect 9318 11516 9331 11540
rect 9355 11521 9540 11540
rect 9564 11521 9677 11545
rect 9355 11516 9677 11521
rect 9318 11512 9677 11516
rect 9744 11542 9955 11548
rect 9744 11540 9905 11542
rect 9744 11520 9755 11540
rect 9775 11520 9905 11540
rect 9744 11513 9905 11520
rect 9744 11512 9785 11513
rect 9220 11486 9256 11511
rect 9068 11459 9105 11460
rect 9164 11459 9201 11460
rect 9220 11459 9227 11486
rect 8968 11450 9106 11459
rect 8968 11430 9077 11450
rect 9097 11430 9106 11450
rect 8968 11423 9106 11430
rect 9164 11456 9227 11459
rect 9248 11459 9256 11486
rect 9275 11459 9312 11460
rect 9248 11456 9312 11459
rect 9164 11450 9312 11456
rect 9164 11430 9173 11450
rect 9193 11430 9283 11450
rect 9303 11430 9312 11450
rect 8968 11421 9064 11423
rect 9164 11420 9312 11430
rect 9371 11450 9408 11460
rect 9483 11459 9520 11460
rect 9464 11457 9520 11459
rect 9371 11430 9379 11450
rect 9399 11430 9408 11450
rect 9220 11419 9256 11420
rect 9068 11288 9105 11289
rect 9371 11288 9408 11430
rect 9433 11450 9520 11457
rect 9433 11447 9491 11450
rect 9433 11427 9438 11447
rect 9459 11430 9491 11447
rect 9511 11430 9520 11450
rect 9459 11427 9520 11430
rect 9433 11420 9520 11427
rect 9579 11450 9616 11460
rect 9579 11430 9587 11450
rect 9607 11430 9616 11450
rect 9433 11419 9464 11420
rect 9579 11351 9616 11430
rect 9646 11459 9677 11512
rect 9890 11505 9905 11513
rect 9945 11505 9955 11542
rect 9890 11496 9955 11505
rect 10103 11503 10168 11524
rect 10103 11485 10128 11503
rect 10146 11485 10168 11503
rect 9696 11459 9733 11460
rect 9646 11450 9733 11459
rect 9646 11430 9704 11450
rect 9724 11430 9733 11450
rect 9646 11420 9733 11430
rect 9792 11450 9829 11460
rect 9792 11430 9800 11450
rect 9820 11430 9829 11450
rect 9646 11419 9677 11420
rect 9641 11351 9751 11364
rect 9792 11351 9829 11430
rect 10103 11409 10168 11485
rect 9579 11349 9829 11351
rect 9579 11346 9680 11349
rect 9579 11327 9644 11346
rect 9641 11319 9644 11327
rect 9673 11319 9680 11346
rect 9708 11322 9718 11349
rect 9747 11327 9829 11349
rect 9852 11374 10169 11409
rect 9747 11322 9751 11327
rect 9708 11319 9751 11322
rect 9641 11305 9751 11319
rect 9067 11287 9408 11288
rect 8992 11285 9408 11287
rect 9852 11285 9892 11374
rect 10103 11347 10168 11374
rect 10103 11329 10126 11347
rect 10144 11329 10168 11347
rect 10103 11309 10168 11329
rect 8989 11282 9892 11285
rect 8989 11262 8995 11282
rect 9015 11262 9892 11282
rect 8989 11258 9892 11262
rect 9852 11255 9892 11258
rect 10104 11248 10169 11269
rect 8322 11240 8983 11241
rect 8322 11233 9256 11240
rect 8322 11232 9228 11233
rect 8322 11212 9173 11232
rect 9205 11213 9228 11232
rect 9253 11213 9256 11233
rect 9205 11212 9256 11213
rect 8322 11205 9256 11212
rect 7921 11163 8089 11164
rect 8324 11163 8363 11205
rect 9152 11203 9256 11205
rect 9221 11201 9256 11203
rect 10104 11230 10128 11248
rect 10146 11230 10169 11248
rect 10104 11183 10169 11230
rect 7921 11137 8365 11163
rect 7921 11135 8089 11137
rect 7921 10784 7948 11135
rect 8324 11131 8365 11137
rect 7988 10924 8052 10936
rect 8328 10932 8365 11131
rect 8827 11158 8899 11175
rect 8827 11119 8835 11158
rect 8880 11119 8899 11158
rect 8593 11021 8704 11036
rect 8593 11019 8635 11021
rect 8593 10999 8600 11019
rect 8619 10999 8635 11019
rect 8593 10991 8635 10999
rect 8663 11019 8704 11021
rect 8663 10999 8677 11019
rect 8696 10999 8704 11019
rect 8663 10991 8704 10999
rect 8593 10985 8704 10991
rect 8536 10963 8785 10985
rect 8536 10932 8573 10963
rect 8749 10961 8785 10963
rect 8749 10932 8786 10961
rect 7988 10923 8023 10924
rect 7965 10918 8023 10923
rect 7965 10898 7968 10918
rect 7988 10904 8023 10918
rect 8043 10904 8052 10924
rect 7988 10896 8052 10904
rect 8014 10895 8052 10896
rect 8015 10894 8052 10895
rect 8118 10928 8154 10929
rect 8226 10928 8262 10929
rect 8118 10920 8262 10928
rect 8118 10900 8126 10920
rect 8146 10900 8234 10920
rect 8254 10900 8262 10920
rect 8118 10894 8262 10900
rect 8328 10924 8366 10932
rect 8434 10928 8470 10929
rect 8328 10904 8337 10924
rect 8357 10904 8366 10924
rect 8328 10895 8366 10904
rect 8385 10921 8470 10928
rect 8385 10901 8392 10921
rect 8413 10920 8470 10921
rect 8413 10901 8442 10920
rect 8385 10900 8442 10901
rect 8462 10900 8470 10920
rect 8328 10894 8365 10895
rect 8385 10894 8470 10900
rect 8536 10924 8574 10932
rect 8647 10928 8683 10929
rect 8536 10904 8545 10924
rect 8565 10904 8574 10924
rect 8536 10895 8574 10904
rect 8598 10920 8683 10928
rect 8598 10900 8655 10920
rect 8675 10900 8683 10920
rect 8536 10894 8573 10895
rect 8598 10894 8683 10900
rect 8749 10924 8787 10932
rect 8749 10904 8758 10924
rect 8778 10904 8787 10924
rect 8749 10895 8787 10904
rect 8827 10909 8899 11119
rect 8969 11153 10169 11183
rect 8969 11152 9413 11153
rect 8969 11150 9137 11152
rect 8827 10895 8910 10909
rect 8749 10894 8786 10895
rect 8172 10873 8208 10894
rect 8598 10873 8629 10894
rect 8827 10873 8844 10895
rect 8005 10869 8105 10873
rect 8005 10865 8067 10869
rect 8005 10839 8012 10865
rect 8038 10843 8067 10865
rect 8093 10843 8105 10869
rect 8038 10839 8105 10843
rect 8005 10836 8105 10839
rect 8173 10836 8208 10873
rect 8270 10870 8629 10873
rect 8270 10865 8492 10870
rect 8270 10841 8283 10865
rect 8307 10846 8492 10865
rect 8516 10846 8629 10870
rect 8307 10841 8629 10846
rect 8270 10837 8629 10841
rect 8696 10865 8844 10873
rect 8696 10845 8707 10865
rect 8727 10862 8844 10865
rect 8897 10862 8910 10895
rect 8727 10845 8910 10862
rect 8696 10838 8910 10845
rect 8696 10837 8737 10838
rect 8827 10837 8910 10838
rect 8172 10811 8208 10836
rect 8020 10784 8057 10785
rect 8116 10784 8153 10785
rect 8172 10784 8179 10811
rect 7920 10775 8058 10784
rect 7920 10755 8029 10775
rect 8049 10755 8058 10775
rect 7920 10748 8058 10755
rect 8116 10781 8179 10784
rect 8200 10784 8208 10811
rect 8227 10784 8264 10785
rect 8200 10781 8264 10784
rect 8116 10775 8264 10781
rect 8116 10755 8125 10775
rect 8145 10755 8235 10775
rect 8255 10755 8264 10775
rect 7920 10746 8016 10748
rect 8116 10745 8264 10755
rect 8323 10775 8360 10785
rect 8435 10784 8472 10785
rect 8416 10782 8472 10784
rect 8323 10755 8331 10775
rect 8351 10755 8360 10775
rect 8172 10744 8208 10745
rect 8020 10613 8057 10614
rect 8323 10613 8360 10755
rect 8385 10775 8472 10782
rect 8385 10772 8443 10775
rect 8385 10752 8390 10772
rect 8411 10755 8443 10772
rect 8463 10755 8472 10775
rect 8411 10752 8472 10755
rect 8385 10745 8472 10752
rect 8531 10775 8568 10785
rect 8531 10755 8539 10775
rect 8559 10755 8568 10775
rect 8385 10744 8416 10745
rect 8531 10676 8568 10755
rect 8598 10784 8629 10837
rect 8835 10804 8849 10837
rect 8902 10804 8910 10837
rect 8835 10798 8910 10804
rect 8835 10793 8905 10798
rect 8648 10784 8685 10785
rect 8598 10775 8685 10784
rect 8598 10755 8656 10775
rect 8676 10755 8685 10775
rect 8598 10745 8685 10755
rect 8744 10775 8781 10785
rect 8969 10780 8996 11150
rect 9036 10920 9100 10932
rect 9376 10928 9413 11152
rect 9884 11133 9948 11135
rect 9880 11121 9948 11133
rect 9880 11088 9891 11121
rect 9931 11088 9948 11121
rect 9880 11078 9948 11088
rect 9641 11017 9752 11032
rect 9641 11015 9683 11017
rect 9641 10995 9648 11015
rect 9667 10995 9683 11015
rect 9641 10987 9683 10995
rect 9711 11015 9752 11017
rect 9711 10995 9725 11015
rect 9744 10995 9752 11015
rect 9711 10987 9752 10995
rect 9641 10981 9752 10987
rect 9584 10959 9833 10981
rect 9584 10928 9621 10959
rect 9797 10957 9833 10959
rect 9797 10928 9834 10957
rect 9036 10919 9071 10920
rect 9013 10914 9071 10919
rect 9013 10894 9016 10914
rect 9036 10900 9071 10914
rect 9091 10900 9100 10920
rect 9036 10892 9100 10900
rect 9062 10891 9100 10892
rect 9063 10890 9100 10891
rect 9166 10924 9202 10925
rect 9274 10924 9310 10925
rect 9166 10916 9310 10924
rect 9166 10896 9174 10916
rect 9194 10896 9282 10916
rect 9302 10896 9310 10916
rect 9166 10890 9310 10896
rect 9376 10920 9414 10928
rect 9482 10924 9518 10925
rect 9376 10900 9385 10920
rect 9405 10900 9414 10920
rect 9376 10891 9414 10900
rect 9433 10917 9518 10924
rect 9433 10897 9440 10917
rect 9461 10916 9518 10917
rect 9461 10897 9490 10916
rect 9433 10896 9490 10897
rect 9510 10896 9518 10916
rect 9376 10890 9413 10891
rect 9433 10890 9518 10896
rect 9584 10920 9622 10928
rect 9695 10924 9731 10925
rect 9584 10900 9593 10920
rect 9613 10900 9622 10920
rect 9584 10891 9622 10900
rect 9646 10916 9731 10924
rect 9646 10896 9703 10916
rect 9723 10896 9731 10916
rect 9584 10890 9621 10891
rect 9646 10890 9731 10896
rect 9797 10920 9835 10928
rect 9797 10900 9806 10920
rect 9826 10900 9835 10920
rect 9797 10891 9835 10900
rect 9884 10894 9948 11078
rect 10104 10952 10169 11153
rect 10104 10934 10126 10952
rect 10144 10934 10169 10952
rect 10104 10915 10169 10934
rect 9797 10890 9834 10891
rect 9220 10869 9256 10890
rect 9646 10869 9677 10890
rect 9884 10885 9892 10894
rect 9881 10869 9892 10885
rect 9053 10865 9153 10869
rect 9053 10861 9115 10865
rect 9053 10835 9060 10861
rect 9086 10839 9115 10861
rect 9141 10839 9153 10865
rect 9086 10835 9153 10839
rect 9053 10832 9153 10835
rect 9221 10832 9256 10869
rect 9318 10866 9677 10869
rect 9318 10861 9540 10866
rect 9318 10837 9331 10861
rect 9355 10842 9540 10861
rect 9564 10842 9677 10866
rect 9355 10837 9677 10842
rect 9318 10833 9677 10837
rect 9744 10861 9892 10869
rect 9744 10841 9755 10861
rect 9775 10852 9892 10861
rect 9941 10885 9948 10894
rect 9941 10852 9949 10885
rect 9775 10841 9949 10852
rect 9744 10834 9949 10841
rect 9744 10833 9785 10834
rect 9220 10807 9256 10832
rect 9068 10780 9105 10781
rect 9164 10780 9201 10781
rect 9220 10780 9227 10807
rect 8744 10755 8752 10775
rect 8772 10755 8781 10775
rect 8598 10744 8629 10745
rect 8593 10676 8703 10689
rect 8744 10676 8781 10755
rect 8968 10771 9106 10780
rect 8968 10751 9077 10771
rect 9097 10751 9106 10771
rect 8968 10744 9106 10751
rect 9164 10777 9227 10780
rect 9248 10780 9256 10807
rect 9275 10780 9312 10781
rect 9248 10777 9312 10780
rect 9164 10771 9312 10777
rect 9164 10751 9173 10771
rect 9193 10751 9283 10771
rect 9303 10751 9312 10771
rect 8968 10742 9064 10744
rect 9164 10741 9312 10751
rect 9371 10771 9408 10781
rect 9483 10780 9520 10781
rect 9464 10778 9520 10780
rect 9371 10751 9379 10771
rect 9399 10751 9408 10771
rect 9220 10740 9256 10741
rect 8531 10674 8781 10676
rect 8531 10671 8632 10674
rect 8531 10652 8596 10671
rect 8593 10644 8596 10652
rect 8625 10644 8632 10671
rect 8660 10647 8670 10674
rect 8699 10652 8781 10674
rect 8699 10647 8703 10652
rect 8660 10644 8703 10647
rect 8593 10630 8703 10644
rect 8019 10612 8360 10613
rect 7944 10607 8360 10612
rect 9068 10609 9105 10610
rect 9371 10609 9408 10751
rect 9433 10771 9520 10778
rect 9433 10768 9491 10771
rect 9433 10748 9438 10768
rect 9459 10751 9491 10768
rect 9511 10751 9520 10771
rect 9459 10748 9520 10751
rect 9433 10741 9520 10748
rect 9579 10771 9616 10781
rect 9579 10751 9587 10771
rect 9607 10751 9616 10771
rect 9433 10740 9464 10741
rect 9579 10672 9616 10751
rect 9646 10780 9677 10833
rect 9881 10831 9949 10834
rect 9881 10789 9893 10831
rect 9942 10789 9949 10831
rect 9696 10780 9733 10781
rect 9646 10771 9733 10780
rect 9646 10751 9704 10771
rect 9724 10751 9733 10771
rect 9646 10741 9733 10751
rect 9792 10771 9829 10781
rect 9881 10776 9949 10789
rect 10104 10853 10169 10870
rect 10104 10835 10128 10853
rect 10146 10835 10169 10853
rect 9792 10751 9800 10771
rect 9820 10751 9829 10771
rect 9646 10740 9677 10741
rect 9641 10672 9751 10685
rect 9792 10672 9829 10751
rect 10104 10696 10169 10835
rect 10104 10690 10126 10696
rect 9579 10670 9829 10672
rect 9579 10667 9680 10670
rect 9579 10648 9644 10667
rect 9641 10640 9644 10648
rect 9673 10640 9680 10667
rect 9708 10643 9718 10670
rect 9747 10648 9829 10670
rect 9858 10678 10126 10690
rect 10144 10678 10169 10696
rect 9858 10655 10169 10678
rect 9858 10654 9913 10655
rect 9747 10643 9751 10648
rect 9708 10640 9751 10643
rect 9641 10626 9751 10640
rect 9067 10608 9408 10609
rect 7944 10587 7947 10607
rect 7967 10587 8360 10607
rect 8992 10607 9408 10608
rect 9858 10607 9901 10654
rect 8992 10603 9901 10607
rect 8311 10554 8356 10587
rect 8992 10583 8995 10603
rect 9015 10583 9901 10603
rect 9369 10578 9901 10583
rect 10109 10597 10168 10619
rect 10109 10579 10128 10597
rect 10146 10579 10168 10597
rect 9157 10554 9256 10556
rect 8311 10544 9256 10554
rect 6868 10524 6927 10534
rect 6868 10496 6881 10524
rect 6909 10496 6927 10524
rect 8311 10518 9179 10544
rect 8312 10517 9179 10518
rect 9157 10506 9179 10517
rect 9204 10509 9223 10544
rect 9248 10509 9256 10544
rect 9204 10506 9256 10509
rect 10109 10508 10168 10579
rect 9157 10498 9256 10506
rect 9183 10497 9255 10498
rect 6868 10447 6927 10496
rect 8837 10471 8904 10490
rect 8837 10450 8854 10471
rect 6474 10312 6642 10313
rect 6878 10312 6925 10447
rect 6474 10286 6925 10312
rect 6474 10284 6642 10286
rect 6474 10017 6501 10284
rect 6878 10280 6925 10286
rect 8835 10405 8854 10450
rect 8884 10450 8904 10471
rect 8884 10405 8905 10450
rect 9374 10447 9415 10449
rect 9646 10447 9750 10449
rect 10106 10447 10170 10508
rect 6541 10157 6605 10169
rect 6881 10165 6918 10280
rect 7146 10254 7257 10269
rect 7146 10252 7188 10254
rect 7146 10232 7153 10252
rect 7172 10232 7188 10252
rect 7146 10224 7188 10232
rect 7216 10252 7257 10254
rect 7216 10232 7230 10252
rect 7249 10232 7257 10252
rect 7216 10224 7257 10232
rect 7146 10218 7257 10224
rect 7089 10196 7338 10218
rect 8835 10197 8905 10405
rect 8967 10412 10170 10447
rect 8967 10398 8995 10412
rect 8969 10267 8995 10398
rect 9374 10409 10170 10412
rect 7089 10165 7126 10196
rect 7302 10194 7338 10196
rect 7302 10165 7339 10194
rect 6541 10156 6576 10157
rect 6518 10151 6576 10156
rect 6518 10131 6521 10151
rect 6541 10137 6576 10151
rect 6596 10137 6605 10157
rect 6541 10129 6605 10137
rect 6567 10128 6605 10129
rect 6568 10127 6605 10128
rect 6671 10161 6707 10162
rect 6779 10161 6815 10162
rect 6671 10153 6815 10161
rect 6671 10133 6679 10153
rect 6699 10133 6787 10153
rect 6807 10133 6815 10153
rect 6671 10127 6815 10133
rect 6881 10157 6919 10165
rect 6987 10161 7023 10162
rect 6881 10137 6890 10157
rect 6910 10137 6919 10157
rect 6881 10128 6919 10137
rect 6938 10154 7023 10161
rect 6938 10134 6945 10154
rect 6966 10153 7023 10154
rect 6966 10134 6995 10153
rect 6938 10133 6995 10134
rect 7015 10133 7023 10153
rect 6881 10127 6918 10128
rect 6938 10127 7023 10133
rect 7089 10157 7127 10165
rect 7200 10161 7236 10162
rect 7089 10137 7098 10157
rect 7118 10137 7127 10157
rect 7089 10128 7127 10137
rect 7151 10153 7236 10161
rect 7151 10133 7208 10153
rect 7228 10133 7236 10153
rect 7089 10127 7126 10128
rect 7151 10127 7236 10133
rect 7302 10157 7340 10165
rect 7302 10137 7311 10157
rect 7331 10137 7340 10157
rect 7302 10128 7340 10137
rect 8827 10146 8907 10197
rect 7302 10127 7339 10128
rect 6725 10106 6761 10127
rect 7151 10106 7182 10127
rect 7362 10112 7419 10120
rect 7362 10106 7370 10112
rect 6558 10102 6658 10106
rect 6558 10098 6620 10102
rect 6558 10072 6565 10098
rect 6591 10076 6620 10098
rect 6646 10076 6658 10102
rect 6591 10072 6658 10076
rect 6558 10069 6658 10072
rect 6726 10069 6761 10106
rect 6823 10103 7182 10106
rect 6823 10098 7045 10103
rect 6823 10074 6836 10098
rect 6860 10079 7045 10098
rect 7069 10079 7182 10103
rect 6860 10074 7182 10079
rect 6823 10070 7182 10074
rect 7249 10098 7370 10106
rect 7249 10078 7260 10098
rect 7280 10089 7370 10098
rect 7396 10089 7419 10112
rect 7280 10078 7419 10089
rect 7249 10076 7419 10078
rect 7722 10105 7794 10125
rect 7722 10082 7750 10105
rect 7776 10082 7794 10105
rect 7249 10071 7370 10076
rect 7249 10070 7290 10071
rect 6725 10044 6761 10069
rect 6573 10017 6610 10018
rect 6669 10017 6706 10018
rect 6725 10017 6732 10044
rect 6473 10008 6611 10017
rect 6473 9988 6582 10008
rect 6602 9988 6611 10008
rect 6473 9981 6611 9988
rect 6669 10014 6732 10017
rect 6753 10017 6761 10044
rect 6780 10017 6817 10018
rect 6753 10014 6817 10017
rect 6669 10008 6817 10014
rect 6669 9988 6678 10008
rect 6698 9988 6788 10008
rect 6808 9988 6817 10008
rect 6473 9979 6569 9981
rect 6669 9978 6817 9988
rect 6876 10008 6913 10018
rect 6988 10017 7025 10018
rect 6969 10015 7025 10017
rect 6876 9988 6884 10008
rect 6904 9988 6913 10008
rect 6725 9977 6761 9978
rect 6573 9846 6610 9847
rect 6876 9846 6913 9988
rect 6938 10008 7025 10015
rect 6938 10005 6996 10008
rect 6938 9985 6943 10005
rect 6964 9988 6996 10005
rect 7016 9988 7025 10008
rect 6964 9985 7025 9988
rect 6938 9978 7025 9985
rect 7084 10008 7121 10018
rect 7084 9988 7092 10008
rect 7112 9988 7121 10008
rect 6938 9977 6969 9978
rect 7084 9909 7121 9988
rect 7151 10017 7182 10070
rect 7722 10020 7794 10082
rect 8827 10120 8843 10146
rect 8883 10120 8907 10146
rect 8827 10101 8907 10120
rect 8827 10075 8846 10101
rect 8886 10075 8907 10101
rect 8827 10048 8907 10075
rect 8827 10022 8850 10048
rect 8890 10022 8907 10048
rect 7201 10017 7238 10018
rect 7151 10008 7238 10017
rect 7151 9988 7209 10008
rect 7229 9988 7238 10008
rect 7151 9978 7238 9988
rect 7297 10008 7334 10018
rect 7297 9988 7305 10008
rect 7325 9988 7334 10008
rect 7151 9977 7182 9978
rect 7146 9909 7256 9922
rect 7297 9909 7334 9988
rect 7084 9907 7334 9909
rect 7084 9904 7185 9907
rect 7084 9885 7149 9904
rect 7146 9877 7149 9885
rect 7178 9877 7185 9904
rect 7213 9880 7223 9907
rect 7252 9885 7334 9907
rect 7252 9880 7256 9885
rect 7213 9877 7256 9880
rect 7146 9863 7256 9877
rect 6572 9845 6913 9846
rect 6497 9840 6913 9845
rect 6497 9820 6500 9840
rect 6520 9820 6914 9840
rect 6723 9787 6760 9797
rect 6723 9750 6732 9787
rect 6749 9750 6760 9787
rect 6723 9729 6760 9750
rect 6432 8790 6600 8791
rect 6729 8790 6758 9729
rect 6871 9115 6914 9820
rect 7726 9469 7788 10020
rect 8827 10011 8907 10022
rect 8969 10012 8996 10267
rect 9374 10259 9415 10409
rect 9646 10403 9750 10409
rect 10106 10406 10170 10409
rect 9841 10347 9962 10365
rect 9841 10345 9912 10347
rect 9841 10304 9856 10345
rect 9893 10306 9912 10345
rect 9949 10306 9962 10347
rect 9893 10304 9962 10306
rect 9841 10294 9962 10304
rect 9036 10152 9100 10164
rect 9376 10160 9413 10259
rect 9641 10249 9752 10262
rect 9641 10247 9683 10249
rect 9641 10227 9648 10247
rect 9667 10227 9683 10247
rect 9641 10219 9683 10227
rect 9711 10247 9752 10249
rect 9711 10227 9725 10247
rect 9744 10227 9752 10247
rect 9711 10219 9752 10227
rect 9641 10213 9752 10219
rect 9584 10191 9833 10213
rect 9584 10160 9621 10191
rect 9797 10189 9833 10191
rect 9797 10160 9834 10189
rect 9036 10151 9071 10152
rect 9013 10146 9071 10151
rect 9013 10126 9016 10146
rect 9036 10132 9071 10146
rect 9091 10132 9100 10152
rect 9036 10124 9100 10132
rect 9062 10123 9100 10124
rect 9063 10122 9100 10123
rect 9166 10156 9202 10157
rect 9274 10156 9310 10157
rect 9166 10148 9310 10156
rect 9166 10128 9174 10148
rect 9194 10128 9282 10148
rect 9302 10128 9310 10148
rect 9166 10122 9310 10128
rect 9376 10152 9414 10160
rect 9482 10156 9518 10157
rect 9376 10132 9385 10152
rect 9405 10132 9414 10152
rect 9376 10123 9414 10132
rect 9433 10149 9518 10156
rect 9433 10129 9440 10149
rect 9461 10148 9518 10149
rect 9461 10129 9490 10148
rect 9433 10128 9490 10129
rect 9510 10128 9518 10148
rect 9376 10122 9413 10123
rect 9433 10122 9518 10128
rect 9584 10152 9622 10160
rect 9695 10156 9731 10157
rect 9584 10132 9593 10152
rect 9613 10132 9622 10152
rect 9584 10123 9622 10132
rect 9646 10148 9731 10156
rect 9646 10128 9703 10148
rect 9723 10128 9731 10148
rect 9584 10122 9621 10123
rect 9646 10122 9731 10128
rect 9797 10152 9835 10160
rect 9797 10132 9806 10152
rect 9826 10132 9835 10152
rect 9890 10142 9955 10294
rect 10108 10268 10163 10406
rect 9797 10123 9835 10132
rect 9888 10135 9955 10142
rect 9797 10122 9834 10123
rect 9220 10101 9256 10122
rect 9646 10101 9677 10122
rect 9888 10114 9905 10135
rect 9941 10114 9955 10135
rect 10107 10155 10163 10268
rect 10107 10137 10126 10155
rect 10144 10137 10163 10155
rect 10107 10117 10163 10137
rect 9888 10101 9955 10114
rect 9053 10097 9153 10101
rect 9053 10093 9115 10097
rect 9053 10067 9060 10093
rect 9086 10071 9115 10093
rect 9141 10071 9153 10097
rect 9086 10067 9153 10071
rect 9053 10064 9153 10067
rect 9221 10064 9256 10101
rect 9318 10098 9677 10101
rect 9318 10093 9540 10098
rect 9318 10069 9331 10093
rect 9355 10074 9540 10093
rect 9564 10074 9677 10098
rect 9355 10069 9677 10074
rect 9318 10065 9677 10069
rect 9744 10095 9955 10101
rect 9744 10093 9905 10095
rect 9744 10073 9755 10093
rect 9775 10073 9905 10093
rect 9744 10066 9905 10073
rect 9744 10065 9785 10066
rect 9220 10039 9256 10064
rect 9068 10012 9105 10013
rect 9164 10012 9201 10013
rect 9220 10012 9227 10039
rect 8968 10003 9106 10012
rect 8968 9983 9077 10003
rect 9097 9983 9106 10003
rect 8968 9976 9106 9983
rect 9164 10009 9227 10012
rect 9248 10012 9256 10039
rect 9275 10012 9312 10013
rect 9248 10009 9312 10012
rect 9164 10003 9312 10009
rect 9164 9983 9173 10003
rect 9193 9983 9283 10003
rect 9303 9983 9312 10003
rect 8968 9974 9064 9976
rect 9164 9973 9312 9983
rect 9371 10003 9408 10013
rect 9483 10012 9520 10013
rect 9464 10010 9520 10012
rect 9371 9983 9379 10003
rect 9399 9983 9408 10003
rect 9220 9972 9256 9973
rect 9068 9841 9105 9842
rect 9371 9841 9408 9983
rect 9433 10003 9520 10010
rect 9433 10000 9491 10003
rect 9433 9980 9438 10000
rect 9459 9983 9491 10000
rect 9511 9983 9520 10003
rect 9459 9980 9520 9983
rect 9433 9973 9520 9980
rect 9579 10003 9616 10013
rect 9579 9983 9587 10003
rect 9607 9983 9616 10003
rect 9433 9972 9464 9973
rect 9579 9904 9616 9983
rect 9646 10012 9677 10065
rect 9890 10058 9905 10066
rect 9945 10058 9955 10095
rect 9890 10049 9955 10058
rect 10103 10056 10168 10077
rect 10103 10038 10128 10056
rect 10146 10038 10168 10056
rect 9696 10012 9733 10013
rect 9646 10003 9733 10012
rect 9646 9983 9704 10003
rect 9724 9983 9733 10003
rect 9646 9973 9733 9983
rect 9792 10003 9829 10013
rect 9792 9983 9800 10003
rect 9820 9983 9829 10003
rect 9646 9972 9677 9973
rect 9641 9904 9751 9917
rect 9792 9904 9829 9983
rect 10103 9962 10168 10038
rect 9579 9902 9829 9904
rect 9579 9899 9680 9902
rect 9579 9880 9644 9899
rect 9641 9872 9644 9880
rect 9673 9872 9680 9899
rect 9708 9875 9718 9902
rect 9747 9880 9829 9902
rect 9852 9927 10169 9962
rect 9747 9875 9751 9880
rect 9708 9872 9751 9875
rect 9641 9858 9751 9872
rect 9067 9840 9408 9841
rect 8992 9838 9408 9840
rect 9852 9838 9892 9927
rect 10103 9900 10168 9927
rect 10103 9882 10126 9900
rect 10144 9882 10168 9900
rect 10103 9862 10168 9882
rect 8989 9835 9892 9838
rect 8989 9815 8995 9835
rect 9015 9815 9892 9835
rect 8989 9811 9892 9815
rect 9852 9808 9892 9811
rect 10104 9801 10169 9822
rect 8322 9793 8983 9794
rect 8322 9786 9256 9793
rect 8322 9785 9228 9786
rect 8322 9765 9173 9785
rect 9205 9766 9228 9785
rect 9253 9766 9256 9786
rect 9205 9765 9256 9766
rect 8322 9758 9256 9765
rect 7921 9716 8089 9717
rect 8324 9716 8363 9758
rect 9152 9756 9256 9758
rect 9221 9754 9256 9756
rect 10104 9783 10128 9801
rect 10146 9783 10169 9801
rect 10104 9736 10169 9783
rect 7921 9690 8365 9716
rect 7921 9688 8089 9690
rect 7723 9385 7792 9469
rect 6872 9107 6914 9115
rect 6872 9096 6917 9107
rect 6872 9058 6882 9096
rect 6907 9058 6917 9096
rect 6872 9049 6917 9058
rect 7721 8906 7792 9385
rect 7921 9337 7948 9688
rect 8324 9684 8365 9690
rect 7988 9477 8052 9489
rect 8328 9485 8365 9684
rect 8827 9711 8899 9728
rect 8827 9672 8835 9711
rect 8880 9672 8899 9711
rect 8593 9574 8704 9589
rect 8593 9572 8635 9574
rect 8593 9552 8600 9572
rect 8619 9552 8635 9572
rect 8593 9544 8635 9552
rect 8663 9572 8704 9574
rect 8663 9552 8677 9572
rect 8696 9552 8704 9572
rect 8663 9544 8704 9552
rect 8593 9538 8704 9544
rect 8536 9516 8785 9538
rect 8536 9485 8573 9516
rect 8749 9514 8785 9516
rect 8749 9485 8786 9514
rect 7988 9476 8023 9477
rect 7965 9471 8023 9476
rect 7965 9451 7968 9471
rect 7988 9457 8023 9471
rect 8043 9457 8052 9477
rect 7988 9449 8052 9457
rect 8014 9448 8052 9449
rect 8015 9447 8052 9448
rect 8118 9481 8154 9482
rect 8226 9481 8262 9482
rect 8118 9473 8262 9481
rect 8118 9453 8126 9473
rect 8146 9453 8234 9473
rect 8254 9453 8262 9473
rect 8118 9447 8262 9453
rect 8328 9477 8366 9485
rect 8434 9481 8470 9482
rect 8328 9457 8337 9477
rect 8357 9457 8366 9477
rect 8328 9448 8366 9457
rect 8385 9474 8470 9481
rect 8385 9454 8392 9474
rect 8413 9473 8470 9474
rect 8413 9454 8442 9473
rect 8385 9453 8442 9454
rect 8462 9453 8470 9473
rect 8328 9447 8365 9448
rect 8385 9447 8470 9453
rect 8536 9477 8574 9485
rect 8647 9481 8683 9482
rect 8536 9457 8545 9477
rect 8565 9457 8574 9477
rect 8536 9448 8574 9457
rect 8598 9473 8683 9481
rect 8598 9453 8655 9473
rect 8675 9453 8683 9473
rect 8536 9447 8573 9448
rect 8598 9447 8683 9453
rect 8749 9477 8787 9485
rect 8749 9457 8758 9477
rect 8778 9457 8787 9477
rect 8749 9448 8787 9457
rect 8827 9462 8899 9672
rect 8969 9706 10169 9736
rect 8969 9705 9413 9706
rect 8969 9703 9137 9705
rect 8827 9448 8910 9462
rect 8749 9447 8786 9448
rect 8172 9426 8208 9447
rect 8598 9426 8629 9447
rect 8827 9426 8844 9448
rect 8005 9422 8105 9426
rect 8005 9418 8067 9422
rect 8005 9392 8012 9418
rect 8038 9396 8067 9418
rect 8093 9396 8105 9422
rect 8038 9392 8105 9396
rect 8005 9389 8105 9392
rect 8173 9389 8208 9426
rect 8270 9423 8629 9426
rect 8270 9418 8492 9423
rect 8270 9394 8283 9418
rect 8307 9399 8492 9418
rect 8516 9399 8629 9423
rect 8307 9394 8629 9399
rect 8270 9390 8629 9394
rect 8696 9418 8844 9426
rect 8696 9398 8707 9418
rect 8727 9415 8844 9418
rect 8897 9415 8910 9448
rect 8727 9398 8910 9415
rect 8696 9391 8910 9398
rect 8696 9390 8737 9391
rect 8827 9390 8910 9391
rect 8172 9364 8208 9389
rect 8020 9337 8057 9338
rect 8116 9337 8153 9338
rect 8172 9337 8179 9364
rect 7920 9328 8058 9337
rect 7920 9308 8029 9328
rect 8049 9308 8058 9328
rect 7920 9301 8058 9308
rect 8116 9334 8179 9337
rect 8200 9337 8208 9364
rect 8227 9337 8264 9338
rect 8200 9334 8264 9337
rect 8116 9328 8264 9334
rect 8116 9308 8125 9328
rect 8145 9308 8235 9328
rect 8255 9308 8264 9328
rect 7920 9299 8016 9301
rect 8116 9298 8264 9308
rect 8323 9328 8360 9338
rect 8435 9337 8472 9338
rect 8416 9335 8472 9337
rect 8323 9308 8331 9328
rect 8351 9308 8360 9328
rect 8172 9297 8208 9298
rect 8020 9166 8057 9167
rect 8323 9166 8360 9308
rect 8385 9328 8472 9335
rect 8385 9325 8443 9328
rect 8385 9305 8390 9325
rect 8411 9308 8443 9325
rect 8463 9308 8472 9328
rect 8411 9305 8472 9308
rect 8385 9298 8472 9305
rect 8531 9328 8568 9338
rect 8531 9308 8539 9328
rect 8559 9308 8568 9328
rect 8385 9297 8416 9298
rect 8531 9229 8568 9308
rect 8598 9337 8629 9390
rect 8835 9357 8849 9390
rect 8902 9357 8910 9390
rect 8835 9351 8910 9357
rect 8835 9346 8905 9351
rect 8648 9337 8685 9338
rect 8598 9328 8685 9337
rect 8598 9308 8656 9328
rect 8676 9308 8685 9328
rect 8598 9298 8685 9308
rect 8744 9328 8781 9338
rect 8969 9333 8996 9703
rect 9036 9473 9100 9485
rect 9376 9481 9413 9705
rect 9884 9686 9948 9688
rect 9880 9674 9948 9686
rect 9880 9641 9891 9674
rect 9931 9641 9948 9674
rect 9880 9631 9948 9641
rect 9641 9570 9752 9585
rect 9641 9568 9683 9570
rect 9641 9548 9648 9568
rect 9667 9548 9683 9568
rect 9641 9540 9683 9548
rect 9711 9568 9752 9570
rect 9711 9548 9725 9568
rect 9744 9548 9752 9568
rect 9711 9540 9752 9548
rect 9641 9534 9752 9540
rect 9584 9512 9833 9534
rect 9584 9481 9621 9512
rect 9797 9510 9833 9512
rect 9797 9481 9834 9510
rect 9036 9472 9071 9473
rect 9013 9467 9071 9472
rect 9013 9447 9016 9467
rect 9036 9453 9071 9467
rect 9091 9453 9100 9473
rect 9036 9445 9100 9453
rect 9062 9444 9100 9445
rect 9063 9443 9100 9444
rect 9166 9477 9202 9478
rect 9274 9477 9310 9478
rect 9166 9469 9310 9477
rect 9166 9449 9174 9469
rect 9194 9449 9282 9469
rect 9302 9449 9310 9469
rect 9166 9443 9310 9449
rect 9376 9473 9414 9481
rect 9482 9477 9518 9478
rect 9376 9453 9385 9473
rect 9405 9453 9414 9473
rect 9376 9444 9414 9453
rect 9433 9470 9518 9477
rect 9433 9450 9440 9470
rect 9461 9469 9518 9470
rect 9461 9450 9490 9469
rect 9433 9449 9490 9450
rect 9510 9449 9518 9469
rect 9376 9443 9413 9444
rect 9433 9443 9518 9449
rect 9584 9473 9622 9481
rect 9695 9477 9731 9478
rect 9584 9453 9593 9473
rect 9613 9453 9622 9473
rect 9584 9444 9622 9453
rect 9646 9469 9731 9477
rect 9646 9449 9703 9469
rect 9723 9449 9731 9469
rect 9584 9443 9621 9444
rect 9646 9443 9731 9449
rect 9797 9473 9835 9481
rect 9797 9453 9806 9473
rect 9826 9453 9835 9473
rect 9797 9444 9835 9453
rect 9884 9447 9948 9631
rect 10104 9505 10169 9706
rect 10104 9487 10126 9505
rect 10144 9487 10169 9505
rect 10104 9468 10169 9487
rect 9797 9443 9834 9444
rect 9220 9422 9256 9443
rect 9646 9422 9677 9443
rect 9884 9438 9892 9447
rect 9881 9422 9892 9438
rect 9053 9418 9153 9422
rect 9053 9414 9115 9418
rect 9053 9388 9060 9414
rect 9086 9392 9115 9414
rect 9141 9392 9153 9418
rect 9086 9388 9153 9392
rect 9053 9385 9153 9388
rect 9221 9385 9256 9422
rect 9318 9419 9677 9422
rect 9318 9414 9540 9419
rect 9318 9390 9331 9414
rect 9355 9395 9540 9414
rect 9564 9395 9677 9419
rect 9355 9390 9677 9395
rect 9318 9386 9677 9390
rect 9744 9414 9892 9422
rect 9744 9394 9755 9414
rect 9775 9405 9892 9414
rect 9941 9438 9948 9447
rect 9941 9405 9949 9438
rect 9775 9394 9949 9405
rect 9744 9387 9949 9394
rect 9744 9386 9785 9387
rect 9220 9360 9256 9385
rect 9068 9333 9105 9334
rect 9164 9333 9201 9334
rect 9220 9333 9227 9360
rect 8744 9308 8752 9328
rect 8772 9308 8781 9328
rect 8598 9297 8629 9298
rect 8593 9229 8703 9242
rect 8744 9229 8781 9308
rect 8968 9324 9106 9333
rect 8968 9304 9077 9324
rect 9097 9304 9106 9324
rect 8968 9297 9106 9304
rect 9164 9330 9227 9333
rect 9248 9333 9256 9360
rect 9275 9333 9312 9334
rect 9248 9330 9312 9333
rect 9164 9324 9312 9330
rect 9164 9304 9173 9324
rect 9193 9304 9283 9324
rect 9303 9304 9312 9324
rect 8968 9295 9064 9297
rect 9164 9294 9312 9304
rect 9371 9324 9408 9334
rect 9483 9333 9520 9334
rect 9464 9331 9520 9333
rect 9371 9304 9379 9324
rect 9399 9304 9408 9324
rect 9220 9293 9256 9294
rect 8531 9227 8781 9229
rect 8531 9224 8632 9227
rect 8531 9205 8596 9224
rect 8593 9197 8596 9205
rect 8625 9197 8632 9224
rect 8660 9200 8670 9227
rect 8699 9205 8781 9227
rect 8699 9200 8703 9205
rect 8660 9197 8703 9200
rect 8593 9183 8703 9197
rect 8019 9165 8360 9166
rect 7944 9160 8360 9165
rect 9068 9162 9105 9163
rect 9371 9162 9408 9304
rect 9433 9324 9520 9331
rect 9433 9321 9491 9324
rect 9433 9301 9438 9321
rect 9459 9304 9491 9321
rect 9511 9304 9520 9324
rect 9459 9301 9520 9304
rect 9433 9294 9520 9301
rect 9579 9324 9616 9334
rect 9579 9304 9587 9324
rect 9607 9304 9616 9324
rect 9433 9293 9464 9294
rect 9579 9225 9616 9304
rect 9646 9333 9677 9386
rect 9881 9384 9949 9387
rect 9881 9342 9893 9384
rect 9942 9342 9949 9384
rect 9696 9333 9733 9334
rect 9646 9324 9733 9333
rect 9646 9304 9704 9324
rect 9724 9304 9733 9324
rect 9646 9294 9733 9304
rect 9792 9324 9829 9334
rect 9881 9329 9949 9342
rect 10104 9406 10169 9423
rect 10104 9388 10128 9406
rect 10146 9388 10169 9406
rect 9792 9304 9800 9324
rect 9820 9304 9829 9324
rect 9646 9293 9677 9294
rect 9641 9225 9751 9238
rect 9792 9225 9829 9304
rect 10104 9249 10169 9388
rect 10104 9243 10126 9249
rect 9579 9223 9829 9225
rect 9579 9220 9680 9223
rect 9579 9201 9644 9220
rect 9641 9193 9644 9201
rect 9673 9193 9680 9220
rect 9708 9196 9718 9223
rect 9747 9201 9829 9223
rect 9858 9231 10126 9243
rect 10144 9231 10169 9249
rect 9858 9208 10169 9231
rect 9858 9207 9913 9208
rect 9747 9196 9751 9201
rect 9708 9193 9751 9196
rect 9641 9179 9751 9193
rect 9067 9161 9408 9162
rect 7944 9140 7947 9160
rect 7967 9140 8360 9160
rect 8992 9160 9408 9161
rect 9858 9160 9901 9207
rect 8992 9156 9901 9160
rect 8311 9107 8356 9140
rect 8992 9136 8995 9156
rect 9015 9136 9901 9156
rect 9369 9131 9901 9136
rect 10109 9150 10168 9172
rect 10109 9132 10128 9150
rect 10146 9132 10168 9150
rect 9157 9107 9256 9109
rect 8311 9097 9256 9107
rect 8311 9071 9179 9097
rect 8312 9070 9179 9071
rect 9157 9059 9179 9070
rect 9204 9062 9223 9097
rect 9248 9062 9256 9097
rect 9204 9059 9256 9062
rect 9157 9051 9256 9059
rect 9183 9050 9255 9051
rect 10109 9002 10168 9132
rect 8831 8972 8907 8996
rect 8831 8906 8843 8972
rect 8897 8906 8907 8972
rect 9375 8927 9416 8929
rect 9647 8927 9751 8929
rect 10109 8927 10170 9002
rect 7721 8856 7793 8906
rect 6432 8764 6876 8790
rect 6432 8762 6600 8764
rect 6432 8495 6459 8762
rect 6729 8760 6758 8764
rect 6499 8635 6563 8647
rect 6839 8643 6876 8764
rect 7104 8732 7215 8747
rect 7104 8730 7146 8732
rect 7104 8710 7111 8730
rect 7130 8710 7146 8730
rect 7104 8702 7146 8710
rect 7174 8730 7215 8732
rect 7174 8710 7188 8730
rect 7207 8710 7215 8730
rect 7174 8702 7215 8710
rect 7104 8696 7215 8702
rect 7047 8674 7296 8696
rect 7047 8643 7084 8674
rect 7260 8672 7296 8674
rect 7260 8643 7297 8672
rect 6499 8634 6534 8635
rect 6476 8629 6534 8634
rect 6476 8609 6479 8629
rect 6499 8615 6534 8629
rect 6554 8615 6563 8635
rect 6499 8607 6563 8615
rect 6525 8606 6563 8607
rect 6526 8605 6563 8606
rect 6629 8639 6665 8640
rect 6737 8639 6773 8640
rect 6629 8631 6773 8639
rect 6629 8611 6637 8631
rect 6657 8611 6745 8631
rect 6765 8611 6773 8631
rect 6629 8605 6773 8611
rect 6839 8635 6877 8643
rect 6945 8639 6981 8640
rect 6839 8615 6848 8635
rect 6868 8615 6877 8635
rect 6839 8606 6877 8615
rect 6896 8632 6981 8639
rect 6896 8612 6903 8632
rect 6924 8631 6981 8632
rect 6924 8612 6953 8631
rect 6896 8611 6953 8612
rect 6973 8611 6981 8631
rect 6839 8605 6876 8606
rect 6896 8605 6981 8611
rect 7047 8635 7085 8643
rect 7158 8639 7194 8640
rect 7047 8615 7056 8635
rect 7076 8615 7085 8635
rect 7047 8606 7085 8615
rect 7109 8631 7194 8639
rect 7109 8611 7166 8631
rect 7186 8611 7194 8631
rect 7047 8605 7084 8606
rect 7109 8605 7194 8611
rect 7260 8635 7298 8643
rect 7260 8615 7269 8635
rect 7289 8615 7298 8635
rect 7260 8606 7298 8615
rect 7260 8605 7297 8606
rect 6683 8584 6719 8605
rect 7109 8584 7140 8605
rect 7290 8584 7624 8588
rect 6516 8580 6616 8584
rect 6516 8576 6578 8580
rect 6516 8550 6523 8576
rect 6549 8554 6578 8576
rect 6604 8554 6616 8580
rect 6549 8550 6616 8554
rect 6516 8547 6616 8550
rect 6684 8547 6719 8584
rect 6781 8581 7140 8584
rect 6781 8576 7003 8581
rect 6781 8552 6794 8576
rect 6818 8557 7003 8576
rect 7027 8557 7140 8581
rect 6818 8552 7140 8557
rect 6781 8548 7140 8552
rect 7207 8576 7624 8584
rect 7207 8556 7218 8576
rect 7238 8556 7624 8576
rect 7207 8549 7624 8556
rect 7207 8548 7248 8549
rect 7290 8548 7624 8549
rect 6683 8522 6719 8547
rect 6531 8495 6568 8496
rect 6627 8495 6664 8496
rect 6683 8495 6690 8522
rect 6431 8486 6569 8495
rect 6431 8466 6540 8486
rect 6560 8466 6569 8486
rect 6431 8459 6569 8466
rect 6627 8492 6690 8495
rect 6711 8495 6719 8522
rect 6738 8495 6775 8496
rect 6711 8492 6775 8495
rect 6627 8486 6775 8492
rect 6627 8466 6636 8486
rect 6656 8466 6746 8486
rect 6766 8466 6775 8486
rect 6431 8457 6527 8459
rect 6627 8456 6775 8466
rect 6834 8486 6871 8496
rect 6946 8495 6983 8496
rect 6927 8493 6983 8495
rect 6834 8466 6842 8486
rect 6862 8466 6871 8486
rect 6683 8455 6719 8456
rect 6531 8324 6568 8325
rect 6834 8324 6871 8466
rect 6896 8486 6983 8493
rect 6896 8483 6954 8486
rect 6896 8463 6901 8483
rect 6922 8466 6954 8483
rect 6974 8466 6983 8486
rect 6922 8463 6983 8466
rect 6896 8456 6983 8463
rect 7042 8486 7079 8496
rect 7042 8466 7050 8486
rect 7070 8466 7079 8486
rect 6896 8455 6927 8456
rect 7042 8387 7079 8466
rect 7109 8495 7140 8548
rect 7159 8495 7196 8496
rect 7109 8486 7196 8495
rect 7109 8466 7167 8486
rect 7187 8466 7196 8486
rect 7109 8456 7196 8466
rect 7255 8486 7292 8496
rect 7255 8466 7263 8486
rect 7283 8466 7292 8486
rect 7109 8455 7140 8456
rect 7104 8387 7214 8400
rect 7255 8387 7292 8466
rect 7042 8385 7292 8387
rect 7042 8382 7143 8385
rect 7042 8363 7107 8382
rect 7104 8355 7107 8363
rect 7136 8355 7143 8382
rect 7171 8358 7181 8385
rect 7210 8363 7292 8385
rect 7210 8358 7214 8363
rect 7171 8355 7214 8358
rect 7104 8341 7214 8355
rect 6530 8323 6871 8324
rect 6455 8318 6871 8323
rect 6455 8298 6458 8318
rect 6478 8298 6871 8318
rect 6764 7933 6795 8298
rect 6682 7904 6795 7933
rect 6683 7604 6719 7904
rect 7543 7799 7624 8548
rect 7723 7947 7793 8856
rect 8831 8886 8907 8906
rect 8831 8849 8848 8886
rect 8892 8849 8907 8886
rect 8968 8892 10170 8927
rect 8968 8878 8996 8892
rect 8831 8833 8907 8849
rect 8836 8677 8906 8833
rect 8970 8747 8996 8878
rect 9375 8889 10170 8892
rect 8828 8626 8908 8677
rect 8828 8600 8844 8626
rect 8884 8600 8908 8626
rect 8828 8581 8908 8600
rect 8828 8555 8847 8581
rect 8887 8555 8908 8581
rect 8828 8528 8908 8555
rect 8828 8502 8851 8528
rect 8891 8502 8908 8528
rect 8828 8491 8908 8502
rect 8970 8492 8997 8747
rect 9375 8739 9416 8889
rect 10109 8877 10170 8889
rect 9842 8827 9963 8845
rect 9842 8825 9913 8827
rect 9842 8784 9857 8825
rect 9894 8786 9913 8825
rect 9950 8786 9963 8827
rect 9894 8784 9963 8786
rect 9842 8774 9963 8784
rect 9647 8744 9751 8753
rect 9037 8632 9101 8644
rect 9377 8640 9414 8739
rect 9642 8729 9753 8744
rect 9642 8727 9684 8729
rect 9642 8707 9649 8727
rect 9668 8707 9684 8727
rect 9642 8699 9684 8707
rect 9712 8727 9753 8729
rect 9712 8707 9726 8727
rect 9745 8707 9753 8727
rect 9712 8699 9753 8707
rect 9642 8693 9753 8699
rect 9585 8671 9834 8693
rect 9585 8640 9622 8671
rect 9798 8669 9834 8671
rect 9798 8640 9835 8669
rect 9037 8631 9072 8632
rect 9014 8626 9072 8631
rect 9014 8606 9017 8626
rect 9037 8612 9072 8626
rect 9092 8612 9101 8632
rect 9037 8604 9101 8612
rect 9063 8603 9101 8604
rect 9064 8602 9101 8603
rect 9167 8636 9203 8637
rect 9275 8636 9311 8637
rect 9167 8628 9311 8636
rect 9167 8608 9175 8628
rect 9195 8608 9283 8628
rect 9303 8608 9311 8628
rect 9167 8602 9311 8608
rect 9377 8632 9415 8640
rect 9483 8636 9519 8637
rect 9377 8612 9386 8632
rect 9406 8612 9415 8632
rect 9377 8603 9415 8612
rect 9434 8629 9519 8636
rect 9434 8609 9441 8629
rect 9462 8628 9519 8629
rect 9462 8609 9491 8628
rect 9434 8608 9491 8609
rect 9511 8608 9519 8628
rect 9377 8602 9414 8603
rect 9434 8602 9519 8608
rect 9585 8632 9623 8640
rect 9696 8636 9732 8637
rect 9585 8612 9594 8632
rect 9614 8612 9623 8632
rect 9585 8603 9623 8612
rect 9647 8628 9732 8636
rect 9647 8608 9704 8628
rect 9724 8608 9732 8628
rect 9585 8602 9622 8603
rect 9647 8602 9732 8608
rect 9798 8632 9836 8640
rect 9798 8612 9807 8632
rect 9827 8612 9836 8632
rect 9891 8622 9956 8774
rect 10109 8748 10164 8877
rect 9798 8603 9836 8612
rect 9889 8615 9956 8622
rect 9798 8602 9835 8603
rect 9221 8581 9257 8602
rect 9647 8581 9678 8602
rect 9889 8594 9906 8615
rect 9942 8594 9956 8615
rect 10108 8635 10164 8748
rect 10108 8617 10127 8635
rect 10145 8617 10164 8635
rect 10108 8597 10164 8617
rect 9889 8581 9956 8594
rect 9054 8577 9154 8581
rect 9054 8573 9116 8577
rect 9054 8547 9061 8573
rect 9087 8551 9116 8573
rect 9142 8551 9154 8577
rect 9087 8547 9154 8551
rect 9054 8544 9154 8547
rect 9222 8544 9257 8581
rect 9319 8578 9678 8581
rect 9319 8573 9541 8578
rect 9319 8549 9332 8573
rect 9356 8554 9541 8573
rect 9565 8554 9678 8578
rect 9356 8549 9678 8554
rect 9319 8545 9678 8549
rect 9745 8575 9956 8581
rect 9745 8573 9906 8575
rect 9745 8553 9756 8573
rect 9776 8553 9906 8573
rect 9745 8546 9906 8553
rect 9745 8545 9786 8546
rect 9221 8519 9257 8544
rect 9069 8492 9106 8493
rect 9165 8492 9202 8493
rect 9221 8492 9228 8519
rect 8969 8483 9107 8492
rect 8969 8463 9078 8483
rect 9098 8463 9107 8483
rect 8969 8456 9107 8463
rect 9165 8489 9228 8492
rect 9249 8492 9257 8519
rect 9276 8492 9313 8493
rect 9249 8489 9313 8492
rect 9165 8483 9313 8489
rect 9165 8463 9174 8483
rect 9194 8463 9284 8483
rect 9304 8463 9313 8483
rect 8969 8454 9065 8456
rect 9165 8453 9313 8463
rect 9372 8483 9409 8493
rect 9484 8492 9521 8493
rect 9465 8490 9521 8492
rect 9372 8463 9380 8483
rect 9400 8463 9409 8483
rect 9221 8452 9257 8453
rect 9069 8321 9106 8322
rect 9372 8321 9409 8463
rect 9434 8483 9521 8490
rect 9434 8480 9492 8483
rect 9434 8460 9439 8480
rect 9460 8463 9492 8480
rect 9512 8463 9521 8483
rect 9460 8460 9521 8463
rect 9434 8453 9521 8460
rect 9580 8483 9617 8493
rect 9580 8463 9588 8483
rect 9608 8463 9617 8483
rect 9434 8452 9465 8453
rect 9580 8384 9617 8463
rect 9647 8492 9678 8545
rect 9891 8538 9906 8546
rect 9946 8538 9956 8575
rect 9891 8529 9956 8538
rect 10104 8536 10169 8557
rect 10104 8518 10129 8536
rect 10147 8518 10169 8536
rect 9697 8492 9734 8493
rect 9647 8483 9734 8492
rect 9647 8463 9705 8483
rect 9725 8463 9734 8483
rect 9647 8453 9734 8463
rect 9793 8483 9830 8493
rect 9793 8463 9801 8483
rect 9821 8463 9830 8483
rect 9647 8452 9678 8453
rect 9642 8384 9752 8397
rect 9793 8384 9830 8463
rect 10104 8442 10169 8518
rect 9580 8382 9830 8384
rect 9580 8379 9681 8382
rect 9580 8360 9645 8379
rect 9642 8352 9645 8360
rect 9674 8352 9681 8379
rect 9709 8355 9719 8382
rect 9748 8360 9830 8382
rect 9853 8407 10170 8442
rect 9748 8355 9752 8360
rect 9709 8352 9752 8355
rect 9642 8338 9752 8352
rect 9068 8320 9409 8321
rect 8993 8318 9409 8320
rect 9853 8318 9893 8407
rect 10104 8380 10169 8407
rect 10104 8362 10127 8380
rect 10145 8362 10169 8380
rect 10104 8342 10169 8362
rect 8990 8315 9893 8318
rect 8990 8295 8996 8315
rect 9016 8295 9893 8315
rect 8990 8291 9893 8295
rect 9853 8288 9893 8291
rect 10105 8281 10170 8302
rect 8323 8273 8984 8274
rect 8323 8266 9257 8273
rect 8323 8265 9229 8266
rect 8323 8245 9174 8265
rect 9206 8246 9229 8265
rect 9254 8246 9257 8266
rect 9206 8245 9257 8246
rect 8323 8238 9257 8245
rect 7922 8196 8090 8197
rect 8325 8196 8364 8238
rect 9153 8236 9257 8238
rect 9222 8234 9257 8236
rect 10105 8263 10129 8281
rect 10147 8263 10170 8281
rect 10105 8216 10170 8263
rect 7922 8170 8366 8196
rect 7922 8168 8090 8170
rect 6683 7581 6687 7604
rect 6711 7581 6719 7604
rect 6883 7582 6982 7586
rect 6683 7560 6719 7581
rect 6683 7537 6687 7560
rect 6711 7537 6719 7560
rect 6683 7533 6719 7537
rect 6879 7576 6982 7582
rect 6879 7538 6905 7576
rect 6930 7541 6949 7576
rect 6974 7541 6982 7576
rect 6930 7538 6982 7541
rect 6879 7530 6982 7538
rect 6879 7529 6981 7530
rect 6475 7451 6643 7452
rect 6879 7451 6926 7529
rect 6475 7425 6926 7451
rect 6475 7423 6643 7425
rect 6475 7050 6502 7423
rect 6672 7375 6758 7384
rect 6672 7357 6691 7375
rect 6743 7357 6758 7375
rect 6672 7353 6758 7357
rect 6542 7190 6606 7202
rect 6542 7189 6577 7190
rect 6519 7184 6577 7189
rect 6519 7164 6522 7184
rect 6542 7170 6577 7184
rect 6597 7170 6606 7190
rect 6542 7162 6606 7170
rect 6568 7161 6606 7162
rect 6569 7160 6606 7161
rect 6672 7194 6708 7195
rect 6728 7194 6758 7353
rect 6879 7313 6926 7425
rect 6882 7198 6919 7313
rect 7147 7287 7258 7302
rect 7147 7285 7189 7287
rect 7147 7265 7154 7285
rect 7173 7265 7189 7285
rect 7147 7257 7189 7265
rect 7217 7285 7258 7287
rect 7217 7265 7231 7285
rect 7250 7265 7258 7285
rect 7217 7257 7258 7265
rect 7147 7251 7258 7257
rect 7090 7229 7339 7251
rect 7090 7198 7127 7229
rect 7303 7227 7339 7229
rect 7303 7198 7340 7227
rect 7544 7214 7623 7799
rect 7720 7347 7799 7947
rect 7922 7817 7949 8168
rect 8325 8164 8366 8170
rect 7989 7957 8053 7969
rect 8329 7965 8366 8164
rect 8828 8191 8900 8208
rect 8828 8152 8836 8191
rect 8881 8152 8900 8191
rect 8594 8054 8705 8069
rect 8594 8052 8636 8054
rect 8594 8032 8601 8052
rect 8620 8032 8636 8052
rect 8594 8024 8636 8032
rect 8664 8052 8705 8054
rect 8664 8032 8678 8052
rect 8697 8032 8705 8052
rect 8664 8024 8705 8032
rect 8594 8018 8705 8024
rect 8537 7996 8786 8018
rect 8537 7965 8574 7996
rect 8750 7994 8786 7996
rect 8750 7965 8787 7994
rect 7989 7956 8024 7957
rect 7966 7951 8024 7956
rect 7966 7931 7969 7951
rect 7989 7937 8024 7951
rect 8044 7937 8053 7957
rect 7989 7929 8053 7937
rect 8015 7928 8053 7929
rect 8016 7927 8053 7928
rect 8119 7961 8155 7962
rect 8227 7961 8263 7962
rect 8119 7953 8263 7961
rect 8119 7933 8127 7953
rect 8147 7933 8235 7953
rect 8255 7933 8263 7953
rect 8119 7927 8263 7933
rect 8329 7957 8367 7965
rect 8435 7961 8471 7962
rect 8329 7937 8338 7957
rect 8358 7937 8367 7957
rect 8329 7928 8367 7937
rect 8386 7954 8471 7961
rect 8386 7934 8393 7954
rect 8414 7953 8471 7954
rect 8414 7934 8443 7953
rect 8386 7933 8443 7934
rect 8463 7933 8471 7953
rect 8329 7927 8366 7928
rect 8386 7927 8471 7933
rect 8537 7957 8575 7965
rect 8648 7961 8684 7962
rect 8537 7937 8546 7957
rect 8566 7937 8575 7957
rect 8537 7928 8575 7937
rect 8599 7953 8684 7961
rect 8599 7933 8656 7953
rect 8676 7933 8684 7953
rect 8537 7927 8574 7928
rect 8599 7927 8684 7933
rect 8750 7957 8788 7965
rect 8750 7937 8759 7957
rect 8779 7937 8788 7957
rect 8750 7928 8788 7937
rect 8828 7942 8900 8152
rect 8970 8186 10170 8216
rect 8970 8185 9414 8186
rect 8970 8183 9138 8185
rect 8828 7928 8911 7942
rect 8750 7927 8787 7928
rect 8173 7906 8209 7927
rect 8599 7906 8630 7927
rect 8828 7906 8845 7928
rect 8006 7902 8106 7906
rect 8006 7898 8068 7902
rect 8006 7872 8013 7898
rect 8039 7876 8068 7898
rect 8094 7876 8106 7902
rect 8039 7872 8106 7876
rect 8006 7869 8106 7872
rect 8174 7869 8209 7906
rect 8271 7903 8630 7906
rect 8271 7898 8493 7903
rect 8271 7874 8284 7898
rect 8308 7879 8493 7898
rect 8517 7879 8630 7903
rect 8308 7874 8630 7879
rect 8271 7870 8630 7874
rect 8697 7898 8845 7906
rect 8697 7878 8708 7898
rect 8728 7895 8845 7898
rect 8898 7895 8911 7928
rect 8728 7878 8911 7895
rect 8697 7871 8911 7878
rect 8697 7870 8738 7871
rect 8828 7870 8911 7871
rect 8173 7844 8209 7869
rect 8021 7817 8058 7818
rect 8117 7817 8154 7818
rect 8173 7817 8180 7844
rect 7921 7808 8059 7817
rect 7921 7788 8030 7808
rect 8050 7788 8059 7808
rect 7921 7781 8059 7788
rect 8117 7814 8180 7817
rect 8201 7817 8209 7844
rect 8228 7817 8265 7818
rect 8201 7814 8265 7817
rect 8117 7808 8265 7814
rect 8117 7788 8126 7808
rect 8146 7788 8236 7808
rect 8256 7788 8265 7808
rect 7921 7779 8017 7781
rect 8117 7778 8265 7788
rect 8324 7808 8361 7818
rect 8436 7817 8473 7818
rect 8417 7815 8473 7817
rect 8324 7788 8332 7808
rect 8352 7788 8361 7808
rect 8173 7777 8209 7778
rect 8021 7646 8058 7647
rect 8324 7646 8361 7788
rect 8386 7808 8473 7815
rect 8386 7805 8444 7808
rect 8386 7785 8391 7805
rect 8412 7788 8444 7805
rect 8464 7788 8473 7808
rect 8412 7785 8473 7788
rect 8386 7778 8473 7785
rect 8532 7808 8569 7818
rect 8532 7788 8540 7808
rect 8560 7788 8569 7808
rect 8386 7777 8417 7778
rect 8532 7709 8569 7788
rect 8599 7817 8630 7870
rect 8836 7837 8850 7870
rect 8903 7837 8911 7870
rect 8836 7831 8911 7837
rect 8836 7826 8906 7831
rect 8649 7817 8686 7818
rect 8599 7808 8686 7817
rect 8599 7788 8657 7808
rect 8677 7788 8686 7808
rect 8599 7778 8686 7788
rect 8745 7808 8782 7818
rect 8970 7813 8997 8183
rect 9037 7953 9101 7965
rect 9377 7961 9414 8185
rect 9885 8166 9949 8168
rect 9881 8154 9949 8166
rect 9881 8121 9892 8154
rect 9932 8121 9949 8154
rect 9881 8111 9949 8121
rect 9642 8050 9753 8065
rect 9642 8048 9684 8050
rect 9642 8028 9649 8048
rect 9668 8028 9684 8048
rect 9642 8020 9684 8028
rect 9712 8048 9753 8050
rect 9712 8028 9726 8048
rect 9745 8028 9753 8048
rect 9712 8020 9753 8028
rect 9642 8014 9753 8020
rect 9585 7992 9834 8014
rect 9585 7961 9622 7992
rect 9798 7990 9834 7992
rect 9798 7961 9835 7990
rect 9037 7952 9072 7953
rect 9014 7947 9072 7952
rect 9014 7927 9017 7947
rect 9037 7933 9072 7947
rect 9092 7933 9101 7953
rect 9037 7925 9101 7933
rect 9063 7924 9101 7925
rect 9064 7923 9101 7924
rect 9167 7957 9203 7958
rect 9275 7957 9311 7958
rect 9167 7949 9311 7957
rect 9167 7929 9175 7949
rect 9195 7929 9283 7949
rect 9303 7929 9311 7949
rect 9167 7923 9311 7929
rect 9377 7953 9415 7961
rect 9483 7957 9519 7958
rect 9377 7933 9386 7953
rect 9406 7933 9415 7953
rect 9377 7924 9415 7933
rect 9434 7950 9519 7957
rect 9434 7930 9441 7950
rect 9462 7949 9519 7950
rect 9462 7930 9491 7949
rect 9434 7929 9491 7930
rect 9511 7929 9519 7949
rect 9377 7923 9414 7924
rect 9434 7923 9519 7929
rect 9585 7953 9623 7961
rect 9696 7957 9732 7958
rect 9585 7933 9594 7953
rect 9614 7933 9623 7953
rect 9585 7924 9623 7933
rect 9647 7949 9732 7957
rect 9647 7929 9704 7949
rect 9724 7929 9732 7949
rect 9585 7923 9622 7924
rect 9647 7923 9732 7929
rect 9798 7953 9836 7961
rect 9798 7933 9807 7953
rect 9827 7933 9836 7953
rect 9798 7924 9836 7933
rect 9885 7927 9949 8111
rect 10105 7985 10170 8186
rect 10105 7967 10127 7985
rect 10145 7967 10170 7985
rect 10105 7948 10170 7967
rect 9798 7923 9835 7924
rect 9221 7902 9257 7923
rect 9647 7902 9678 7923
rect 9885 7918 9893 7927
rect 9882 7902 9893 7918
rect 9054 7898 9154 7902
rect 9054 7894 9116 7898
rect 9054 7868 9061 7894
rect 9087 7872 9116 7894
rect 9142 7872 9154 7898
rect 9087 7868 9154 7872
rect 9054 7865 9154 7868
rect 9222 7865 9257 7902
rect 9319 7899 9678 7902
rect 9319 7894 9541 7899
rect 9319 7870 9332 7894
rect 9356 7875 9541 7894
rect 9565 7875 9678 7899
rect 9356 7870 9678 7875
rect 9319 7866 9678 7870
rect 9745 7894 9893 7902
rect 9745 7874 9756 7894
rect 9776 7885 9893 7894
rect 9942 7918 9949 7927
rect 9942 7885 9950 7918
rect 9776 7874 9950 7885
rect 9745 7867 9950 7874
rect 9745 7866 9786 7867
rect 9221 7840 9257 7865
rect 9069 7813 9106 7814
rect 9165 7813 9202 7814
rect 9221 7813 9228 7840
rect 8745 7788 8753 7808
rect 8773 7788 8782 7808
rect 8599 7777 8630 7778
rect 8594 7709 8704 7722
rect 8745 7709 8782 7788
rect 8969 7804 9107 7813
rect 8969 7784 9078 7804
rect 9098 7784 9107 7804
rect 8969 7777 9107 7784
rect 9165 7810 9228 7813
rect 9249 7813 9257 7840
rect 9276 7813 9313 7814
rect 9249 7810 9313 7813
rect 9165 7804 9313 7810
rect 9165 7784 9174 7804
rect 9194 7784 9284 7804
rect 9304 7784 9313 7804
rect 8969 7775 9065 7777
rect 9165 7774 9313 7784
rect 9372 7804 9409 7814
rect 9484 7813 9521 7814
rect 9465 7811 9521 7813
rect 9372 7784 9380 7804
rect 9400 7784 9409 7804
rect 9221 7773 9257 7774
rect 8532 7707 8782 7709
rect 8532 7704 8633 7707
rect 8532 7685 8597 7704
rect 8594 7677 8597 7685
rect 8626 7677 8633 7704
rect 8661 7680 8671 7707
rect 8700 7685 8782 7707
rect 8700 7680 8704 7685
rect 8661 7677 8704 7680
rect 8594 7663 8704 7677
rect 8020 7645 8361 7646
rect 7945 7640 8361 7645
rect 9069 7642 9106 7643
rect 9372 7642 9409 7784
rect 9434 7804 9521 7811
rect 9434 7801 9492 7804
rect 9434 7781 9439 7801
rect 9460 7784 9492 7801
rect 9512 7784 9521 7804
rect 9460 7781 9521 7784
rect 9434 7774 9521 7781
rect 9580 7804 9617 7814
rect 9580 7784 9588 7804
rect 9608 7784 9617 7804
rect 9434 7773 9465 7774
rect 9580 7705 9617 7784
rect 9647 7813 9678 7866
rect 9882 7864 9950 7867
rect 9882 7822 9894 7864
rect 9943 7822 9950 7864
rect 9697 7813 9734 7814
rect 9647 7804 9734 7813
rect 9647 7784 9705 7804
rect 9725 7784 9734 7804
rect 9647 7774 9734 7784
rect 9793 7804 9830 7814
rect 9882 7809 9950 7822
rect 10105 7886 10170 7903
rect 10105 7868 10129 7886
rect 10147 7868 10170 7886
rect 9793 7784 9801 7804
rect 9821 7784 9830 7804
rect 9647 7773 9678 7774
rect 9642 7705 9752 7718
rect 9793 7705 9830 7784
rect 10105 7729 10170 7868
rect 10105 7723 10127 7729
rect 9580 7703 9830 7705
rect 9580 7700 9681 7703
rect 9580 7681 9645 7700
rect 9642 7673 9645 7681
rect 9674 7673 9681 7700
rect 9709 7676 9719 7703
rect 9748 7681 9830 7703
rect 9859 7711 10127 7723
rect 10145 7711 10170 7729
rect 9859 7688 10170 7711
rect 9859 7687 9914 7688
rect 9748 7676 9752 7681
rect 9709 7673 9752 7676
rect 9642 7659 9752 7673
rect 9068 7641 9409 7642
rect 7945 7620 7948 7640
rect 7968 7620 8361 7640
rect 8993 7640 9409 7641
rect 9859 7640 9902 7687
rect 8993 7636 9902 7640
rect 8312 7587 8357 7620
rect 8993 7616 8996 7636
rect 9016 7616 9902 7636
rect 9370 7611 9902 7616
rect 10110 7630 10169 7652
rect 10110 7612 10129 7630
rect 10147 7612 10169 7630
rect 9158 7587 9257 7589
rect 8312 7577 9257 7587
rect 8312 7551 9180 7577
rect 8313 7550 9180 7551
rect 9158 7539 9180 7550
rect 9205 7542 9224 7577
rect 9249 7542 9257 7577
rect 9205 7539 9257 7542
rect 10110 7541 10169 7612
rect 9158 7531 9257 7539
rect 9184 7530 9256 7531
rect 8838 7504 8905 7523
rect 8838 7483 8855 7504
rect 7719 7305 7799 7347
rect 8836 7438 8855 7483
rect 8885 7483 8905 7504
rect 8885 7438 8906 7483
rect 9375 7480 9416 7482
rect 9647 7480 9751 7482
rect 10107 7480 10171 7541
rect 6780 7194 6816 7195
rect 6672 7186 6816 7194
rect 6672 7166 6680 7186
rect 6700 7166 6788 7186
rect 6808 7166 6816 7186
rect 6672 7160 6816 7166
rect 6882 7190 6920 7198
rect 6988 7194 7024 7195
rect 6882 7170 6891 7190
rect 6911 7170 6920 7190
rect 6882 7161 6920 7170
rect 6939 7187 7024 7194
rect 6939 7167 6946 7187
rect 6967 7186 7024 7187
rect 6967 7167 6996 7186
rect 6939 7166 6996 7167
rect 7016 7166 7024 7186
rect 6882 7160 6919 7161
rect 6939 7160 7024 7166
rect 7090 7190 7128 7198
rect 7201 7194 7237 7195
rect 7090 7170 7099 7190
rect 7119 7170 7128 7190
rect 7090 7161 7128 7170
rect 7152 7186 7237 7194
rect 7152 7166 7209 7186
rect 7229 7166 7237 7186
rect 7090 7160 7127 7161
rect 7152 7160 7237 7166
rect 7303 7190 7341 7198
rect 7303 7170 7312 7190
rect 7332 7170 7341 7190
rect 7303 7161 7341 7170
rect 7541 7178 7627 7214
rect 7303 7160 7340 7161
rect 6726 7139 6762 7160
rect 7152 7139 7183 7160
rect 7379 7139 7425 7143
rect 6559 7135 6659 7139
rect 6559 7131 6621 7135
rect 6559 7105 6566 7131
rect 6592 7109 6621 7131
rect 6647 7109 6659 7135
rect 6592 7105 6659 7109
rect 6559 7102 6659 7105
rect 6727 7102 6762 7139
rect 6824 7136 7183 7139
rect 6824 7131 7046 7136
rect 6824 7107 6837 7131
rect 6861 7112 7046 7131
rect 7070 7112 7183 7136
rect 6861 7107 7183 7112
rect 6824 7103 7183 7107
rect 7250 7131 7425 7139
rect 7250 7111 7261 7131
rect 7281 7111 7425 7131
rect 7541 7137 7558 7178
rect 7612 7137 7627 7178
rect 7541 7118 7627 7137
rect 7250 7104 7425 7111
rect 7250 7103 7291 7104
rect 6726 7077 6762 7102
rect 6574 7050 6611 7051
rect 6670 7050 6707 7051
rect 6726 7050 6733 7077
rect 6474 7041 6612 7050
rect 6474 7021 6583 7041
rect 6603 7021 6612 7041
rect 6474 7014 6612 7021
rect 6670 7047 6733 7050
rect 6754 7050 6762 7077
rect 6781 7050 6818 7051
rect 6754 7047 6818 7050
rect 6670 7041 6818 7047
rect 6670 7021 6679 7041
rect 6699 7021 6789 7041
rect 6809 7021 6818 7041
rect 6474 7012 6570 7014
rect 6670 7011 6818 7021
rect 6877 7041 6914 7051
rect 6989 7050 7026 7051
rect 6970 7048 7026 7050
rect 6877 7021 6885 7041
rect 6905 7021 6914 7041
rect 6726 7010 6762 7011
rect 6574 6879 6611 6880
rect 6877 6879 6914 7021
rect 6939 7041 7026 7048
rect 6939 7038 6997 7041
rect 6939 7018 6944 7038
rect 6965 7021 6997 7038
rect 7017 7021 7026 7041
rect 6965 7018 7026 7021
rect 6939 7011 7026 7018
rect 7085 7041 7122 7051
rect 7085 7021 7093 7041
rect 7113 7021 7122 7041
rect 6939 7010 6970 7011
rect 7085 6942 7122 7021
rect 7152 7050 7183 7103
rect 7202 7050 7239 7051
rect 7152 7041 7239 7050
rect 7152 7021 7210 7041
rect 7230 7021 7239 7041
rect 7152 7011 7239 7021
rect 7298 7041 7335 7051
rect 7298 7021 7306 7041
rect 7326 7021 7335 7041
rect 7152 7010 7183 7011
rect 7147 6942 7257 6955
rect 7298 6942 7335 7021
rect 7379 7021 7425 7104
rect 7719 7021 7794 7305
rect 8836 7230 8906 7438
rect 8968 7445 10171 7480
rect 8968 7431 8996 7445
rect 8970 7300 8996 7431
rect 9375 7442 10171 7445
rect 8828 7179 8908 7230
rect 8828 7153 8844 7179
rect 8884 7153 8908 7179
rect 8828 7134 8908 7153
rect 8828 7108 8847 7134
rect 8887 7108 8908 7134
rect 8828 7081 8908 7108
rect 8828 7055 8851 7081
rect 8891 7055 8908 7081
rect 8828 7044 8908 7055
rect 8970 7045 8997 7300
rect 9375 7292 9416 7442
rect 9647 7436 9751 7442
rect 10107 7439 10171 7442
rect 9842 7380 9963 7398
rect 9842 7378 9913 7380
rect 9842 7337 9857 7378
rect 9894 7339 9913 7378
rect 9950 7339 9963 7380
rect 9894 7337 9963 7339
rect 9842 7327 9963 7337
rect 9037 7185 9101 7197
rect 9377 7193 9414 7292
rect 9642 7282 9753 7295
rect 9642 7280 9684 7282
rect 9642 7260 9649 7280
rect 9668 7260 9684 7280
rect 9642 7252 9684 7260
rect 9712 7280 9753 7282
rect 9712 7260 9726 7280
rect 9745 7260 9753 7280
rect 9712 7252 9753 7260
rect 9642 7246 9753 7252
rect 9585 7224 9834 7246
rect 9585 7193 9622 7224
rect 9798 7222 9834 7224
rect 9798 7193 9835 7222
rect 9037 7184 9072 7185
rect 9014 7179 9072 7184
rect 9014 7159 9017 7179
rect 9037 7165 9072 7179
rect 9092 7165 9101 7185
rect 9037 7157 9101 7165
rect 9063 7156 9101 7157
rect 9064 7155 9101 7156
rect 9167 7189 9203 7190
rect 9275 7189 9311 7190
rect 9167 7181 9311 7189
rect 9167 7161 9175 7181
rect 9195 7161 9283 7181
rect 9303 7161 9311 7181
rect 9167 7155 9311 7161
rect 9377 7185 9415 7193
rect 9483 7189 9519 7190
rect 9377 7165 9386 7185
rect 9406 7165 9415 7185
rect 9377 7156 9415 7165
rect 9434 7182 9519 7189
rect 9434 7162 9441 7182
rect 9462 7181 9519 7182
rect 9462 7162 9491 7181
rect 9434 7161 9491 7162
rect 9511 7161 9519 7181
rect 9377 7155 9414 7156
rect 9434 7155 9519 7161
rect 9585 7185 9623 7193
rect 9696 7189 9732 7190
rect 9585 7165 9594 7185
rect 9614 7165 9623 7185
rect 9585 7156 9623 7165
rect 9647 7181 9732 7189
rect 9647 7161 9704 7181
rect 9724 7161 9732 7181
rect 9585 7155 9622 7156
rect 9647 7155 9732 7161
rect 9798 7185 9836 7193
rect 9798 7165 9807 7185
rect 9827 7165 9836 7185
rect 9891 7175 9956 7327
rect 10109 7301 10164 7439
rect 9798 7156 9836 7165
rect 9889 7168 9956 7175
rect 9798 7155 9835 7156
rect 9221 7134 9257 7155
rect 9647 7134 9678 7155
rect 9889 7147 9906 7168
rect 9942 7147 9956 7168
rect 10108 7188 10164 7301
rect 10108 7170 10127 7188
rect 10145 7170 10164 7188
rect 10108 7150 10164 7170
rect 9889 7134 9956 7147
rect 9054 7130 9154 7134
rect 9054 7126 9116 7130
rect 9054 7100 9061 7126
rect 9087 7104 9116 7126
rect 9142 7104 9154 7130
rect 9087 7100 9154 7104
rect 9054 7097 9154 7100
rect 9222 7097 9257 7134
rect 9319 7131 9678 7134
rect 9319 7126 9541 7131
rect 9319 7102 9332 7126
rect 9356 7107 9541 7126
rect 9565 7107 9678 7131
rect 9356 7102 9678 7107
rect 9319 7098 9678 7102
rect 9745 7128 9956 7134
rect 9745 7126 9906 7128
rect 9745 7106 9756 7126
rect 9776 7106 9906 7126
rect 9745 7099 9906 7106
rect 9745 7098 9786 7099
rect 9221 7072 9257 7097
rect 9069 7045 9106 7046
rect 9165 7045 9202 7046
rect 9221 7045 9228 7072
rect 7379 6986 7794 7021
rect 8969 7036 9107 7045
rect 8969 7016 9078 7036
rect 9098 7016 9107 7036
rect 8969 7009 9107 7016
rect 9165 7042 9228 7045
rect 9249 7045 9257 7072
rect 9276 7045 9313 7046
rect 9249 7042 9313 7045
rect 9165 7036 9313 7042
rect 9165 7016 9174 7036
rect 9194 7016 9284 7036
rect 9304 7016 9313 7036
rect 8969 7007 9065 7009
rect 9165 7006 9313 7016
rect 9372 7036 9409 7046
rect 9484 7045 9521 7046
rect 9465 7043 9521 7045
rect 9372 7016 9380 7036
rect 9400 7016 9409 7036
rect 9221 7005 9257 7006
rect 7379 6985 7425 6986
rect 7085 6940 7335 6942
rect 7085 6937 7186 6940
rect 7085 6918 7150 6937
rect 7147 6910 7150 6918
rect 7179 6910 7186 6937
rect 7214 6913 7224 6940
rect 7253 6918 7335 6940
rect 7719 6934 7794 6986
rect 7253 6913 7257 6918
rect 7214 6910 7257 6913
rect 7147 6896 7257 6910
rect 6573 6878 6914 6879
rect 6498 6873 6914 6878
rect 6498 6853 6501 6873
rect 6521 6853 6915 6873
rect 5555 6206 6361 6281
rect 4794 6162 4803 6196
rect 4832 6195 5242 6196
rect 4832 6162 4849 6195
rect 5074 6194 5242 6195
rect 4794 6136 4849 6162
rect 4794 6102 4802 6136
rect 4831 6102 4849 6136
rect 4794 6090 4849 6102
rect 2990 6045 3074 6066
rect 2990 6017 3018 6045
rect 3062 6017 3074 6045
rect 2804 5966 2878 5994
rect 2804 5918 2827 5966
rect 2864 5918 2878 5966
rect 2990 5988 3074 6017
rect 2990 5960 3015 5988
rect 3059 5960 3074 5988
rect 2990 5935 3074 5960
rect 5130 5949 5218 5953
rect 2804 5909 2878 5918
rect 437 5859 503 5907
rect 2814 5905 2878 5909
rect 5130 5932 5394 5949
rect 5130 5878 5310 5932
rect 5373 5878 5394 5932
rect 3027 5868 3738 5870
rect 2400 5867 3738 5868
rect 1350 5866 1422 5867
rect 437 5785 496 5859
rect 1349 5858 1448 5866
rect 1349 5855 1401 5858
rect 1349 5820 1357 5855
rect 1382 5820 1401 5855
rect 1426 5847 1448 5858
rect 2399 5859 3738 5867
rect 2399 5856 2451 5859
rect 1426 5846 2293 5847
rect 1426 5820 2294 5846
rect 1349 5810 2294 5820
rect 1349 5808 1448 5810
rect 437 5767 459 5785
rect 477 5767 496 5785
rect 437 5745 496 5767
rect 704 5781 1236 5786
rect 704 5761 1590 5781
rect 1610 5761 1613 5781
rect 2249 5777 2294 5810
rect 2399 5821 2407 5856
rect 2432 5821 2451 5856
rect 2476 5821 3738 5859
rect 2399 5812 3738 5821
rect 2399 5809 2488 5812
rect 3027 5810 3738 5812
rect 5130 5861 5394 5878
rect 704 5757 1613 5761
rect 704 5710 747 5757
rect 1197 5756 1613 5757
rect 2245 5757 2638 5777
rect 2658 5757 2661 5777
rect 1197 5755 1538 5756
rect 854 5724 964 5738
rect 854 5721 897 5724
rect 854 5716 858 5721
rect 692 5709 747 5710
rect 436 5686 747 5709
rect 436 5668 461 5686
rect 479 5674 747 5686
rect 776 5694 858 5716
rect 887 5694 897 5721
rect 925 5697 932 5724
rect 961 5716 964 5724
rect 961 5697 1026 5716
rect 925 5694 1026 5697
rect 776 5692 1026 5694
rect 479 5668 501 5674
rect 436 5529 501 5668
rect 776 5613 813 5692
rect 854 5679 964 5692
rect 928 5623 959 5624
rect 776 5593 785 5613
rect 805 5593 813 5613
rect 436 5511 459 5529
rect 477 5511 501 5529
rect 436 5494 501 5511
rect 656 5575 724 5588
rect 776 5583 813 5593
rect 872 5613 959 5623
rect 872 5593 881 5613
rect 901 5593 959 5613
rect 872 5584 959 5593
rect 872 5583 909 5584
rect 656 5533 663 5575
rect 712 5533 724 5575
rect 656 5530 724 5533
rect 928 5531 959 5584
rect 989 5613 1026 5692
rect 1141 5623 1172 5624
rect 989 5593 998 5613
rect 1018 5593 1026 5613
rect 989 5583 1026 5593
rect 1085 5616 1172 5623
rect 1085 5613 1146 5616
rect 1085 5593 1094 5613
rect 1114 5596 1146 5613
rect 1167 5596 1172 5616
rect 1114 5593 1172 5596
rect 1085 5586 1172 5593
rect 1197 5613 1234 5755
rect 1500 5754 1537 5755
rect 2245 5752 2661 5757
rect 2245 5751 2586 5752
rect 1902 5720 2012 5734
rect 1902 5717 1945 5720
rect 1902 5712 1906 5717
rect 1824 5690 1906 5712
rect 1935 5690 1945 5717
rect 1973 5693 1980 5720
rect 2009 5712 2012 5720
rect 2009 5693 2074 5712
rect 1973 5690 2074 5693
rect 1824 5688 2074 5690
rect 1349 5623 1385 5624
rect 1197 5593 1206 5613
rect 1226 5593 1234 5613
rect 1085 5584 1141 5586
rect 1085 5583 1122 5584
rect 1197 5583 1234 5593
rect 1293 5613 1441 5623
rect 1541 5620 1637 5622
rect 1293 5593 1302 5613
rect 1322 5593 1412 5613
rect 1432 5593 1441 5613
rect 1293 5587 1441 5593
rect 1293 5584 1357 5587
rect 1293 5583 1330 5584
rect 1349 5557 1357 5584
rect 1378 5584 1441 5587
rect 1499 5613 1637 5620
rect 1499 5593 1508 5613
rect 1528 5593 1637 5613
rect 1499 5584 1637 5593
rect 1824 5609 1861 5688
rect 1902 5675 2012 5688
rect 1976 5619 2007 5620
rect 1824 5589 1833 5609
rect 1853 5589 1861 5609
rect 1378 5557 1385 5584
rect 1404 5583 1441 5584
rect 1500 5583 1537 5584
rect 1349 5532 1385 5557
rect 820 5530 861 5531
rect 656 5523 861 5530
rect 656 5512 830 5523
rect 656 5479 664 5512
rect 657 5470 664 5479
rect 713 5503 830 5512
rect 850 5503 861 5523
rect 713 5495 861 5503
rect 928 5527 1287 5531
rect 928 5522 1250 5527
rect 928 5498 1041 5522
rect 1065 5503 1250 5522
rect 1274 5503 1287 5527
rect 1065 5498 1287 5503
rect 928 5495 1287 5498
rect 1349 5495 1384 5532
rect 1452 5529 1552 5532
rect 1452 5525 1519 5529
rect 1452 5499 1464 5525
rect 1490 5503 1519 5525
rect 1545 5503 1552 5529
rect 1490 5499 1552 5503
rect 1452 5495 1552 5499
rect 713 5479 724 5495
rect 713 5470 721 5479
rect 928 5474 959 5495
rect 1349 5474 1385 5495
rect 771 5473 808 5474
rect 436 5430 501 5449
rect 436 5412 461 5430
rect 479 5412 501 5430
rect 436 5211 501 5412
rect 657 5286 721 5470
rect 770 5464 808 5473
rect 770 5444 779 5464
rect 799 5444 808 5464
rect 770 5436 808 5444
rect 874 5468 959 5474
rect 984 5473 1021 5474
rect 874 5448 882 5468
rect 902 5448 959 5468
rect 874 5440 959 5448
rect 983 5464 1021 5473
rect 983 5444 992 5464
rect 1012 5444 1021 5464
rect 874 5439 910 5440
rect 983 5436 1021 5444
rect 1087 5468 1172 5474
rect 1192 5473 1229 5474
rect 1087 5448 1095 5468
rect 1115 5467 1172 5468
rect 1115 5448 1144 5467
rect 1087 5447 1144 5448
rect 1165 5447 1172 5467
rect 1087 5440 1172 5447
rect 1191 5464 1229 5473
rect 1191 5444 1200 5464
rect 1220 5444 1229 5464
rect 1087 5439 1123 5440
rect 1191 5436 1229 5444
rect 1295 5468 1439 5474
rect 1295 5448 1303 5468
rect 1323 5448 1411 5468
rect 1431 5448 1439 5468
rect 1295 5440 1439 5448
rect 1295 5439 1331 5440
rect 1403 5439 1439 5440
rect 1505 5473 1542 5474
rect 1505 5472 1543 5473
rect 1505 5464 1569 5472
rect 1505 5444 1514 5464
rect 1534 5450 1569 5464
rect 1589 5450 1592 5470
rect 1534 5445 1592 5450
rect 1534 5444 1569 5445
rect 771 5407 808 5436
rect 772 5405 808 5407
rect 984 5405 1021 5436
rect 772 5383 1021 5405
rect 853 5377 964 5383
rect 853 5369 894 5377
rect 853 5349 861 5369
rect 880 5349 894 5369
rect 853 5347 894 5349
rect 922 5369 964 5377
rect 922 5349 938 5369
rect 957 5349 964 5369
rect 922 5347 964 5349
rect 853 5332 964 5347
rect 657 5276 725 5286
rect 657 5243 674 5276
rect 714 5243 725 5276
rect 657 5231 725 5243
rect 657 5229 721 5231
rect 1192 5212 1229 5436
rect 1505 5432 1569 5444
rect 1609 5214 1636 5584
rect 1824 5579 1861 5589
rect 1920 5609 2007 5619
rect 1920 5589 1929 5609
rect 1949 5589 2007 5609
rect 1920 5580 2007 5589
rect 1920 5579 1957 5580
rect 1700 5566 1770 5571
rect 1695 5560 1770 5566
rect 1695 5527 1703 5560
rect 1756 5527 1770 5560
rect 1976 5527 2007 5580
rect 2037 5609 2074 5688
rect 2189 5619 2220 5620
rect 2037 5589 2046 5609
rect 2066 5589 2074 5609
rect 2037 5579 2074 5589
rect 2133 5612 2220 5619
rect 2133 5609 2194 5612
rect 2133 5589 2142 5609
rect 2162 5592 2194 5609
rect 2215 5592 2220 5612
rect 2162 5589 2220 5592
rect 2133 5582 2220 5589
rect 2245 5609 2282 5751
rect 2548 5750 2585 5751
rect 2397 5619 2433 5620
rect 2245 5589 2254 5609
rect 2274 5589 2282 5609
rect 2133 5580 2189 5582
rect 2133 5579 2170 5580
rect 2245 5579 2282 5589
rect 2341 5609 2489 5619
rect 2589 5616 2685 5618
rect 2341 5589 2350 5609
rect 2370 5589 2460 5609
rect 2480 5589 2489 5609
rect 2341 5583 2489 5589
rect 2341 5580 2405 5583
rect 2341 5579 2378 5580
rect 2397 5553 2405 5580
rect 2426 5580 2489 5583
rect 2547 5609 2685 5616
rect 2547 5589 2556 5609
rect 2576 5589 2685 5609
rect 2547 5580 2685 5589
rect 2426 5553 2433 5580
rect 2452 5579 2489 5580
rect 2548 5579 2585 5580
rect 2397 5528 2433 5553
rect 1695 5526 1778 5527
rect 1868 5526 1909 5527
rect 1695 5519 1909 5526
rect 1695 5502 1878 5519
rect 1695 5469 1708 5502
rect 1761 5499 1878 5502
rect 1898 5499 1909 5519
rect 1761 5491 1909 5499
rect 1976 5523 2335 5527
rect 1976 5518 2298 5523
rect 1976 5494 2089 5518
rect 2113 5499 2298 5518
rect 2322 5499 2335 5523
rect 2113 5494 2335 5499
rect 1976 5491 2335 5494
rect 2397 5491 2432 5528
rect 2500 5525 2600 5528
rect 2500 5521 2567 5525
rect 2500 5495 2512 5521
rect 2538 5499 2567 5521
rect 2593 5499 2600 5525
rect 2538 5495 2600 5499
rect 2500 5491 2600 5495
rect 1761 5469 1778 5491
rect 1976 5470 2007 5491
rect 2397 5470 2433 5491
rect 1819 5469 1856 5470
rect 1695 5455 1778 5469
rect 1468 5212 1636 5214
rect 1192 5211 1636 5212
rect 436 5181 1636 5211
rect 1706 5245 1778 5455
rect 1818 5460 1856 5469
rect 1818 5440 1827 5460
rect 1847 5440 1856 5460
rect 1818 5432 1856 5440
rect 1922 5464 2007 5470
rect 2032 5469 2069 5470
rect 1922 5444 1930 5464
rect 1950 5444 2007 5464
rect 1922 5436 2007 5444
rect 2031 5460 2069 5469
rect 2031 5440 2040 5460
rect 2060 5440 2069 5460
rect 1922 5435 1958 5436
rect 2031 5432 2069 5440
rect 2135 5464 2220 5470
rect 2240 5469 2277 5470
rect 2135 5444 2143 5464
rect 2163 5463 2220 5464
rect 2163 5444 2192 5463
rect 2135 5443 2192 5444
rect 2213 5443 2220 5463
rect 2135 5436 2220 5443
rect 2239 5460 2277 5469
rect 2239 5440 2248 5460
rect 2268 5440 2277 5460
rect 2135 5435 2171 5436
rect 2239 5432 2277 5440
rect 2343 5464 2487 5470
rect 2343 5444 2351 5464
rect 2371 5444 2459 5464
rect 2479 5444 2487 5464
rect 2343 5436 2487 5444
rect 2343 5435 2379 5436
rect 2451 5435 2487 5436
rect 2553 5469 2590 5470
rect 2553 5468 2591 5469
rect 2553 5460 2617 5468
rect 2553 5440 2562 5460
rect 2582 5446 2617 5460
rect 2637 5446 2640 5466
rect 2582 5441 2640 5446
rect 2582 5440 2617 5441
rect 1819 5403 1856 5432
rect 1820 5401 1856 5403
rect 2032 5401 2069 5432
rect 1820 5379 2069 5401
rect 1901 5373 2012 5379
rect 1901 5365 1942 5373
rect 1901 5345 1909 5365
rect 1928 5345 1942 5365
rect 1901 5343 1942 5345
rect 1970 5365 2012 5373
rect 1970 5345 1986 5365
rect 2005 5345 2012 5365
rect 1970 5343 2012 5345
rect 1901 5328 2012 5343
rect 1706 5206 1725 5245
rect 1770 5206 1778 5245
rect 1706 5189 1778 5206
rect 2240 5233 2277 5432
rect 2553 5428 2617 5440
rect 2240 5227 2281 5233
rect 2657 5229 2684 5580
rect 2979 5567 3074 5593
rect 2815 5545 2879 5564
rect 2815 5506 2828 5545
rect 2862 5506 2879 5545
rect 2815 5487 2879 5506
rect 2516 5227 2684 5229
rect 2240 5201 2684 5227
rect 436 5134 501 5181
rect 436 5116 459 5134
rect 477 5116 501 5134
rect 1349 5161 1384 5163
rect 1349 5159 1453 5161
rect 2242 5159 2281 5201
rect 2516 5200 2684 5201
rect 1349 5152 2283 5159
rect 1349 5151 1400 5152
rect 1349 5131 1352 5151
rect 1377 5132 1400 5151
rect 1432 5132 2283 5152
rect 1377 5131 2283 5132
rect 1349 5124 2283 5131
rect 1622 5123 2283 5124
rect 436 5095 501 5116
rect 713 5106 753 5109
rect 713 5102 1616 5106
rect 713 5082 1590 5102
rect 1610 5082 1616 5102
rect 713 5079 1616 5082
rect 437 5035 502 5055
rect 437 5017 461 5035
rect 479 5017 502 5035
rect 437 4990 502 5017
rect 713 4990 753 5079
rect 1197 5077 1613 5079
rect 1197 5076 1538 5077
rect 854 5045 964 5059
rect 854 5042 897 5045
rect 854 5037 858 5042
rect 436 4955 753 4990
rect 776 5015 858 5037
rect 887 5015 897 5042
rect 925 5018 932 5045
rect 961 5037 964 5045
rect 961 5018 1026 5037
rect 925 5015 1026 5018
rect 776 5013 1026 5015
rect 437 4879 502 4955
rect 776 4934 813 5013
rect 854 5000 964 5013
rect 928 4944 959 4945
rect 776 4914 785 4934
rect 805 4914 813 4934
rect 776 4904 813 4914
rect 872 4934 959 4944
rect 872 4914 881 4934
rect 901 4914 959 4934
rect 872 4905 959 4914
rect 872 4904 909 4905
rect 437 4861 459 4879
rect 477 4861 502 4879
rect 437 4840 502 4861
rect 650 4859 715 4868
rect 650 4822 660 4859
rect 700 4851 715 4859
rect 928 4852 959 4905
rect 989 4934 1026 5013
rect 1141 4944 1172 4945
rect 989 4914 998 4934
rect 1018 4914 1026 4934
rect 989 4904 1026 4914
rect 1085 4937 1172 4944
rect 1085 4934 1146 4937
rect 1085 4914 1094 4934
rect 1114 4917 1146 4934
rect 1167 4917 1172 4937
rect 1114 4914 1172 4917
rect 1085 4907 1172 4914
rect 1197 4934 1234 5076
rect 1500 5075 1537 5076
rect 2817 5016 2879 5487
rect 2979 5526 3005 5567
rect 3041 5526 3074 5567
rect 2979 5230 3074 5526
rect 2979 5186 2994 5230
rect 3054 5186 3074 5230
rect 2979 5166 3074 5186
rect 3691 5097 3734 5810
rect 3691 5077 4085 5097
rect 4105 5077 4108 5097
rect 3692 5072 4108 5077
rect 3692 5071 4033 5072
rect 3349 5040 3459 5054
rect 3349 5037 3392 5040
rect 3349 5032 3353 5037
rect 2812 4964 2887 5016
rect 3271 5010 3353 5032
rect 3382 5010 3392 5037
rect 3420 5013 3427 5040
rect 3456 5032 3459 5040
rect 3456 5013 3521 5032
rect 3420 5010 3521 5013
rect 3271 5008 3521 5010
rect 3181 4964 3227 4965
rect 1349 4944 1385 4945
rect 1197 4914 1206 4934
rect 1226 4914 1234 4934
rect 1085 4905 1141 4907
rect 1085 4904 1122 4905
rect 1197 4904 1234 4914
rect 1293 4934 1441 4944
rect 1541 4941 1637 4943
rect 1293 4914 1302 4934
rect 1322 4914 1412 4934
rect 1432 4914 1441 4934
rect 1293 4908 1441 4914
rect 1293 4905 1357 4908
rect 1293 4904 1330 4905
rect 1349 4878 1357 4905
rect 1378 4905 1441 4908
rect 1499 4934 1637 4941
rect 1499 4914 1508 4934
rect 1528 4914 1637 4934
rect 1499 4905 1637 4914
rect 2812 4929 3227 4964
rect 1378 4878 1385 4905
rect 1404 4904 1441 4905
rect 1500 4904 1537 4905
rect 1349 4853 1385 4878
rect 820 4851 861 4852
rect 700 4844 861 4851
rect 700 4824 830 4844
rect 850 4824 861 4844
rect 700 4822 861 4824
rect 650 4816 861 4822
rect 928 4848 1287 4852
rect 928 4843 1250 4848
rect 928 4819 1041 4843
rect 1065 4824 1250 4843
rect 1274 4824 1287 4848
rect 1065 4819 1287 4824
rect 928 4816 1287 4819
rect 1349 4816 1384 4853
rect 1452 4850 1552 4853
rect 1452 4846 1519 4850
rect 1452 4820 1464 4846
rect 1490 4824 1519 4846
rect 1545 4824 1552 4850
rect 1490 4820 1552 4824
rect 1452 4816 1552 4820
rect 650 4803 717 4816
rect 442 4780 498 4800
rect 442 4762 461 4780
rect 479 4762 498 4780
rect 442 4649 498 4762
rect 650 4782 664 4803
rect 700 4782 717 4803
rect 928 4795 959 4816
rect 1349 4795 1385 4816
rect 771 4794 808 4795
rect 650 4775 717 4782
rect 770 4785 808 4794
rect 442 4511 497 4649
rect 650 4623 715 4775
rect 770 4765 779 4785
rect 799 4765 808 4785
rect 770 4757 808 4765
rect 874 4789 959 4795
rect 984 4794 1021 4795
rect 874 4769 882 4789
rect 902 4769 959 4789
rect 874 4761 959 4769
rect 983 4785 1021 4794
rect 983 4765 992 4785
rect 1012 4765 1021 4785
rect 874 4760 910 4761
rect 983 4757 1021 4765
rect 1087 4789 1172 4795
rect 1192 4794 1229 4795
rect 1087 4769 1095 4789
rect 1115 4788 1172 4789
rect 1115 4769 1144 4788
rect 1087 4768 1144 4769
rect 1165 4768 1172 4788
rect 1087 4761 1172 4768
rect 1191 4785 1229 4794
rect 1191 4765 1200 4785
rect 1220 4765 1229 4785
rect 1087 4760 1123 4761
rect 1191 4757 1229 4765
rect 1295 4789 1439 4795
rect 1295 4769 1303 4789
rect 1323 4769 1411 4789
rect 1431 4769 1439 4789
rect 1295 4761 1439 4769
rect 1295 4760 1331 4761
rect 1403 4760 1439 4761
rect 1505 4794 1542 4795
rect 1505 4793 1543 4794
rect 1505 4785 1569 4793
rect 1505 4765 1514 4785
rect 1534 4771 1569 4785
rect 1589 4771 1592 4791
rect 1534 4766 1592 4771
rect 1534 4765 1569 4766
rect 771 4728 808 4757
rect 772 4726 808 4728
rect 984 4726 1021 4757
rect 772 4704 1021 4726
rect 853 4698 964 4704
rect 853 4690 894 4698
rect 853 4670 861 4690
rect 880 4670 894 4690
rect 853 4668 894 4670
rect 922 4690 964 4698
rect 922 4670 938 4690
rect 957 4670 964 4690
rect 922 4668 964 4670
rect 853 4655 964 4668
rect 1192 4658 1229 4757
rect 1505 4753 1569 4765
rect 643 4613 764 4623
rect 643 4611 712 4613
rect 643 4570 656 4611
rect 693 4572 712 4611
rect 749 4572 764 4613
rect 693 4570 764 4572
rect 643 4552 764 4570
rect 435 4508 499 4511
rect 855 4508 959 4514
rect 1190 4508 1231 4658
rect 1609 4650 1636 4905
rect 1698 4895 1778 4906
rect 1698 4869 1715 4895
rect 1755 4869 1778 4895
rect 1698 4842 1778 4869
rect 1698 4816 1719 4842
rect 1759 4816 1778 4842
rect 1698 4797 1778 4816
rect 1698 4771 1722 4797
rect 1762 4771 1778 4797
rect 1698 4720 1778 4771
rect 435 4505 1231 4508
rect 1610 4519 1636 4650
rect 1610 4505 1638 4519
rect 435 4470 1638 4505
rect 1700 4512 1770 4720
rect 2812 4645 2887 4929
rect 3181 4846 3227 4929
rect 3271 4929 3308 5008
rect 3349 4995 3459 5008
rect 3423 4939 3454 4940
rect 3271 4909 3280 4929
rect 3300 4909 3308 4929
rect 3271 4899 3308 4909
rect 3367 4929 3454 4939
rect 3367 4909 3376 4929
rect 3396 4909 3454 4929
rect 3367 4900 3454 4909
rect 3367 4899 3404 4900
rect 3423 4847 3454 4900
rect 3484 4929 3521 5008
rect 3636 4939 3667 4940
rect 3484 4909 3493 4929
rect 3513 4909 3521 4929
rect 3484 4899 3521 4909
rect 3580 4932 3667 4939
rect 3580 4929 3641 4932
rect 3580 4909 3589 4929
rect 3609 4912 3641 4929
rect 3662 4912 3667 4932
rect 3609 4909 3667 4912
rect 3580 4902 3667 4909
rect 3692 4929 3729 5071
rect 3995 5070 4032 5071
rect 3844 4939 3880 4940
rect 3692 4909 3701 4929
rect 3721 4909 3729 4929
rect 3580 4900 3636 4902
rect 3580 4899 3617 4900
rect 3692 4899 3729 4909
rect 3788 4929 3936 4939
rect 4036 4936 4132 4938
rect 3788 4909 3797 4929
rect 3817 4909 3907 4929
rect 3927 4909 3936 4929
rect 3788 4903 3936 4909
rect 3788 4900 3852 4903
rect 3788 4899 3825 4900
rect 3844 4873 3852 4900
rect 3873 4900 3936 4903
rect 3994 4929 4132 4936
rect 3994 4909 4003 4929
rect 4023 4909 4132 4929
rect 3994 4900 4132 4909
rect 3873 4873 3880 4900
rect 3899 4899 3936 4900
rect 3995 4899 4032 4900
rect 3844 4848 3880 4873
rect 3315 4846 3356 4847
rect 3181 4839 3356 4846
rect 2979 4813 3065 4832
rect 2979 4772 2994 4813
rect 3048 4772 3065 4813
rect 3181 4819 3325 4839
rect 3345 4819 3356 4839
rect 3181 4811 3356 4819
rect 3423 4843 3782 4847
rect 3423 4838 3745 4843
rect 3423 4814 3536 4838
rect 3560 4819 3745 4838
rect 3769 4819 3782 4843
rect 3560 4814 3782 4819
rect 3423 4811 3782 4814
rect 3844 4811 3879 4848
rect 3947 4845 4047 4848
rect 3947 4841 4014 4845
rect 3947 4815 3959 4841
rect 3985 4819 4014 4841
rect 4040 4819 4047 4845
rect 3985 4815 4047 4819
rect 3947 4811 4047 4815
rect 3181 4807 3227 4811
rect 3423 4790 3454 4811
rect 3844 4790 3880 4811
rect 3266 4789 3303 4790
rect 2979 4736 3065 4772
rect 3265 4780 3303 4789
rect 3265 4760 3274 4780
rect 3294 4760 3303 4780
rect 3265 4752 3303 4760
rect 3369 4784 3454 4790
rect 3479 4789 3516 4790
rect 3369 4764 3377 4784
rect 3397 4764 3454 4784
rect 3369 4756 3454 4764
rect 3478 4780 3516 4789
rect 3478 4760 3487 4780
rect 3507 4760 3516 4780
rect 3369 4755 3405 4756
rect 3478 4752 3516 4760
rect 3582 4784 3667 4790
rect 3687 4789 3724 4790
rect 3582 4764 3590 4784
rect 3610 4783 3667 4784
rect 3610 4764 3639 4783
rect 3582 4763 3639 4764
rect 3660 4763 3667 4783
rect 3582 4756 3667 4763
rect 3686 4780 3724 4789
rect 3686 4760 3695 4780
rect 3715 4760 3724 4780
rect 3582 4755 3618 4756
rect 3686 4752 3724 4760
rect 3790 4784 3934 4790
rect 3790 4764 3798 4784
rect 3818 4764 3906 4784
rect 3926 4764 3934 4784
rect 3790 4756 3934 4764
rect 3790 4755 3826 4756
rect 435 4409 499 4470
rect 855 4468 959 4470
rect 1190 4468 1231 4470
rect 1700 4467 1721 4512
rect 1701 4446 1721 4467
rect 1751 4467 1770 4512
rect 2807 4603 2887 4645
rect 1751 4446 1768 4467
rect 1701 4427 1768 4446
rect 1350 4419 1422 4420
rect 1349 4411 1448 4419
rect 437 4338 496 4409
rect 1349 4408 1401 4411
rect 1349 4373 1357 4408
rect 1382 4373 1401 4408
rect 1426 4400 1448 4411
rect 1426 4399 2293 4400
rect 1426 4373 2294 4399
rect 1349 4363 2294 4373
rect 1349 4361 1448 4363
rect 437 4320 459 4338
rect 477 4320 496 4338
rect 437 4298 496 4320
rect 704 4334 1236 4339
rect 704 4314 1590 4334
rect 1610 4314 1613 4334
rect 2249 4330 2294 4363
rect 704 4310 1613 4314
rect 704 4263 747 4310
rect 1197 4309 1613 4310
rect 2245 4310 2638 4330
rect 2658 4310 2661 4330
rect 1197 4308 1538 4309
rect 854 4277 964 4291
rect 854 4274 897 4277
rect 854 4269 858 4274
rect 692 4262 747 4263
rect 436 4239 747 4262
rect 436 4221 461 4239
rect 479 4227 747 4239
rect 776 4247 858 4269
rect 887 4247 897 4274
rect 925 4250 932 4277
rect 961 4269 964 4277
rect 961 4250 1026 4269
rect 925 4247 1026 4250
rect 776 4245 1026 4247
rect 479 4221 501 4227
rect 436 4082 501 4221
rect 776 4166 813 4245
rect 854 4232 964 4245
rect 928 4176 959 4177
rect 776 4146 785 4166
rect 805 4146 813 4166
rect 436 4064 459 4082
rect 477 4064 501 4082
rect 436 4047 501 4064
rect 656 4128 724 4141
rect 776 4136 813 4146
rect 872 4166 959 4176
rect 872 4146 881 4166
rect 901 4146 959 4166
rect 872 4137 959 4146
rect 872 4136 909 4137
rect 656 4086 663 4128
rect 712 4086 724 4128
rect 656 4083 724 4086
rect 928 4084 959 4137
rect 989 4166 1026 4245
rect 1141 4176 1172 4177
rect 989 4146 998 4166
rect 1018 4146 1026 4166
rect 989 4136 1026 4146
rect 1085 4169 1172 4176
rect 1085 4166 1146 4169
rect 1085 4146 1094 4166
rect 1114 4149 1146 4166
rect 1167 4149 1172 4169
rect 1114 4146 1172 4149
rect 1085 4139 1172 4146
rect 1197 4166 1234 4308
rect 1500 4307 1537 4308
rect 2245 4305 2661 4310
rect 2245 4304 2586 4305
rect 1902 4273 2012 4287
rect 1902 4270 1945 4273
rect 1902 4265 1906 4270
rect 1824 4243 1906 4265
rect 1935 4243 1945 4270
rect 1973 4246 1980 4273
rect 2009 4265 2012 4273
rect 2009 4246 2074 4265
rect 1973 4243 2074 4246
rect 1824 4241 2074 4243
rect 1349 4176 1385 4177
rect 1197 4146 1206 4166
rect 1226 4146 1234 4166
rect 1085 4137 1141 4139
rect 1085 4136 1122 4137
rect 1197 4136 1234 4146
rect 1293 4166 1441 4176
rect 1541 4173 1637 4175
rect 1293 4146 1302 4166
rect 1322 4146 1412 4166
rect 1432 4146 1441 4166
rect 1293 4140 1441 4146
rect 1293 4137 1357 4140
rect 1293 4136 1330 4137
rect 1349 4110 1357 4137
rect 1378 4137 1441 4140
rect 1499 4166 1637 4173
rect 1499 4146 1508 4166
rect 1528 4146 1637 4166
rect 1499 4137 1637 4146
rect 1824 4162 1861 4241
rect 1902 4228 2012 4241
rect 1976 4172 2007 4173
rect 1824 4142 1833 4162
rect 1853 4142 1861 4162
rect 1378 4110 1385 4137
rect 1404 4136 1441 4137
rect 1500 4136 1537 4137
rect 1349 4085 1385 4110
rect 820 4083 861 4084
rect 656 4076 861 4083
rect 656 4065 830 4076
rect 656 4032 664 4065
rect 657 4023 664 4032
rect 713 4056 830 4065
rect 850 4056 861 4076
rect 713 4048 861 4056
rect 928 4080 1287 4084
rect 928 4075 1250 4080
rect 928 4051 1041 4075
rect 1065 4056 1250 4075
rect 1274 4056 1287 4080
rect 1065 4051 1287 4056
rect 928 4048 1287 4051
rect 1349 4048 1384 4085
rect 1452 4082 1552 4085
rect 1452 4078 1519 4082
rect 1452 4052 1464 4078
rect 1490 4056 1519 4078
rect 1545 4056 1552 4082
rect 1490 4052 1552 4056
rect 1452 4048 1552 4052
rect 713 4032 724 4048
rect 713 4023 721 4032
rect 928 4027 959 4048
rect 1349 4027 1385 4048
rect 771 4026 808 4027
rect 436 3983 501 4002
rect 436 3965 461 3983
rect 479 3965 501 3983
rect 436 3764 501 3965
rect 657 3839 721 4023
rect 770 4017 808 4026
rect 770 3997 779 4017
rect 799 3997 808 4017
rect 770 3989 808 3997
rect 874 4021 959 4027
rect 984 4026 1021 4027
rect 874 4001 882 4021
rect 902 4001 959 4021
rect 874 3993 959 4001
rect 983 4017 1021 4026
rect 983 3997 992 4017
rect 1012 3997 1021 4017
rect 874 3992 910 3993
rect 983 3989 1021 3997
rect 1087 4021 1172 4027
rect 1192 4026 1229 4027
rect 1087 4001 1095 4021
rect 1115 4020 1172 4021
rect 1115 4001 1144 4020
rect 1087 4000 1144 4001
rect 1165 4000 1172 4020
rect 1087 3993 1172 4000
rect 1191 4017 1229 4026
rect 1191 3997 1200 4017
rect 1220 3997 1229 4017
rect 1087 3992 1123 3993
rect 1191 3989 1229 3997
rect 1295 4021 1439 4027
rect 1295 4001 1303 4021
rect 1323 4001 1411 4021
rect 1431 4001 1439 4021
rect 1295 3993 1439 4001
rect 1295 3992 1331 3993
rect 1403 3992 1439 3993
rect 1505 4026 1542 4027
rect 1505 4025 1543 4026
rect 1505 4017 1569 4025
rect 1505 3997 1514 4017
rect 1534 4003 1569 4017
rect 1589 4003 1592 4023
rect 1534 3998 1592 4003
rect 1534 3997 1569 3998
rect 771 3960 808 3989
rect 772 3958 808 3960
rect 984 3958 1021 3989
rect 772 3936 1021 3958
rect 853 3930 964 3936
rect 853 3922 894 3930
rect 853 3902 861 3922
rect 880 3902 894 3922
rect 853 3900 894 3902
rect 922 3922 964 3930
rect 922 3902 938 3922
rect 957 3902 964 3922
rect 922 3900 964 3902
rect 853 3885 964 3900
rect 657 3829 725 3839
rect 657 3796 674 3829
rect 714 3796 725 3829
rect 657 3784 725 3796
rect 657 3782 721 3784
rect 1192 3765 1229 3989
rect 1505 3985 1569 3997
rect 1609 3767 1636 4137
rect 1824 4132 1861 4142
rect 1920 4162 2007 4172
rect 1920 4142 1929 4162
rect 1949 4142 2007 4162
rect 1920 4133 2007 4142
rect 1920 4132 1957 4133
rect 1700 4119 1770 4124
rect 1695 4113 1770 4119
rect 1695 4080 1703 4113
rect 1756 4080 1770 4113
rect 1976 4080 2007 4133
rect 2037 4162 2074 4241
rect 2189 4172 2220 4173
rect 2037 4142 2046 4162
rect 2066 4142 2074 4162
rect 2037 4132 2074 4142
rect 2133 4165 2220 4172
rect 2133 4162 2194 4165
rect 2133 4142 2142 4162
rect 2162 4145 2194 4162
rect 2215 4145 2220 4165
rect 2162 4142 2220 4145
rect 2133 4135 2220 4142
rect 2245 4162 2282 4304
rect 2548 4303 2585 4304
rect 2397 4172 2433 4173
rect 2245 4142 2254 4162
rect 2274 4142 2282 4162
rect 2133 4133 2189 4135
rect 2133 4132 2170 4133
rect 2245 4132 2282 4142
rect 2341 4162 2489 4172
rect 2589 4169 2685 4171
rect 2341 4142 2350 4162
rect 2370 4142 2460 4162
rect 2480 4142 2489 4162
rect 2341 4136 2489 4142
rect 2341 4133 2405 4136
rect 2341 4132 2378 4133
rect 2397 4106 2405 4133
rect 2426 4133 2489 4136
rect 2547 4162 2685 4169
rect 2547 4142 2556 4162
rect 2576 4142 2685 4162
rect 2547 4133 2685 4142
rect 2426 4106 2433 4133
rect 2452 4132 2489 4133
rect 2548 4132 2585 4133
rect 2397 4081 2433 4106
rect 1695 4079 1778 4080
rect 1868 4079 1909 4080
rect 1695 4072 1909 4079
rect 1695 4055 1878 4072
rect 1695 4022 1708 4055
rect 1761 4052 1878 4055
rect 1898 4052 1909 4072
rect 1761 4044 1909 4052
rect 1976 4076 2335 4080
rect 1976 4071 2298 4076
rect 1976 4047 2089 4071
rect 2113 4052 2298 4071
rect 2322 4052 2335 4076
rect 2113 4047 2335 4052
rect 1976 4044 2335 4047
rect 2397 4044 2432 4081
rect 2500 4078 2600 4081
rect 2500 4074 2567 4078
rect 2500 4048 2512 4074
rect 2538 4052 2567 4074
rect 2593 4052 2600 4078
rect 2538 4048 2600 4052
rect 2500 4044 2600 4048
rect 1761 4022 1778 4044
rect 1976 4023 2007 4044
rect 2397 4023 2433 4044
rect 1819 4022 1856 4023
rect 1695 4008 1778 4022
rect 1468 3765 1636 3767
rect 1192 3764 1636 3765
rect 436 3734 1636 3764
rect 1706 3798 1778 4008
rect 1818 4013 1856 4022
rect 1818 3993 1827 4013
rect 1847 3993 1856 4013
rect 1818 3985 1856 3993
rect 1922 4017 2007 4023
rect 2032 4022 2069 4023
rect 1922 3997 1930 4017
rect 1950 3997 2007 4017
rect 1922 3989 2007 3997
rect 2031 4013 2069 4022
rect 2031 3993 2040 4013
rect 2060 3993 2069 4013
rect 1922 3988 1958 3989
rect 2031 3985 2069 3993
rect 2135 4017 2220 4023
rect 2240 4022 2277 4023
rect 2135 3997 2143 4017
rect 2163 4016 2220 4017
rect 2163 3997 2192 4016
rect 2135 3996 2192 3997
rect 2213 3996 2220 4016
rect 2135 3989 2220 3996
rect 2239 4013 2277 4022
rect 2239 3993 2248 4013
rect 2268 3993 2277 4013
rect 2135 3988 2171 3989
rect 2239 3985 2277 3993
rect 2343 4017 2487 4023
rect 2343 3997 2351 4017
rect 2371 3997 2459 4017
rect 2479 3997 2487 4017
rect 2343 3989 2487 3997
rect 2343 3988 2379 3989
rect 2451 3988 2487 3989
rect 2553 4022 2590 4023
rect 2553 4021 2591 4022
rect 2553 4013 2617 4021
rect 2553 3993 2562 4013
rect 2582 3999 2617 4013
rect 2637 3999 2640 4019
rect 2582 3994 2640 3999
rect 2582 3993 2617 3994
rect 1819 3956 1856 3985
rect 1820 3954 1856 3956
rect 2032 3954 2069 3985
rect 1820 3932 2069 3954
rect 1901 3926 2012 3932
rect 1901 3918 1942 3926
rect 1901 3898 1909 3918
rect 1928 3898 1942 3918
rect 1901 3896 1942 3898
rect 1970 3918 2012 3926
rect 1970 3898 1986 3918
rect 2005 3898 2012 3918
rect 1970 3896 2012 3898
rect 1901 3881 2012 3896
rect 1706 3759 1725 3798
rect 1770 3759 1778 3798
rect 1706 3742 1778 3759
rect 2240 3786 2277 3985
rect 2553 3981 2617 3993
rect 2240 3780 2281 3786
rect 2657 3782 2684 4133
rect 2807 4003 2886 4603
rect 2983 4151 3062 4736
rect 3266 4723 3303 4752
rect 3267 4721 3303 4723
rect 3479 4721 3516 4752
rect 3267 4699 3516 4721
rect 3348 4693 3459 4699
rect 3348 4685 3389 4693
rect 3348 4665 3356 4685
rect 3375 4665 3389 4685
rect 3348 4663 3389 4665
rect 3417 4685 3459 4693
rect 3417 4665 3433 4685
rect 3452 4665 3459 4685
rect 3417 4663 3459 4665
rect 3348 4648 3459 4663
rect 3687 4637 3724 4752
rect 3680 4525 3727 4637
rect 3848 4597 3878 4756
rect 3898 4755 3934 4756
rect 4000 4789 4037 4790
rect 4000 4788 4038 4789
rect 4000 4780 4064 4788
rect 4000 4760 4009 4780
rect 4029 4766 4064 4780
rect 4084 4766 4087 4786
rect 4029 4761 4087 4766
rect 4029 4760 4064 4761
rect 4000 4748 4064 4760
rect 3848 4593 3934 4597
rect 3848 4575 3863 4593
rect 3915 4575 3934 4593
rect 3848 4566 3934 4575
rect 4104 4527 4131 4900
rect 3963 4525 4131 4527
rect 3680 4499 4131 4525
rect 3680 4421 3727 4499
rect 3963 4498 4131 4499
rect 3625 4420 3727 4421
rect 3624 4412 3727 4420
rect 3624 4409 3676 4412
rect 3624 4374 3632 4409
rect 3657 4374 3676 4409
rect 3701 4374 3727 4412
rect 3624 4368 3727 4374
rect 3887 4413 3923 4417
rect 3887 4390 3895 4413
rect 3919 4390 3923 4413
rect 3887 4369 3923 4390
rect 3624 4364 3723 4368
rect 3887 4346 3895 4369
rect 3919 4346 3923 4369
rect 2516 3780 2684 3782
rect 2240 3754 2684 3780
rect 436 3687 501 3734
rect 436 3669 459 3687
rect 477 3669 501 3687
rect 1349 3714 1384 3716
rect 1349 3712 1453 3714
rect 2242 3712 2281 3754
rect 2516 3753 2684 3754
rect 1349 3705 2283 3712
rect 1349 3704 1400 3705
rect 1349 3684 1352 3704
rect 1377 3685 1400 3704
rect 1432 3685 2283 3705
rect 1377 3684 2283 3685
rect 1349 3677 2283 3684
rect 1622 3676 2283 3677
rect 436 3648 501 3669
rect 713 3659 753 3662
rect 713 3655 1616 3659
rect 713 3635 1590 3655
rect 1610 3635 1616 3655
rect 713 3632 1616 3635
rect 437 3588 502 3608
rect 437 3570 461 3588
rect 479 3570 502 3588
rect 437 3543 502 3570
rect 713 3543 753 3632
rect 1197 3630 1613 3632
rect 1197 3629 1538 3630
rect 854 3598 964 3612
rect 854 3595 897 3598
rect 854 3590 858 3595
rect 436 3508 753 3543
rect 776 3568 858 3590
rect 887 3568 897 3595
rect 925 3571 932 3598
rect 961 3590 964 3598
rect 961 3571 1026 3590
rect 925 3568 1026 3571
rect 776 3566 1026 3568
rect 437 3432 502 3508
rect 776 3487 813 3566
rect 854 3553 964 3566
rect 928 3497 959 3498
rect 776 3467 785 3487
rect 805 3467 813 3487
rect 776 3457 813 3467
rect 872 3487 959 3497
rect 872 3467 881 3487
rect 901 3467 959 3487
rect 872 3458 959 3467
rect 872 3457 909 3458
rect 437 3414 459 3432
rect 477 3414 502 3432
rect 437 3393 502 3414
rect 650 3412 715 3421
rect 650 3375 660 3412
rect 700 3404 715 3412
rect 928 3405 959 3458
rect 989 3487 1026 3566
rect 1141 3497 1172 3498
rect 989 3467 998 3487
rect 1018 3467 1026 3487
rect 989 3457 1026 3467
rect 1085 3490 1172 3497
rect 1085 3487 1146 3490
rect 1085 3467 1094 3487
rect 1114 3470 1146 3487
rect 1167 3470 1172 3490
rect 1114 3467 1172 3470
rect 1085 3460 1172 3467
rect 1197 3487 1234 3629
rect 1500 3628 1537 3629
rect 1349 3497 1385 3498
rect 1197 3467 1206 3487
rect 1226 3467 1234 3487
rect 1085 3458 1141 3460
rect 1085 3457 1122 3458
rect 1197 3457 1234 3467
rect 1293 3487 1441 3497
rect 1541 3494 1637 3496
rect 1293 3467 1302 3487
rect 1322 3467 1412 3487
rect 1432 3467 1441 3487
rect 1293 3461 1441 3467
rect 1293 3458 1357 3461
rect 1293 3457 1330 3458
rect 1349 3431 1357 3458
rect 1378 3458 1441 3461
rect 1499 3487 1637 3494
rect 1499 3467 1508 3487
rect 1528 3467 1637 3487
rect 1499 3458 1637 3467
rect 1378 3431 1385 3458
rect 1404 3457 1441 3458
rect 1500 3457 1537 3458
rect 1349 3406 1385 3431
rect 820 3404 861 3405
rect 700 3397 861 3404
rect 700 3377 830 3397
rect 850 3377 861 3397
rect 700 3375 861 3377
rect 650 3369 861 3375
rect 928 3401 1287 3405
rect 928 3396 1250 3401
rect 928 3372 1041 3396
rect 1065 3377 1250 3396
rect 1274 3377 1287 3401
rect 1065 3372 1287 3377
rect 928 3369 1287 3372
rect 1349 3369 1384 3406
rect 1452 3403 1552 3406
rect 1452 3399 1519 3403
rect 1452 3373 1464 3399
rect 1490 3377 1519 3399
rect 1545 3377 1552 3403
rect 1490 3373 1552 3377
rect 1452 3369 1552 3373
rect 650 3356 717 3369
rect 442 3333 498 3353
rect 442 3315 461 3333
rect 479 3315 498 3333
rect 442 3202 498 3315
rect 650 3335 664 3356
rect 700 3335 717 3356
rect 928 3348 959 3369
rect 1349 3348 1385 3369
rect 771 3347 808 3348
rect 650 3328 717 3335
rect 770 3338 808 3347
rect 442 3073 497 3202
rect 650 3176 715 3328
rect 770 3318 779 3338
rect 799 3318 808 3338
rect 770 3310 808 3318
rect 874 3342 959 3348
rect 984 3347 1021 3348
rect 874 3322 882 3342
rect 902 3322 959 3342
rect 874 3314 959 3322
rect 983 3338 1021 3347
rect 983 3318 992 3338
rect 1012 3318 1021 3338
rect 874 3313 910 3314
rect 983 3310 1021 3318
rect 1087 3342 1172 3348
rect 1192 3347 1229 3348
rect 1087 3322 1095 3342
rect 1115 3341 1172 3342
rect 1115 3322 1144 3341
rect 1087 3321 1144 3322
rect 1165 3321 1172 3341
rect 1087 3314 1172 3321
rect 1191 3338 1229 3347
rect 1191 3318 1200 3338
rect 1220 3318 1229 3338
rect 1087 3313 1123 3314
rect 1191 3310 1229 3318
rect 1295 3342 1439 3348
rect 1295 3322 1303 3342
rect 1323 3322 1411 3342
rect 1431 3322 1439 3342
rect 1295 3314 1439 3322
rect 1295 3313 1331 3314
rect 1403 3313 1439 3314
rect 1505 3347 1542 3348
rect 1505 3346 1543 3347
rect 1505 3338 1569 3346
rect 1505 3318 1514 3338
rect 1534 3324 1569 3338
rect 1589 3324 1592 3344
rect 1534 3319 1592 3324
rect 1534 3318 1569 3319
rect 771 3281 808 3310
rect 772 3279 808 3281
rect 984 3279 1021 3310
rect 772 3257 1021 3279
rect 853 3251 964 3257
rect 853 3243 894 3251
rect 853 3223 861 3243
rect 880 3223 894 3243
rect 853 3221 894 3223
rect 922 3243 964 3251
rect 922 3223 938 3243
rect 957 3223 964 3243
rect 922 3221 964 3223
rect 853 3206 964 3221
rect 1192 3211 1229 3310
rect 1505 3306 1569 3318
rect 855 3197 959 3206
rect 643 3166 764 3176
rect 643 3164 712 3166
rect 643 3123 656 3164
rect 693 3125 712 3164
rect 749 3125 764 3166
rect 693 3123 764 3125
rect 643 3105 764 3123
rect 436 3061 497 3073
rect 1190 3061 1231 3211
rect 1609 3203 1636 3458
rect 1698 3448 1778 3459
rect 1698 3422 1715 3448
rect 1755 3422 1778 3448
rect 1698 3395 1778 3422
rect 1698 3369 1719 3395
rect 1759 3369 1778 3395
rect 1698 3350 1778 3369
rect 1698 3324 1722 3350
rect 1762 3324 1778 3350
rect 1698 3273 1778 3324
rect 436 3058 1231 3061
rect 1610 3072 1636 3203
rect 1700 3117 1770 3273
rect 1699 3101 1775 3117
rect 1610 3058 1638 3072
rect 436 3023 1638 3058
rect 1699 3064 1714 3101
rect 1758 3064 1775 3101
rect 1699 3044 1775 3064
rect 2813 3094 2883 4003
rect 2982 3482 3063 4151
rect 3887 4046 3923 4346
rect 3811 4017 3924 4046
rect 3811 3652 3842 4017
rect 3735 3632 4128 3652
rect 4148 3632 4151 3652
rect 3735 3627 4151 3632
rect 3735 3626 4076 3627
rect 3392 3595 3502 3609
rect 3392 3592 3435 3595
rect 3392 3587 3396 3592
rect 3314 3565 3396 3587
rect 3425 3565 3435 3592
rect 3463 3568 3470 3595
rect 3499 3587 3502 3595
rect 3499 3568 3564 3587
rect 3463 3565 3564 3568
rect 3314 3563 3564 3565
rect 3314 3484 3351 3563
rect 3392 3550 3502 3563
rect 3466 3494 3497 3495
rect 2976 3402 3075 3482
rect 3314 3464 3323 3484
rect 3343 3464 3351 3484
rect 3314 3454 3351 3464
rect 3410 3484 3497 3494
rect 3410 3464 3419 3484
rect 3439 3464 3497 3484
rect 3410 3455 3497 3464
rect 3410 3454 3447 3455
rect 3466 3402 3497 3455
rect 3527 3484 3564 3563
rect 3679 3494 3710 3495
rect 3527 3464 3536 3484
rect 3556 3464 3564 3484
rect 3527 3454 3564 3464
rect 3623 3487 3710 3494
rect 3623 3484 3684 3487
rect 3623 3464 3632 3484
rect 3652 3467 3684 3484
rect 3705 3467 3710 3487
rect 3652 3464 3710 3467
rect 3623 3457 3710 3464
rect 3735 3484 3772 3626
rect 4038 3625 4075 3626
rect 3887 3494 3923 3495
rect 3735 3464 3744 3484
rect 3764 3464 3772 3484
rect 3623 3455 3679 3457
rect 3623 3454 3660 3455
rect 3735 3454 3772 3464
rect 3831 3484 3979 3494
rect 4079 3491 4175 3493
rect 3831 3464 3840 3484
rect 3860 3464 3950 3484
rect 3970 3464 3979 3484
rect 3831 3458 3979 3464
rect 3831 3455 3895 3458
rect 3831 3454 3868 3455
rect 3887 3428 3895 3455
rect 3916 3455 3979 3458
rect 4037 3484 4175 3491
rect 4037 3464 4046 3484
rect 4066 3464 4175 3484
rect 4037 3455 4175 3464
rect 3916 3428 3923 3455
rect 3942 3454 3979 3455
rect 4038 3454 4075 3455
rect 3887 3403 3923 3428
rect 2976 3401 3316 3402
rect 3358 3401 3399 3402
rect 2976 3394 3399 3401
rect 2976 3374 3368 3394
rect 3388 3374 3399 3394
rect 2976 3366 3399 3374
rect 3466 3398 3825 3402
rect 3466 3393 3788 3398
rect 3466 3369 3579 3393
rect 3603 3374 3788 3393
rect 3812 3374 3825 3398
rect 3603 3369 3825 3374
rect 3466 3366 3825 3369
rect 3887 3366 3922 3403
rect 3990 3400 4090 3403
rect 3990 3396 4057 3400
rect 3990 3370 4002 3396
rect 4028 3374 4057 3396
rect 4083 3374 4090 3400
rect 4028 3370 4090 3374
rect 3990 3366 4090 3370
rect 2976 3362 3316 3366
rect 2813 3044 2885 3094
rect 436 2948 497 3023
rect 855 3021 959 3023
rect 1190 3021 1231 3023
rect 1699 2978 1709 3044
rect 1763 2978 1775 3044
rect 1699 2954 1775 2978
rect 438 2818 497 2948
rect 1351 2899 1423 2900
rect 1350 2891 1449 2899
rect 1350 2888 1402 2891
rect 1350 2853 1358 2888
rect 1383 2853 1402 2888
rect 1427 2880 1449 2891
rect 1427 2879 2294 2880
rect 1427 2853 2295 2879
rect 1350 2843 2295 2853
rect 1350 2841 1449 2843
rect 438 2800 460 2818
rect 478 2800 497 2818
rect 438 2778 497 2800
rect 705 2814 1237 2819
rect 705 2794 1591 2814
rect 1611 2794 1614 2814
rect 2250 2810 2295 2843
rect 705 2790 1614 2794
rect 705 2743 748 2790
rect 1198 2789 1614 2790
rect 2246 2790 2639 2810
rect 2659 2790 2662 2810
rect 1198 2788 1539 2789
rect 855 2757 965 2771
rect 855 2754 898 2757
rect 855 2749 859 2754
rect 693 2742 748 2743
rect 437 2719 748 2742
rect 437 2701 462 2719
rect 480 2707 748 2719
rect 777 2727 859 2749
rect 888 2727 898 2754
rect 926 2730 933 2757
rect 962 2749 965 2757
rect 962 2730 1027 2749
rect 926 2727 1027 2730
rect 777 2725 1027 2727
rect 480 2701 502 2707
rect 437 2562 502 2701
rect 777 2646 814 2725
rect 855 2712 965 2725
rect 929 2656 960 2657
rect 777 2626 786 2646
rect 806 2626 814 2646
rect 437 2544 460 2562
rect 478 2544 502 2562
rect 437 2527 502 2544
rect 657 2608 725 2621
rect 777 2616 814 2626
rect 873 2646 960 2656
rect 873 2626 882 2646
rect 902 2626 960 2646
rect 873 2617 960 2626
rect 873 2616 910 2617
rect 657 2566 664 2608
rect 713 2566 725 2608
rect 657 2563 725 2566
rect 929 2564 960 2617
rect 990 2646 1027 2725
rect 1142 2656 1173 2657
rect 990 2626 999 2646
rect 1019 2626 1027 2646
rect 990 2616 1027 2626
rect 1086 2649 1173 2656
rect 1086 2646 1147 2649
rect 1086 2626 1095 2646
rect 1115 2629 1147 2646
rect 1168 2629 1173 2649
rect 1115 2626 1173 2629
rect 1086 2619 1173 2626
rect 1198 2646 1235 2788
rect 1501 2787 1538 2788
rect 2246 2785 2662 2790
rect 2246 2784 2587 2785
rect 1903 2753 2013 2767
rect 1903 2750 1946 2753
rect 1903 2745 1907 2750
rect 1825 2723 1907 2745
rect 1936 2723 1946 2750
rect 1974 2726 1981 2753
rect 2010 2745 2013 2753
rect 2010 2726 2075 2745
rect 1974 2723 2075 2726
rect 1825 2721 2075 2723
rect 1350 2656 1386 2657
rect 1198 2626 1207 2646
rect 1227 2626 1235 2646
rect 1086 2617 1142 2619
rect 1086 2616 1123 2617
rect 1198 2616 1235 2626
rect 1294 2646 1442 2656
rect 1542 2653 1638 2655
rect 1294 2626 1303 2646
rect 1323 2626 1413 2646
rect 1433 2626 1442 2646
rect 1294 2620 1442 2626
rect 1294 2617 1358 2620
rect 1294 2616 1331 2617
rect 1350 2590 1358 2617
rect 1379 2617 1442 2620
rect 1500 2646 1638 2653
rect 1500 2626 1509 2646
rect 1529 2626 1638 2646
rect 1500 2617 1638 2626
rect 1825 2642 1862 2721
rect 1903 2708 2013 2721
rect 1977 2652 2008 2653
rect 1825 2622 1834 2642
rect 1854 2622 1862 2642
rect 1379 2590 1386 2617
rect 1405 2616 1442 2617
rect 1501 2616 1538 2617
rect 1350 2565 1386 2590
rect 821 2563 862 2564
rect 657 2556 862 2563
rect 657 2545 831 2556
rect 657 2512 665 2545
rect 658 2503 665 2512
rect 714 2536 831 2545
rect 851 2536 862 2556
rect 714 2528 862 2536
rect 929 2560 1288 2564
rect 929 2555 1251 2560
rect 929 2531 1042 2555
rect 1066 2536 1251 2555
rect 1275 2536 1288 2560
rect 1066 2531 1288 2536
rect 929 2528 1288 2531
rect 1350 2528 1385 2565
rect 1453 2562 1553 2565
rect 1453 2558 1520 2562
rect 1453 2532 1465 2558
rect 1491 2536 1520 2558
rect 1546 2536 1553 2562
rect 1491 2532 1553 2536
rect 1453 2528 1553 2532
rect 714 2512 725 2528
rect 714 2503 722 2512
rect 929 2507 960 2528
rect 1350 2507 1386 2528
rect 772 2506 809 2507
rect 437 2463 502 2482
rect 437 2445 462 2463
rect 480 2445 502 2463
rect 437 2244 502 2445
rect 658 2319 722 2503
rect 771 2497 809 2506
rect 771 2477 780 2497
rect 800 2477 809 2497
rect 771 2469 809 2477
rect 875 2501 960 2507
rect 985 2506 1022 2507
rect 875 2481 883 2501
rect 903 2481 960 2501
rect 875 2473 960 2481
rect 984 2497 1022 2506
rect 984 2477 993 2497
rect 1013 2477 1022 2497
rect 875 2472 911 2473
rect 984 2469 1022 2477
rect 1088 2501 1173 2507
rect 1193 2506 1230 2507
rect 1088 2481 1096 2501
rect 1116 2500 1173 2501
rect 1116 2481 1145 2500
rect 1088 2480 1145 2481
rect 1166 2480 1173 2500
rect 1088 2473 1173 2480
rect 1192 2497 1230 2506
rect 1192 2477 1201 2497
rect 1221 2477 1230 2497
rect 1088 2472 1124 2473
rect 1192 2469 1230 2477
rect 1296 2501 1440 2507
rect 1296 2481 1304 2501
rect 1324 2481 1412 2501
rect 1432 2481 1440 2501
rect 1296 2473 1440 2481
rect 1296 2472 1332 2473
rect 1404 2472 1440 2473
rect 1506 2506 1543 2507
rect 1506 2505 1544 2506
rect 1506 2497 1570 2505
rect 1506 2477 1515 2497
rect 1535 2483 1570 2497
rect 1590 2483 1593 2503
rect 1535 2478 1593 2483
rect 1535 2477 1570 2478
rect 772 2440 809 2469
rect 773 2438 809 2440
rect 985 2438 1022 2469
rect 773 2416 1022 2438
rect 854 2410 965 2416
rect 854 2402 895 2410
rect 854 2382 862 2402
rect 881 2382 895 2402
rect 854 2380 895 2382
rect 923 2402 965 2410
rect 923 2382 939 2402
rect 958 2382 965 2402
rect 923 2380 965 2382
rect 854 2365 965 2380
rect 658 2309 726 2319
rect 658 2276 675 2309
rect 715 2276 726 2309
rect 658 2264 726 2276
rect 658 2262 722 2264
rect 1193 2245 1230 2469
rect 1506 2465 1570 2477
rect 1610 2247 1637 2617
rect 1825 2612 1862 2622
rect 1921 2642 2008 2652
rect 1921 2622 1930 2642
rect 1950 2622 2008 2642
rect 1921 2613 2008 2622
rect 1921 2612 1958 2613
rect 1701 2599 1771 2604
rect 1696 2593 1771 2599
rect 1696 2560 1704 2593
rect 1757 2560 1771 2593
rect 1977 2560 2008 2613
rect 2038 2642 2075 2721
rect 2190 2652 2221 2653
rect 2038 2622 2047 2642
rect 2067 2622 2075 2642
rect 2038 2612 2075 2622
rect 2134 2645 2221 2652
rect 2134 2642 2195 2645
rect 2134 2622 2143 2642
rect 2163 2625 2195 2642
rect 2216 2625 2221 2645
rect 2163 2622 2221 2625
rect 2134 2615 2221 2622
rect 2246 2642 2283 2784
rect 2549 2783 2586 2784
rect 2398 2652 2434 2653
rect 2246 2622 2255 2642
rect 2275 2622 2283 2642
rect 2134 2613 2190 2615
rect 2134 2612 2171 2613
rect 2246 2612 2283 2622
rect 2342 2642 2490 2652
rect 2590 2649 2686 2651
rect 2342 2622 2351 2642
rect 2371 2622 2461 2642
rect 2481 2622 2490 2642
rect 2342 2616 2490 2622
rect 2342 2613 2406 2616
rect 2342 2612 2379 2613
rect 2398 2586 2406 2613
rect 2427 2613 2490 2616
rect 2548 2642 2686 2649
rect 2548 2622 2557 2642
rect 2577 2622 2686 2642
rect 2548 2613 2686 2622
rect 2427 2586 2434 2613
rect 2453 2612 2490 2613
rect 2549 2612 2586 2613
rect 2398 2561 2434 2586
rect 1696 2559 1779 2560
rect 1869 2559 1910 2560
rect 1696 2552 1910 2559
rect 1696 2535 1879 2552
rect 1696 2502 1709 2535
rect 1762 2532 1879 2535
rect 1899 2532 1910 2552
rect 1762 2524 1910 2532
rect 1977 2556 2336 2560
rect 1977 2551 2299 2556
rect 1977 2527 2090 2551
rect 2114 2532 2299 2551
rect 2323 2532 2336 2556
rect 2114 2527 2336 2532
rect 1977 2524 2336 2527
rect 2398 2524 2433 2561
rect 2501 2558 2601 2561
rect 2501 2554 2568 2558
rect 2501 2528 2513 2554
rect 2539 2532 2568 2554
rect 2594 2532 2601 2558
rect 2539 2528 2601 2532
rect 2501 2524 2601 2528
rect 1762 2502 1779 2524
rect 1977 2503 2008 2524
rect 2398 2503 2434 2524
rect 1820 2502 1857 2503
rect 1696 2488 1779 2502
rect 1469 2245 1637 2247
rect 1193 2244 1637 2245
rect 437 2214 1637 2244
rect 1707 2278 1779 2488
rect 1819 2493 1857 2502
rect 1819 2473 1828 2493
rect 1848 2473 1857 2493
rect 1819 2465 1857 2473
rect 1923 2497 2008 2503
rect 2033 2502 2070 2503
rect 1923 2477 1931 2497
rect 1951 2477 2008 2497
rect 1923 2469 2008 2477
rect 2032 2493 2070 2502
rect 2032 2473 2041 2493
rect 2061 2473 2070 2493
rect 1923 2468 1959 2469
rect 2032 2465 2070 2473
rect 2136 2497 2221 2503
rect 2241 2502 2278 2503
rect 2136 2477 2144 2497
rect 2164 2496 2221 2497
rect 2164 2477 2193 2496
rect 2136 2476 2193 2477
rect 2214 2476 2221 2496
rect 2136 2469 2221 2476
rect 2240 2493 2278 2502
rect 2240 2473 2249 2493
rect 2269 2473 2278 2493
rect 2136 2468 2172 2469
rect 2240 2465 2278 2473
rect 2344 2497 2488 2503
rect 2344 2477 2352 2497
rect 2372 2477 2460 2497
rect 2480 2477 2488 2497
rect 2344 2469 2488 2477
rect 2344 2468 2380 2469
rect 2452 2468 2488 2469
rect 2554 2502 2591 2503
rect 2554 2501 2592 2502
rect 2554 2493 2618 2501
rect 2554 2473 2563 2493
rect 2583 2479 2618 2493
rect 2638 2479 2641 2499
rect 2583 2474 2641 2479
rect 2583 2473 2618 2474
rect 1820 2436 1857 2465
rect 1821 2434 1857 2436
rect 2033 2434 2070 2465
rect 1821 2412 2070 2434
rect 1902 2406 2013 2412
rect 1902 2398 1943 2406
rect 1902 2378 1910 2398
rect 1929 2378 1943 2398
rect 1902 2376 1943 2378
rect 1971 2398 2013 2406
rect 1971 2378 1987 2398
rect 2006 2378 2013 2398
rect 1971 2376 2013 2378
rect 1902 2361 2013 2376
rect 1707 2239 1726 2278
rect 1771 2239 1779 2278
rect 1707 2222 1779 2239
rect 2241 2266 2278 2465
rect 2554 2461 2618 2473
rect 2241 2260 2282 2266
rect 2658 2262 2685 2613
rect 2814 2565 2885 3044
rect 2814 2481 2883 2565
rect 2517 2260 2685 2262
rect 2241 2234 2685 2260
rect 437 2167 502 2214
rect 437 2149 460 2167
rect 478 2149 502 2167
rect 1350 2194 1385 2196
rect 1350 2192 1454 2194
rect 2243 2192 2282 2234
rect 2517 2233 2685 2234
rect 1350 2185 2284 2192
rect 1350 2184 1401 2185
rect 1350 2164 1353 2184
rect 1378 2165 1401 2184
rect 1433 2165 2284 2185
rect 1378 2164 2284 2165
rect 1350 2157 2284 2164
rect 1623 2156 2284 2157
rect 437 2128 502 2149
rect 714 2139 754 2142
rect 714 2135 1617 2139
rect 714 2115 1591 2135
rect 1611 2115 1617 2135
rect 714 2112 1617 2115
rect 438 2068 503 2088
rect 438 2050 462 2068
rect 480 2050 503 2068
rect 438 2023 503 2050
rect 714 2023 754 2112
rect 1198 2110 1614 2112
rect 1198 2109 1539 2110
rect 855 2078 965 2092
rect 855 2075 898 2078
rect 855 2070 859 2075
rect 437 1988 754 2023
rect 777 2048 859 2070
rect 888 2048 898 2075
rect 926 2051 933 2078
rect 962 2070 965 2078
rect 962 2051 1027 2070
rect 926 2048 1027 2051
rect 777 2046 1027 2048
rect 438 1912 503 1988
rect 777 1967 814 2046
rect 855 2033 965 2046
rect 929 1977 960 1978
rect 777 1947 786 1967
rect 806 1947 814 1967
rect 777 1937 814 1947
rect 873 1967 960 1977
rect 873 1947 882 1967
rect 902 1947 960 1967
rect 873 1938 960 1947
rect 873 1937 910 1938
rect 438 1894 460 1912
rect 478 1894 503 1912
rect 438 1873 503 1894
rect 651 1892 716 1901
rect 651 1855 661 1892
rect 701 1884 716 1892
rect 929 1885 960 1938
rect 990 1967 1027 2046
rect 1142 1977 1173 1978
rect 990 1947 999 1967
rect 1019 1947 1027 1967
rect 990 1937 1027 1947
rect 1086 1970 1173 1977
rect 1086 1967 1147 1970
rect 1086 1947 1095 1967
rect 1115 1950 1147 1967
rect 1168 1950 1173 1970
rect 1115 1947 1173 1950
rect 1086 1940 1173 1947
rect 1198 1967 1235 2109
rect 1501 2108 1538 2109
rect 1350 1977 1386 1978
rect 1198 1947 1207 1967
rect 1227 1947 1235 1967
rect 1086 1938 1142 1940
rect 1086 1937 1123 1938
rect 1198 1937 1235 1947
rect 1294 1967 1442 1977
rect 1542 1974 1638 1976
rect 1294 1947 1303 1967
rect 1323 1947 1413 1967
rect 1433 1947 1442 1967
rect 1294 1941 1442 1947
rect 1294 1938 1358 1941
rect 1294 1937 1331 1938
rect 1350 1911 1358 1938
rect 1379 1938 1442 1941
rect 1500 1967 1638 1974
rect 2818 1969 2880 2481
rect 1500 1947 1509 1967
rect 1529 1947 1638 1967
rect 1500 1938 1638 1947
rect 1379 1911 1386 1938
rect 1405 1937 1442 1938
rect 1501 1937 1538 1938
rect 1350 1886 1386 1911
rect 821 1884 862 1885
rect 701 1877 862 1884
rect 701 1857 831 1877
rect 851 1857 862 1877
rect 701 1855 862 1857
rect 651 1849 862 1855
rect 929 1881 1288 1885
rect 929 1876 1251 1881
rect 929 1852 1042 1876
rect 1066 1857 1251 1876
rect 1275 1857 1288 1881
rect 1066 1852 1288 1857
rect 929 1849 1288 1852
rect 1350 1849 1385 1886
rect 1453 1883 1553 1886
rect 1453 1879 1520 1883
rect 1453 1853 1465 1879
rect 1491 1857 1520 1879
rect 1546 1857 1553 1883
rect 1491 1853 1553 1857
rect 1453 1849 1553 1853
rect 651 1836 718 1849
rect 443 1813 499 1833
rect 443 1795 462 1813
rect 480 1795 499 1813
rect 443 1682 499 1795
rect 651 1815 665 1836
rect 701 1815 718 1836
rect 929 1828 960 1849
rect 1350 1828 1386 1849
rect 772 1827 809 1828
rect 651 1808 718 1815
rect 771 1818 809 1827
rect 443 1544 498 1682
rect 651 1656 716 1808
rect 771 1798 780 1818
rect 800 1798 809 1818
rect 771 1790 809 1798
rect 875 1822 960 1828
rect 985 1827 1022 1828
rect 875 1802 883 1822
rect 903 1802 960 1822
rect 875 1794 960 1802
rect 984 1818 1022 1827
rect 984 1798 993 1818
rect 1013 1798 1022 1818
rect 875 1793 911 1794
rect 984 1790 1022 1798
rect 1088 1822 1173 1828
rect 1193 1827 1230 1828
rect 1088 1802 1096 1822
rect 1116 1821 1173 1822
rect 1116 1802 1145 1821
rect 1088 1801 1145 1802
rect 1166 1801 1173 1821
rect 1088 1794 1173 1801
rect 1192 1818 1230 1827
rect 1192 1798 1201 1818
rect 1221 1798 1230 1818
rect 1088 1793 1124 1794
rect 1192 1790 1230 1798
rect 1296 1822 1440 1828
rect 1296 1802 1304 1822
rect 1324 1802 1412 1822
rect 1432 1802 1440 1822
rect 1296 1794 1440 1802
rect 1296 1793 1332 1794
rect 1404 1793 1440 1794
rect 1506 1827 1543 1828
rect 1506 1826 1544 1827
rect 1506 1818 1570 1826
rect 1506 1798 1515 1818
rect 1535 1804 1570 1818
rect 1590 1804 1593 1824
rect 1535 1799 1593 1804
rect 1535 1798 1570 1799
rect 772 1761 809 1790
rect 773 1759 809 1761
rect 985 1759 1022 1790
rect 773 1737 1022 1759
rect 854 1731 965 1737
rect 854 1723 895 1731
rect 854 1703 862 1723
rect 881 1703 895 1723
rect 854 1701 895 1703
rect 923 1723 965 1731
rect 923 1703 939 1723
rect 958 1703 965 1723
rect 923 1701 965 1703
rect 854 1688 965 1701
rect 1193 1691 1230 1790
rect 1506 1786 1570 1798
rect 644 1646 765 1656
rect 644 1644 713 1646
rect 644 1603 657 1644
rect 694 1605 713 1644
rect 750 1605 765 1646
rect 694 1603 765 1605
rect 644 1585 765 1603
rect 436 1541 500 1544
rect 856 1541 960 1547
rect 1191 1541 1232 1691
rect 1610 1683 1637 1938
rect 1699 1928 1779 1939
rect 1699 1902 1716 1928
rect 1756 1902 1779 1928
rect 1699 1875 1779 1902
rect 2822 1930 2880 1969
rect 2822 1895 2884 1930
rect 1699 1849 1720 1875
rect 1760 1849 1779 1875
rect 1699 1830 1779 1849
rect 1699 1804 1723 1830
rect 1763 1804 1779 1830
rect 1699 1753 1779 1804
rect 2771 1868 2884 1895
rect 2771 1866 2830 1868
rect 2771 1835 2785 1866
rect 2810 1845 2830 1866
rect 2856 1845 2884 1868
rect 2810 1835 2884 1845
rect 2771 1825 2884 1835
rect 436 1538 1232 1541
rect 1611 1552 1637 1683
rect 1611 1538 1639 1552
rect 436 1503 1639 1538
rect 1701 1545 1771 1753
rect 436 1442 500 1503
rect 856 1501 960 1503
rect 1191 1501 1232 1503
rect 1701 1500 1722 1545
rect 1702 1479 1722 1500
rect 1752 1500 1771 1545
rect 1752 1479 1769 1500
rect 1702 1460 1769 1479
rect 1351 1452 1423 1453
rect 1350 1444 1449 1452
rect 438 1371 497 1442
rect 1350 1441 1402 1444
rect 1350 1406 1358 1441
rect 1383 1406 1402 1441
rect 1427 1433 1449 1444
rect 1427 1432 2294 1433
rect 1427 1406 2295 1432
rect 1350 1396 2295 1406
rect 1350 1394 1449 1396
rect 438 1353 460 1371
rect 478 1353 497 1371
rect 438 1331 497 1353
rect 705 1367 1237 1372
rect 705 1347 1591 1367
rect 1611 1347 1614 1367
rect 2250 1363 2295 1396
rect 705 1343 1614 1347
rect 705 1296 748 1343
rect 1198 1342 1614 1343
rect 2246 1343 2639 1363
rect 2659 1343 2662 1363
rect 1198 1341 1539 1342
rect 855 1310 965 1324
rect 855 1307 898 1310
rect 855 1302 859 1307
rect 693 1295 748 1296
rect 437 1272 748 1295
rect 437 1254 462 1272
rect 480 1260 748 1272
rect 777 1280 859 1302
rect 888 1280 898 1307
rect 926 1283 933 1310
rect 962 1302 965 1310
rect 962 1283 1027 1302
rect 926 1280 1027 1283
rect 777 1278 1027 1280
rect 480 1254 502 1260
rect 437 1115 502 1254
rect 777 1199 814 1278
rect 855 1265 965 1278
rect 929 1209 960 1210
rect 777 1179 786 1199
rect 806 1179 814 1199
rect 437 1097 460 1115
rect 478 1097 502 1115
rect 437 1080 502 1097
rect 657 1161 725 1174
rect 777 1169 814 1179
rect 873 1199 960 1209
rect 873 1179 882 1199
rect 902 1179 960 1199
rect 873 1170 960 1179
rect 873 1169 910 1170
rect 657 1119 664 1161
rect 713 1119 725 1161
rect 657 1116 725 1119
rect 929 1117 960 1170
rect 990 1199 1027 1278
rect 1142 1209 1173 1210
rect 990 1179 999 1199
rect 1019 1179 1027 1199
rect 990 1169 1027 1179
rect 1086 1202 1173 1209
rect 1086 1199 1147 1202
rect 1086 1179 1095 1199
rect 1115 1182 1147 1199
rect 1168 1182 1173 1202
rect 1115 1179 1173 1182
rect 1086 1172 1173 1179
rect 1198 1199 1235 1341
rect 1501 1340 1538 1341
rect 2246 1338 2662 1343
rect 2246 1337 2587 1338
rect 1903 1306 2013 1320
rect 1903 1303 1946 1306
rect 1903 1298 1907 1303
rect 1825 1276 1907 1298
rect 1936 1276 1946 1303
rect 1974 1279 1981 1306
rect 2010 1298 2013 1306
rect 2010 1279 2075 1298
rect 1974 1276 2075 1279
rect 1825 1274 2075 1276
rect 1350 1209 1386 1210
rect 1198 1179 1207 1199
rect 1227 1179 1235 1199
rect 1086 1170 1142 1172
rect 1086 1169 1123 1170
rect 1198 1169 1235 1179
rect 1294 1199 1442 1209
rect 1542 1206 1638 1208
rect 1294 1179 1303 1199
rect 1323 1179 1413 1199
rect 1433 1179 1442 1199
rect 1294 1173 1442 1179
rect 1294 1170 1358 1173
rect 1294 1169 1331 1170
rect 1350 1143 1358 1170
rect 1379 1170 1442 1173
rect 1500 1199 1638 1206
rect 1500 1179 1509 1199
rect 1529 1179 1638 1199
rect 1500 1170 1638 1179
rect 1825 1195 1862 1274
rect 1903 1261 2013 1274
rect 1977 1205 2008 1206
rect 1825 1175 1834 1195
rect 1854 1175 1862 1195
rect 1379 1143 1386 1170
rect 1405 1169 1442 1170
rect 1501 1169 1538 1170
rect 1350 1118 1386 1143
rect 821 1116 862 1117
rect 657 1109 862 1116
rect 657 1098 831 1109
rect 657 1065 665 1098
rect 658 1056 665 1065
rect 714 1089 831 1098
rect 851 1089 862 1109
rect 714 1081 862 1089
rect 929 1113 1288 1117
rect 929 1108 1251 1113
rect 929 1084 1042 1108
rect 1066 1089 1251 1108
rect 1275 1089 1288 1113
rect 1066 1084 1288 1089
rect 929 1081 1288 1084
rect 1350 1081 1385 1118
rect 1453 1115 1553 1118
rect 1453 1111 1520 1115
rect 1453 1085 1465 1111
rect 1491 1089 1520 1111
rect 1546 1089 1553 1115
rect 1491 1085 1553 1089
rect 1453 1081 1553 1085
rect 714 1065 725 1081
rect 714 1056 722 1065
rect 929 1060 960 1081
rect 1350 1060 1386 1081
rect 772 1059 809 1060
rect 437 1016 502 1035
rect 437 998 462 1016
rect 480 998 502 1016
rect 437 797 502 998
rect 658 872 722 1056
rect 771 1050 809 1059
rect 771 1030 780 1050
rect 800 1030 809 1050
rect 771 1022 809 1030
rect 875 1054 960 1060
rect 985 1059 1022 1060
rect 875 1034 883 1054
rect 903 1034 960 1054
rect 875 1026 960 1034
rect 984 1050 1022 1059
rect 984 1030 993 1050
rect 1013 1030 1022 1050
rect 875 1025 911 1026
rect 984 1022 1022 1030
rect 1088 1054 1173 1060
rect 1193 1059 1230 1060
rect 1088 1034 1096 1054
rect 1116 1053 1173 1054
rect 1116 1034 1145 1053
rect 1088 1033 1145 1034
rect 1166 1033 1173 1053
rect 1088 1026 1173 1033
rect 1192 1050 1230 1059
rect 1192 1030 1201 1050
rect 1221 1030 1230 1050
rect 1088 1025 1124 1026
rect 1192 1022 1230 1030
rect 1296 1054 1440 1060
rect 1296 1034 1304 1054
rect 1324 1034 1412 1054
rect 1432 1034 1440 1054
rect 1296 1026 1440 1034
rect 1296 1025 1332 1026
rect 1404 1025 1440 1026
rect 1506 1059 1543 1060
rect 1506 1058 1544 1059
rect 1506 1050 1570 1058
rect 1506 1030 1515 1050
rect 1535 1036 1570 1050
rect 1590 1036 1593 1056
rect 1535 1031 1593 1036
rect 1535 1030 1570 1031
rect 772 993 809 1022
rect 773 991 809 993
rect 985 991 1022 1022
rect 773 969 1022 991
rect 854 963 965 969
rect 854 955 895 963
rect 854 935 862 955
rect 881 935 895 955
rect 854 933 895 935
rect 923 955 965 963
rect 923 935 939 955
rect 958 935 965 955
rect 923 933 965 935
rect 854 918 965 933
rect 658 862 726 872
rect 658 829 675 862
rect 715 829 726 862
rect 658 817 726 829
rect 658 815 722 817
rect 1193 798 1230 1022
rect 1506 1018 1570 1030
rect 1610 800 1637 1170
rect 1825 1165 1862 1175
rect 1921 1195 2008 1205
rect 1921 1175 1930 1195
rect 1950 1175 2008 1195
rect 1921 1166 2008 1175
rect 1921 1165 1958 1166
rect 1701 1152 1771 1157
rect 1696 1146 1771 1152
rect 1696 1113 1704 1146
rect 1757 1113 1771 1146
rect 1977 1113 2008 1166
rect 2038 1195 2075 1274
rect 2190 1205 2221 1206
rect 2038 1175 2047 1195
rect 2067 1175 2075 1195
rect 2038 1165 2075 1175
rect 2134 1198 2221 1205
rect 2134 1195 2195 1198
rect 2134 1175 2143 1195
rect 2163 1178 2195 1195
rect 2216 1178 2221 1198
rect 2163 1175 2221 1178
rect 2134 1168 2221 1175
rect 2246 1195 2283 1337
rect 2549 1336 2586 1337
rect 2398 1205 2434 1206
rect 2246 1175 2255 1195
rect 2275 1175 2283 1195
rect 2134 1166 2190 1168
rect 2134 1165 2171 1166
rect 2246 1165 2283 1175
rect 2342 1195 2490 1205
rect 2590 1202 2686 1204
rect 2342 1175 2351 1195
rect 2371 1175 2461 1195
rect 2481 1175 2490 1195
rect 2342 1169 2490 1175
rect 2342 1166 2406 1169
rect 2342 1165 2379 1166
rect 2398 1139 2406 1166
rect 2427 1166 2490 1169
rect 2548 1195 2686 1202
rect 2548 1175 2557 1195
rect 2577 1175 2686 1195
rect 2548 1166 2686 1175
rect 2427 1139 2434 1166
rect 2453 1165 2490 1166
rect 2549 1165 2586 1166
rect 2398 1114 2434 1139
rect 1696 1112 1779 1113
rect 1869 1112 1910 1113
rect 1696 1105 1910 1112
rect 1696 1088 1879 1105
rect 1696 1055 1709 1088
rect 1762 1085 1879 1088
rect 1899 1085 1910 1105
rect 1762 1077 1910 1085
rect 1977 1109 2336 1113
rect 1977 1104 2299 1109
rect 1977 1080 2090 1104
rect 2114 1085 2299 1104
rect 2323 1085 2336 1109
rect 2114 1080 2336 1085
rect 1977 1077 2336 1080
rect 2398 1077 2433 1114
rect 2501 1111 2601 1114
rect 2501 1107 2568 1111
rect 2501 1081 2513 1107
rect 2539 1085 2568 1107
rect 2594 1085 2601 1111
rect 2539 1081 2601 1085
rect 2501 1077 2601 1081
rect 1762 1055 1779 1077
rect 1977 1056 2008 1077
rect 2398 1056 2434 1077
rect 1820 1055 1857 1056
rect 1696 1041 1779 1055
rect 1469 798 1637 800
rect 1193 797 1637 798
rect 437 767 1637 797
rect 1707 831 1779 1041
rect 1819 1046 1857 1055
rect 1819 1026 1828 1046
rect 1848 1026 1857 1046
rect 1819 1018 1857 1026
rect 1923 1050 2008 1056
rect 2033 1055 2070 1056
rect 1923 1030 1931 1050
rect 1951 1030 2008 1050
rect 1923 1022 2008 1030
rect 2032 1046 2070 1055
rect 2032 1026 2041 1046
rect 2061 1026 2070 1046
rect 1923 1021 1959 1022
rect 2032 1018 2070 1026
rect 2136 1050 2221 1056
rect 2241 1055 2278 1056
rect 2136 1030 2144 1050
rect 2164 1049 2221 1050
rect 2164 1030 2193 1049
rect 2136 1029 2193 1030
rect 2214 1029 2221 1049
rect 2136 1022 2221 1029
rect 2240 1046 2278 1055
rect 2240 1026 2249 1046
rect 2269 1026 2278 1046
rect 2136 1021 2172 1022
rect 2240 1018 2278 1026
rect 2344 1050 2488 1056
rect 2344 1030 2352 1050
rect 2372 1030 2460 1050
rect 2480 1030 2488 1050
rect 2344 1022 2488 1030
rect 2344 1021 2380 1022
rect 2452 1021 2488 1022
rect 2554 1055 2591 1056
rect 2554 1054 2592 1055
rect 2554 1046 2618 1054
rect 2554 1026 2563 1046
rect 2583 1032 2618 1046
rect 2638 1032 2641 1052
rect 2583 1027 2641 1032
rect 2583 1026 2618 1027
rect 1820 989 1857 1018
rect 1821 987 1857 989
rect 2033 987 2070 1018
rect 1821 965 2070 987
rect 1902 959 2013 965
rect 1902 951 1943 959
rect 1902 931 1910 951
rect 1929 931 1943 951
rect 1902 929 1943 931
rect 1971 951 2013 959
rect 1971 931 1987 951
rect 2006 931 2013 951
rect 1971 929 2013 931
rect 1902 914 2013 929
rect 1707 792 1726 831
rect 1771 792 1779 831
rect 1707 775 1779 792
rect 2241 819 2278 1018
rect 2554 1014 2618 1026
rect 2241 813 2282 819
rect 2658 815 2685 1166
rect 2517 813 2685 815
rect 2241 787 2685 813
rect 437 720 502 767
rect 437 702 460 720
rect 478 702 502 720
rect 1350 747 1385 749
rect 1350 745 1454 747
rect 2243 745 2282 787
rect 2517 786 2685 787
rect 1350 738 2284 745
rect 1350 737 1401 738
rect 1350 717 1353 737
rect 1378 718 1401 737
rect 1433 718 2284 738
rect 1378 717 2284 718
rect 1350 710 2284 717
rect 1623 709 2284 710
rect 437 681 502 702
rect 714 692 754 695
rect 714 688 1617 692
rect 714 668 1591 688
rect 1611 668 1617 688
rect 714 665 1617 668
rect 438 621 503 641
rect 438 603 462 621
rect 480 603 503 621
rect 438 576 503 603
rect 714 576 754 665
rect 1198 663 1614 665
rect 1198 662 1539 663
rect 855 631 965 645
rect 855 628 898 631
rect 855 623 859 628
rect 437 541 754 576
rect 777 601 859 623
rect 888 601 898 628
rect 926 604 933 631
rect 962 623 965 631
rect 962 604 1027 623
rect 926 601 1027 604
rect 777 599 1027 601
rect 438 465 503 541
rect 777 520 814 599
rect 855 586 965 599
rect 929 530 960 531
rect 777 500 786 520
rect 806 500 814 520
rect 777 490 814 500
rect 873 520 960 530
rect 873 500 882 520
rect 902 500 960 520
rect 873 491 960 500
rect 873 490 910 491
rect 438 447 460 465
rect 478 447 503 465
rect 438 426 503 447
rect 651 445 716 454
rect 651 408 661 445
rect 701 437 716 445
rect 929 438 960 491
rect 990 520 1027 599
rect 1142 530 1173 531
rect 990 500 999 520
rect 1019 500 1027 520
rect 990 490 1027 500
rect 1086 523 1173 530
rect 1086 520 1147 523
rect 1086 500 1095 520
rect 1115 503 1147 520
rect 1168 503 1173 523
rect 1115 500 1173 503
rect 1086 493 1173 500
rect 1198 520 1235 662
rect 1501 661 1538 662
rect 1350 530 1386 531
rect 1198 500 1207 520
rect 1227 500 1235 520
rect 1086 491 1142 493
rect 1086 490 1123 491
rect 1198 490 1235 500
rect 1294 520 1442 530
rect 1542 527 1638 529
rect 1294 500 1303 520
rect 1323 500 1413 520
rect 1433 500 1442 520
rect 1294 494 1442 500
rect 1294 491 1358 494
rect 1294 490 1331 491
rect 1350 464 1358 491
rect 1379 491 1442 494
rect 1500 520 1638 527
rect 1500 500 1509 520
rect 1529 500 1638 520
rect 1500 491 1638 500
rect 1379 464 1386 491
rect 1405 490 1442 491
rect 1501 490 1538 491
rect 1350 439 1386 464
rect 821 437 862 438
rect 701 430 862 437
rect 701 410 831 430
rect 851 410 862 430
rect 701 408 862 410
rect 651 402 862 408
rect 929 434 1288 438
rect 929 429 1251 434
rect 929 405 1042 429
rect 1066 410 1251 429
rect 1275 410 1288 434
rect 1066 405 1288 410
rect 929 402 1288 405
rect 1350 402 1385 439
rect 1453 436 1553 439
rect 1453 432 1520 436
rect 1453 406 1465 432
rect 1491 410 1520 432
rect 1546 410 1553 436
rect 1491 406 1553 410
rect 1453 402 1553 406
rect 651 389 718 402
rect 443 366 499 386
rect 443 348 462 366
rect 480 348 499 366
rect 443 313 499 348
rect 405 235 499 313
rect 651 368 665 389
rect 701 368 718 389
rect 929 381 960 402
rect 1350 381 1386 402
rect 772 380 809 381
rect 651 361 718 368
rect 771 371 809 380
rect 405 94 498 235
rect 651 209 716 361
rect 771 351 780 371
rect 800 351 809 371
rect 771 343 809 351
rect 875 375 960 381
rect 985 380 1022 381
rect 875 355 883 375
rect 903 355 960 375
rect 875 347 960 355
rect 984 371 1022 380
rect 984 351 993 371
rect 1013 351 1022 371
rect 875 346 911 347
rect 984 343 1022 351
rect 1088 375 1173 381
rect 1193 380 1230 381
rect 1088 355 1096 375
rect 1116 374 1173 375
rect 1116 355 1145 374
rect 1088 354 1145 355
rect 1166 354 1173 374
rect 1088 347 1173 354
rect 1192 371 1230 380
rect 1192 351 1201 371
rect 1221 351 1230 371
rect 1088 346 1124 347
rect 1192 343 1230 351
rect 1296 375 1440 381
rect 1296 355 1304 375
rect 1324 355 1412 375
rect 1432 355 1440 375
rect 1296 347 1440 355
rect 1296 346 1332 347
rect 1404 346 1440 347
rect 1506 380 1543 381
rect 1506 379 1544 380
rect 1506 371 1570 379
rect 1506 351 1515 371
rect 1535 357 1570 371
rect 1590 357 1593 377
rect 1535 352 1593 357
rect 1535 351 1570 352
rect 772 314 809 343
rect 773 312 809 314
rect 985 312 1022 343
rect 773 290 1022 312
rect 854 284 965 290
rect 854 276 895 284
rect 854 256 862 276
rect 881 256 895 276
rect 854 254 895 256
rect 923 276 965 284
rect 923 256 939 276
rect 958 256 965 276
rect 923 254 965 256
rect 854 239 965 254
rect 1193 244 1230 343
rect 1506 339 1570 351
rect 1610 300 1637 491
rect 856 230 960 239
rect 644 199 765 209
rect 644 197 713 199
rect 644 156 657 197
rect 694 158 713 197
rect 750 158 765 199
rect 694 156 765 158
rect 644 138 765 156
rect 856 94 960 103
rect 1191 94 1232 244
rect 405 92 1232 94
rect 413 91 1232 92
rect 1611 210 1636 300
rect 2771 268 2870 1825
rect 2976 461 3075 3362
rect 3466 3345 3497 3366
rect 3887 3345 3923 3366
rect 3309 3344 3346 3345
rect 3308 3335 3346 3344
rect 3308 3315 3317 3335
rect 3337 3315 3346 3335
rect 3308 3307 3346 3315
rect 3412 3339 3497 3345
rect 3522 3344 3559 3345
rect 3412 3319 3420 3339
rect 3440 3319 3497 3339
rect 3412 3311 3497 3319
rect 3521 3335 3559 3344
rect 3521 3315 3530 3335
rect 3550 3315 3559 3335
rect 3412 3310 3448 3311
rect 3521 3307 3559 3315
rect 3625 3339 3710 3345
rect 3730 3344 3767 3345
rect 3625 3319 3633 3339
rect 3653 3338 3710 3339
rect 3653 3319 3682 3338
rect 3625 3318 3682 3319
rect 3703 3318 3710 3338
rect 3625 3311 3710 3318
rect 3729 3335 3767 3344
rect 3729 3315 3738 3335
rect 3758 3315 3767 3335
rect 3625 3310 3661 3311
rect 3729 3307 3767 3315
rect 3833 3339 3977 3345
rect 3833 3319 3841 3339
rect 3861 3319 3949 3339
rect 3969 3319 3977 3339
rect 3833 3311 3977 3319
rect 3833 3310 3869 3311
rect 3941 3310 3977 3311
rect 4043 3344 4080 3345
rect 4043 3343 4081 3344
rect 4043 3335 4107 3343
rect 4043 3315 4052 3335
rect 4072 3321 4107 3335
rect 4127 3321 4130 3341
rect 4072 3316 4130 3321
rect 4072 3315 4107 3316
rect 3309 3278 3346 3307
rect 3310 3276 3346 3278
rect 3522 3276 3559 3307
rect 3310 3254 3559 3276
rect 3391 3248 3502 3254
rect 3391 3240 3432 3248
rect 3391 3220 3399 3240
rect 3418 3220 3432 3240
rect 3391 3218 3432 3220
rect 3460 3240 3502 3248
rect 3460 3220 3476 3240
rect 3495 3220 3502 3240
rect 3460 3218 3502 3220
rect 3391 3203 3502 3218
rect 3730 3186 3767 3307
rect 4043 3303 4107 3315
rect 3848 3186 3877 3190
rect 4147 3188 4174 3455
rect 4006 3186 4174 3188
rect 3730 3160 4174 3186
rect 3689 2892 3734 2901
rect 3689 2854 3699 2892
rect 3724 2854 3734 2892
rect 3689 2843 3734 2854
rect 3692 2835 3734 2843
rect 3692 2130 3735 2835
rect 3848 2221 3877 3160
rect 4006 3159 4174 3160
rect 4578 3010 4662 3014
rect 5130 3010 5218 5861
rect 5757 5848 5812 5860
rect 5757 5814 5775 5848
rect 5804 5814 5812 5848
rect 5757 5788 5812 5814
rect 5364 5755 5532 5756
rect 5757 5755 5774 5788
rect 5364 5754 5774 5755
rect 5803 5754 5812 5788
rect 5364 5729 5812 5754
rect 5364 5727 5532 5729
rect 5364 5460 5391 5727
rect 5757 5723 5812 5729
rect 5431 5600 5495 5612
rect 5771 5608 5808 5723
rect 6036 5697 6147 5712
rect 6036 5695 6078 5697
rect 6036 5675 6043 5695
rect 6062 5675 6078 5695
rect 6036 5667 6078 5675
rect 6106 5695 6147 5697
rect 6106 5675 6120 5695
rect 6139 5675 6147 5695
rect 6106 5667 6147 5675
rect 6036 5661 6147 5667
rect 5979 5639 6228 5661
rect 5979 5608 6016 5639
rect 6192 5637 6228 5639
rect 6192 5608 6229 5637
rect 5431 5599 5466 5600
rect 5408 5594 5466 5599
rect 5408 5574 5411 5594
rect 5431 5580 5466 5594
rect 5486 5580 5495 5600
rect 5431 5572 5495 5580
rect 5457 5571 5495 5572
rect 5458 5570 5495 5571
rect 5561 5604 5597 5605
rect 5669 5604 5705 5605
rect 5561 5596 5705 5604
rect 5561 5576 5569 5596
rect 5589 5576 5677 5596
rect 5697 5576 5705 5596
rect 5561 5570 5705 5576
rect 5771 5600 5809 5608
rect 5877 5604 5913 5605
rect 5771 5580 5780 5600
rect 5800 5580 5809 5600
rect 5771 5571 5809 5580
rect 5828 5597 5913 5604
rect 5828 5577 5835 5597
rect 5856 5596 5913 5597
rect 5856 5577 5885 5596
rect 5828 5576 5885 5577
rect 5905 5576 5913 5596
rect 5771 5570 5808 5571
rect 5828 5570 5913 5576
rect 5979 5600 6017 5608
rect 6090 5604 6126 5605
rect 5979 5580 5988 5600
rect 6008 5580 6017 5600
rect 5979 5571 6017 5580
rect 6041 5596 6126 5604
rect 6041 5576 6098 5596
rect 6118 5576 6126 5596
rect 5979 5570 6016 5571
rect 6041 5570 6126 5576
rect 6192 5600 6230 5608
rect 6192 5580 6201 5600
rect 6221 5580 6230 5600
rect 6192 5571 6230 5580
rect 6192 5570 6229 5571
rect 5615 5549 5651 5570
rect 6041 5549 6072 5570
rect 6286 5553 6357 6206
rect 6872 6140 6915 6853
rect 7532 6764 7627 6784
rect 7532 6720 7552 6764
rect 7612 6720 7627 6764
rect 7532 6424 7627 6720
rect 7532 6383 7565 6424
rect 7601 6383 7627 6424
rect 7727 6463 7789 6934
rect 9069 6874 9106 6875
rect 9372 6874 9409 7016
rect 9434 7036 9521 7043
rect 9434 7033 9492 7036
rect 9434 7013 9439 7033
rect 9460 7016 9492 7033
rect 9512 7016 9521 7036
rect 9460 7013 9521 7016
rect 9434 7006 9521 7013
rect 9580 7036 9617 7046
rect 9580 7016 9588 7036
rect 9608 7016 9617 7036
rect 9434 7005 9465 7006
rect 9580 6937 9617 7016
rect 9647 7045 9678 7098
rect 9891 7091 9906 7099
rect 9946 7091 9956 7128
rect 9891 7082 9956 7091
rect 10104 7089 10169 7110
rect 10104 7071 10129 7089
rect 10147 7071 10169 7089
rect 9697 7045 9734 7046
rect 9647 7036 9734 7045
rect 9647 7016 9705 7036
rect 9725 7016 9734 7036
rect 9647 7006 9734 7016
rect 9793 7036 9830 7046
rect 9793 7016 9801 7036
rect 9821 7016 9830 7036
rect 9647 7005 9678 7006
rect 9642 6937 9752 6950
rect 9793 6937 9830 7016
rect 10104 6995 10169 7071
rect 9580 6935 9830 6937
rect 9580 6932 9681 6935
rect 9580 6913 9645 6932
rect 9642 6905 9645 6913
rect 9674 6905 9681 6932
rect 9709 6908 9719 6935
rect 9748 6913 9830 6935
rect 9853 6960 10170 6995
rect 9748 6908 9752 6913
rect 9709 6905 9752 6908
rect 9642 6891 9752 6905
rect 9068 6873 9409 6874
rect 8993 6871 9409 6873
rect 9853 6871 9893 6960
rect 10104 6933 10169 6960
rect 10104 6915 10127 6933
rect 10145 6915 10169 6933
rect 10104 6895 10169 6915
rect 8990 6868 9893 6871
rect 8990 6848 8996 6868
rect 9016 6848 9893 6868
rect 8990 6844 9893 6848
rect 9853 6841 9893 6844
rect 10105 6834 10170 6855
rect 8323 6826 8984 6827
rect 8323 6819 9257 6826
rect 8323 6818 9229 6819
rect 8323 6798 9174 6818
rect 9206 6799 9229 6818
rect 9254 6799 9257 6819
rect 9206 6798 9257 6799
rect 8323 6791 9257 6798
rect 7922 6749 8090 6750
rect 8325 6749 8364 6791
rect 9153 6789 9257 6791
rect 9222 6787 9257 6789
rect 10105 6816 10129 6834
rect 10147 6816 10170 6834
rect 10105 6769 10170 6816
rect 7922 6723 8366 6749
rect 7922 6721 8090 6723
rect 7727 6444 7791 6463
rect 7727 6405 7744 6444
rect 7778 6405 7791 6444
rect 7727 6386 7791 6405
rect 7532 6357 7627 6383
rect 7922 6370 7949 6721
rect 8325 6717 8366 6723
rect 7989 6510 8053 6522
rect 8329 6518 8366 6717
rect 8828 6744 8900 6761
rect 8828 6705 8836 6744
rect 8881 6705 8900 6744
rect 8594 6607 8705 6622
rect 8594 6605 8636 6607
rect 8594 6585 8601 6605
rect 8620 6585 8636 6605
rect 8594 6577 8636 6585
rect 8664 6605 8705 6607
rect 8664 6585 8678 6605
rect 8697 6585 8705 6605
rect 8664 6577 8705 6585
rect 8594 6571 8705 6577
rect 8537 6549 8786 6571
rect 8537 6518 8574 6549
rect 8750 6547 8786 6549
rect 8750 6518 8787 6547
rect 7989 6509 8024 6510
rect 7966 6504 8024 6509
rect 7966 6484 7969 6504
rect 7989 6490 8024 6504
rect 8044 6490 8053 6510
rect 7989 6482 8053 6490
rect 8015 6481 8053 6482
rect 8016 6480 8053 6481
rect 8119 6514 8155 6515
rect 8227 6514 8263 6515
rect 8119 6506 8263 6514
rect 8119 6486 8127 6506
rect 8147 6486 8235 6506
rect 8255 6486 8263 6506
rect 8119 6480 8263 6486
rect 8329 6510 8367 6518
rect 8435 6514 8471 6515
rect 8329 6490 8338 6510
rect 8358 6490 8367 6510
rect 8329 6481 8367 6490
rect 8386 6507 8471 6514
rect 8386 6487 8393 6507
rect 8414 6506 8471 6507
rect 8414 6487 8443 6506
rect 8386 6486 8443 6487
rect 8463 6486 8471 6506
rect 8329 6480 8366 6481
rect 8386 6480 8471 6486
rect 8537 6510 8575 6518
rect 8648 6514 8684 6515
rect 8537 6490 8546 6510
rect 8566 6490 8575 6510
rect 8537 6481 8575 6490
rect 8599 6506 8684 6514
rect 8599 6486 8656 6506
rect 8676 6486 8684 6506
rect 8537 6480 8574 6481
rect 8599 6480 8684 6486
rect 8750 6510 8788 6518
rect 8750 6490 8759 6510
rect 8779 6490 8788 6510
rect 8750 6481 8788 6490
rect 8828 6495 8900 6705
rect 8970 6739 10170 6769
rect 8970 6738 9414 6739
rect 8970 6736 9138 6738
rect 8828 6481 8911 6495
rect 8750 6480 8787 6481
rect 8173 6459 8209 6480
rect 8599 6459 8630 6480
rect 8828 6459 8845 6481
rect 8006 6455 8106 6459
rect 8006 6451 8068 6455
rect 8006 6425 8013 6451
rect 8039 6429 8068 6451
rect 8094 6429 8106 6455
rect 8039 6425 8106 6429
rect 8006 6422 8106 6425
rect 8174 6422 8209 6459
rect 8271 6456 8630 6459
rect 8271 6451 8493 6456
rect 8271 6427 8284 6451
rect 8308 6432 8493 6451
rect 8517 6432 8630 6456
rect 8308 6427 8630 6432
rect 8271 6423 8630 6427
rect 8697 6451 8845 6459
rect 8697 6431 8708 6451
rect 8728 6448 8845 6451
rect 8898 6448 8911 6481
rect 8728 6431 8911 6448
rect 8697 6424 8911 6431
rect 8697 6423 8738 6424
rect 8828 6423 8911 6424
rect 8173 6397 8209 6422
rect 8021 6370 8058 6371
rect 8117 6370 8154 6371
rect 8173 6370 8180 6397
rect 7921 6361 8059 6370
rect 7921 6341 8030 6361
rect 8050 6341 8059 6361
rect 7921 6334 8059 6341
rect 8117 6367 8180 6370
rect 8201 6370 8209 6397
rect 8228 6370 8265 6371
rect 8201 6367 8265 6370
rect 8117 6361 8265 6367
rect 8117 6341 8126 6361
rect 8146 6341 8236 6361
rect 8256 6341 8265 6361
rect 7921 6332 8017 6334
rect 8117 6331 8265 6341
rect 8324 6361 8361 6371
rect 8436 6370 8473 6371
rect 8417 6368 8473 6370
rect 8324 6341 8332 6361
rect 8352 6341 8361 6361
rect 8173 6330 8209 6331
rect 8021 6199 8058 6200
rect 8324 6199 8361 6341
rect 8386 6361 8473 6368
rect 8386 6358 8444 6361
rect 8386 6338 8391 6358
rect 8412 6341 8444 6358
rect 8464 6341 8473 6361
rect 8412 6338 8473 6341
rect 8386 6331 8473 6338
rect 8532 6361 8569 6371
rect 8532 6341 8540 6361
rect 8560 6341 8569 6361
rect 8386 6330 8417 6331
rect 8532 6262 8569 6341
rect 8599 6370 8630 6423
rect 8836 6390 8850 6423
rect 8903 6390 8911 6423
rect 8836 6384 8911 6390
rect 8836 6379 8906 6384
rect 8649 6370 8686 6371
rect 8599 6361 8686 6370
rect 8599 6341 8657 6361
rect 8677 6341 8686 6361
rect 8599 6331 8686 6341
rect 8745 6361 8782 6371
rect 8970 6366 8997 6736
rect 9037 6506 9101 6518
rect 9377 6514 9414 6738
rect 9885 6719 9949 6721
rect 9881 6707 9949 6719
rect 9881 6674 9892 6707
rect 9932 6674 9949 6707
rect 9881 6664 9949 6674
rect 9642 6603 9753 6618
rect 9642 6601 9684 6603
rect 9642 6581 9649 6601
rect 9668 6581 9684 6601
rect 9642 6573 9684 6581
rect 9712 6601 9753 6603
rect 9712 6581 9726 6601
rect 9745 6581 9753 6601
rect 9712 6573 9753 6581
rect 9642 6567 9753 6573
rect 9585 6545 9834 6567
rect 9585 6514 9622 6545
rect 9798 6543 9834 6545
rect 9798 6514 9835 6543
rect 9037 6505 9072 6506
rect 9014 6500 9072 6505
rect 9014 6480 9017 6500
rect 9037 6486 9072 6500
rect 9092 6486 9101 6506
rect 9037 6478 9101 6486
rect 9063 6477 9101 6478
rect 9064 6476 9101 6477
rect 9167 6510 9203 6511
rect 9275 6510 9311 6511
rect 9167 6502 9311 6510
rect 9167 6482 9175 6502
rect 9195 6482 9283 6502
rect 9303 6482 9311 6502
rect 9167 6476 9311 6482
rect 9377 6506 9415 6514
rect 9483 6510 9519 6511
rect 9377 6486 9386 6506
rect 9406 6486 9415 6506
rect 9377 6477 9415 6486
rect 9434 6503 9519 6510
rect 9434 6483 9441 6503
rect 9462 6502 9519 6503
rect 9462 6483 9491 6502
rect 9434 6482 9491 6483
rect 9511 6482 9519 6502
rect 9377 6476 9414 6477
rect 9434 6476 9519 6482
rect 9585 6506 9623 6514
rect 9696 6510 9732 6511
rect 9585 6486 9594 6506
rect 9614 6486 9623 6506
rect 9585 6477 9623 6486
rect 9647 6502 9732 6510
rect 9647 6482 9704 6502
rect 9724 6482 9732 6502
rect 9585 6476 9622 6477
rect 9647 6476 9732 6482
rect 9798 6506 9836 6514
rect 9798 6486 9807 6506
rect 9827 6486 9836 6506
rect 9798 6477 9836 6486
rect 9885 6480 9949 6664
rect 10105 6538 10170 6739
rect 10105 6520 10127 6538
rect 10145 6520 10170 6538
rect 10105 6501 10170 6520
rect 9798 6476 9835 6477
rect 9221 6455 9257 6476
rect 9647 6455 9678 6476
rect 9885 6471 9893 6480
rect 9882 6455 9893 6471
rect 9054 6451 9154 6455
rect 9054 6447 9116 6451
rect 9054 6421 9061 6447
rect 9087 6425 9116 6447
rect 9142 6425 9154 6451
rect 9087 6421 9154 6425
rect 9054 6418 9154 6421
rect 9222 6418 9257 6455
rect 9319 6452 9678 6455
rect 9319 6447 9541 6452
rect 9319 6423 9332 6447
rect 9356 6428 9541 6447
rect 9565 6428 9678 6452
rect 9356 6423 9678 6428
rect 9319 6419 9678 6423
rect 9745 6447 9893 6455
rect 9745 6427 9756 6447
rect 9776 6438 9893 6447
rect 9942 6471 9949 6480
rect 9942 6438 9950 6471
rect 9776 6427 9950 6438
rect 9745 6420 9950 6427
rect 9745 6419 9786 6420
rect 9221 6393 9257 6418
rect 9069 6366 9106 6367
rect 9165 6366 9202 6367
rect 9221 6366 9228 6393
rect 8745 6341 8753 6361
rect 8773 6341 8782 6361
rect 8599 6330 8630 6331
rect 8594 6262 8704 6275
rect 8745 6262 8782 6341
rect 8969 6357 9107 6366
rect 8969 6337 9078 6357
rect 9098 6337 9107 6357
rect 8969 6330 9107 6337
rect 9165 6363 9228 6366
rect 9249 6366 9257 6393
rect 9276 6366 9313 6367
rect 9249 6363 9313 6366
rect 9165 6357 9313 6363
rect 9165 6337 9174 6357
rect 9194 6337 9284 6357
rect 9304 6337 9313 6357
rect 8969 6328 9065 6330
rect 9165 6327 9313 6337
rect 9372 6357 9409 6367
rect 9484 6366 9521 6367
rect 9465 6364 9521 6366
rect 9372 6337 9380 6357
rect 9400 6337 9409 6357
rect 9221 6326 9257 6327
rect 8532 6260 8782 6262
rect 8532 6257 8633 6260
rect 8532 6238 8597 6257
rect 8594 6230 8597 6238
rect 8626 6230 8633 6257
rect 8661 6233 8671 6260
rect 8700 6238 8782 6260
rect 8700 6233 8704 6238
rect 8661 6230 8704 6233
rect 8594 6216 8704 6230
rect 8020 6198 8361 6199
rect 7945 6193 8361 6198
rect 9069 6195 9106 6196
rect 9372 6195 9409 6337
rect 9434 6357 9521 6364
rect 9434 6354 9492 6357
rect 9434 6334 9439 6354
rect 9460 6337 9492 6354
rect 9512 6337 9521 6357
rect 9460 6334 9521 6337
rect 9434 6327 9521 6334
rect 9580 6357 9617 6367
rect 9580 6337 9588 6357
rect 9608 6337 9617 6357
rect 9434 6326 9465 6327
rect 9580 6258 9617 6337
rect 9647 6366 9678 6419
rect 9882 6417 9950 6420
rect 9882 6375 9894 6417
rect 9943 6375 9950 6417
rect 9697 6366 9734 6367
rect 9647 6357 9734 6366
rect 9647 6337 9705 6357
rect 9725 6337 9734 6357
rect 9647 6327 9734 6337
rect 9793 6357 9830 6367
rect 9882 6362 9950 6375
rect 10105 6439 10170 6456
rect 10105 6421 10129 6439
rect 10147 6421 10170 6439
rect 9793 6337 9801 6357
rect 9821 6337 9830 6357
rect 9647 6326 9678 6327
rect 9642 6258 9752 6271
rect 9793 6258 9830 6337
rect 10105 6282 10170 6421
rect 10105 6276 10127 6282
rect 9580 6256 9830 6258
rect 9580 6253 9681 6256
rect 9580 6234 9645 6253
rect 9642 6226 9645 6234
rect 9674 6226 9681 6253
rect 9709 6229 9719 6256
rect 9748 6234 9830 6256
rect 9859 6264 10127 6276
rect 10145 6264 10170 6282
rect 9859 6241 10170 6264
rect 9859 6240 9914 6241
rect 9748 6229 9752 6234
rect 9709 6226 9752 6229
rect 9642 6212 9752 6226
rect 9068 6194 9409 6195
rect 7945 6173 7948 6193
rect 7968 6173 8361 6193
rect 8993 6193 9409 6194
rect 9859 6193 9902 6240
rect 8993 6189 9902 6193
rect 6868 6138 7579 6140
rect 8118 6138 8207 6141
rect 6868 6129 8207 6138
rect 6868 6091 8130 6129
rect 8155 6094 8174 6129
rect 8199 6094 8207 6129
rect 8312 6140 8357 6173
rect 8993 6169 8996 6189
rect 9016 6169 9902 6189
rect 9370 6164 9902 6169
rect 10110 6183 10169 6205
rect 10110 6165 10129 6183
rect 10147 6165 10169 6183
rect 9158 6140 9257 6142
rect 8312 6130 9257 6140
rect 8312 6104 9180 6130
rect 8313 6103 9180 6104
rect 8155 6091 8207 6094
rect 6868 6083 8207 6091
rect 9158 6092 9180 6103
rect 9205 6095 9224 6130
rect 9249 6095 9257 6130
rect 9205 6092 9257 6095
rect 9158 6084 9257 6092
rect 10110 6091 10169 6165
rect 9184 6083 9256 6084
rect 6868 6082 8206 6083
rect 6868 6080 7579 6082
rect 7728 6041 7792 6045
rect 10103 6043 10169 6091
rect 7728 6032 7802 6041
rect 6243 5549 6357 5553
rect 5448 5545 5548 5549
rect 5448 5541 5510 5545
rect 5448 5515 5455 5541
rect 5481 5519 5510 5541
rect 5536 5519 5548 5545
rect 5481 5515 5548 5519
rect 5448 5512 5548 5515
rect 5616 5512 5651 5549
rect 5713 5546 6072 5549
rect 5713 5541 5935 5546
rect 5713 5517 5726 5541
rect 5750 5522 5935 5541
rect 5959 5522 6072 5546
rect 5750 5517 6072 5522
rect 5713 5513 6072 5517
rect 6139 5546 6357 5549
rect 6139 5545 6322 5546
rect 6139 5541 6265 5545
rect 6139 5521 6150 5541
rect 6170 5521 6265 5541
rect 6289 5522 6322 5545
rect 6346 5522 6357 5546
rect 6289 5521 6357 5522
rect 6139 5514 6357 5521
rect 6139 5513 6180 5514
rect 5615 5487 5651 5512
rect 5463 5460 5500 5461
rect 5559 5460 5596 5461
rect 5615 5460 5622 5487
rect 5363 5451 5501 5460
rect 5363 5431 5472 5451
rect 5492 5431 5501 5451
rect 5363 5424 5501 5431
rect 5559 5457 5622 5460
rect 5643 5460 5651 5487
rect 5670 5460 5707 5461
rect 5643 5457 5707 5460
rect 5559 5451 5707 5457
rect 5559 5431 5568 5451
rect 5588 5431 5678 5451
rect 5698 5431 5707 5451
rect 5363 5422 5459 5424
rect 5559 5421 5707 5431
rect 5766 5451 5803 5461
rect 5878 5460 5915 5461
rect 5859 5458 5915 5460
rect 5766 5431 5774 5451
rect 5794 5431 5803 5451
rect 5615 5420 5651 5421
rect 5463 5289 5500 5290
rect 5766 5289 5803 5431
rect 5828 5451 5915 5458
rect 5828 5448 5886 5451
rect 5828 5428 5833 5448
rect 5854 5431 5886 5448
rect 5906 5431 5915 5451
rect 5854 5428 5915 5431
rect 5828 5421 5915 5428
rect 5974 5451 6011 5461
rect 5974 5431 5982 5451
rect 6002 5431 6011 5451
rect 5828 5420 5859 5421
rect 5974 5352 6011 5431
rect 6041 5460 6072 5513
rect 6243 5511 6357 5514
rect 6286 5479 6357 5511
rect 7532 5990 7616 6015
rect 7532 5962 7547 5990
rect 7591 5962 7616 5990
rect 7532 5933 7616 5962
rect 7728 5984 7742 6032
rect 7779 5984 7802 6032
rect 7728 5956 7802 5984
rect 7532 5905 7544 5933
rect 7588 5905 7616 5933
rect 7532 5884 7616 5905
rect 6091 5460 6128 5461
rect 6041 5451 6128 5460
rect 6041 5431 6099 5451
rect 6119 5431 6128 5451
rect 6041 5421 6128 5431
rect 6187 5451 6224 5461
rect 6187 5431 6195 5451
rect 6215 5431 6224 5451
rect 6041 5420 6072 5421
rect 6036 5352 6146 5365
rect 6187 5352 6224 5431
rect 5974 5350 6224 5352
rect 5974 5347 6075 5350
rect 5974 5328 6039 5347
rect 6036 5320 6039 5328
rect 6068 5320 6075 5347
rect 6103 5323 6113 5350
rect 6142 5328 6224 5350
rect 6142 5323 6146 5328
rect 6103 5320 6146 5323
rect 6036 5306 6146 5320
rect 5462 5288 5803 5289
rect 5387 5285 5803 5288
rect 5387 5283 5810 5285
rect 5387 5263 5390 5283
rect 5410 5263 5810 5283
rect 4578 2922 5218 3010
rect 4578 2571 4662 2922
rect 5144 2891 5188 2897
rect 5144 2865 5152 2891
rect 5177 2865 5188 2891
rect 5144 2816 5188 2865
rect 5144 2796 5541 2816
rect 5561 2796 5564 2816
rect 5144 2791 5564 2796
rect 5144 2790 5489 2791
rect 5144 2786 5188 2790
rect 5451 2789 5488 2790
rect 4805 2759 4915 2773
rect 4805 2756 4848 2759
rect 4805 2751 4809 2756
rect 4727 2729 4809 2751
rect 4838 2729 4848 2756
rect 4876 2732 4883 2759
rect 4912 2751 4915 2759
rect 4912 2732 4977 2751
rect 4876 2729 4977 2732
rect 4727 2727 4977 2729
rect 4727 2648 4764 2727
rect 4805 2714 4915 2727
rect 4879 2658 4910 2659
rect 4727 2628 4736 2648
rect 4756 2628 4764 2648
rect 4727 2618 4764 2628
rect 4823 2648 4910 2658
rect 4823 2628 4832 2648
rect 4852 2628 4910 2648
rect 4823 2619 4910 2628
rect 4823 2618 4860 2619
rect 4578 2565 4687 2571
rect 4879 2566 4910 2619
rect 4940 2648 4977 2727
rect 5092 2658 5123 2659
rect 4940 2628 4949 2648
rect 4969 2628 4977 2648
rect 4940 2618 4977 2628
rect 5036 2651 5123 2658
rect 5036 2648 5097 2651
rect 5036 2628 5045 2648
rect 5065 2631 5097 2648
rect 5118 2631 5123 2651
rect 5065 2628 5123 2631
rect 5036 2621 5123 2628
rect 5148 2648 5185 2786
rect 5300 2658 5336 2659
rect 5148 2628 5157 2648
rect 5177 2628 5185 2648
rect 5036 2619 5092 2621
rect 5036 2618 5073 2619
rect 5148 2618 5185 2628
rect 5244 2648 5392 2658
rect 5492 2655 5588 2657
rect 5244 2628 5253 2648
rect 5273 2628 5363 2648
rect 5383 2628 5392 2648
rect 5244 2622 5392 2628
rect 5244 2619 5308 2622
rect 5244 2618 5281 2619
rect 5300 2592 5308 2619
rect 5329 2619 5392 2622
rect 5450 2648 5588 2655
rect 5450 2628 5459 2648
rect 5479 2628 5588 2648
rect 5450 2619 5588 2628
rect 5329 2592 5336 2619
rect 5355 2618 5392 2619
rect 5451 2618 5488 2619
rect 5300 2567 5336 2592
rect 4771 2565 4812 2566
rect 4578 2558 4812 2565
rect 4578 2538 4781 2558
rect 4801 2538 4812 2558
rect 4578 2530 4812 2538
rect 4879 2562 5238 2566
rect 4879 2557 5201 2562
rect 4879 2533 4992 2557
rect 5016 2538 5201 2557
rect 5225 2538 5238 2562
rect 5016 2533 5238 2538
rect 4879 2530 5238 2533
rect 5300 2530 5335 2567
rect 5403 2564 5503 2567
rect 5403 2560 5470 2564
rect 5403 2534 5415 2560
rect 5441 2538 5470 2560
rect 5496 2538 5503 2564
rect 5441 2534 5503 2538
rect 5403 2530 5503 2534
rect 4578 2512 4687 2530
rect 4879 2509 4910 2530
rect 5300 2509 5336 2530
rect 4722 2508 4759 2509
rect 4721 2499 4759 2508
rect 4721 2479 4730 2499
rect 4750 2479 4759 2499
rect 4721 2471 4759 2479
rect 4825 2503 4910 2509
rect 4935 2508 4972 2509
rect 4825 2483 4833 2503
rect 4853 2483 4910 2503
rect 4825 2475 4910 2483
rect 4934 2499 4972 2508
rect 4934 2479 4943 2499
rect 4963 2479 4972 2499
rect 4825 2474 4861 2475
rect 4934 2471 4972 2479
rect 5038 2503 5123 2509
rect 5143 2508 5180 2509
rect 5038 2483 5046 2503
rect 5066 2502 5123 2503
rect 5066 2483 5095 2502
rect 5038 2482 5095 2483
rect 5116 2482 5123 2502
rect 5038 2475 5123 2482
rect 5142 2499 5180 2508
rect 5142 2479 5151 2499
rect 5171 2479 5180 2499
rect 5038 2474 5074 2475
rect 5142 2471 5180 2479
rect 5246 2504 5390 2509
rect 5246 2503 5299 2504
rect 5246 2483 5254 2503
rect 5274 2484 5299 2503
rect 5332 2503 5390 2504
rect 5332 2484 5362 2503
rect 5274 2483 5362 2484
rect 5382 2483 5390 2503
rect 5246 2475 5390 2483
rect 5246 2474 5282 2475
rect 5354 2474 5390 2475
rect 5456 2508 5493 2509
rect 5456 2507 5494 2508
rect 5456 2499 5520 2507
rect 5456 2479 5465 2499
rect 5485 2485 5520 2499
rect 5540 2485 5543 2505
rect 5485 2480 5543 2485
rect 5485 2479 5520 2480
rect 4722 2442 4759 2471
rect 4723 2440 4759 2442
rect 4935 2440 4972 2471
rect 4723 2418 4972 2440
rect 4804 2412 4915 2418
rect 4804 2404 4845 2412
rect 4804 2384 4812 2404
rect 4831 2384 4845 2404
rect 4804 2382 4845 2384
rect 4873 2404 4915 2412
rect 4873 2384 4889 2404
rect 4908 2384 4915 2404
rect 4873 2382 4915 2384
rect 4804 2367 4915 2382
rect 5143 2350 5180 2471
rect 5456 2467 5520 2479
rect 5560 2356 5587 2619
rect 5614 2365 5650 2372
rect 5614 2356 5620 2365
rect 5538 2352 5620 2356
rect 5419 2350 5620 2352
rect 5143 2327 5620 2350
rect 5643 2327 5650 2365
rect 5143 2324 5650 2327
rect 5419 2323 5587 2324
rect 5614 2321 5650 2324
rect 5732 2223 5810 5263
rect 6866 4516 6925 4526
rect 6866 4488 6879 4516
rect 6907 4488 6925 4516
rect 6866 4439 6925 4488
rect 6472 4304 6640 4305
rect 6876 4304 6923 4439
rect 6472 4278 6923 4304
rect 6472 4276 6640 4278
rect 6472 4009 6499 4276
rect 6876 4272 6923 4278
rect 6539 4149 6603 4161
rect 6879 4157 6916 4272
rect 7144 4246 7255 4261
rect 7144 4244 7186 4246
rect 7144 4224 7151 4244
rect 7170 4224 7186 4244
rect 7144 4216 7186 4224
rect 7214 4244 7255 4246
rect 7214 4224 7228 4244
rect 7247 4224 7255 4244
rect 7214 4216 7255 4224
rect 7144 4210 7255 4216
rect 7087 4188 7336 4210
rect 7087 4157 7124 4188
rect 7300 4186 7336 4188
rect 7300 4157 7337 4186
rect 6539 4148 6574 4149
rect 6516 4143 6574 4148
rect 6516 4123 6519 4143
rect 6539 4129 6574 4143
rect 6594 4129 6603 4149
rect 6539 4121 6603 4129
rect 6565 4120 6603 4121
rect 6566 4119 6603 4120
rect 6669 4153 6705 4154
rect 6777 4153 6813 4154
rect 6669 4145 6813 4153
rect 6669 4125 6677 4145
rect 6697 4125 6785 4145
rect 6805 4125 6813 4145
rect 6669 4119 6813 4125
rect 6879 4149 6917 4157
rect 6985 4153 7021 4154
rect 6879 4129 6888 4149
rect 6908 4129 6917 4149
rect 6879 4120 6917 4129
rect 6936 4146 7021 4153
rect 6936 4126 6943 4146
rect 6964 4145 7021 4146
rect 6964 4126 6993 4145
rect 6936 4125 6993 4126
rect 7013 4125 7021 4145
rect 6879 4119 6916 4120
rect 6936 4119 7021 4125
rect 7087 4149 7125 4157
rect 7198 4153 7234 4154
rect 7087 4129 7096 4149
rect 7116 4129 7125 4149
rect 7087 4120 7125 4129
rect 7149 4145 7234 4153
rect 7149 4125 7206 4145
rect 7226 4125 7234 4145
rect 7087 4119 7124 4120
rect 7149 4119 7234 4125
rect 7300 4149 7338 4157
rect 7300 4129 7309 4149
rect 7329 4129 7338 4149
rect 7300 4120 7338 4129
rect 7300 4119 7337 4120
rect 6723 4098 6759 4119
rect 7149 4098 7180 4119
rect 7360 4104 7417 4112
rect 7360 4098 7368 4104
rect 6556 4094 6656 4098
rect 6556 4090 6618 4094
rect 6556 4064 6563 4090
rect 6589 4068 6618 4090
rect 6644 4068 6656 4094
rect 6589 4064 6656 4068
rect 6556 4061 6656 4064
rect 6724 4061 6759 4098
rect 6821 4095 7180 4098
rect 6821 4090 7043 4095
rect 6821 4066 6834 4090
rect 6858 4071 7043 4090
rect 7067 4071 7180 4095
rect 6858 4066 7180 4071
rect 6821 4062 7180 4066
rect 7247 4090 7368 4098
rect 7247 4070 7258 4090
rect 7278 4081 7368 4090
rect 7394 4081 7417 4104
rect 7278 4070 7417 4081
rect 7247 4068 7417 4070
rect 7247 4063 7368 4068
rect 7247 4062 7288 4063
rect 6723 4036 6759 4061
rect 6571 4009 6608 4010
rect 6667 4009 6704 4010
rect 6723 4009 6730 4036
rect 6471 4000 6609 4009
rect 6471 3980 6580 4000
rect 6600 3980 6609 4000
rect 6471 3973 6609 3980
rect 6667 4006 6730 4009
rect 6751 4009 6759 4036
rect 6778 4009 6815 4010
rect 6751 4006 6815 4009
rect 6667 4000 6815 4006
rect 6667 3980 6676 4000
rect 6696 3980 6786 4000
rect 6806 3980 6815 4000
rect 6471 3971 6567 3973
rect 6667 3970 6815 3980
rect 6874 4000 6911 4010
rect 6986 4009 7023 4010
rect 6967 4007 7023 4009
rect 6874 3980 6882 4000
rect 6902 3980 6911 4000
rect 6723 3969 6759 3970
rect 6571 3838 6608 3839
rect 6874 3838 6911 3980
rect 6936 4000 7023 4007
rect 6936 3997 6994 4000
rect 6936 3977 6941 3997
rect 6962 3980 6994 3997
rect 7014 3980 7023 4000
rect 6962 3977 7023 3980
rect 6936 3970 7023 3977
rect 7082 4000 7119 4010
rect 7082 3980 7090 4000
rect 7110 3980 7119 4000
rect 6936 3969 6967 3970
rect 7082 3901 7119 3980
rect 7149 4009 7180 4062
rect 7199 4009 7236 4010
rect 7149 4000 7236 4009
rect 7149 3980 7207 4000
rect 7227 3980 7236 4000
rect 7149 3970 7236 3980
rect 7295 4000 7332 4010
rect 7295 3980 7303 4000
rect 7323 3980 7332 4000
rect 7149 3969 7180 3970
rect 7144 3901 7254 3914
rect 7295 3901 7332 3980
rect 7082 3899 7332 3901
rect 7082 3896 7183 3899
rect 7082 3877 7147 3896
rect 7144 3869 7147 3877
rect 7176 3869 7183 3896
rect 7211 3872 7221 3899
rect 7250 3877 7332 3899
rect 7250 3872 7254 3877
rect 7211 3869 7254 3872
rect 7144 3855 7254 3869
rect 6570 3837 6911 3838
rect 6495 3832 6911 3837
rect 6495 3812 6498 3832
rect 6518 3812 6912 3832
rect 6721 3779 6758 3789
rect 6721 3742 6730 3779
rect 6747 3742 6758 3779
rect 6721 3721 6758 3742
rect 6430 2782 6598 2783
rect 6727 2782 6756 3721
rect 6869 3107 6912 3812
rect 6870 3099 6912 3107
rect 6870 3088 6915 3099
rect 6870 3050 6880 3088
rect 6905 3050 6915 3088
rect 6870 3041 6915 3050
rect 6430 2756 6874 2782
rect 6430 2754 6598 2756
rect 6430 2487 6457 2754
rect 6727 2752 6756 2756
rect 6497 2627 6561 2639
rect 6837 2635 6874 2756
rect 7102 2724 7213 2739
rect 7102 2722 7144 2724
rect 7102 2702 7109 2722
rect 7128 2702 7144 2722
rect 7102 2694 7144 2702
rect 7172 2722 7213 2724
rect 7172 2702 7186 2722
rect 7205 2702 7213 2722
rect 7172 2694 7213 2702
rect 7102 2688 7213 2694
rect 7045 2666 7294 2688
rect 7045 2635 7082 2666
rect 7258 2664 7294 2666
rect 7258 2635 7295 2664
rect 6497 2626 6532 2627
rect 6474 2621 6532 2626
rect 6474 2601 6477 2621
rect 6497 2607 6532 2621
rect 6552 2607 6561 2627
rect 6497 2599 6561 2607
rect 6523 2598 6561 2599
rect 6524 2597 6561 2598
rect 6627 2631 6663 2632
rect 6735 2631 6771 2632
rect 6627 2623 6771 2631
rect 6627 2603 6635 2623
rect 6655 2603 6743 2623
rect 6763 2603 6771 2623
rect 6627 2597 6771 2603
rect 6837 2627 6875 2635
rect 6943 2631 6979 2632
rect 6837 2607 6846 2627
rect 6866 2607 6875 2627
rect 6837 2598 6875 2607
rect 6894 2624 6979 2631
rect 6894 2604 6901 2624
rect 6922 2623 6979 2624
rect 6922 2604 6951 2623
rect 6894 2603 6951 2604
rect 6971 2603 6979 2623
rect 6837 2597 6874 2598
rect 6894 2597 6979 2603
rect 7045 2627 7083 2635
rect 7156 2631 7192 2632
rect 7045 2607 7054 2627
rect 7074 2607 7083 2627
rect 7045 2598 7083 2607
rect 7107 2623 7192 2631
rect 7107 2603 7164 2623
rect 7184 2603 7192 2623
rect 7045 2597 7082 2598
rect 7107 2597 7192 2603
rect 7258 2627 7296 2635
rect 7258 2607 7267 2627
rect 7287 2607 7296 2627
rect 7258 2598 7296 2607
rect 7258 2597 7295 2598
rect 6681 2576 6717 2597
rect 7107 2576 7138 2597
rect 7532 2580 7624 5884
rect 7730 4117 7802 5956
rect 8832 5906 8904 5923
rect 8832 5858 8844 5906
rect 8890 5858 8904 5906
rect 9372 5886 9413 5888
rect 9644 5886 9748 5888
rect 10103 5886 10168 6043
rect 8832 5836 8904 5858
rect 8965 5851 10168 5886
rect 8965 5837 8993 5851
rect 8833 5636 8903 5836
rect 8967 5706 8993 5837
rect 9372 5848 10168 5851
rect 8825 5585 8905 5636
rect 8825 5559 8841 5585
rect 8881 5559 8905 5585
rect 8825 5540 8905 5559
rect 8825 5514 8844 5540
rect 8884 5514 8905 5540
rect 8825 5487 8905 5514
rect 8825 5461 8848 5487
rect 8888 5461 8905 5487
rect 8825 5450 8905 5461
rect 8967 5451 8994 5706
rect 9372 5698 9413 5848
rect 9644 5846 9748 5848
rect 10103 5814 10168 5848
rect 9839 5786 9960 5804
rect 9839 5784 9910 5786
rect 9839 5743 9854 5784
rect 9891 5745 9910 5784
rect 9947 5745 9960 5786
rect 9891 5743 9960 5745
rect 9839 5733 9960 5743
rect 9644 5703 9748 5706
rect 9034 5591 9098 5603
rect 9374 5599 9411 5698
rect 9639 5688 9750 5703
rect 9639 5686 9681 5688
rect 9639 5666 9646 5686
rect 9665 5666 9681 5686
rect 9639 5658 9681 5666
rect 9709 5686 9750 5688
rect 9709 5666 9723 5686
rect 9742 5666 9750 5686
rect 9709 5658 9750 5666
rect 9639 5652 9750 5658
rect 9582 5630 9831 5652
rect 9582 5599 9619 5630
rect 9795 5628 9831 5630
rect 9795 5599 9832 5628
rect 9034 5590 9069 5591
rect 9011 5585 9069 5590
rect 9011 5565 9014 5585
rect 9034 5571 9069 5585
rect 9089 5571 9098 5591
rect 9034 5563 9098 5571
rect 9060 5562 9098 5563
rect 9061 5561 9098 5562
rect 9164 5595 9200 5596
rect 9272 5595 9308 5596
rect 9164 5587 9308 5595
rect 9164 5567 9172 5587
rect 9192 5567 9280 5587
rect 9300 5567 9308 5587
rect 9164 5561 9308 5567
rect 9374 5591 9412 5599
rect 9480 5595 9516 5596
rect 9374 5571 9383 5591
rect 9403 5571 9412 5591
rect 9374 5562 9412 5571
rect 9431 5588 9516 5595
rect 9431 5568 9438 5588
rect 9459 5587 9516 5588
rect 9459 5568 9488 5587
rect 9431 5567 9488 5568
rect 9508 5567 9516 5587
rect 9374 5561 9411 5562
rect 9431 5561 9516 5567
rect 9582 5591 9620 5599
rect 9693 5595 9729 5596
rect 9582 5571 9591 5591
rect 9611 5571 9620 5591
rect 9582 5562 9620 5571
rect 9644 5587 9729 5595
rect 9644 5567 9701 5587
rect 9721 5567 9729 5587
rect 9582 5561 9619 5562
rect 9644 5561 9729 5567
rect 9795 5591 9833 5599
rect 9795 5571 9804 5591
rect 9824 5571 9833 5591
rect 9888 5581 9953 5733
rect 10106 5707 10161 5814
rect 9795 5562 9833 5571
rect 9886 5574 9953 5581
rect 9795 5561 9832 5562
rect 9218 5540 9254 5561
rect 9644 5540 9675 5561
rect 9886 5553 9903 5574
rect 9939 5553 9953 5574
rect 10105 5594 10161 5707
rect 10105 5576 10124 5594
rect 10142 5576 10161 5594
rect 10105 5556 10161 5576
rect 9886 5540 9953 5553
rect 9051 5536 9151 5540
rect 9051 5532 9113 5536
rect 9051 5506 9058 5532
rect 9084 5510 9113 5532
rect 9139 5510 9151 5536
rect 9084 5506 9151 5510
rect 9051 5503 9151 5506
rect 9219 5503 9254 5540
rect 9316 5537 9675 5540
rect 9316 5532 9538 5537
rect 9316 5508 9329 5532
rect 9353 5513 9538 5532
rect 9562 5513 9675 5537
rect 9353 5508 9675 5513
rect 9316 5504 9675 5508
rect 9742 5534 9953 5540
rect 9742 5532 9903 5534
rect 9742 5512 9753 5532
rect 9773 5512 9903 5532
rect 9742 5505 9903 5512
rect 9742 5504 9783 5505
rect 9218 5478 9254 5503
rect 9066 5451 9103 5452
rect 9162 5451 9199 5452
rect 9218 5451 9225 5478
rect 8966 5442 9104 5451
rect 8966 5422 9075 5442
rect 9095 5422 9104 5442
rect 8966 5415 9104 5422
rect 9162 5448 9225 5451
rect 9246 5451 9254 5478
rect 9273 5451 9310 5452
rect 9246 5448 9310 5451
rect 9162 5442 9310 5448
rect 9162 5422 9171 5442
rect 9191 5422 9281 5442
rect 9301 5422 9310 5442
rect 8966 5413 9062 5415
rect 9162 5412 9310 5422
rect 9369 5442 9406 5452
rect 9481 5451 9518 5452
rect 9462 5449 9518 5451
rect 9369 5422 9377 5442
rect 9397 5422 9406 5442
rect 9218 5411 9254 5412
rect 9066 5280 9103 5281
rect 9369 5280 9406 5422
rect 9431 5442 9518 5449
rect 9431 5439 9489 5442
rect 9431 5419 9436 5439
rect 9457 5422 9489 5439
rect 9509 5422 9518 5442
rect 9457 5419 9518 5422
rect 9431 5412 9518 5419
rect 9577 5442 9614 5452
rect 9577 5422 9585 5442
rect 9605 5422 9614 5442
rect 9431 5411 9462 5412
rect 9577 5343 9614 5422
rect 9644 5451 9675 5504
rect 9888 5497 9903 5505
rect 9943 5497 9953 5534
rect 9888 5488 9953 5497
rect 10101 5495 10166 5516
rect 10101 5477 10126 5495
rect 10144 5477 10166 5495
rect 9694 5451 9731 5452
rect 9644 5442 9731 5451
rect 9644 5422 9702 5442
rect 9722 5422 9731 5442
rect 9644 5412 9731 5422
rect 9790 5442 9827 5452
rect 9790 5422 9798 5442
rect 9818 5422 9827 5442
rect 9644 5411 9675 5412
rect 9639 5343 9749 5356
rect 9790 5343 9827 5422
rect 10101 5401 10166 5477
rect 9577 5341 9827 5343
rect 9577 5338 9678 5341
rect 9577 5319 9642 5338
rect 9639 5311 9642 5319
rect 9671 5311 9678 5338
rect 9706 5314 9716 5341
rect 9745 5319 9827 5341
rect 9850 5366 10167 5401
rect 9745 5314 9749 5319
rect 9706 5311 9749 5314
rect 9639 5297 9749 5311
rect 9065 5279 9406 5280
rect 8990 5277 9406 5279
rect 9850 5277 9890 5366
rect 10101 5339 10166 5366
rect 10101 5321 10124 5339
rect 10142 5321 10166 5339
rect 10101 5301 10166 5321
rect 8987 5274 9890 5277
rect 8987 5254 8993 5274
rect 9013 5254 9890 5274
rect 8987 5250 9890 5254
rect 9850 5247 9890 5250
rect 10102 5240 10167 5261
rect 8320 5232 8981 5233
rect 8320 5225 9254 5232
rect 8320 5224 9226 5225
rect 8320 5204 9171 5224
rect 9203 5205 9226 5224
rect 9251 5205 9254 5225
rect 9203 5204 9254 5205
rect 8320 5197 9254 5204
rect 7919 5155 8087 5156
rect 8322 5155 8361 5197
rect 9150 5195 9254 5197
rect 9219 5193 9254 5195
rect 10102 5222 10126 5240
rect 10144 5222 10167 5240
rect 10102 5175 10167 5222
rect 7919 5129 8363 5155
rect 7919 5127 8087 5129
rect 7919 4776 7946 5127
rect 8322 5123 8363 5129
rect 7986 4916 8050 4928
rect 8326 4924 8363 5123
rect 8825 5150 8897 5167
rect 8825 5111 8833 5150
rect 8878 5111 8897 5150
rect 8591 5013 8702 5028
rect 8591 5011 8633 5013
rect 8591 4991 8598 5011
rect 8617 4991 8633 5011
rect 8591 4983 8633 4991
rect 8661 5011 8702 5013
rect 8661 4991 8675 5011
rect 8694 4991 8702 5011
rect 8661 4983 8702 4991
rect 8591 4977 8702 4983
rect 8534 4955 8783 4977
rect 8534 4924 8571 4955
rect 8747 4953 8783 4955
rect 8747 4924 8784 4953
rect 7986 4915 8021 4916
rect 7963 4910 8021 4915
rect 7963 4890 7966 4910
rect 7986 4896 8021 4910
rect 8041 4896 8050 4916
rect 7986 4888 8050 4896
rect 8012 4887 8050 4888
rect 8013 4886 8050 4887
rect 8116 4920 8152 4921
rect 8224 4920 8260 4921
rect 8116 4912 8260 4920
rect 8116 4892 8124 4912
rect 8144 4892 8232 4912
rect 8252 4892 8260 4912
rect 8116 4886 8260 4892
rect 8326 4916 8364 4924
rect 8432 4920 8468 4921
rect 8326 4896 8335 4916
rect 8355 4896 8364 4916
rect 8326 4887 8364 4896
rect 8383 4913 8468 4920
rect 8383 4893 8390 4913
rect 8411 4912 8468 4913
rect 8411 4893 8440 4912
rect 8383 4892 8440 4893
rect 8460 4892 8468 4912
rect 8326 4886 8363 4887
rect 8383 4886 8468 4892
rect 8534 4916 8572 4924
rect 8645 4920 8681 4921
rect 8534 4896 8543 4916
rect 8563 4896 8572 4916
rect 8534 4887 8572 4896
rect 8596 4912 8681 4920
rect 8596 4892 8653 4912
rect 8673 4892 8681 4912
rect 8534 4886 8571 4887
rect 8596 4886 8681 4892
rect 8747 4916 8785 4924
rect 8747 4896 8756 4916
rect 8776 4896 8785 4916
rect 8747 4887 8785 4896
rect 8825 4901 8897 5111
rect 8967 5145 10167 5175
rect 8967 5144 9411 5145
rect 8967 5142 9135 5144
rect 8825 4887 8908 4901
rect 8747 4886 8784 4887
rect 8170 4865 8206 4886
rect 8596 4865 8627 4886
rect 8825 4865 8842 4887
rect 8003 4861 8103 4865
rect 8003 4857 8065 4861
rect 8003 4831 8010 4857
rect 8036 4835 8065 4857
rect 8091 4835 8103 4861
rect 8036 4831 8103 4835
rect 8003 4828 8103 4831
rect 8171 4828 8206 4865
rect 8268 4862 8627 4865
rect 8268 4857 8490 4862
rect 8268 4833 8281 4857
rect 8305 4838 8490 4857
rect 8514 4838 8627 4862
rect 8305 4833 8627 4838
rect 8268 4829 8627 4833
rect 8694 4857 8842 4865
rect 8694 4837 8705 4857
rect 8725 4854 8842 4857
rect 8895 4854 8908 4887
rect 8725 4837 8908 4854
rect 8694 4830 8908 4837
rect 8694 4829 8735 4830
rect 8825 4829 8908 4830
rect 8170 4803 8206 4828
rect 8018 4776 8055 4777
rect 8114 4776 8151 4777
rect 8170 4776 8177 4803
rect 7918 4767 8056 4776
rect 7918 4747 8027 4767
rect 8047 4747 8056 4767
rect 7918 4740 8056 4747
rect 8114 4773 8177 4776
rect 8198 4776 8206 4803
rect 8225 4776 8262 4777
rect 8198 4773 8262 4776
rect 8114 4767 8262 4773
rect 8114 4747 8123 4767
rect 8143 4747 8233 4767
rect 8253 4747 8262 4767
rect 7918 4738 8014 4740
rect 8114 4737 8262 4747
rect 8321 4767 8358 4777
rect 8433 4776 8470 4777
rect 8414 4774 8470 4776
rect 8321 4747 8329 4767
rect 8349 4747 8358 4767
rect 8170 4736 8206 4737
rect 8018 4605 8055 4606
rect 8321 4605 8358 4747
rect 8383 4767 8470 4774
rect 8383 4764 8441 4767
rect 8383 4744 8388 4764
rect 8409 4747 8441 4764
rect 8461 4747 8470 4767
rect 8409 4744 8470 4747
rect 8383 4737 8470 4744
rect 8529 4767 8566 4777
rect 8529 4747 8537 4767
rect 8557 4747 8566 4767
rect 8383 4736 8414 4737
rect 8529 4668 8566 4747
rect 8596 4776 8627 4829
rect 8833 4796 8847 4829
rect 8900 4796 8908 4829
rect 8833 4790 8908 4796
rect 8833 4785 8903 4790
rect 8646 4776 8683 4777
rect 8596 4767 8683 4776
rect 8596 4747 8654 4767
rect 8674 4747 8683 4767
rect 8596 4737 8683 4747
rect 8742 4767 8779 4777
rect 8967 4772 8994 5142
rect 9034 4912 9098 4924
rect 9374 4920 9411 5144
rect 9882 5125 9946 5127
rect 9878 5113 9946 5125
rect 9878 5080 9889 5113
rect 9929 5080 9946 5113
rect 9878 5070 9946 5080
rect 9639 5009 9750 5024
rect 9639 5007 9681 5009
rect 9639 4987 9646 5007
rect 9665 4987 9681 5007
rect 9639 4979 9681 4987
rect 9709 5007 9750 5009
rect 9709 4987 9723 5007
rect 9742 4987 9750 5007
rect 9709 4979 9750 4987
rect 9639 4973 9750 4979
rect 9582 4951 9831 4973
rect 9582 4920 9619 4951
rect 9795 4949 9831 4951
rect 9795 4920 9832 4949
rect 9034 4911 9069 4912
rect 9011 4906 9069 4911
rect 9011 4886 9014 4906
rect 9034 4892 9069 4906
rect 9089 4892 9098 4912
rect 9034 4884 9098 4892
rect 9060 4883 9098 4884
rect 9061 4882 9098 4883
rect 9164 4916 9200 4917
rect 9272 4916 9308 4917
rect 9164 4908 9308 4916
rect 9164 4888 9172 4908
rect 9192 4888 9280 4908
rect 9300 4888 9308 4908
rect 9164 4882 9308 4888
rect 9374 4912 9412 4920
rect 9480 4916 9516 4917
rect 9374 4892 9383 4912
rect 9403 4892 9412 4912
rect 9374 4883 9412 4892
rect 9431 4909 9516 4916
rect 9431 4889 9438 4909
rect 9459 4908 9516 4909
rect 9459 4889 9488 4908
rect 9431 4888 9488 4889
rect 9508 4888 9516 4908
rect 9374 4882 9411 4883
rect 9431 4882 9516 4888
rect 9582 4912 9620 4920
rect 9693 4916 9729 4917
rect 9582 4892 9591 4912
rect 9611 4892 9620 4912
rect 9582 4883 9620 4892
rect 9644 4908 9729 4916
rect 9644 4888 9701 4908
rect 9721 4888 9729 4908
rect 9582 4882 9619 4883
rect 9644 4882 9729 4888
rect 9795 4912 9833 4920
rect 9795 4892 9804 4912
rect 9824 4892 9833 4912
rect 9795 4883 9833 4892
rect 9882 4886 9946 5070
rect 10102 4944 10167 5145
rect 10102 4926 10124 4944
rect 10142 4926 10167 4944
rect 10102 4907 10167 4926
rect 9795 4882 9832 4883
rect 9218 4861 9254 4882
rect 9644 4861 9675 4882
rect 9882 4877 9890 4886
rect 9879 4861 9890 4877
rect 9051 4857 9151 4861
rect 9051 4853 9113 4857
rect 9051 4827 9058 4853
rect 9084 4831 9113 4853
rect 9139 4831 9151 4857
rect 9084 4827 9151 4831
rect 9051 4824 9151 4827
rect 9219 4824 9254 4861
rect 9316 4858 9675 4861
rect 9316 4853 9538 4858
rect 9316 4829 9329 4853
rect 9353 4834 9538 4853
rect 9562 4834 9675 4858
rect 9353 4829 9675 4834
rect 9316 4825 9675 4829
rect 9742 4853 9890 4861
rect 9742 4833 9753 4853
rect 9773 4844 9890 4853
rect 9939 4877 9946 4886
rect 9939 4844 9947 4877
rect 9773 4833 9947 4844
rect 9742 4826 9947 4833
rect 9742 4825 9783 4826
rect 9218 4799 9254 4824
rect 9066 4772 9103 4773
rect 9162 4772 9199 4773
rect 9218 4772 9225 4799
rect 8742 4747 8750 4767
rect 8770 4747 8779 4767
rect 8596 4736 8627 4737
rect 8591 4668 8701 4681
rect 8742 4668 8779 4747
rect 8966 4763 9104 4772
rect 8966 4743 9075 4763
rect 9095 4743 9104 4763
rect 8966 4736 9104 4743
rect 9162 4769 9225 4772
rect 9246 4772 9254 4799
rect 9273 4772 9310 4773
rect 9246 4769 9310 4772
rect 9162 4763 9310 4769
rect 9162 4743 9171 4763
rect 9191 4743 9281 4763
rect 9301 4743 9310 4763
rect 8966 4734 9062 4736
rect 9162 4733 9310 4743
rect 9369 4763 9406 4773
rect 9481 4772 9518 4773
rect 9462 4770 9518 4772
rect 9369 4743 9377 4763
rect 9397 4743 9406 4763
rect 9218 4732 9254 4733
rect 8529 4666 8779 4668
rect 8529 4663 8630 4666
rect 8529 4644 8594 4663
rect 8591 4636 8594 4644
rect 8623 4636 8630 4663
rect 8658 4639 8668 4666
rect 8697 4644 8779 4666
rect 8697 4639 8701 4644
rect 8658 4636 8701 4639
rect 8591 4622 8701 4636
rect 8017 4604 8358 4605
rect 7942 4599 8358 4604
rect 9066 4601 9103 4602
rect 9369 4601 9406 4743
rect 9431 4763 9518 4770
rect 9431 4760 9489 4763
rect 9431 4740 9436 4760
rect 9457 4743 9489 4760
rect 9509 4743 9518 4763
rect 9457 4740 9518 4743
rect 9431 4733 9518 4740
rect 9577 4763 9614 4773
rect 9577 4743 9585 4763
rect 9605 4743 9614 4763
rect 9431 4732 9462 4733
rect 9577 4664 9614 4743
rect 9644 4772 9675 4825
rect 9879 4823 9947 4826
rect 9879 4781 9891 4823
rect 9940 4781 9947 4823
rect 9694 4772 9731 4773
rect 9644 4763 9731 4772
rect 9644 4743 9702 4763
rect 9722 4743 9731 4763
rect 9644 4733 9731 4743
rect 9790 4763 9827 4773
rect 9879 4768 9947 4781
rect 10102 4845 10167 4862
rect 10102 4827 10126 4845
rect 10144 4827 10167 4845
rect 9790 4743 9798 4763
rect 9818 4743 9827 4763
rect 9644 4732 9675 4733
rect 9639 4664 9749 4677
rect 9790 4664 9827 4743
rect 10102 4688 10167 4827
rect 10102 4682 10124 4688
rect 9577 4662 9827 4664
rect 9577 4659 9678 4662
rect 9577 4640 9642 4659
rect 9639 4632 9642 4640
rect 9671 4632 9678 4659
rect 9706 4635 9716 4662
rect 9745 4640 9827 4662
rect 9856 4670 10124 4682
rect 10142 4670 10167 4688
rect 9856 4647 10167 4670
rect 9856 4646 9911 4647
rect 9745 4635 9749 4640
rect 9706 4632 9749 4635
rect 9639 4618 9749 4632
rect 9065 4600 9406 4601
rect 7942 4579 7945 4599
rect 7965 4579 8358 4599
rect 8990 4599 9406 4600
rect 9856 4599 9899 4646
rect 8990 4595 9899 4599
rect 8309 4546 8354 4579
rect 8990 4575 8993 4595
rect 9013 4575 9899 4595
rect 9367 4570 9899 4575
rect 10107 4589 10166 4611
rect 10107 4571 10126 4589
rect 10144 4571 10166 4589
rect 9155 4546 9254 4548
rect 8309 4536 9254 4546
rect 8309 4510 9177 4536
rect 8310 4509 9177 4510
rect 9155 4498 9177 4509
rect 9202 4501 9221 4536
rect 9246 4501 9254 4536
rect 9202 4498 9254 4501
rect 10107 4500 10166 4571
rect 9155 4490 9254 4498
rect 9181 4489 9253 4490
rect 8835 4463 8902 4482
rect 8835 4442 8852 4463
rect 8833 4397 8852 4442
rect 8882 4442 8902 4463
rect 8882 4397 8903 4442
rect 9372 4439 9413 4441
rect 9644 4439 9748 4441
rect 10104 4439 10168 4500
rect 8833 4189 8903 4397
rect 8965 4404 10168 4439
rect 8965 4390 8993 4404
rect 8967 4259 8993 4390
rect 9372 4401 10168 4404
rect 7720 4097 7802 4117
rect 7720 4074 7748 4097
rect 7774 4074 7802 4097
rect 7720 4012 7802 4074
rect 7724 3977 7802 4012
rect 8825 4138 8905 4189
rect 8825 4112 8841 4138
rect 8881 4112 8905 4138
rect 8825 4093 8905 4112
rect 8825 4067 8844 4093
rect 8884 4067 8905 4093
rect 8825 4040 8905 4067
rect 8825 4014 8848 4040
rect 8888 4014 8905 4040
rect 8825 4003 8905 4014
rect 8967 4004 8994 4259
rect 9372 4251 9413 4401
rect 9644 4395 9748 4401
rect 10104 4398 10168 4401
rect 9839 4339 9960 4357
rect 9839 4337 9910 4339
rect 9839 4296 9854 4337
rect 9891 4298 9910 4337
rect 9947 4298 9960 4339
rect 9891 4296 9960 4298
rect 9839 4286 9960 4296
rect 9034 4144 9098 4156
rect 9374 4152 9411 4251
rect 9639 4241 9750 4254
rect 9639 4239 9681 4241
rect 9639 4219 9646 4239
rect 9665 4219 9681 4239
rect 9639 4211 9681 4219
rect 9709 4239 9750 4241
rect 9709 4219 9723 4239
rect 9742 4219 9750 4239
rect 9709 4211 9750 4219
rect 9639 4205 9750 4211
rect 9582 4183 9831 4205
rect 9582 4152 9619 4183
rect 9795 4181 9831 4183
rect 9795 4152 9832 4181
rect 9034 4143 9069 4144
rect 9011 4138 9069 4143
rect 9011 4118 9014 4138
rect 9034 4124 9069 4138
rect 9089 4124 9098 4144
rect 9034 4116 9098 4124
rect 9060 4115 9098 4116
rect 9061 4114 9098 4115
rect 9164 4148 9200 4149
rect 9272 4148 9308 4149
rect 9164 4140 9308 4148
rect 9164 4120 9172 4140
rect 9192 4120 9280 4140
rect 9300 4120 9308 4140
rect 9164 4114 9308 4120
rect 9374 4144 9412 4152
rect 9480 4148 9516 4149
rect 9374 4124 9383 4144
rect 9403 4124 9412 4144
rect 9374 4115 9412 4124
rect 9431 4141 9516 4148
rect 9431 4121 9438 4141
rect 9459 4140 9516 4141
rect 9459 4121 9488 4140
rect 9431 4120 9488 4121
rect 9508 4120 9516 4140
rect 9374 4114 9411 4115
rect 9431 4114 9516 4120
rect 9582 4144 9620 4152
rect 9693 4148 9729 4149
rect 9582 4124 9591 4144
rect 9611 4124 9620 4144
rect 9582 4115 9620 4124
rect 9644 4140 9729 4148
rect 9644 4120 9701 4140
rect 9721 4120 9729 4140
rect 9582 4114 9619 4115
rect 9644 4114 9729 4120
rect 9795 4144 9833 4152
rect 9795 4124 9804 4144
rect 9824 4124 9833 4144
rect 9888 4134 9953 4286
rect 10106 4260 10161 4398
rect 9795 4115 9833 4124
rect 9886 4127 9953 4134
rect 9795 4114 9832 4115
rect 9218 4093 9254 4114
rect 9644 4093 9675 4114
rect 9886 4106 9903 4127
rect 9939 4106 9953 4127
rect 10105 4147 10161 4260
rect 10105 4129 10124 4147
rect 10142 4129 10161 4147
rect 10105 4109 10161 4129
rect 9886 4093 9953 4106
rect 9051 4089 9151 4093
rect 9051 4085 9113 4089
rect 9051 4059 9058 4085
rect 9084 4063 9113 4085
rect 9139 4063 9151 4089
rect 9084 4059 9151 4063
rect 9051 4056 9151 4059
rect 9219 4056 9254 4093
rect 9316 4090 9675 4093
rect 9316 4085 9538 4090
rect 9316 4061 9329 4085
rect 9353 4066 9538 4085
rect 9562 4066 9675 4090
rect 9353 4061 9675 4066
rect 9316 4057 9675 4061
rect 9742 4087 9953 4093
rect 9742 4085 9903 4087
rect 9742 4065 9753 4085
rect 9773 4065 9903 4085
rect 9742 4058 9903 4065
rect 9742 4057 9783 4058
rect 9218 4031 9254 4056
rect 9066 4004 9103 4005
rect 9162 4004 9199 4005
rect 9218 4004 9225 4031
rect 8966 3995 9104 4004
rect 7724 3461 7786 3977
rect 8966 3975 9075 3995
rect 9095 3975 9104 3995
rect 8966 3968 9104 3975
rect 9162 4001 9225 4004
rect 9246 4004 9254 4031
rect 9273 4004 9310 4005
rect 9246 4001 9310 4004
rect 9162 3995 9310 4001
rect 9162 3975 9171 3995
rect 9191 3975 9281 3995
rect 9301 3975 9310 3995
rect 8966 3966 9062 3968
rect 9162 3965 9310 3975
rect 9369 3995 9406 4005
rect 9481 4004 9518 4005
rect 9462 4002 9518 4004
rect 9369 3975 9377 3995
rect 9397 3975 9406 3995
rect 9218 3964 9254 3965
rect 9066 3833 9103 3834
rect 9369 3833 9406 3975
rect 9431 3995 9518 4002
rect 9431 3992 9489 3995
rect 9431 3972 9436 3992
rect 9457 3975 9489 3992
rect 9509 3975 9518 3995
rect 9457 3972 9518 3975
rect 9431 3965 9518 3972
rect 9577 3995 9614 4005
rect 9577 3975 9585 3995
rect 9605 3975 9614 3995
rect 9431 3964 9462 3965
rect 9577 3896 9614 3975
rect 9644 4004 9675 4057
rect 9888 4050 9903 4058
rect 9943 4050 9953 4087
rect 9888 4041 9953 4050
rect 10101 4048 10166 4069
rect 10101 4030 10126 4048
rect 10144 4030 10166 4048
rect 9694 4004 9731 4005
rect 9644 3995 9731 4004
rect 9644 3975 9702 3995
rect 9722 3975 9731 3995
rect 9644 3965 9731 3975
rect 9790 3995 9827 4005
rect 9790 3975 9798 3995
rect 9818 3975 9827 3995
rect 9644 3964 9675 3965
rect 9639 3896 9749 3909
rect 9790 3896 9827 3975
rect 10101 3954 10166 4030
rect 9577 3894 9827 3896
rect 9577 3891 9678 3894
rect 9577 3872 9642 3891
rect 9639 3864 9642 3872
rect 9671 3864 9678 3891
rect 9706 3867 9716 3894
rect 9745 3872 9827 3894
rect 9850 3919 10167 3954
rect 9745 3867 9749 3872
rect 9706 3864 9749 3867
rect 9639 3850 9749 3864
rect 9065 3832 9406 3833
rect 8990 3830 9406 3832
rect 9850 3830 9890 3919
rect 10101 3892 10166 3919
rect 10101 3874 10124 3892
rect 10142 3874 10166 3892
rect 10101 3854 10166 3874
rect 8987 3827 9890 3830
rect 8987 3807 8993 3827
rect 9013 3807 9890 3827
rect 8987 3803 9890 3807
rect 9850 3800 9890 3803
rect 10102 3793 10167 3814
rect 8320 3785 8981 3786
rect 8320 3778 9254 3785
rect 8320 3777 9226 3778
rect 8320 3757 9171 3777
rect 9203 3758 9226 3777
rect 9251 3758 9254 3778
rect 9203 3757 9254 3758
rect 8320 3750 9254 3757
rect 7919 3708 8087 3709
rect 8322 3708 8361 3750
rect 9150 3748 9254 3750
rect 9219 3746 9254 3748
rect 10102 3775 10126 3793
rect 10144 3775 10167 3793
rect 10102 3728 10167 3775
rect 7919 3682 8363 3708
rect 7919 3680 8087 3682
rect 7721 3377 7790 3461
rect 7719 2898 7790 3377
rect 7919 3329 7946 3680
rect 8322 3676 8363 3682
rect 7986 3469 8050 3481
rect 8326 3477 8363 3676
rect 8825 3703 8897 3720
rect 8825 3664 8833 3703
rect 8878 3664 8897 3703
rect 8591 3566 8702 3581
rect 8591 3564 8633 3566
rect 8591 3544 8598 3564
rect 8617 3544 8633 3564
rect 8591 3536 8633 3544
rect 8661 3564 8702 3566
rect 8661 3544 8675 3564
rect 8694 3544 8702 3564
rect 8661 3536 8702 3544
rect 8591 3530 8702 3536
rect 8534 3508 8783 3530
rect 8534 3477 8571 3508
rect 8747 3506 8783 3508
rect 8747 3477 8784 3506
rect 7986 3468 8021 3469
rect 7963 3463 8021 3468
rect 7963 3443 7966 3463
rect 7986 3449 8021 3463
rect 8041 3449 8050 3469
rect 7986 3441 8050 3449
rect 8012 3440 8050 3441
rect 8013 3439 8050 3440
rect 8116 3473 8152 3474
rect 8224 3473 8260 3474
rect 8116 3465 8260 3473
rect 8116 3445 8124 3465
rect 8144 3445 8232 3465
rect 8252 3445 8260 3465
rect 8116 3439 8260 3445
rect 8326 3469 8364 3477
rect 8432 3473 8468 3474
rect 8326 3449 8335 3469
rect 8355 3449 8364 3469
rect 8326 3440 8364 3449
rect 8383 3466 8468 3473
rect 8383 3446 8390 3466
rect 8411 3465 8468 3466
rect 8411 3446 8440 3465
rect 8383 3445 8440 3446
rect 8460 3445 8468 3465
rect 8326 3439 8363 3440
rect 8383 3439 8468 3445
rect 8534 3469 8572 3477
rect 8645 3473 8681 3474
rect 8534 3449 8543 3469
rect 8563 3449 8572 3469
rect 8534 3440 8572 3449
rect 8596 3465 8681 3473
rect 8596 3445 8653 3465
rect 8673 3445 8681 3465
rect 8534 3439 8571 3440
rect 8596 3439 8681 3445
rect 8747 3469 8785 3477
rect 8747 3449 8756 3469
rect 8776 3449 8785 3469
rect 8747 3440 8785 3449
rect 8825 3454 8897 3664
rect 8967 3698 10167 3728
rect 8967 3697 9411 3698
rect 8967 3695 9135 3697
rect 8825 3440 8908 3454
rect 8747 3439 8784 3440
rect 8170 3418 8206 3439
rect 8596 3418 8627 3439
rect 8825 3418 8842 3440
rect 8003 3414 8103 3418
rect 8003 3410 8065 3414
rect 8003 3384 8010 3410
rect 8036 3388 8065 3410
rect 8091 3388 8103 3414
rect 8036 3384 8103 3388
rect 8003 3381 8103 3384
rect 8171 3381 8206 3418
rect 8268 3415 8627 3418
rect 8268 3410 8490 3415
rect 8268 3386 8281 3410
rect 8305 3391 8490 3410
rect 8514 3391 8627 3415
rect 8305 3386 8627 3391
rect 8268 3382 8627 3386
rect 8694 3410 8842 3418
rect 8694 3390 8705 3410
rect 8725 3407 8842 3410
rect 8895 3407 8908 3440
rect 8725 3390 8908 3407
rect 8694 3383 8908 3390
rect 8694 3382 8735 3383
rect 8825 3382 8908 3383
rect 8170 3356 8206 3381
rect 8018 3329 8055 3330
rect 8114 3329 8151 3330
rect 8170 3329 8177 3356
rect 7918 3320 8056 3329
rect 7918 3300 8027 3320
rect 8047 3300 8056 3320
rect 7918 3293 8056 3300
rect 8114 3326 8177 3329
rect 8198 3329 8206 3356
rect 8225 3329 8262 3330
rect 8198 3326 8262 3329
rect 8114 3320 8262 3326
rect 8114 3300 8123 3320
rect 8143 3300 8233 3320
rect 8253 3300 8262 3320
rect 7918 3291 8014 3293
rect 8114 3290 8262 3300
rect 8321 3320 8358 3330
rect 8433 3329 8470 3330
rect 8414 3327 8470 3329
rect 8321 3300 8329 3320
rect 8349 3300 8358 3320
rect 8170 3289 8206 3290
rect 8018 3158 8055 3159
rect 8321 3158 8358 3300
rect 8383 3320 8470 3327
rect 8383 3317 8441 3320
rect 8383 3297 8388 3317
rect 8409 3300 8441 3317
rect 8461 3300 8470 3320
rect 8409 3297 8470 3300
rect 8383 3290 8470 3297
rect 8529 3320 8566 3330
rect 8529 3300 8537 3320
rect 8557 3300 8566 3320
rect 8383 3289 8414 3290
rect 8529 3221 8566 3300
rect 8596 3329 8627 3382
rect 8833 3349 8847 3382
rect 8900 3349 8908 3382
rect 8833 3343 8908 3349
rect 8833 3338 8903 3343
rect 8646 3329 8683 3330
rect 8596 3320 8683 3329
rect 8596 3300 8654 3320
rect 8674 3300 8683 3320
rect 8596 3290 8683 3300
rect 8742 3320 8779 3330
rect 8967 3325 8994 3695
rect 9034 3465 9098 3477
rect 9374 3473 9411 3697
rect 9882 3678 9946 3680
rect 9878 3666 9946 3678
rect 9878 3633 9889 3666
rect 9929 3633 9946 3666
rect 9878 3623 9946 3633
rect 9639 3562 9750 3577
rect 9639 3560 9681 3562
rect 9639 3540 9646 3560
rect 9665 3540 9681 3560
rect 9639 3532 9681 3540
rect 9709 3560 9750 3562
rect 9709 3540 9723 3560
rect 9742 3540 9750 3560
rect 9709 3532 9750 3540
rect 9639 3526 9750 3532
rect 9582 3504 9831 3526
rect 9582 3473 9619 3504
rect 9795 3502 9831 3504
rect 9795 3473 9832 3502
rect 9034 3464 9069 3465
rect 9011 3459 9069 3464
rect 9011 3439 9014 3459
rect 9034 3445 9069 3459
rect 9089 3445 9098 3465
rect 9034 3437 9098 3445
rect 9060 3436 9098 3437
rect 9061 3435 9098 3436
rect 9164 3469 9200 3470
rect 9272 3469 9308 3470
rect 9164 3461 9308 3469
rect 9164 3441 9172 3461
rect 9192 3441 9280 3461
rect 9300 3441 9308 3461
rect 9164 3435 9308 3441
rect 9374 3465 9412 3473
rect 9480 3469 9516 3470
rect 9374 3445 9383 3465
rect 9403 3445 9412 3465
rect 9374 3436 9412 3445
rect 9431 3462 9516 3469
rect 9431 3442 9438 3462
rect 9459 3461 9516 3462
rect 9459 3442 9488 3461
rect 9431 3441 9488 3442
rect 9508 3441 9516 3461
rect 9374 3435 9411 3436
rect 9431 3435 9516 3441
rect 9582 3465 9620 3473
rect 9693 3469 9729 3470
rect 9582 3445 9591 3465
rect 9611 3445 9620 3465
rect 9582 3436 9620 3445
rect 9644 3461 9729 3469
rect 9644 3441 9701 3461
rect 9721 3441 9729 3461
rect 9582 3435 9619 3436
rect 9644 3435 9729 3441
rect 9795 3465 9833 3473
rect 9795 3445 9804 3465
rect 9824 3445 9833 3465
rect 9795 3436 9833 3445
rect 9882 3439 9946 3623
rect 10102 3497 10167 3698
rect 10102 3479 10124 3497
rect 10142 3479 10167 3497
rect 10102 3460 10167 3479
rect 9795 3435 9832 3436
rect 9218 3414 9254 3435
rect 9644 3414 9675 3435
rect 9882 3430 9890 3439
rect 9879 3414 9890 3430
rect 9051 3410 9151 3414
rect 9051 3406 9113 3410
rect 9051 3380 9058 3406
rect 9084 3384 9113 3406
rect 9139 3384 9151 3410
rect 9084 3380 9151 3384
rect 9051 3377 9151 3380
rect 9219 3377 9254 3414
rect 9316 3411 9675 3414
rect 9316 3406 9538 3411
rect 9316 3382 9329 3406
rect 9353 3387 9538 3406
rect 9562 3387 9675 3411
rect 9353 3382 9675 3387
rect 9316 3378 9675 3382
rect 9742 3406 9890 3414
rect 9742 3386 9753 3406
rect 9773 3397 9890 3406
rect 9939 3430 9946 3439
rect 9939 3397 9947 3430
rect 9773 3386 9947 3397
rect 9742 3379 9947 3386
rect 9742 3378 9783 3379
rect 9218 3352 9254 3377
rect 9066 3325 9103 3326
rect 9162 3325 9199 3326
rect 9218 3325 9225 3352
rect 8742 3300 8750 3320
rect 8770 3300 8779 3320
rect 8596 3289 8627 3290
rect 8591 3221 8701 3234
rect 8742 3221 8779 3300
rect 8966 3316 9104 3325
rect 8966 3296 9075 3316
rect 9095 3296 9104 3316
rect 8966 3289 9104 3296
rect 9162 3322 9225 3325
rect 9246 3325 9254 3352
rect 9273 3325 9310 3326
rect 9246 3322 9310 3325
rect 9162 3316 9310 3322
rect 9162 3296 9171 3316
rect 9191 3296 9281 3316
rect 9301 3296 9310 3316
rect 8966 3287 9062 3289
rect 9162 3286 9310 3296
rect 9369 3316 9406 3326
rect 9481 3325 9518 3326
rect 9462 3323 9518 3325
rect 9369 3296 9377 3316
rect 9397 3296 9406 3316
rect 9218 3285 9254 3286
rect 8529 3219 8779 3221
rect 8529 3216 8630 3219
rect 8529 3197 8594 3216
rect 8591 3189 8594 3197
rect 8623 3189 8630 3216
rect 8658 3192 8668 3219
rect 8697 3197 8779 3219
rect 8697 3192 8701 3197
rect 8658 3189 8701 3192
rect 8591 3175 8701 3189
rect 8017 3157 8358 3158
rect 7942 3152 8358 3157
rect 9066 3154 9103 3155
rect 9369 3154 9406 3296
rect 9431 3316 9518 3323
rect 9431 3313 9489 3316
rect 9431 3293 9436 3313
rect 9457 3296 9489 3313
rect 9509 3296 9518 3316
rect 9457 3293 9518 3296
rect 9431 3286 9518 3293
rect 9577 3316 9614 3326
rect 9577 3296 9585 3316
rect 9605 3296 9614 3316
rect 9431 3285 9462 3286
rect 9577 3217 9614 3296
rect 9644 3325 9675 3378
rect 9879 3376 9947 3379
rect 9879 3334 9891 3376
rect 9940 3334 9947 3376
rect 9694 3325 9731 3326
rect 9644 3316 9731 3325
rect 9644 3296 9702 3316
rect 9722 3296 9731 3316
rect 9644 3286 9731 3296
rect 9790 3316 9827 3326
rect 9879 3321 9947 3334
rect 10102 3398 10167 3415
rect 10102 3380 10126 3398
rect 10144 3380 10167 3398
rect 9790 3296 9798 3316
rect 9818 3296 9827 3316
rect 9644 3285 9675 3286
rect 9639 3217 9749 3230
rect 9790 3217 9827 3296
rect 10102 3241 10167 3380
rect 10102 3235 10124 3241
rect 9577 3215 9827 3217
rect 9577 3212 9678 3215
rect 9577 3193 9642 3212
rect 9639 3185 9642 3193
rect 9671 3185 9678 3212
rect 9706 3188 9716 3215
rect 9745 3193 9827 3215
rect 9856 3223 10124 3235
rect 10142 3223 10167 3241
rect 9856 3200 10167 3223
rect 9856 3199 9911 3200
rect 9745 3188 9749 3193
rect 9706 3185 9749 3188
rect 9639 3171 9749 3185
rect 9065 3153 9406 3154
rect 7942 3132 7945 3152
rect 7965 3132 8358 3152
rect 8990 3152 9406 3153
rect 9856 3152 9899 3199
rect 8990 3148 9899 3152
rect 8309 3099 8354 3132
rect 8990 3128 8993 3148
rect 9013 3128 9899 3148
rect 9367 3123 9899 3128
rect 10107 3142 10166 3164
rect 10107 3124 10126 3142
rect 10144 3124 10166 3142
rect 9155 3099 9254 3101
rect 8309 3089 9254 3099
rect 8309 3063 9177 3089
rect 8310 3062 9177 3063
rect 9155 3051 9177 3062
rect 9202 3054 9221 3089
rect 9246 3054 9254 3089
rect 9202 3051 9254 3054
rect 9155 3043 9254 3051
rect 9181 3042 9253 3043
rect 10107 2994 10166 3124
rect 8829 2964 8905 2988
rect 8829 2898 8841 2964
rect 8895 2898 8905 2964
rect 9373 2919 9414 2921
rect 9645 2919 9749 2921
rect 10107 2919 10168 2994
rect 7719 2848 7791 2898
rect 7288 2576 7624 2580
rect 6514 2572 6614 2576
rect 6514 2568 6576 2572
rect 6514 2542 6521 2568
rect 6547 2546 6576 2568
rect 6602 2546 6614 2572
rect 6547 2542 6614 2546
rect 6514 2539 6614 2542
rect 6682 2539 6717 2576
rect 6779 2573 7138 2576
rect 6779 2568 7001 2573
rect 6779 2544 6792 2568
rect 6816 2549 7001 2568
rect 7025 2549 7138 2573
rect 6816 2544 7138 2549
rect 6779 2540 7138 2544
rect 7205 2568 7624 2576
rect 7205 2548 7216 2568
rect 7236 2548 7624 2568
rect 7205 2541 7624 2548
rect 7205 2540 7246 2541
rect 7288 2540 7624 2541
rect 6681 2514 6717 2539
rect 6529 2487 6566 2488
rect 6625 2487 6662 2488
rect 6681 2487 6688 2514
rect 6429 2478 6567 2487
rect 6429 2458 6538 2478
rect 6558 2458 6567 2478
rect 6429 2451 6567 2458
rect 6625 2484 6688 2487
rect 6709 2487 6717 2514
rect 6736 2487 6773 2488
rect 6709 2484 6773 2487
rect 6625 2478 6773 2484
rect 6625 2458 6634 2478
rect 6654 2458 6744 2478
rect 6764 2458 6773 2478
rect 6429 2449 6525 2451
rect 6625 2448 6773 2458
rect 6832 2478 6869 2488
rect 6944 2487 6981 2488
rect 6925 2485 6981 2487
rect 6832 2458 6840 2478
rect 6860 2458 6869 2478
rect 6681 2447 6717 2448
rect 6529 2316 6566 2317
rect 6832 2316 6869 2458
rect 6894 2478 6981 2485
rect 6894 2475 6952 2478
rect 6894 2455 6899 2475
rect 6920 2458 6952 2475
rect 6972 2458 6981 2478
rect 6920 2455 6981 2458
rect 6894 2448 6981 2455
rect 7040 2478 7077 2488
rect 7040 2458 7048 2478
rect 7068 2458 7077 2478
rect 6894 2447 6925 2448
rect 7040 2379 7077 2458
rect 7107 2487 7138 2540
rect 7532 2504 7624 2540
rect 7157 2487 7194 2488
rect 7107 2478 7194 2487
rect 7107 2458 7165 2478
rect 7185 2458 7194 2478
rect 7107 2448 7194 2458
rect 7253 2478 7290 2488
rect 7253 2458 7261 2478
rect 7281 2458 7290 2478
rect 7107 2447 7138 2448
rect 7102 2379 7212 2392
rect 7253 2379 7290 2458
rect 7040 2377 7290 2379
rect 7040 2374 7141 2377
rect 7040 2355 7105 2374
rect 7102 2347 7105 2355
rect 7134 2347 7141 2374
rect 7169 2350 7179 2377
rect 7208 2355 7290 2377
rect 7208 2350 7212 2355
rect 7169 2347 7212 2350
rect 7102 2333 7212 2347
rect 6528 2315 6869 2316
rect 6453 2310 6869 2315
rect 6453 2290 6456 2310
rect 6476 2290 6869 2310
rect 6613 2246 6718 2249
rect 6612 2223 6718 2246
rect 5732 2221 6233 2223
rect 6374 2221 6723 2223
rect 3846 2200 3883 2221
rect 3846 2163 3857 2200
rect 3874 2163 3883 2200
rect 5732 2215 6723 2221
rect 5732 2210 6684 2215
rect 5732 2189 6643 2210
rect 6663 2194 6684 2210
rect 6704 2194 6723 2215
rect 6663 2189 6723 2194
rect 5732 2164 6723 2189
rect 6208 2163 6390 2164
rect 3846 2153 3883 2163
rect 3692 2110 4086 2130
rect 4106 2110 4109 2130
rect 3693 2105 4109 2110
rect 3693 2104 4034 2105
rect 3350 2073 3460 2087
rect 3350 2070 3393 2073
rect 3350 2065 3354 2070
rect 3272 2043 3354 2065
rect 3383 2043 3393 2070
rect 3421 2046 3428 2073
rect 3457 2065 3460 2073
rect 3457 2046 3522 2065
rect 3421 2043 3522 2046
rect 3272 2041 3522 2043
rect 3272 1962 3309 2041
rect 3350 2028 3460 2041
rect 3424 1972 3455 1973
rect 3272 1942 3281 1962
rect 3301 1942 3309 1962
rect 3272 1932 3309 1942
rect 3368 1962 3455 1972
rect 3368 1942 3377 1962
rect 3397 1942 3455 1962
rect 3368 1933 3455 1942
rect 3368 1932 3405 1933
rect 3424 1880 3455 1933
rect 3485 1962 3522 2041
rect 3637 1972 3668 1973
rect 3485 1942 3494 1962
rect 3514 1942 3522 1962
rect 3485 1932 3522 1942
rect 3581 1965 3668 1972
rect 3581 1962 3642 1965
rect 3581 1942 3590 1962
rect 3610 1945 3642 1962
rect 3663 1945 3668 1965
rect 3610 1942 3668 1945
rect 3581 1935 3668 1942
rect 3693 1962 3730 2104
rect 3996 2103 4033 2104
rect 3845 1972 3881 1973
rect 3693 1942 3702 1962
rect 3722 1942 3730 1962
rect 3581 1933 3637 1935
rect 3581 1932 3618 1933
rect 3693 1932 3730 1942
rect 3789 1962 3937 1972
rect 4037 1969 4133 1971
rect 3789 1942 3798 1962
rect 3818 1942 3908 1962
rect 3928 1942 3937 1962
rect 3789 1936 3937 1942
rect 3789 1933 3853 1936
rect 3789 1932 3826 1933
rect 3845 1906 3853 1933
rect 3874 1933 3937 1936
rect 3995 1962 4133 1969
rect 3995 1942 4004 1962
rect 4024 1942 4133 1962
rect 3995 1933 4133 1942
rect 6762 1934 6793 2290
rect 3874 1906 3881 1933
rect 3900 1932 3937 1933
rect 3996 1932 4033 1933
rect 3845 1881 3881 1906
rect 3316 1879 3357 1880
rect 3236 1874 3357 1879
rect 3187 1872 3357 1874
rect 3187 1861 3326 1872
rect 3187 1838 3210 1861
rect 3236 1852 3326 1861
rect 3346 1852 3357 1872
rect 3236 1844 3357 1852
rect 3424 1876 3783 1880
rect 3424 1871 3746 1876
rect 3424 1847 3537 1871
rect 3561 1852 3746 1871
rect 3770 1852 3783 1876
rect 3561 1847 3783 1852
rect 3424 1844 3783 1847
rect 3845 1844 3880 1881
rect 3948 1878 4048 1881
rect 3948 1874 4015 1878
rect 3948 1848 3960 1874
rect 3986 1852 4015 1874
rect 4041 1852 4048 1878
rect 3986 1848 4048 1852
rect 3948 1844 4048 1848
rect 3236 1838 3244 1844
rect 3187 1830 3244 1838
rect 3424 1823 3455 1844
rect 3845 1823 3881 1844
rect 3267 1822 3304 1823
rect 3266 1813 3304 1822
rect 3266 1793 3275 1813
rect 3295 1793 3304 1813
rect 3266 1785 3304 1793
rect 3370 1817 3455 1823
rect 3480 1822 3517 1823
rect 3370 1797 3378 1817
rect 3398 1797 3455 1817
rect 3370 1789 3455 1797
rect 3479 1813 3517 1822
rect 3479 1793 3488 1813
rect 3508 1793 3517 1813
rect 3370 1788 3406 1789
rect 3479 1785 3517 1793
rect 3583 1817 3668 1823
rect 3688 1822 3725 1823
rect 3583 1797 3591 1817
rect 3611 1816 3668 1817
rect 3611 1797 3640 1816
rect 3583 1796 3640 1797
rect 3661 1796 3668 1816
rect 3583 1789 3668 1796
rect 3687 1813 3725 1822
rect 3687 1793 3696 1813
rect 3716 1793 3725 1813
rect 3583 1788 3619 1789
rect 3687 1785 3725 1793
rect 3791 1817 3935 1823
rect 3791 1797 3799 1817
rect 3819 1797 3907 1817
rect 3927 1797 3935 1817
rect 3791 1789 3935 1797
rect 3791 1788 3827 1789
rect 3899 1788 3935 1789
rect 4001 1822 4038 1823
rect 4001 1821 4039 1822
rect 4001 1813 4065 1821
rect 4001 1793 4010 1813
rect 4030 1799 4065 1813
rect 4085 1799 4088 1819
rect 4030 1794 4088 1799
rect 4030 1793 4065 1794
rect 3267 1756 3304 1785
rect 3268 1754 3304 1756
rect 3480 1754 3517 1785
rect 3268 1732 3517 1754
rect 3349 1726 3460 1732
rect 3349 1718 3390 1726
rect 3349 1698 3357 1718
rect 3376 1698 3390 1718
rect 3349 1696 3390 1698
rect 3418 1718 3460 1726
rect 3418 1698 3434 1718
rect 3453 1698 3460 1718
rect 3418 1696 3460 1698
rect 3349 1681 3460 1696
rect 3688 1670 3725 1785
rect 4001 1781 4065 1793
rect 3681 1664 3728 1670
rect 4105 1666 4132 1933
rect 6680 1905 6793 1934
rect 3964 1664 4132 1666
rect 3681 1638 4132 1664
rect 3681 1503 3728 1638
rect 3964 1637 4132 1638
rect 6681 1596 6717 1905
rect 7541 1791 7622 2504
rect 7721 1939 7791 2848
rect 8829 2878 8905 2898
rect 8829 2841 8846 2878
rect 8890 2841 8905 2878
rect 8966 2884 10168 2919
rect 8966 2870 8994 2884
rect 8829 2825 8905 2841
rect 8834 2669 8904 2825
rect 8968 2739 8994 2870
rect 9373 2881 10168 2884
rect 8826 2618 8906 2669
rect 8826 2592 8842 2618
rect 8882 2592 8906 2618
rect 8826 2573 8906 2592
rect 8826 2547 8845 2573
rect 8885 2547 8906 2573
rect 8826 2520 8906 2547
rect 8826 2494 8849 2520
rect 8889 2494 8906 2520
rect 8826 2483 8906 2494
rect 8968 2484 8995 2739
rect 9373 2731 9414 2881
rect 10107 2869 10168 2881
rect 9840 2819 9961 2837
rect 9840 2817 9911 2819
rect 9840 2776 9855 2817
rect 9892 2778 9911 2817
rect 9948 2778 9961 2819
rect 9892 2776 9961 2778
rect 9840 2766 9961 2776
rect 9645 2736 9749 2745
rect 9035 2624 9099 2636
rect 9375 2632 9412 2731
rect 9640 2721 9751 2736
rect 9640 2719 9682 2721
rect 9640 2699 9647 2719
rect 9666 2699 9682 2719
rect 9640 2691 9682 2699
rect 9710 2719 9751 2721
rect 9710 2699 9724 2719
rect 9743 2699 9751 2719
rect 9710 2691 9751 2699
rect 9640 2685 9751 2691
rect 9583 2663 9832 2685
rect 9583 2632 9620 2663
rect 9796 2661 9832 2663
rect 9796 2632 9833 2661
rect 9035 2623 9070 2624
rect 9012 2618 9070 2623
rect 9012 2598 9015 2618
rect 9035 2604 9070 2618
rect 9090 2604 9099 2624
rect 9035 2596 9099 2604
rect 9061 2595 9099 2596
rect 9062 2594 9099 2595
rect 9165 2628 9201 2629
rect 9273 2628 9309 2629
rect 9165 2620 9309 2628
rect 9165 2600 9173 2620
rect 9193 2600 9281 2620
rect 9301 2600 9309 2620
rect 9165 2594 9309 2600
rect 9375 2624 9413 2632
rect 9481 2628 9517 2629
rect 9375 2604 9384 2624
rect 9404 2604 9413 2624
rect 9375 2595 9413 2604
rect 9432 2621 9517 2628
rect 9432 2601 9439 2621
rect 9460 2620 9517 2621
rect 9460 2601 9489 2620
rect 9432 2600 9489 2601
rect 9509 2600 9517 2620
rect 9375 2594 9412 2595
rect 9432 2594 9517 2600
rect 9583 2624 9621 2632
rect 9694 2628 9730 2629
rect 9583 2604 9592 2624
rect 9612 2604 9621 2624
rect 9583 2595 9621 2604
rect 9645 2620 9730 2628
rect 9645 2600 9702 2620
rect 9722 2600 9730 2620
rect 9583 2594 9620 2595
rect 9645 2594 9730 2600
rect 9796 2624 9834 2632
rect 9796 2604 9805 2624
rect 9825 2604 9834 2624
rect 9889 2614 9954 2766
rect 10107 2740 10162 2869
rect 9796 2595 9834 2604
rect 9887 2607 9954 2614
rect 9796 2594 9833 2595
rect 9219 2573 9255 2594
rect 9645 2573 9676 2594
rect 9887 2586 9904 2607
rect 9940 2586 9954 2607
rect 10106 2627 10162 2740
rect 10106 2609 10125 2627
rect 10143 2609 10162 2627
rect 10106 2589 10162 2609
rect 9887 2573 9954 2586
rect 9052 2569 9152 2573
rect 9052 2565 9114 2569
rect 9052 2539 9059 2565
rect 9085 2543 9114 2565
rect 9140 2543 9152 2569
rect 9085 2539 9152 2543
rect 9052 2536 9152 2539
rect 9220 2536 9255 2573
rect 9317 2570 9676 2573
rect 9317 2565 9539 2570
rect 9317 2541 9330 2565
rect 9354 2546 9539 2565
rect 9563 2546 9676 2570
rect 9354 2541 9676 2546
rect 9317 2537 9676 2541
rect 9743 2567 9954 2573
rect 9743 2565 9904 2567
rect 9743 2545 9754 2565
rect 9774 2545 9904 2565
rect 9743 2538 9904 2545
rect 9743 2537 9784 2538
rect 9219 2511 9255 2536
rect 9067 2484 9104 2485
rect 9163 2484 9200 2485
rect 9219 2484 9226 2511
rect 8967 2475 9105 2484
rect 8967 2455 9076 2475
rect 9096 2455 9105 2475
rect 8967 2448 9105 2455
rect 9163 2481 9226 2484
rect 9247 2484 9255 2511
rect 9274 2484 9311 2485
rect 9247 2481 9311 2484
rect 9163 2475 9311 2481
rect 9163 2455 9172 2475
rect 9192 2455 9282 2475
rect 9302 2455 9311 2475
rect 8967 2446 9063 2448
rect 9163 2445 9311 2455
rect 9370 2475 9407 2485
rect 9482 2484 9519 2485
rect 9463 2482 9519 2484
rect 9370 2455 9378 2475
rect 9398 2455 9407 2475
rect 9219 2444 9255 2445
rect 9067 2313 9104 2314
rect 9370 2313 9407 2455
rect 9432 2475 9519 2482
rect 9432 2472 9490 2475
rect 9432 2452 9437 2472
rect 9458 2455 9490 2472
rect 9510 2455 9519 2475
rect 9458 2452 9519 2455
rect 9432 2445 9519 2452
rect 9578 2475 9615 2485
rect 9578 2455 9586 2475
rect 9606 2455 9615 2475
rect 9432 2444 9463 2445
rect 9578 2376 9615 2455
rect 9645 2484 9676 2537
rect 9889 2530 9904 2538
rect 9944 2530 9954 2567
rect 9889 2521 9954 2530
rect 10102 2528 10167 2549
rect 10102 2510 10127 2528
rect 10145 2510 10167 2528
rect 9695 2484 9732 2485
rect 9645 2475 9732 2484
rect 9645 2455 9703 2475
rect 9723 2455 9732 2475
rect 9645 2445 9732 2455
rect 9791 2475 9828 2485
rect 9791 2455 9799 2475
rect 9819 2455 9828 2475
rect 9645 2444 9676 2445
rect 9640 2376 9750 2389
rect 9791 2376 9828 2455
rect 10102 2434 10167 2510
rect 9578 2374 9828 2376
rect 9578 2371 9679 2374
rect 9578 2352 9643 2371
rect 9640 2344 9643 2352
rect 9672 2344 9679 2371
rect 9707 2347 9717 2374
rect 9746 2352 9828 2374
rect 9851 2399 10168 2434
rect 9746 2347 9750 2352
rect 9707 2344 9750 2347
rect 9640 2330 9750 2344
rect 9066 2312 9407 2313
rect 8991 2310 9407 2312
rect 9851 2310 9891 2399
rect 10102 2372 10167 2399
rect 10102 2354 10125 2372
rect 10143 2354 10167 2372
rect 10102 2334 10167 2354
rect 8988 2307 9891 2310
rect 8988 2287 8994 2307
rect 9014 2287 9891 2307
rect 8988 2283 9891 2287
rect 9851 2280 9891 2283
rect 10103 2273 10168 2294
rect 8321 2265 8982 2266
rect 8321 2258 9255 2265
rect 8321 2257 9227 2258
rect 8321 2237 9172 2257
rect 9204 2238 9227 2257
rect 9252 2238 9255 2258
rect 9204 2237 9255 2238
rect 8321 2230 9255 2237
rect 7920 2188 8088 2189
rect 8323 2188 8362 2230
rect 9151 2228 9255 2230
rect 9220 2226 9255 2228
rect 10103 2255 10127 2273
rect 10145 2255 10168 2273
rect 10103 2208 10168 2255
rect 7920 2162 8364 2188
rect 7920 2160 8088 2162
rect 6681 1573 6685 1596
rect 6709 1573 6717 1596
rect 6881 1574 6980 1578
rect 6681 1552 6717 1573
rect 6681 1529 6685 1552
rect 6709 1529 6717 1552
rect 6681 1525 6717 1529
rect 6877 1568 6980 1574
rect 6877 1530 6903 1568
rect 6928 1533 6947 1568
rect 6972 1533 6980 1568
rect 6928 1530 6980 1533
rect 6877 1522 6980 1530
rect 6877 1521 6979 1522
rect 3679 1454 3738 1503
rect 3679 1426 3697 1454
rect 3725 1426 3738 1454
rect 3679 1416 3738 1426
rect 6473 1443 6641 1444
rect 6877 1443 6924 1521
rect 6473 1417 6924 1443
rect 6473 1415 6641 1417
rect 6473 1042 6500 1415
rect 6670 1367 6756 1376
rect 6670 1349 6689 1367
rect 6741 1349 6756 1367
rect 6670 1345 6756 1349
rect 6540 1182 6604 1194
rect 6540 1181 6575 1182
rect 6517 1176 6575 1181
rect 6517 1156 6520 1176
rect 6540 1162 6575 1176
rect 6595 1162 6604 1182
rect 6540 1154 6604 1162
rect 6566 1153 6604 1154
rect 6567 1152 6604 1153
rect 6670 1186 6706 1187
rect 6726 1186 6756 1345
rect 6877 1305 6924 1417
rect 6880 1190 6917 1305
rect 7145 1279 7256 1294
rect 7145 1277 7187 1279
rect 7145 1257 7152 1277
rect 7171 1257 7187 1277
rect 7145 1249 7187 1257
rect 7215 1277 7256 1279
rect 7215 1257 7229 1277
rect 7248 1257 7256 1277
rect 7215 1249 7256 1257
rect 7145 1243 7256 1249
rect 7088 1221 7337 1243
rect 7088 1190 7125 1221
rect 7301 1219 7337 1221
rect 7301 1190 7338 1219
rect 7542 1206 7621 1791
rect 7718 1339 7797 1939
rect 7920 1809 7947 2160
rect 8323 2156 8364 2162
rect 7987 1949 8051 1961
rect 8327 1957 8364 2156
rect 8826 2183 8898 2200
rect 8826 2144 8834 2183
rect 8879 2144 8898 2183
rect 8592 2046 8703 2061
rect 8592 2044 8634 2046
rect 8592 2024 8599 2044
rect 8618 2024 8634 2044
rect 8592 2016 8634 2024
rect 8662 2044 8703 2046
rect 8662 2024 8676 2044
rect 8695 2024 8703 2044
rect 8662 2016 8703 2024
rect 8592 2010 8703 2016
rect 8535 1988 8784 2010
rect 8535 1957 8572 1988
rect 8748 1986 8784 1988
rect 8748 1957 8785 1986
rect 7987 1948 8022 1949
rect 7964 1943 8022 1948
rect 7964 1923 7967 1943
rect 7987 1929 8022 1943
rect 8042 1929 8051 1949
rect 7987 1921 8051 1929
rect 8013 1920 8051 1921
rect 8014 1919 8051 1920
rect 8117 1953 8153 1954
rect 8225 1953 8261 1954
rect 8117 1945 8261 1953
rect 8117 1925 8125 1945
rect 8145 1925 8233 1945
rect 8253 1925 8261 1945
rect 8117 1919 8261 1925
rect 8327 1949 8365 1957
rect 8433 1953 8469 1954
rect 8327 1929 8336 1949
rect 8356 1929 8365 1949
rect 8327 1920 8365 1929
rect 8384 1946 8469 1953
rect 8384 1926 8391 1946
rect 8412 1945 8469 1946
rect 8412 1926 8441 1945
rect 8384 1925 8441 1926
rect 8461 1925 8469 1945
rect 8327 1919 8364 1920
rect 8384 1919 8469 1925
rect 8535 1949 8573 1957
rect 8646 1953 8682 1954
rect 8535 1929 8544 1949
rect 8564 1929 8573 1949
rect 8535 1920 8573 1929
rect 8597 1945 8682 1953
rect 8597 1925 8654 1945
rect 8674 1925 8682 1945
rect 8535 1919 8572 1920
rect 8597 1919 8682 1925
rect 8748 1949 8786 1957
rect 8748 1929 8757 1949
rect 8777 1929 8786 1949
rect 8748 1920 8786 1929
rect 8826 1934 8898 2144
rect 8968 2178 10168 2208
rect 8968 2177 9412 2178
rect 8968 2175 9136 2177
rect 8826 1920 8909 1934
rect 8748 1919 8785 1920
rect 8171 1898 8207 1919
rect 8597 1898 8628 1919
rect 8826 1898 8843 1920
rect 8004 1894 8104 1898
rect 8004 1890 8066 1894
rect 8004 1864 8011 1890
rect 8037 1868 8066 1890
rect 8092 1868 8104 1894
rect 8037 1864 8104 1868
rect 8004 1861 8104 1864
rect 8172 1861 8207 1898
rect 8269 1895 8628 1898
rect 8269 1890 8491 1895
rect 8269 1866 8282 1890
rect 8306 1871 8491 1890
rect 8515 1871 8628 1895
rect 8306 1866 8628 1871
rect 8269 1862 8628 1866
rect 8695 1890 8843 1898
rect 8695 1870 8706 1890
rect 8726 1887 8843 1890
rect 8896 1887 8909 1920
rect 8726 1870 8909 1887
rect 8695 1863 8909 1870
rect 8695 1862 8736 1863
rect 8826 1862 8909 1863
rect 8171 1836 8207 1861
rect 8019 1809 8056 1810
rect 8115 1809 8152 1810
rect 8171 1809 8178 1836
rect 7919 1800 8057 1809
rect 7919 1780 8028 1800
rect 8048 1780 8057 1800
rect 7919 1773 8057 1780
rect 8115 1806 8178 1809
rect 8199 1809 8207 1836
rect 8226 1809 8263 1810
rect 8199 1806 8263 1809
rect 8115 1800 8263 1806
rect 8115 1780 8124 1800
rect 8144 1780 8234 1800
rect 8254 1780 8263 1800
rect 7919 1771 8015 1773
rect 8115 1770 8263 1780
rect 8322 1800 8359 1810
rect 8434 1809 8471 1810
rect 8415 1807 8471 1809
rect 8322 1780 8330 1800
rect 8350 1780 8359 1800
rect 8171 1769 8207 1770
rect 8019 1638 8056 1639
rect 8322 1638 8359 1780
rect 8384 1800 8471 1807
rect 8384 1797 8442 1800
rect 8384 1777 8389 1797
rect 8410 1780 8442 1797
rect 8462 1780 8471 1800
rect 8410 1777 8471 1780
rect 8384 1770 8471 1777
rect 8530 1800 8567 1810
rect 8530 1780 8538 1800
rect 8558 1780 8567 1800
rect 8384 1769 8415 1770
rect 8530 1701 8567 1780
rect 8597 1809 8628 1862
rect 8834 1829 8848 1862
rect 8901 1829 8909 1862
rect 8834 1823 8909 1829
rect 8834 1818 8904 1823
rect 8647 1809 8684 1810
rect 8597 1800 8684 1809
rect 8597 1780 8655 1800
rect 8675 1780 8684 1800
rect 8597 1770 8684 1780
rect 8743 1800 8780 1810
rect 8968 1805 8995 2175
rect 9035 1945 9099 1957
rect 9375 1953 9412 2177
rect 9883 2158 9947 2160
rect 9879 2146 9947 2158
rect 9879 2113 9890 2146
rect 9930 2113 9947 2146
rect 9879 2103 9947 2113
rect 9640 2042 9751 2057
rect 9640 2040 9682 2042
rect 9640 2020 9647 2040
rect 9666 2020 9682 2040
rect 9640 2012 9682 2020
rect 9710 2040 9751 2042
rect 9710 2020 9724 2040
rect 9743 2020 9751 2040
rect 9710 2012 9751 2020
rect 9640 2006 9751 2012
rect 9583 1984 9832 2006
rect 9583 1953 9620 1984
rect 9796 1982 9832 1984
rect 9796 1953 9833 1982
rect 9035 1944 9070 1945
rect 9012 1939 9070 1944
rect 9012 1919 9015 1939
rect 9035 1925 9070 1939
rect 9090 1925 9099 1945
rect 9035 1917 9099 1925
rect 9061 1916 9099 1917
rect 9062 1915 9099 1916
rect 9165 1949 9201 1950
rect 9273 1949 9309 1950
rect 9165 1941 9309 1949
rect 9165 1921 9173 1941
rect 9193 1921 9281 1941
rect 9301 1921 9309 1941
rect 9165 1915 9309 1921
rect 9375 1945 9413 1953
rect 9481 1949 9517 1950
rect 9375 1925 9384 1945
rect 9404 1925 9413 1945
rect 9375 1916 9413 1925
rect 9432 1942 9517 1949
rect 9432 1922 9439 1942
rect 9460 1941 9517 1942
rect 9460 1922 9489 1941
rect 9432 1921 9489 1922
rect 9509 1921 9517 1941
rect 9375 1915 9412 1916
rect 9432 1915 9517 1921
rect 9583 1945 9621 1953
rect 9694 1949 9730 1950
rect 9583 1925 9592 1945
rect 9612 1925 9621 1945
rect 9583 1916 9621 1925
rect 9645 1941 9730 1949
rect 9645 1921 9702 1941
rect 9722 1921 9730 1941
rect 9583 1915 9620 1916
rect 9645 1915 9730 1921
rect 9796 1945 9834 1953
rect 9796 1925 9805 1945
rect 9825 1925 9834 1945
rect 9796 1916 9834 1925
rect 9883 1919 9947 2103
rect 10103 1977 10168 2178
rect 10103 1959 10125 1977
rect 10143 1959 10168 1977
rect 10103 1940 10168 1959
rect 9796 1915 9833 1916
rect 9219 1894 9255 1915
rect 9645 1894 9676 1915
rect 9883 1910 9891 1919
rect 9880 1894 9891 1910
rect 9052 1890 9152 1894
rect 9052 1886 9114 1890
rect 9052 1860 9059 1886
rect 9085 1864 9114 1886
rect 9140 1864 9152 1890
rect 9085 1860 9152 1864
rect 9052 1857 9152 1860
rect 9220 1857 9255 1894
rect 9317 1891 9676 1894
rect 9317 1886 9539 1891
rect 9317 1862 9330 1886
rect 9354 1867 9539 1886
rect 9563 1867 9676 1891
rect 9354 1862 9676 1867
rect 9317 1858 9676 1862
rect 9743 1886 9891 1894
rect 9743 1866 9754 1886
rect 9774 1877 9891 1886
rect 9940 1910 9947 1919
rect 9940 1877 9948 1910
rect 9774 1866 9948 1877
rect 9743 1859 9948 1866
rect 9743 1858 9784 1859
rect 9219 1832 9255 1857
rect 9067 1805 9104 1806
rect 9163 1805 9200 1806
rect 9219 1805 9226 1832
rect 8743 1780 8751 1800
rect 8771 1780 8780 1800
rect 8597 1769 8628 1770
rect 8592 1701 8702 1714
rect 8743 1701 8780 1780
rect 8967 1796 9105 1805
rect 8967 1776 9076 1796
rect 9096 1776 9105 1796
rect 8967 1769 9105 1776
rect 9163 1802 9226 1805
rect 9247 1805 9255 1832
rect 9274 1805 9311 1806
rect 9247 1802 9311 1805
rect 9163 1796 9311 1802
rect 9163 1776 9172 1796
rect 9192 1776 9282 1796
rect 9302 1776 9311 1796
rect 8967 1767 9063 1769
rect 9163 1766 9311 1776
rect 9370 1796 9407 1806
rect 9482 1805 9519 1806
rect 9463 1803 9519 1805
rect 9370 1776 9378 1796
rect 9398 1776 9407 1796
rect 9219 1765 9255 1766
rect 8530 1699 8780 1701
rect 8530 1696 8631 1699
rect 8530 1677 8595 1696
rect 8592 1669 8595 1677
rect 8624 1669 8631 1696
rect 8659 1672 8669 1699
rect 8698 1677 8780 1699
rect 8698 1672 8702 1677
rect 8659 1669 8702 1672
rect 8592 1655 8702 1669
rect 8018 1637 8359 1638
rect 7943 1632 8359 1637
rect 9067 1634 9104 1635
rect 9370 1634 9407 1776
rect 9432 1796 9519 1803
rect 9432 1793 9490 1796
rect 9432 1773 9437 1793
rect 9458 1776 9490 1793
rect 9510 1776 9519 1796
rect 9458 1773 9519 1776
rect 9432 1766 9519 1773
rect 9578 1796 9615 1806
rect 9578 1776 9586 1796
rect 9606 1776 9615 1796
rect 9432 1765 9463 1766
rect 9578 1697 9615 1776
rect 9645 1805 9676 1858
rect 9880 1856 9948 1859
rect 9880 1814 9892 1856
rect 9941 1814 9948 1856
rect 9695 1805 9732 1806
rect 9645 1796 9732 1805
rect 9645 1776 9703 1796
rect 9723 1776 9732 1796
rect 9645 1766 9732 1776
rect 9791 1796 9828 1806
rect 9880 1801 9948 1814
rect 10103 1878 10168 1895
rect 10103 1860 10127 1878
rect 10145 1860 10168 1878
rect 9791 1776 9799 1796
rect 9819 1776 9828 1796
rect 9645 1765 9676 1766
rect 9640 1697 9750 1710
rect 9791 1697 9828 1776
rect 10103 1721 10168 1860
rect 10103 1715 10125 1721
rect 9578 1695 9828 1697
rect 9578 1692 9679 1695
rect 9578 1673 9643 1692
rect 9640 1665 9643 1673
rect 9672 1665 9679 1692
rect 9707 1668 9717 1695
rect 9746 1673 9828 1695
rect 9857 1703 10125 1715
rect 10143 1703 10168 1721
rect 9857 1680 10168 1703
rect 9857 1679 9912 1680
rect 9746 1668 9750 1673
rect 9707 1665 9750 1668
rect 9640 1651 9750 1665
rect 9066 1633 9407 1634
rect 7943 1612 7946 1632
rect 7966 1612 8359 1632
rect 8991 1632 9407 1633
rect 9857 1632 9900 1679
rect 8991 1628 9900 1632
rect 8310 1579 8355 1612
rect 8991 1608 8994 1628
rect 9014 1608 9900 1628
rect 9368 1603 9900 1608
rect 10108 1622 10167 1644
rect 10108 1604 10127 1622
rect 10145 1604 10167 1622
rect 9156 1579 9255 1581
rect 8310 1569 9255 1579
rect 8310 1543 9178 1569
rect 8311 1542 9178 1543
rect 9156 1531 9178 1542
rect 9203 1534 9222 1569
rect 9247 1534 9255 1569
rect 9203 1531 9255 1534
rect 10108 1533 10167 1604
rect 9156 1523 9255 1531
rect 9182 1522 9254 1523
rect 8836 1496 8903 1515
rect 8836 1475 8853 1496
rect 7717 1297 7797 1339
rect 8834 1430 8853 1475
rect 8883 1475 8903 1496
rect 8883 1430 8904 1475
rect 9373 1472 9414 1474
rect 9645 1472 9749 1474
rect 10105 1472 10169 1533
rect 6778 1186 6814 1187
rect 6670 1178 6814 1186
rect 6670 1158 6678 1178
rect 6698 1158 6786 1178
rect 6806 1158 6814 1178
rect 6670 1152 6814 1158
rect 6880 1182 6918 1190
rect 6986 1186 7022 1187
rect 6880 1162 6889 1182
rect 6909 1162 6918 1182
rect 6880 1153 6918 1162
rect 6937 1179 7022 1186
rect 6937 1159 6944 1179
rect 6965 1178 7022 1179
rect 6965 1159 6994 1178
rect 6937 1158 6994 1159
rect 7014 1158 7022 1178
rect 6880 1152 6917 1153
rect 6937 1152 7022 1158
rect 7088 1182 7126 1190
rect 7199 1186 7235 1187
rect 7088 1162 7097 1182
rect 7117 1162 7126 1182
rect 7088 1153 7126 1162
rect 7150 1178 7235 1186
rect 7150 1158 7207 1178
rect 7227 1158 7235 1178
rect 7088 1152 7125 1153
rect 7150 1152 7235 1158
rect 7301 1182 7339 1190
rect 7301 1162 7310 1182
rect 7330 1162 7339 1182
rect 7301 1153 7339 1162
rect 7539 1170 7625 1206
rect 7301 1152 7338 1153
rect 6724 1131 6760 1152
rect 7150 1131 7181 1152
rect 7377 1131 7423 1135
rect 6557 1127 6657 1131
rect 6557 1123 6619 1127
rect 6557 1097 6564 1123
rect 6590 1101 6619 1123
rect 6645 1101 6657 1127
rect 6590 1097 6657 1101
rect 6557 1094 6657 1097
rect 6725 1094 6760 1131
rect 6822 1128 7181 1131
rect 6822 1123 7044 1128
rect 6822 1099 6835 1123
rect 6859 1104 7044 1123
rect 7068 1104 7181 1128
rect 6859 1099 7181 1104
rect 6822 1095 7181 1099
rect 7248 1123 7423 1131
rect 7248 1103 7259 1123
rect 7279 1103 7423 1123
rect 7539 1129 7556 1170
rect 7610 1129 7625 1170
rect 7539 1110 7625 1129
rect 7248 1096 7423 1103
rect 7248 1095 7289 1096
rect 6724 1069 6760 1094
rect 6572 1042 6609 1043
rect 6668 1042 6705 1043
rect 6724 1042 6731 1069
rect 6472 1033 6610 1042
rect 6472 1013 6581 1033
rect 6601 1013 6610 1033
rect 6472 1006 6610 1013
rect 6668 1039 6731 1042
rect 6752 1042 6760 1069
rect 6779 1042 6816 1043
rect 6752 1039 6816 1042
rect 6668 1033 6816 1039
rect 6668 1013 6677 1033
rect 6697 1013 6787 1033
rect 6807 1013 6816 1033
rect 6472 1004 6568 1006
rect 6668 1003 6816 1013
rect 6875 1033 6912 1043
rect 6987 1042 7024 1043
rect 6968 1040 7024 1042
rect 6875 1013 6883 1033
rect 6903 1013 6912 1033
rect 6724 1002 6760 1003
rect 6572 871 6609 872
rect 6875 871 6912 1013
rect 6937 1033 7024 1040
rect 6937 1030 6995 1033
rect 6937 1010 6942 1030
rect 6963 1013 6995 1030
rect 7015 1013 7024 1033
rect 6963 1010 7024 1013
rect 6937 1003 7024 1010
rect 7083 1033 7120 1043
rect 7083 1013 7091 1033
rect 7111 1013 7120 1033
rect 6937 1002 6968 1003
rect 7083 934 7120 1013
rect 7150 1042 7181 1095
rect 7200 1042 7237 1043
rect 7150 1033 7237 1042
rect 7150 1013 7208 1033
rect 7228 1013 7237 1033
rect 7150 1003 7237 1013
rect 7296 1033 7333 1043
rect 7296 1013 7304 1033
rect 7324 1013 7333 1033
rect 7150 1002 7181 1003
rect 7145 934 7255 947
rect 7296 934 7333 1013
rect 7377 1013 7423 1096
rect 7717 1013 7792 1297
rect 8834 1222 8904 1430
rect 8966 1437 10169 1472
rect 8966 1423 8994 1437
rect 8968 1292 8994 1423
rect 9373 1434 10169 1437
rect 8826 1171 8906 1222
rect 8826 1145 8842 1171
rect 8882 1145 8906 1171
rect 8826 1126 8906 1145
rect 8826 1100 8845 1126
rect 8885 1100 8906 1126
rect 8826 1073 8906 1100
rect 8826 1047 8849 1073
rect 8889 1047 8906 1073
rect 8826 1036 8906 1047
rect 8968 1037 8995 1292
rect 9373 1284 9414 1434
rect 9645 1428 9749 1434
rect 10105 1431 10169 1434
rect 9840 1372 9961 1390
rect 9840 1370 9911 1372
rect 9840 1329 9855 1370
rect 9892 1331 9911 1370
rect 9948 1331 9961 1372
rect 9892 1329 9961 1331
rect 9840 1319 9961 1329
rect 9035 1177 9099 1189
rect 9375 1185 9412 1284
rect 9640 1274 9751 1287
rect 9640 1272 9682 1274
rect 9640 1252 9647 1272
rect 9666 1252 9682 1272
rect 9640 1244 9682 1252
rect 9710 1272 9751 1274
rect 9710 1252 9724 1272
rect 9743 1252 9751 1272
rect 9710 1244 9751 1252
rect 9640 1238 9751 1244
rect 9583 1216 9832 1238
rect 9583 1185 9620 1216
rect 9796 1214 9832 1216
rect 9796 1185 9833 1214
rect 9035 1176 9070 1177
rect 9012 1171 9070 1176
rect 9012 1151 9015 1171
rect 9035 1157 9070 1171
rect 9090 1157 9099 1177
rect 9035 1149 9099 1157
rect 9061 1148 9099 1149
rect 9062 1147 9099 1148
rect 9165 1181 9201 1182
rect 9273 1181 9309 1182
rect 9165 1173 9309 1181
rect 9165 1153 9173 1173
rect 9193 1153 9281 1173
rect 9301 1153 9309 1173
rect 9165 1147 9309 1153
rect 9375 1177 9413 1185
rect 9481 1181 9517 1182
rect 9375 1157 9384 1177
rect 9404 1157 9413 1177
rect 9375 1148 9413 1157
rect 9432 1174 9517 1181
rect 9432 1154 9439 1174
rect 9460 1173 9517 1174
rect 9460 1154 9489 1173
rect 9432 1153 9489 1154
rect 9509 1153 9517 1173
rect 9375 1147 9412 1148
rect 9432 1147 9517 1153
rect 9583 1177 9621 1185
rect 9694 1181 9730 1182
rect 9583 1157 9592 1177
rect 9612 1157 9621 1177
rect 9583 1148 9621 1157
rect 9645 1173 9730 1181
rect 9645 1153 9702 1173
rect 9722 1153 9730 1173
rect 9583 1147 9620 1148
rect 9645 1147 9730 1153
rect 9796 1177 9834 1185
rect 9796 1157 9805 1177
rect 9825 1157 9834 1177
rect 9889 1167 9954 1319
rect 10107 1293 10162 1431
rect 9796 1148 9834 1157
rect 9887 1160 9954 1167
rect 9796 1147 9833 1148
rect 9219 1126 9255 1147
rect 9645 1126 9676 1147
rect 9887 1139 9904 1160
rect 9940 1139 9954 1160
rect 10106 1180 10162 1293
rect 10106 1162 10125 1180
rect 10143 1162 10162 1180
rect 10106 1142 10162 1162
rect 9887 1126 9954 1139
rect 9052 1122 9152 1126
rect 9052 1118 9114 1122
rect 9052 1092 9059 1118
rect 9085 1096 9114 1118
rect 9140 1096 9152 1122
rect 9085 1092 9152 1096
rect 9052 1089 9152 1092
rect 9220 1089 9255 1126
rect 9317 1123 9676 1126
rect 9317 1118 9539 1123
rect 9317 1094 9330 1118
rect 9354 1099 9539 1118
rect 9563 1099 9676 1123
rect 9354 1094 9676 1099
rect 9317 1090 9676 1094
rect 9743 1120 9954 1126
rect 9743 1118 9904 1120
rect 9743 1098 9754 1118
rect 9774 1098 9904 1118
rect 9743 1091 9904 1098
rect 9743 1090 9784 1091
rect 9219 1064 9255 1089
rect 9067 1037 9104 1038
rect 9163 1037 9200 1038
rect 9219 1037 9226 1064
rect 7377 978 7792 1013
rect 8967 1028 9105 1037
rect 8967 1008 9076 1028
rect 9096 1008 9105 1028
rect 8967 1001 9105 1008
rect 9163 1034 9226 1037
rect 9247 1037 9255 1064
rect 9274 1037 9311 1038
rect 9247 1034 9311 1037
rect 9163 1028 9311 1034
rect 9163 1008 9172 1028
rect 9192 1008 9282 1028
rect 9302 1008 9311 1028
rect 8967 999 9063 1001
rect 9163 998 9311 1008
rect 9370 1028 9407 1038
rect 9482 1037 9519 1038
rect 9463 1035 9519 1037
rect 9370 1008 9378 1028
rect 9398 1008 9407 1028
rect 9219 997 9255 998
rect 7377 977 7423 978
rect 7083 932 7333 934
rect 7083 929 7184 932
rect 7083 910 7148 929
rect 7145 902 7148 910
rect 7177 902 7184 929
rect 7212 905 7222 932
rect 7251 910 7333 932
rect 7717 926 7792 978
rect 7251 905 7255 910
rect 7212 902 7255 905
rect 7145 888 7255 902
rect 6571 870 6912 871
rect 6496 865 6912 870
rect 6496 845 6499 865
rect 6519 845 6913 865
rect 2976 436 6044 461
rect 2976 371 5839 436
rect 5970 371 6044 436
rect 2976 354 6044 371
rect 6870 341 6913 845
rect 7530 756 7625 776
rect 7530 712 7550 756
rect 7610 712 7625 756
rect 7530 416 7625 712
rect 7530 375 7563 416
rect 7599 375 7625 416
rect 7725 455 7787 926
rect 9067 866 9104 867
rect 9370 866 9407 1008
rect 9432 1028 9519 1035
rect 9432 1025 9490 1028
rect 9432 1005 9437 1025
rect 9458 1008 9490 1025
rect 9510 1008 9519 1028
rect 9458 1005 9519 1008
rect 9432 998 9519 1005
rect 9578 1028 9615 1038
rect 9578 1008 9586 1028
rect 9606 1008 9615 1028
rect 9432 997 9463 998
rect 9578 929 9615 1008
rect 9645 1037 9676 1090
rect 9889 1083 9904 1091
rect 9944 1083 9954 1120
rect 9889 1074 9954 1083
rect 10102 1081 10167 1102
rect 10102 1063 10127 1081
rect 10145 1063 10167 1081
rect 9695 1037 9732 1038
rect 9645 1028 9732 1037
rect 9645 1008 9703 1028
rect 9723 1008 9732 1028
rect 9645 998 9732 1008
rect 9791 1028 9828 1038
rect 9791 1008 9799 1028
rect 9819 1008 9828 1028
rect 9645 997 9676 998
rect 9640 929 9750 942
rect 9791 929 9828 1008
rect 10102 987 10167 1063
rect 9578 927 9828 929
rect 9578 924 9679 927
rect 9578 905 9643 924
rect 9640 897 9643 905
rect 9672 897 9679 924
rect 9707 900 9717 927
rect 9746 905 9828 927
rect 9851 952 10168 987
rect 9746 900 9750 905
rect 9707 897 9750 900
rect 9640 883 9750 897
rect 9066 865 9407 866
rect 8991 863 9407 865
rect 9851 863 9891 952
rect 10102 925 10167 952
rect 10102 907 10125 925
rect 10143 907 10167 925
rect 10102 887 10167 907
rect 8988 860 9891 863
rect 8988 840 8994 860
rect 9014 840 9891 860
rect 8988 836 9891 840
rect 9851 833 9891 836
rect 10103 826 10168 847
rect 8321 818 8982 819
rect 8321 811 9255 818
rect 8321 810 9227 811
rect 8321 790 9172 810
rect 9204 791 9227 810
rect 9252 791 9255 811
rect 9204 790 9255 791
rect 8321 783 9255 790
rect 7920 741 8088 742
rect 8323 741 8362 783
rect 9151 781 9255 783
rect 9220 779 9255 781
rect 10103 808 10127 826
rect 10145 808 10168 826
rect 10103 761 10168 808
rect 7920 715 8364 741
rect 7920 713 8088 715
rect 7725 436 7789 455
rect 7725 397 7742 436
rect 7776 397 7789 436
rect 7725 378 7789 397
rect 7530 349 7625 375
rect 7920 362 7947 713
rect 8323 709 8364 715
rect 7987 502 8051 514
rect 8327 510 8364 709
rect 8826 736 8898 753
rect 8826 697 8834 736
rect 8879 697 8898 736
rect 8592 599 8703 614
rect 8592 597 8634 599
rect 8592 577 8599 597
rect 8618 577 8634 597
rect 8592 569 8634 577
rect 8662 597 8703 599
rect 8662 577 8676 597
rect 8695 577 8703 597
rect 8662 569 8703 577
rect 8592 563 8703 569
rect 8535 541 8784 563
rect 8535 510 8572 541
rect 8748 539 8784 541
rect 8748 510 8785 539
rect 7987 501 8022 502
rect 7964 496 8022 501
rect 7964 476 7967 496
rect 7987 482 8022 496
rect 8042 482 8051 502
rect 7987 474 8051 482
rect 8013 473 8051 474
rect 8014 472 8051 473
rect 8117 506 8153 507
rect 8225 506 8261 507
rect 8117 498 8261 506
rect 8117 478 8125 498
rect 8145 478 8233 498
rect 8253 478 8261 498
rect 8117 472 8261 478
rect 8327 502 8365 510
rect 8433 506 8469 507
rect 8327 482 8336 502
rect 8356 482 8365 502
rect 8327 473 8365 482
rect 8384 499 8469 506
rect 8384 479 8391 499
rect 8412 498 8469 499
rect 8412 479 8441 498
rect 8384 478 8441 479
rect 8461 478 8469 498
rect 8327 472 8364 473
rect 8384 472 8469 478
rect 8535 502 8573 510
rect 8646 506 8682 507
rect 8535 482 8544 502
rect 8564 482 8573 502
rect 8535 473 8573 482
rect 8597 498 8682 506
rect 8597 478 8654 498
rect 8674 478 8682 498
rect 8535 472 8572 473
rect 8597 472 8682 478
rect 8748 502 8786 510
rect 8748 482 8757 502
rect 8777 482 8786 502
rect 8748 473 8786 482
rect 8826 487 8898 697
rect 8968 731 10168 761
rect 8968 730 9412 731
rect 8968 728 9136 730
rect 8826 473 8909 487
rect 8748 472 8785 473
rect 8171 451 8207 472
rect 8597 451 8628 472
rect 8826 451 8843 473
rect 8004 447 8104 451
rect 8004 443 8066 447
rect 8004 417 8011 443
rect 8037 421 8066 443
rect 8092 421 8104 447
rect 8037 417 8104 421
rect 8004 414 8104 417
rect 8172 414 8207 451
rect 8269 448 8628 451
rect 8269 443 8491 448
rect 8269 419 8282 443
rect 8306 424 8491 443
rect 8515 424 8628 448
rect 8306 419 8628 424
rect 8269 415 8628 419
rect 8695 443 8843 451
rect 8695 423 8706 443
rect 8726 440 8843 443
rect 8896 440 8909 473
rect 8726 423 8909 440
rect 8695 416 8909 423
rect 8695 415 8736 416
rect 8826 415 8909 416
rect 8171 389 8207 414
rect 8019 362 8056 363
rect 8115 362 8152 363
rect 8171 362 8178 389
rect 7919 353 8057 362
rect 2731 255 2888 268
rect 2731 251 2892 255
rect 1611 105 1637 210
rect 2731 144 2772 251
rect 2872 144 2892 251
rect 2731 115 2892 144
rect 6868 132 6917 341
rect 7919 333 8028 353
rect 8048 333 8057 353
rect 7919 326 8057 333
rect 8115 359 8178 362
rect 8199 362 8207 389
rect 8226 362 8263 363
rect 8199 359 8263 362
rect 8115 353 8263 359
rect 8115 333 8124 353
rect 8144 333 8234 353
rect 8254 333 8263 353
rect 7919 324 8015 326
rect 8115 323 8263 333
rect 8322 353 8359 363
rect 8434 362 8471 363
rect 8415 360 8471 362
rect 8322 333 8330 353
rect 8350 333 8359 353
rect 8171 322 8207 323
rect 8019 191 8056 192
rect 8322 191 8359 333
rect 8384 353 8471 360
rect 8384 350 8442 353
rect 8384 330 8389 350
rect 8410 333 8442 350
rect 8462 333 8471 353
rect 8410 330 8471 333
rect 8384 323 8471 330
rect 8530 353 8567 363
rect 8530 333 8538 353
rect 8558 333 8567 353
rect 8384 322 8415 323
rect 8530 254 8567 333
rect 8597 362 8628 415
rect 8834 382 8848 415
rect 8901 382 8909 415
rect 8834 376 8909 382
rect 8834 371 8904 376
rect 8647 362 8684 363
rect 8597 353 8684 362
rect 8597 333 8655 353
rect 8675 333 8684 353
rect 8597 323 8684 333
rect 8743 353 8780 363
rect 8968 358 8995 728
rect 9035 498 9099 510
rect 9375 506 9412 730
rect 9883 711 9947 713
rect 9879 699 9947 711
rect 9879 666 9890 699
rect 9930 666 9947 699
rect 9879 656 9947 666
rect 9640 595 9751 610
rect 9640 593 9682 595
rect 9640 573 9647 593
rect 9666 573 9682 593
rect 9640 565 9682 573
rect 9710 593 9751 595
rect 9710 573 9724 593
rect 9743 573 9751 593
rect 9710 565 9751 573
rect 9640 559 9751 565
rect 9583 537 9832 559
rect 9583 506 9620 537
rect 9796 535 9832 537
rect 9796 506 9833 535
rect 9035 497 9070 498
rect 9012 492 9070 497
rect 9012 472 9015 492
rect 9035 478 9070 492
rect 9090 478 9099 498
rect 9035 470 9099 478
rect 9061 469 9099 470
rect 9062 468 9099 469
rect 9165 502 9201 503
rect 9273 502 9309 503
rect 9165 494 9309 502
rect 9165 474 9173 494
rect 9193 474 9281 494
rect 9301 474 9309 494
rect 9165 468 9309 474
rect 9375 498 9413 506
rect 9481 502 9517 503
rect 9375 478 9384 498
rect 9404 478 9413 498
rect 9375 469 9413 478
rect 9432 495 9517 502
rect 9432 475 9439 495
rect 9460 494 9517 495
rect 9460 475 9489 494
rect 9432 474 9489 475
rect 9509 474 9517 494
rect 9375 468 9412 469
rect 9432 468 9517 474
rect 9583 498 9621 506
rect 9694 502 9730 503
rect 9583 478 9592 498
rect 9612 478 9621 498
rect 9583 469 9621 478
rect 9645 494 9730 502
rect 9645 474 9702 494
rect 9722 474 9730 494
rect 9583 468 9620 469
rect 9645 468 9730 474
rect 9796 498 9834 506
rect 9796 478 9805 498
rect 9825 478 9834 498
rect 9796 469 9834 478
rect 9883 472 9947 656
rect 10103 530 10168 731
rect 10103 512 10125 530
rect 10143 512 10168 530
rect 10103 493 10168 512
rect 9796 468 9833 469
rect 9219 447 9255 468
rect 9645 447 9676 468
rect 9883 463 9891 472
rect 9880 447 9891 463
rect 9052 443 9152 447
rect 9052 439 9114 443
rect 9052 413 9059 439
rect 9085 417 9114 439
rect 9140 417 9152 443
rect 9085 413 9152 417
rect 9052 410 9152 413
rect 9220 410 9255 447
rect 9317 444 9676 447
rect 9317 439 9539 444
rect 9317 415 9330 439
rect 9354 420 9539 439
rect 9563 420 9676 444
rect 9354 415 9676 420
rect 9317 411 9676 415
rect 9743 439 9891 447
rect 9743 419 9754 439
rect 9774 430 9891 439
rect 9940 463 9947 472
rect 9940 430 9948 463
rect 9774 419 9948 430
rect 9743 412 9948 419
rect 9743 411 9784 412
rect 9219 385 9255 410
rect 9067 358 9104 359
rect 9163 358 9200 359
rect 9219 358 9226 385
rect 8743 333 8751 353
rect 8771 333 8780 353
rect 8597 322 8628 323
rect 8592 254 8702 267
rect 8743 254 8780 333
rect 8967 349 9105 358
rect 8967 329 9076 349
rect 9096 329 9105 349
rect 8967 322 9105 329
rect 9163 355 9226 358
rect 9247 358 9255 385
rect 9274 358 9311 359
rect 9247 355 9311 358
rect 9163 349 9311 355
rect 9163 329 9172 349
rect 9192 329 9282 349
rect 9302 329 9311 349
rect 8967 320 9063 322
rect 9163 319 9311 329
rect 9370 349 9407 359
rect 9482 358 9519 359
rect 9463 356 9519 358
rect 9370 329 9378 349
rect 9398 329 9407 349
rect 9219 318 9255 319
rect 8530 252 8780 254
rect 8530 249 8631 252
rect 8530 230 8595 249
rect 8592 222 8595 230
rect 8624 222 8631 249
rect 8659 225 8669 252
rect 8698 230 8780 252
rect 8698 225 8702 230
rect 8659 222 8702 225
rect 8592 208 8702 222
rect 8018 190 8359 191
rect 7943 185 8359 190
rect 9067 187 9104 188
rect 9370 187 9407 329
rect 9432 349 9519 356
rect 9432 346 9490 349
rect 9432 326 9437 346
rect 9458 329 9490 346
rect 9510 329 9519 349
rect 9458 326 9519 329
rect 9432 319 9519 326
rect 9578 349 9615 359
rect 9578 329 9586 349
rect 9606 329 9615 349
rect 9432 318 9463 319
rect 9578 250 9615 329
rect 9645 358 9676 411
rect 9880 409 9948 412
rect 9880 367 9892 409
rect 9941 367 9948 409
rect 9695 358 9732 359
rect 9645 349 9732 358
rect 9645 329 9703 349
rect 9723 329 9732 349
rect 9645 319 9732 329
rect 9791 349 9828 359
rect 9880 354 9948 367
rect 10103 431 10168 448
rect 10103 413 10127 431
rect 10145 413 10168 431
rect 9791 329 9799 349
rect 9819 329 9828 349
rect 9645 318 9676 319
rect 9640 250 9750 263
rect 9791 250 9828 329
rect 10103 274 10168 413
rect 10103 268 10125 274
rect 9578 248 9828 250
rect 9578 245 9679 248
rect 9578 226 9643 245
rect 9640 218 9643 226
rect 9672 218 9679 245
rect 9707 221 9717 248
rect 9746 226 9828 248
rect 9857 256 10125 268
rect 10143 256 10168 274
rect 9857 233 10168 256
rect 9857 232 9912 233
rect 9746 221 9750 226
rect 9707 218 9750 221
rect 9640 204 9750 218
rect 9066 186 9407 187
rect 7943 165 7946 185
rect 7966 165 8359 185
rect 8991 185 9407 186
rect 9857 185 9900 232
rect 8991 181 9900 185
rect 1611 91 1639 105
rect 2735 102 2892 115
rect 6866 130 7683 132
rect 8116 130 8205 133
rect 6866 121 8205 130
rect 413 56 1639 91
rect 6866 83 8128 121
rect 8153 86 8172 121
rect 8197 86 8205 121
rect 8310 132 8355 165
rect 8991 161 8994 181
rect 9014 161 9900 181
rect 9368 156 9900 161
rect 10108 175 10167 197
rect 10108 157 10127 175
rect 10145 157 10167 175
rect 9156 132 9255 134
rect 8310 122 9255 132
rect 8310 96 9178 122
rect 8311 95 9178 96
rect 8153 83 8205 86
rect 6866 75 8205 83
rect 9156 84 9178 95
rect 9203 87 9222 122
rect 9247 87 9255 122
rect 9203 84 9255 87
rect 9156 76 9255 84
rect 9182 75 9254 76
rect 6866 74 8204 75
rect 6866 72 7683 74
rect 7457 68 7683 72
rect 413 -20 498 56
rect 856 54 960 56
rect 1191 54 1232 56
rect 10108 -20 10167 157
rect 413 -93 10181 -20
rect 427 -108 10181 -93
rect 7496 -113 7650 -108
<< viali >>
rect 2829 12119 2866 12167
rect 1359 11828 1384 11863
rect 1403 11828 1428 11866
rect 1592 11769 1612 11789
rect 2409 11829 2434 11864
rect 2453 11829 2478 11867
rect 2640 11765 2660 11785
rect 860 11702 889 11729
rect 934 11705 963 11732
rect 665 11541 714 11583
rect 1148 11604 1169 11624
rect 1908 11698 1937 11725
rect 1982 11701 2011 11728
rect 1359 11565 1380 11595
rect 666 11478 715 11520
rect 1521 11511 1547 11537
rect 1146 11455 1167 11475
rect 1571 11458 1591 11478
rect 863 11357 882 11377
rect 940 11357 959 11377
rect 676 11251 716 11284
rect 1705 11535 1758 11568
rect 2196 11600 2217 11620
rect 2407 11561 2428 11591
rect 1710 11477 1763 11510
rect 2569 11507 2595 11533
rect 2194 11451 2215 11471
rect 2619 11454 2639 11474
rect 1911 11353 1930 11373
rect 1988 11353 2007 11373
rect 1727 11214 1772 11253
rect 2830 11514 2864 11553
rect 1354 11139 1379 11159
rect 1402 11140 1434 11160
rect 1592 11090 1612 11110
rect 860 11023 889 11050
rect 934 11026 963 11053
rect 662 10830 702 10867
rect 1148 10925 1169 10945
rect 3007 11534 3043 11575
rect 2996 11194 3056 11238
rect 5579 11641 5665 11708
rect 4087 11085 4107 11105
rect 3355 11018 3384 11045
rect 3429 11021 3458 11048
rect 1359 10886 1380 10916
rect 1521 10832 1547 10858
rect 666 10790 702 10811
rect 1146 10776 1167 10796
rect 1571 10779 1591 10799
rect 863 10678 882 10698
rect 940 10678 959 10698
rect 658 10578 695 10619
rect 714 10580 751 10621
rect 1717 10877 1757 10903
rect 1721 10824 1761 10850
rect 1724 10779 1764 10805
rect 3643 10920 3664 10940
rect 3854 10881 3875 10911
rect 2996 10780 3050 10821
rect 4016 10827 4042 10853
rect 3641 10771 3662 10791
rect 1723 10454 1753 10520
rect 1359 10381 1384 10416
rect 1403 10381 1428 10419
rect 1592 10322 1612 10342
rect 2640 10318 2660 10338
rect 860 10255 889 10282
rect 934 10258 963 10285
rect 665 10094 714 10136
rect 1148 10157 1169 10177
rect 1908 10251 1937 10278
rect 1982 10254 2011 10281
rect 1359 10118 1380 10148
rect 666 10031 715 10073
rect 1521 10064 1547 10090
rect 1146 10008 1167 10028
rect 1571 10011 1591 10031
rect 863 9910 882 9930
rect 940 9910 959 9930
rect 676 9804 716 9837
rect 1705 10088 1758 10121
rect 2196 10153 2217 10173
rect 2407 10114 2428 10144
rect 1710 10030 1763 10063
rect 2569 10060 2595 10086
rect 2194 10004 2215 10024
rect 2619 10007 2639 10027
rect 1911 9906 1930 9926
rect 1988 9906 2007 9926
rect 1727 9767 1772 9806
rect 3358 10673 3377 10693
rect 3435 10673 3454 10693
rect 4066 10774 4086 10794
rect 3865 10583 3917 10601
rect 3634 10382 3659 10417
rect 3678 10382 3703 10420
rect 3897 10398 3921 10421
rect 3897 10354 3921 10377
rect 1354 9692 1379 9712
rect 1402 9693 1434 9713
rect 1592 9643 1612 9663
rect 860 9576 889 9603
rect 934 9579 963 9606
rect 662 9383 702 9420
rect 1148 9478 1169 9498
rect 1359 9439 1380 9469
rect 1521 9385 1547 9411
rect 666 9343 702 9364
rect 1146 9329 1167 9349
rect 1571 9332 1591 9352
rect 863 9231 882 9251
rect 940 9231 959 9251
rect 658 9131 695 9172
rect 714 9133 751 9174
rect 1717 9430 1757 9456
rect 1721 9377 1761 9403
rect 1724 9332 1764 9358
rect 1716 9072 1760 9109
rect 3902 9735 3922 9756
rect 3943 9740 3963 9761
rect 4130 9640 4150 9660
rect 3398 9573 3427 9600
rect 3472 9576 3501 9603
rect 3686 9475 3707 9495
rect 3897 9436 3918 9466
rect 4059 9382 4085 9408
rect 1711 8986 1765 9052
rect 1360 8861 1385 8896
rect 1404 8861 1429 8899
rect 1593 8802 1613 8822
rect 2641 8798 2661 8818
rect 861 8735 890 8762
rect 935 8738 964 8765
rect 666 8574 715 8616
rect 1149 8637 1170 8657
rect 1909 8731 1938 8758
rect 1983 8734 2012 8761
rect 1360 8598 1381 8628
rect 667 8511 716 8553
rect 1522 8544 1548 8570
rect 1147 8488 1168 8508
rect 1572 8491 1592 8511
rect 864 8390 883 8410
rect 941 8390 960 8410
rect 677 8284 717 8317
rect 1706 8568 1759 8601
rect 2197 8633 2218 8653
rect 2408 8594 2429 8624
rect 1711 8510 1764 8543
rect 2570 8540 2596 8566
rect 2195 8484 2216 8504
rect 2620 8487 2640 8507
rect 1912 8386 1931 8406
rect 1989 8386 2008 8406
rect 1728 8247 1773 8286
rect 1355 8172 1380 8192
rect 1403 8173 1435 8193
rect 1593 8123 1613 8143
rect 861 8056 890 8083
rect 935 8059 964 8086
rect 663 7863 703 7900
rect 1149 7958 1170 7978
rect 1360 7919 1381 7949
rect 1522 7865 1548 7891
rect 667 7823 703 7844
rect 1147 7809 1168 7829
rect 1572 7812 1592 7832
rect 864 7711 883 7731
rect 941 7711 960 7731
rect 659 7611 696 7652
rect 715 7613 752 7654
rect 1718 7910 1758 7936
rect 1722 7857 1762 7883
rect 1725 7812 1765 7838
rect 2832 7853 2858 7876
rect 1724 7487 1754 7553
rect 1360 7414 1385 7449
rect 1404 7414 1429 7452
rect 1593 7355 1613 7375
rect 2641 7351 2661 7371
rect 861 7288 890 7315
rect 935 7291 964 7318
rect 666 7127 715 7169
rect 1149 7190 1170 7210
rect 1909 7284 1938 7311
rect 1983 7287 2012 7314
rect 1360 7151 1381 7181
rect 667 7064 716 7106
rect 1522 7097 1548 7123
rect 1147 7041 1168 7061
rect 1572 7044 1592 7064
rect 864 6943 883 6963
rect 941 6943 960 6963
rect 677 6837 717 6870
rect 1706 7121 1759 7154
rect 2197 7186 2218 7206
rect 2408 7147 2429 7177
rect 1711 7063 1764 7096
rect 2570 7093 2596 7119
rect 2195 7037 2216 7057
rect 2620 7040 2640 7060
rect 1912 6939 1931 6959
rect 1989 6939 2008 6959
rect 1728 6800 1773 6839
rect 1355 6725 1380 6745
rect 1403 6726 1435 6746
rect 1593 6676 1613 6696
rect 861 6609 890 6636
rect 935 6612 964 6639
rect 663 6416 703 6453
rect 1149 6511 1170 6531
rect 1360 6472 1381 6502
rect 1522 6418 1548 6444
rect 667 6376 703 6397
rect 1147 6362 1168 6382
rect 1572 6365 1592 6385
rect 864 6264 883 6284
rect 941 6264 960 6284
rect 659 6164 696 6205
rect 715 6166 752 6207
rect 1718 6463 1758 6489
rect 1722 6410 1762 6436
rect 1725 6365 1765 6391
rect 1716 6044 1762 6092
rect 3684 9326 3705 9346
rect 4109 9329 4129 9349
rect 3401 9228 3420 9248
rect 3478 9228 3497 9248
rect 3701 8862 3726 8900
rect 3859 8171 3876 8208
rect 4088 8118 4108 8138
rect 3356 8051 3385 8078
rect 3430 8054 3459 8081
rect 3644 7953 3665 7973
rect 3855 7914 3876 7944
rect 3212 7846 3238 7869
rect 4017 7860 4043 7886
rect 3642 7804 3663 7824
rect 4067 7807 4087 7827
rect 3359 7706 3378 7726
rect 3436 7706 3455 7726
rect 3699 7434 3727 7462
rect 5196 6667 5216 6687
rect 4464 6600 4493 6627
rect 4538 6603 4567 6630
rect 4752 6502 4773 6522
rect 4963 6463 4984 6493
rect 4260 6404 4284 6428
rect 4317 6405 4341 6429
rect 5125 6409 5151 6435
rect 4750 6353 4771 6373
rect 4963 6351 4987 6373
rect 5175 6356 5195 6376
rect 4467 6255 4486 6275
rect 4544 6255 4563 6275
rect 8843 11567 8883 11593
rect 8846 11522 8886 11548
rect 8850 11469 8890 11495
rect 9856 11751 9893 11792
rect 9912 11753 9949 11794
rect 9648 11674 9667 11694
rect 9725 11674 9744 11694
rect 9016 11573 9036 11593
rect 9440 11576 9461 11596
rect 9905 11561 9941 11582
rect 9060 11514 9086 11540
rect 9227 11456 9248 11486
rect 9438 11427 9459 11447
rect 9905 11505 9945 11542
rect 9644 11319 9673 11346
rect 9718 11322 9747 11349
rect 8995 11262 9015 11282
rect 9173 11212 9205 11232
rect 9228 11213 9253 11233
rect 8835 11119 8880 11158
rect 8600 10999 8619 11019
rect 8677 10999 8696 11019
rect 7968 10898 7988 10918
rect 8392 10901 8413 10921
rect 8012 10839 8038 10865
rect 8844 10862 8897 10895
rect 8179 10781 8200 10811
rect 8390 10752 8411 10772
rect 8849 10804 8902 10837
rect 9891 11088 9931 11121
rect 9648 10995 9667 11015
rect 9725 10995 9744 11015
rect 9016 10894 9036 10914
rect 9440 10897 9461 10917
rect 9060 10835 9086 10861
rect 9892 10852 9941 10894
rect 9227 10777 9248 10807
rect 8596 10644 8625 10671
rect 8670 10647 8699 10674
rect 9438 10748 9459 10768
rect 9893 10789 9942 10831
rect 9644 10640 9673 10667
rect 9718 10643 9747 10670
rect 7947 10587 7967 10607
rect 8995 10583 9015 10603
rect 6881 10496 6909 10524
rect 9179 10506 9204 10544
rect 9223 10509 9248 10544
rect 8854 10405 8884 10471
rect 7153 10232 7172 10252
rect 7230 10232 7249 10252
rect 6521 10131 6541 10151
rect 6945 10134 6966 10154
rect 6565 10072 6591 10098
rect 7370 10089 7396 10112
rect 7750 10082 7776 10105
rect 6732 10014 6753 10044
rect 6943 9985 6964 10005
rect 8843 10120 8883 10146
rect 8846 10075 8886 10101
rect 8850 10022 8890 10048
rect 7149 9877 7178 9904
rect 7223 9880 7252 9907
rect 6500 9820 6520 9840
rect 6732 9750 6749 9787
rect 9856 10304 9893 10345
rect 9912 10306 9949 10347
rect 9648 10227 9667 10247
rect 9725 10227 9744 10247
rect 9016 10126 9036 10146
rect 9440 10129 9461 10149
rect 9905 10114 9941 10135
rect 9060 10067 9086 10093
rect 9227 10009 9248 10039
rect 9438 9980 9459 10000
rect 9905 10058 9945 10095
rect 9644 9872 9673 9899
rect 9718 9875 9747 9902
rect 8995 9815 9015 9835
rect 9173 9765 9205 9785
rect 9228 9766 9253 9786
rect 6882 9058 6907 9096
rect 8835 9672 8880 9711
rect 8600 9552 8619 9572
rect 8677 9552 8696 9572
rect 7968 9451 7988 9471
rect 8392 9454 8413 9474
rect 8012 9392 8038 9418
rect 8844 9415 8897 9448
rect 8179 9334 8200 9364
rect 8390 9305 8411 9325
rect 8849 9357 8902 9390
rect 9891 9641 9931 9674
rect 9648 9548 9667 9568
rect 9725 9548 9744 9568
rect 9016 9447 9036 9467
rect 9440 9450 9461 9470
rect 9060 9388 9086 9414
rect 9892 9405 9941 9447
rect 9227 9330 9248 9360
rect 8596 9197 8625 9224
rect 8670 9200 8699 9227
rect 9438 9301 9459 9321
rect 9893 9342 9942 9384
rect 9644 9193 9673 9220
rect 9718 9196 9747 9223
rect 7947 9140 7967 9160
rect 8995 9136 9015 9156
rect 9179 9059 9204 9097
rect 9223 9062 9248 9097
rect 8843 8906 8897 8972
rect 7111 8710 7130 8730
rect 7188 8710 7207 8730
rect 6479 8609 6499 8629
rect 6903 8612 6924 8632
rect 6523 8550 6549 8576
rect 6690 8492 6711 8522
rect 6901 8463 6922 8483
rect 7107 8355 7136 8382
rect 7181 8358 7210 8385
rect 6458 8298 6478 8318
rect 8848 8849 8892 8886
rect 8844 8600 8884 8626
rect 8847 8555 8887 8581
rect 8851 8502 8891 8528
rect 9857 8784 9894 8825
rect 9913 8786 9950 8827
rect 9649 8707 9668 8727
rect 9726 8707 9745 8727
rect 9017 8606 9037 8626
rect 9441 8609 9462 8629
rect 9906 8594 9942 8615
rect 9061 8547 9087 8573
rect 9228 8489 9249 8519
rect 9439 8460 9460 8480
rect 9906 8538 9946 8575
rect 9645 8352 9674 8379
rect 9719 8355 9748 8382
rect 8996 8295 9016 8315
rect 9174 8245 9206 8265
rect 9229 8246 9254 8266
rect 6687 7581 6711 7604
rect 6687 7537 6711 7560
rect 6905 7538 6930 7576
rect 6949 7541 6974 7576
rect 6691 7357 6743 7375
rect 6522 7164 6542 7184
rect 7154 7265 7173 7285
rect 7231 7265 7250 7285
rect 8836 8152 8881 8191
rect 8601 8032 8620 8052
rect 8678 8032 8697 8052
rect 7969 7931 7989 7951
rect 8393 7934 8414 7954
rect 8013 7872 8039 7898
rect 8845 7895 8898 7928
rect 8180 7814 8201 7844
rect 8391 7785 8412 7805
rect 8850 7837 8903 7870
rect 9892 8121 9932 8154
rect 9649 8028 9668 8048
rect 9726 8028 9745 8048
rect 9017 7927 9037 7947
rect 9441 7930 9462 7950
rect 9061 7868 9087 7894
rect 9893 7885 9942 7927
rect 9228 7810 9249 7840
rect 8597 7677 8626 7704
rect 8671 7680 8700 7707
rect 9439 7781 9460 7801
rect 9894 7822 9943 7864
rect 9645 7673 9674 7700
rect 9719 7676 9748 7703
rect 7948 7620 7968 7640
rect 8996 7616 9016 7636
rect 9180 7539 9205 7577
rect 9224 7542 9249 7577
rect 8855 7438 8885 7504
rect 6946 7167 6967 7187
rect 6566 7105 6592 7131
rect 7558 7137 7612 7178
rect 6733 7047 6754 7077
rect 6944 7018 6965 7038
rect 8844 7153 8884 7179
rect 8847 7108 8887 7134
rect 8851 7055 8891 7081
rect 9857 7337 9894 7378
rect 9913 7339 9950 7380
rect 9649 7260 9668 7280
rect 9726 7260 9745 7280
rect 9017 7159 9037 7179
rect 9441 7162 9462 7182
rect 9906 7147 9942 7168
rect 9061 7100 9087 7126
rect 9228 7042 9249 7072
rect 7150 6910 7179 6937
rect 7224 6913 7253 6940
rect 6501 6853 6521 6873
rect 4803 6162 4832 6196
rect 4802 6102 4831 6136
rect 3018 6017 3062 6045
rect 2827 5918 2864 5966
rect 3015 5960 3059 5988
rect 5310 5878 5373 5932
rect 1357 5820 1382 5855
rect 1401 5820 1426 5858
rect 1590 5761 1610 5781
rect 2407 5821 2432 5856
rect 2451 5821 2476 5859
rect 2638 5757 2658 5777
rect 858 5694 887 5721
rect 932 5697 961 5724
rect 663 5533 712 5575
rect 1146 5596 1167 5616
rect 1906 5690 1935 5717
rect 1980 5693 2009 5720
rect 1357 5557 1378 5587
rect 664 5470 713 5512
rect 1519 5503 1545 5529
rect 1144 5447 1165 5467
rect 1569 5450 1589 5470
rect 861 5349 880 5369
rect 938 5349 957 5369
rect 674 5243 714 5276
rect 1703 5527 1756 5560
rect 2194 5592 2215 5612
rect 2405 5553 2426 5583
rect 1708 5469 1761 5502
rect 2567 5499 2593 5525
rect 2192 5443 2213 5463
rect 2617 5446 2637 5466
rect 1909 5345 1928 5365
rect 1986 5345 2005 5365
rect 1725 5206 1770 5245
rect 2828 5506 2862 5545
rect 1352 5131 1377 5151
rect 1400 5132 1432 5152
rect 1590 5082 1610 5102
rect 858 5015 887 5042
rect 932 5018 961 5045
rect 660 4822 700 4859
rect 1146 4917 1167 4937
rect 3005 5526 3041 5567
rect 2994 5186 3054 5230
rect 4085 5077 4105 5097
rect 3353 5010 3382 5037
rect 3427 5013 3456 5040
rect 1357 4878 1378 4908
rect 1519 4824 1545 4850
rect 664 4782 700 4803
rect 1144 4768 1165 4788
rect 1569 4771 1589 4791
rect 861 4670 880 4690
rect 938 4670 957 4690
rect 656 4570 693 4611
rect 712 4572 749 4613
rect 1715 4869 1755 4895
rect 1719 4816 1759 4842
rect 1722 4771 1762 4797
rect 3641 4912 3662 4932
rect 3852 4873 3873 4903
rect 2994 4772 3048 4813
rect 4014 4819 4040 4845
rect 3639 4763 3660 4783
rect 1721 4446 1751 4512
rect 1357 4373 1382 4408
rect 1401 4373 1426 4411
rect 1590 4314 1610 4334
rect 2638 4310 2658 4330
rect 858 4247 887 4274
rect 932 4250 961 4277
rect 663 4086 712 4128
rect 1146 4149 1167 4169
rect 1906 4243 1935 4270
rect 1980 4246 2009 4273
rect 1357 4110 1378 4140
rect 664 4023 713 4065
rect 1519 4056 1545 4082
rect 1144 4000 1165 4020
rect 1569 4003 1589 4023
rect 861 3902 880 3922
rect 938 3902 957 3922
rect 674 3796 714 3829
rect 1703 4080 1756 4113
rect 2194 4145 2215 4165
rect 2405 4106 2426 4136
rect 1708 4022 1761 4055
rect 2567 4052 2593 4078
rect 2192 3996 2213 4016
rect 2617 3999 2637 4019
rect 1909 3898 1928 3918
rect 1986 3898 2005 3918
rect 1725 3759 1770 3798
rect 3356 4665 3375 4685
rect 3433 4665 3452 4685
rect 4064 4766 4084 4786
rect 3863 4575 3915 4593
rect 3632 4374 3657 4409
rect 3676 4374 3701 4412
rect 3895 4390 3919 4413
rect 3895 4346 3919 4369
rect 1352 3684 1377 3704
rect 1400 3685 1432 3705
rect 1590 3635 1610 3655
rect 858 3568 887 3595
rect 932 3571 961 3598
rect 660 3375 700 3412
rect 1146 3470 1167 3490
rect 1357 3431 1378 3461
rect 1519 3377 1545 3403
rect 664 3335 700 3356
rect 1144 3321 1165 3341
rect 1569 3324 1589 3344
rect 861 3223 880 3243
rect 938 3223 957 3243
rect 656 3123 693 3164
rect 712 3125 749 3166
rect 1715 3422 1755 3448
rect 1719 3369 1759 3395
rect 1722 3324 1762 3350
rect 1714 3064 1758 3101
rect 4128 3632 4148 3652
rect 3396 3565 3425 3592
rect 3470 3568 3499 3595
rect 3684 3467 3705 3487
rect 3895 3428 3916 3458
rect 4057 3374 4083 3400
rect 1709 2978 1763 3044
rect 1358 2853 1383 2888
rect 1402 2853 1427 2891
rect 1591 2794 1611 2814
rect 2639 2790 2659 2810
rect 859 2727 888 2754
rect 933 2730 962 2757
rect 664 2566 713 2608
rect 1147 2629 1168 2649
rect 1907 2723 1936 2750
rect 1981 2726 2010 2753
rect 1358 2590 1379 2620
rect 665 2503 714 2545
rect 1520 2536 1546 2562
rect 1145 2480 1166 2500
rect 1570 2483 1590 2503
rect 862 2382 881 2402
rect 939 2382 958 2402
rect 675 2276 715 2309
rect 1704 2560 1757 2593
rect 2195 2625 2216 2645
rect 2406 2586 2427 2616
rect 1709 2502 1762 2535
rect 2568 2532 2594 2558
rect 2193 2476 2214 2496
rect 2618 2479 2638 2499
rect 1910 2378 1929 2398
rect 1987 2378 2006 2398
rect 1726 2239 1771 2278
rect 1353 2164 1378 2184
rect 1401 2165 1433 2185
rect 1591 2115 1611 2135
rect 859 2048 888 2075
rect 933 2051 962 2078
rect 661 1855 701 1892
rect 1147 1950 1168 1970
rect 1358 1911 1379 1941
rect 1520 1857 1546 1883
rect 665 1815 701 1836
rect 1145 1801 1166 1821
rect 1570 1804 1590 1824
rect 862 1703 881 1723
rect 939 1703 958 1723
rect 657 1603 694 1644
rect 713 1605 750 1646
rect 1716 1902 1756 1928
rect 1720 1849 1760 1875
rect 1723 1804 1763 1830
rect 2785 1835 2810 1866
rect 2830 1845 2856 1868
rect 1722 1479 1752 1545
rect 1358 1406 1383 1441
rect 1402 1406 1427 1444
rect 1591 1347 1611 1367
rect 2639 1343 2659 1363
rect 859 1280 888 1307
rect 933 1283 962 1310
rect 664 1119 713 1161
rect 1147 1182 1168 1202
rect 1907 1276 1936 1303
rect 1981 1279 2010 1306
rect 1358 1143 1379 1173
rect 665 1056 714 1098
rect 1520 1089 1546 1115
rect 1145 1033 1166 1053
rect 1570 1036 1590 1056
rect 862 935 881 955
rect 939 935 958 955
rect 675 829 715 862
rect 1704 1113 1757 1146
rect 2195 1178 2216 1198
rect 2406 1139 2427 1169
rect 1709 1055 1762 1088
rect 2568 1085 2594 1111
rect 2193 1029 2214 1049
rect 2618 1032 2638 1052
rect 1910 931 1929 951
rect 1987 931 2006 951
rect 1726 792 1771 831
rect 1353 717 1378 737
rect 1401 718 1433 738
rect 1591 668 1611 688
rect 859 601 888 628
rect 933 604 962 631
rect 661 408 701 445
rect 1147 503 1168 523
rect 1358 464 1379 494
rect 1520 410 1546 436
rect 665 368 701 389
rect 1145 354 1166 374
rect 1570 357 1590 377
rect 862 256 881 276
rect 939 256 958 276
rect 657 156 694 197
rect 713 158 750 199
rect 3682 3318 3703 3338
rect 4107 3321 4127 3341
rect 3399 3220 3418 3240
rect 3476 3220 3495 3240
rect 3699 2854 3724 2892
rect 5775 5814 5804 5848
rect 5774 5754 5803 5788
rect 6043 5675 6062 5695
rect 6120 5675 6139 5695
rect 5411 5574 5431 5594
rect 5835 5577 5856 5597
rect 7552 6720 7612 6764
rect 7565 6383 7601 6424
rect 9439 7013 9460 7033
rect 9906 7091 9946 7128
rect 9645 6905 9674 6932
rect 9719 6908 9748 6935
rect 8996 6848 9016 6868
rect 9174 6798 9206 6818
rect 9229 6799 9254 6819
rect 7744 6405 7778 6444
rect 8836 6705 8881 6744
rect 8601 6585 8620 6605
rect 8678 6585 8697 6605
rect 7969 6484 7989 6504
rect 8393 6487 8414 6507
rect 8013 6425 8039 6451
rect 8845 6448 8898 6481
rect 8180 6367 8201 6397
rect 8391 6338 8412 6358
rect 8850 6390 8903 6423
rect 9892 6674 9932 6707
rect 9649 6581 9668 6601
rect 9726 6581 9745 6601
rect 9017 6480 9037 6500
rect 9441 6483 9462 6503
rect 9061 6421 9087 6447
rect 9893 6438 9942 6480
rect 9228 6363 9249 6393
rect 8597 6230 8626 6257
rect 8671 6233 8700 6260
rect 9439 6334 9460 6354
rect 9894 6375 9943 6417
rect 9645 6226 9674 6253
rect 9719 6229 9748 6256
rect 7948 6173 7968 6193
rect 8130 6091 8155 6129
rect 8174 6094 8199 6129
rect 8996 6169 9016 6189
rect 9180 6092 9205 6130
rect 9224 6095 9249 6130
rect 5455 5515 5481 5541
rect 6265 5521 6289 5545
rect 6322 5522 6346 5546
rect 5622 5457 5643 5487
rect 5833 5428 5854 5448
rect 7547 5962 7591 5990
rect 7742 5984 7779 6032
rect 7544 5905 7588 5933
rect 6039 5320 6068 5347
rect 6113 5323 6142 5350
rect 5390 5263 5410 5283
rect 5152 2865 5177 2891
rect 5541 2796 5561 2816
rect 4809 2729 4838 2756
rect 4883 2732 4912 2759
rect 5097 2631 5118 2651
rect 5308 2592 5329 2622
rect 5470 2538 5496 2564
rect 5095 2482 5116 2502
rect 5299 2484 5332 2504
rect 5520 2485 5540 2505
rect 4812 2384 4831 2404
rect 4889 2384 4908 2404
rect 5620 2327 5643 2365
rect 6879 4488 6907 4516
rect 7151 4224 7170 4244
rect 7228 4224 7247 4244
rect 6519 4123 6539 4143
rect 6943 4126 6964 4146
rect 6563 4064 6589 4090
rect 7368 4081 7394 4104
rect 6730 4006 6751 4036
rect 6941 3977 6962 3997
rect 7147 3869 7176 3896
rect 7221 3872 7250 3899
rect 6498 3812 6518 3832
rect 6730 3742 6747 3779
rect 6880 3050 6905 3088
rect 7109 2702 7128 2722
rect 7186 2702 7205 2722
rect 6477 2601 6497 2621
rect 6901 2604 6922 2624
rect 8844 5858 8890 5906
rect 8841 5559 8881 5585
rect 8844 5514 8884 5540
rect 8848 5461 8888 5487
rect 9854 5743 9891 5784
rect 9910 5745 9947 5786
rect 9646 5666 9665 5686
rect 9723 5666 9742 5686
rect 9014 5565 9034 5585
rect 9438 5568 9459 5588
rect 9903 5553 9939 5574
rect 9058 5506 9084 5532
rect 9225 5448 9246 5478
rect 9436 5419 9457 5439
rect 9903 5497 9943 5534
rect 9642 5311 9671 5338
rect 9716 5314 9745 5341
rect 8993 5254 9013 5274
rect 9171 5204 9203 5224
rect 9226 5205 9251 5225
rect 8833 5111 8878 5150
rect 8598 4991 8617 5011
rect 8675 4991 8694 5011
rect 7966 4890 7986 4910
rect 8390 4893 8411 4913
rect 8010 4831 8036 4857
rect 8842 4854 8895 4887
rect 8177 4773 8198 4803
rect 8388 4744 8409 4764
rect 8847 4796 8900 4829
rect 9889 5080 9929 5113
rect 9646 4987 9665 5007
rect 9723 4987 9742 5007
rect 9014 4886 9034 4906
rect 9438 4889 9459 4909
rect 9058 4827 9084 4853
rect 9890 4844 9939 4886
rect 9225 4769 9246 4799
rect 8594 4636 8623 4663
rect 8668 4639 8697 4666
rect 9436 4740 9457 4760
rect 9891 4781 9940 4823
rect 9642 4632 9671 4659
rect 9716 4635 9745 4662
rect 7945 4579 7965 4599
rect 8993 4575 9013 4595
rect 9177 4498 9202 4536
rect 9221 4501 9246 4536
rect 8852 4397 8882 4463
rect 7748 4074 7774 4097
rect 8841 4112 8881 4138
rect 8844 4067 8884 4093
rect 8848 4014 8888 4040
rect 9854 4296 9891 4337
rect 9910 4298 9947 4339
rect 9646 4219 9665 4239
rect 9723 4219 9742 4239
rect 9014 4118 9034 4138
rect 9438 4121 9459 4141
rect 9903 4106 9939 4127
rect 9058 4059 9084 4085
rect 9225 4001 9246 4031
rect 9436 3972 9457 3992
rect 9903 4050 9943 4087
rect 9642 3864 9671 3891
rect 9716 3867 9745 3894
rect 8993 3807 9013 3827
rect 9171 3757 9203 3777
rect 9226 3758 9251 3778
rect 8833 3664 8878 3703
rect 8598 3544 8617 3564
rect 8675 3544 8694 3564
rect 7966 3443 7986 3463
rect 8390 3446 8411 3466
rect 8010 3384 8036 3410
rect 8842 3407 8895 3440
rect 8177 3326 8198 3356
rect 8388 3297 8409 3317
rect 8847 3349 8900 3382
rect 9889 3633 9929 3666
rect 9646 3540 9665 3560
rect 9723 3540 9742 3560
rect 9014 3439 9034 3459
rect 9438 3442 9459 3462
rect 9058 3380 9084 3406
rect 9890 3397 9939 3439
rect 9225 3322 9246 3352
rect 8594 3189 8623 3216
rect 8668 3192 8697 3219
rect 9436 3293 9457 3313
rect 9891 3334 9940 3376
rect 9642 3185 9671 3212
rect 9716 3188 9745 3215
rect 7945 3132 7965 3152
rect 8993 3128 9013 3148
rect 9177 3051 9202 3089
rect 9221 3054 9246 3089
rect 8841 2898 8895 2964
rect 6521 2542 6547 2568
rect 6688 2484 6709 2514
rect 6899 2455 6920 2475
rect 7105 2347 7134 2374
rect 7179 2350 7208 2377
rect 6456 2290 6476 2310
rect 3857 2163 3874 2200
rect 6643 2189 6663 2210
rect 6684 2194 6704 2215
rect 4086 2110 4106 2130
rect 3354 2043 3383 2070
rect 3428 2046 3457 2073
rect 3642 1945 3663 1965
rect 3853 1906 3874 1936
rect 3210 1838 3236 1861
rect 4015 1852 4041 1878
rect 3640 1796 3661 1816
rect 4065 1799 4085 1819
rect 3357 1698 3376 1718
rect 3434 1698 3453 1718
rect 8846 2841 8890 2878
rect 8842 2592 8882 2618
rect 8845 2547 8885 2573
rect 8849 2494 8889 2520
rect 9855 2776 9892 2817
rect 9911 2778 9948 2819
rect 9647 2699 9666 2719
rect 9724 2699 9743 2719
rect 9015 2598 9035 2618
rect 9439 2601 9460 2621
rect 9904 2586 9940 2607
rect 9059 2539 9085 2565
rect 9226 2481 9247 2511
rect 9437 2452 9458 2472
rect 9904 2530 9944 2567
rect 9643 2344 9672 2371
rect 9717 2347 9746 2374
rect 8994 2287 9014 2307
rect 9172 2237 9204 2257
rect 9227 2238 9252 2258
rect 6685 1573 6709 1596
rect 6685 1529 6709 1552
rect 6903 1530 6928 1568
rect 6947 1533 6972 1568
rect 3697 1426 3725 1454
rect 6689 1349 6741 1367
rect 6520 1156 6540 1176
rect 7152 1257 7171 1277
rect 7229 1257 7248 1277
rect 8834 2144 8879 2183
rect 8599 2024 8618 2044
rect 8676 2024 8695 2044
rect 7967 1923 7987 1943
rect 8391 1926 8412 1946
rect 8011 1864 8037 1890
rect 8843 1887 8896 1920
rect 8178 1806 8199 1836
rect 8389 1777 8410 1797
rect 8848 1829 8901 1862
rect 9890 2113 9930 2146
rect 9647 2020 9666 2040
rect 9724 2020 9743 2040
rect 9015 1919 9035 1939
rect 9439 1922 9460 1942
rect 9059 1860 9085 1886
rect 9891 1877 9940 1919
rect 9226 1802 9247 1832
rect 8595 1669 8624 1696
rect 8669 1672 8698 1699
rect 9437 1773 9458 1793
rect 9892 1814 9941 1856
rect 9643 1665 9672 1692
rect 9717 1668 9746 1695
rect 7946 1612 7966 1632
rect 8994 1608 9014 1628
rect 9178 1531 9203 1569
rect 9222 1534 9247 1569
rect 8853 1430 8883 1496
rect 6944 1159 6965 1179
rect 6564 1097 6590 1123
rect 7556 1129 7610 1170
rect 6731 1039 6752 1069
rect 6942 1010 6963 1030
rect 8842 1145 8882 1171
rect 8845 1100 8885 1126
rect 8849 1047 8889 1073
rect 9855 1329 9892 1370
rect 9911 1331 9948 1372
rect 9647 1252 9666 1272
rect 9724 1252 9743 1272
rect 9015 1151 9035 1171
rect 9439 1154 9460 1174
rect 9904 1139 9940 1160
rect 9059 1092 9085 1118
rect 9226 1034 9247 1064
rect 7148 902 7177 929
rect 7222 905 7251 932
rect 6499 845 6519 865
rect 5839 371 5970 436
rect 7550 712 7610 756
rect 7563 375 7599 416
rect 9437 1005 9458 1025
rect 9904 1083 9944 1120
rect 9643 897 9672 924
rect 9717 900 9746 927
rect 8994 840 9014 860
rect 9172 790 9204 810
rect 9227 791 9252 811
rect 7742 397 7776 436
rect 8834 697 8879 736
rect 8599 577 8618 597
rect 8676 577 8695 597
rect 7967 476 7987 496
rect 8391 479 8412 499
rect 8011 417 8037 443
rect 8843 440 8896 473
rect 2772 144 2872 251
rect 8178 359 8199 389
rect 8389 330 8410 350
rect 8848 382 8901 415
rect 9890 666 9930 699
rect 9647 573 9666 593
rect 9724 573 9743 593
rect 9015 472 9035 492
rect 9439 475 9460 495
rect 9059 413 9085 439
rect 9891 430 9940 472
rect 9226 355 9247 385
rect 8595 222 8624 249
rect 8669 225 8698 252
rect 9437 326 9458 346
rect 9892 367 9941 409
rect 9643 218 9672 245
rect 9717 221 9746 248
rect 7946 165 7966 185
rect 8128 83 8153 121
rect 8172 86 8197 121
rect 8994 161 9014 181
rect 9178 84 9203 122
rect 9222 87 9247 122
<< metal1 >>
rect 177 11395 284 12185
rect 656 11583 728 12176
rect 1352 11874 1424 11875
rect 1351 11866 1450 11874
rect 1351 11863 1403 11866
rect 1351 11828 1359 11863
rect 1384 11828 1403 11863
rect 1428 11828 1450 11866
rect 1351 11816 1450 11828
rect 1352 11797 1420 11816
rect 1353 11794 1386 11797
rect 1588 11794 1620 11795
rect 763 11733 966 11746
rect 763 11700 787 11733
rect 823 11732 966 11733
rect 823 11729 934 11732
rect 823 11702 860 11729
rect 889 11705 934 11729
rect 963 11705 966 11732
rect 889 11702 966 11705
rect 823 11700 966 11702
rect 763 11687 966 11700
rect 763 11686 864 11687
rect 656 11541 665 11583
rect 714 11541 728 11583
rect 656 11520 728 11541
rect 656 11478 666 11520
rect 715 11478 728 11520
rect 656 11460 728 11478
rect 1141 11624 1173 11631
rect 1141 11604 1148 11624
rect 1169 11604 1173 11624
rect 1141 11539 1173 11604
rect 1353 11595 1384 11794
rect 1585 11789 1620 11794
rect 1585 11769 1592 11789
rect 1612 11769 1620 11789
rect 1585 11761 1620 11769
rect 1353 11565 1359 11595
rect 1380 11565 1384 11595
rect 1353 11557 1384 11565
rect 1511 11539 1551 11540
rect 1141 11537 1553 11539
rect 1141 11511 1521 11537
rect 1547 11511 1553 11537
rect 1141 11503 1553 11511
rect 1141 11475 1173 11503
rect 1586 11483 1620 11761
rect 1702 11574 1772 12177
rect 2816 12167 2881 12202
rect 2816 12163 2829 12167
rect 2817 12119 2829 12163
rect 2866 12163 2881 12167
rect 2866 12119 2879 12163
rect 2402 11875 2474 11876
rect 2401 11867 2490 11875
rect 2401 11864 2453 11867
rect 2401 11829 2409 11864
rect 2434 11829 2453 11864
rect 2478 11829 2490 11867
rect 2401 11817 2490 11829
rect 2401 11816 2470 11817
rect 2401 11798 2437 11816
rect 1811 11729 2014 11742
rect 1811 11696 1835 11729
rect 1871 11728 2014 11729
rect 1871 11725 1982 11728
rect 1871 11698 1908 11725
rect 1937 11701 1982 11725
rect 2011 11701 2014 11728
rect 1937 11698 2014 11701
rect 1871 11696 2014 11698
rect 1811 11683 2014 11696
rect 1811 11682 1912 11683
rect 1141 11455 1146 11475
rect 1167 11455 1173 11475
rect 1141 11448 1173 11455
rect 1564 11478 1620 11483
rect 1564 11458 1571 11478
rect 1591 11458 1620 11478
rect 1697 11568 1772 11574
rect 1697 11535 1705 11568
rect 1758 11535 1772 11568
rect 1697 11510 1772 11535
rect 1697 11477 1710 11510
rect 1763 11477 1772 11510
rect 1697 11468 1772 11477
rect 2189 11620 2221 11627
rect 2189 11600 2196 11620
rect 2217 11600 2221 11620
rect 2189 11535 2221 11600
rect 2401 11591 2432 11798
rect 2636 11790 2668 11791
rect 2633 11785 2668 11790
rect 2633 11765 2640 11785
rect 2660 11765 2668 11785
rect 2633 11757 2668 11765
rect 2401 11561 2407 11591
rect 2428 11561 2432 11591
rect 2401 11553 2432 11561
rect 2559 11535 2599 11536
rect 2189 11533 2601 11535
rect 2189 11507 2569 11533
rect 2595 11507 2601 11533
rect 2189 11499 2601 11507
rect 2189 11471 2221 11499
rect 2634 11479 2668 11757
rect 2817 11572 2879 12119
rect 2986 11575 3068 12197
rect 4253 11724 4302 12237
rect 9891 11812 9956 11950
rect 9841 11794 9962 11812
rect 9841 11792 9912 11794
rect 9841 11751 9856 11792
rect 9893 11753 9912 11792
rect 9949 11753 9962 11794
rect 9893 11751 9962 11753
rect 9841 11741 9962 11751
rect 5547 11736 5685 11740
rect 5185 11724 5685 11736
rect 4243 11708 5685 11724
rect 4243 11641 5579 11708
rect 5665 11641 5685 11708
rect 6357 11712 7835 11714
rect 10323 11712 10430 11912
rect 6357 11694 10432 11712
rect 6357 11674 9648 11694
rect 9667 11674 9725 11694
rect 9744 11674 10432 11694
rect 6357 11656 10432 11674
rect 7790 11655 7997 11656
rect 9641 11652 9752 11656
rect 4243 11625 5685 11641
rect 2817 11553 2881 11572
rect 2817 11514 2830 11553
rect 2864 11514 2881 11553
rect 2817 11495 2881 11514
rect 2986 11534 3007 11575
rect 3043 11534 3068 11575
rect 2986 11505 3068 11534
rect 1697 11463 1755 11468
rect 1564 11451 1620 11458
rect 2189 11451 2194 11471
rect 2215 11451 2221 11471
rect 1564 11450 1599 11451
rect 2189 11444 2221 11451
rect 2612 11474 2668 11479
rect 2612 11454 2619 11474
rect 2639 11454 2668 11474
rect 2612 11447 2668 11454
rect 2612 11446 2647 11447
rect 855 11395 966 11399
rect 2638 11395 3751 11396
rect 177 11377 3751 11395
rect 177 11357 863 11377
rect 882 11357 940 11377
rect 959 11373 3751 11377
rect 959 11357 1911 11373
rect 177 11353 1911 11357
rect 1930 11353 1988 11373
rect 2007 11353 3751 11373
rect 177 11339 3751 11353
rect 177 10716 284 11339
rect 1903 11336 2014 11339
rect 663 11290 727 11294
rect 659 11284 727 11290
rect 659 11251 676 11284
rect 716 11251 727 11284
rect 659 11239 727 11251
rect 1710 11253 1775 11275
rect 659 11237 716 11239
rect 663 10876 714 11237
rect 1710 11214 1727 11253
rect 1772 11214 1775 11253
rect 1351 11169 1386 11171
rect 1351 11160 1455 11169
rect 1351 11159 1402 11160
rect 1351 11139 1354 11159
rect 1379 11140 1402 11159
rect 1434 11140 1455 11160
rect 1379 11139 1455 11140
rect 1351 11132 1455 11139
rect 1351 11120 1386 11132
rect 763 11054 966 11067
rect 763 11021 787 11054
rect 823 11053 966 11054
rect 823 11050 934 11053
rect 823 11023 860 11050
rect 889 11026 934 11050
rect 963 11026 966 11053
rect 889 11023 966 11026
rect 823 11021 966 11023
rect 763 11008 966 11021
rect 763 11007 864 11008
rect 1141 10945 1173 10952
rect 1141 10925 1148 10945
rect 1169 10925 1173 10945
rect 652 10867 717 10876
rect 652 10830 662 10867
rect 702 10833 717 10867
rect 1141 10860 1173 10925
rect 1353 10916 1384 11120
rect 1588 11115 1620 11116
rect 1585 11110 1620 11115
rect 1585 11090 1592 11110
rect 1612 11090 1620 11110
rect 1585 11082 1620 11090
rect 1353 10886 1359 10916
rect 1380 10886 1384 10916
rect 1353 10878 1384 10886
rect 1511 10860 1551 10861
rect 1141 10858 1553 10860
rect 702 10830 719 10833
rect 652 10811 719 10830
rect 652 10790 666 10811
rect 702 10790 719 10811
rect 652 10783 719 10790
rect 1141 10832 1521 10858
rect 1547 10832 1553 10858
rect 1141 10824 1553 10832
rect 1141 10796 1173 10824
rect 1586 10804 1620 11082
rect 1710 10914 1775 11214
rect 2981 11238 3074 11253
rect 2981 11194 2996 11238
rect 3056 11194 3074 11238
rect 1141 10776 1146 10796
rect 1167 10776 1173 10796
rect 1141 10769 1173 10776
rect 1564 10799 1620 10804
rect 1564 10779 1571 10799
rect 1591 10779 1620 10799
rect 1564 10772 1620 10779
rect 1700 10903 1780 10914
rect 1700 10877 1717 10903
rect 1757 10877 1780 10903
rect 1700 10850 1780 10877
rect 1700 10824 1721 10850
rect 1761 10824 1780 10850
rect 1700 10805 1780 10824
rect 1700 10779 1724 10805
rect 1764 10779 1780 10805
rect 1564 10771 1599 10772
rect 1700 10767 1780 10779
rect 2981 10821 3074 11194
rect 3258 11049 3461 11062
rect 3258 11016 3282 11049
rect 3318 11048 3461 11049
rect 3318 11045 3429 11048
rect 3318 11018 3355 11045
rect 3384 11021 3429 11045
rect 3458 11021 3461 11048
rect 3384 11018 3461 11021
rect 3318 11016 3461 11018
rect 3258 11003 3461 11016
rect 3258 11002 3359 11003
rect 2981 10780 2996 10821
rect 3050 10780 3074 10821
rect 2981 10773 3074 10780
rect 3636 10940 3668 10947
rect 3636 10920 3643 10940
rect 3664 10920 3668 10940
rect 3636 10855 3668 10920
rect 3848 10911 3879 11112
rect 4083 11110 4115 11111
rect 4080 11105 4115 11110
rect 4080 11085 4087 11105
rect 4107 11085 4115 11105
rect 4080 11077 4115 11085
rect 3848 10881 3854 10911
rect 3875 10881 3879 10911
rect 3848 10873 3879 10881
rect 4006 10855 4046 10856
rect 3636 10853 4048 10855
rect 3636 10827 4016 10853
rect 4042 10827 4048 10853
rect 3636 10819 4048 10827
rect 3636 10791 3668 10819
rect 4081 10799 4115 11077
rect 3636 10771 3641 10791
rect 3662 10771 3668 10791
rect 3636 10764 3668 10771
rect 4059 10794 4115 10799
rect 4059 10774 4066 10794
rect 4086 10774 4115 10794
rect 4059 10767 4115 10774
rect 4059 10766 4094 10767
rect 855 10716 966 10720
rect 2597 10716 4146 10719
rect 175 10698 4146 10716
rect 175 10678 863 10698
rect 882 10678 940 10698
rect 959 10693 4146 10698
rect 959 10678 3358 10693
rect 175 10673 3358 10678
rect 3377 10673 3435 10693
rect 3454 10673 4146 10693
rect 175 10663 4146 10673
rect 175 10660 800 10663
rect 987 10660 4146 10663
rect 177 10432 284 10660
rect 2597 10659 4146 10660
rect 3350 10656 3461 10659
rect 645 10621 766 10631
rect 645 10619 714 10621
rect 645 10578 658 10619
rect 695 10580 714 10619
rect 751 10580 766 10621
rect 695 10578 766 10580
rect 645 10560 766 10578
rect 3850 10601 3936 10605
rect 3850 10583 3865 10601
rect 3917 10583 3936 10601
rect 3850 10574 3936 10583
rect 651 10458 730 10560
rect 1703 10520 1770 10539
rect 1703 10500 1723 10520
rect 177 10377 285 10432
rect 652 10377 730 10458
rect 1702 10454 1723 10500
rect 1753 10500 1770 10520
rect 1753 10470 1772 10500
rect 1753 10454 1773 10470
rect 1702 10438 1773 10454
rect 1352 10427 1424 10428
rect 1351 10419 1450 10427
rect 1351 10416 1403 10419
rect 1351 10381 1359 10416
rect 1384 10381 1403 10416
rect 1428 10381 1450 10419
rect 177 9948 284 10377
rect 656 10136 728 10377
rect 1351 10369 1450 10381
rect 1352 10350 1420 10369
rect 1353 10347 1386 10350
rect 1588 10347 1620 10348
rect 763 10286 966 10299
rect 763 10253 787 10286
rect 823 10285 966 10286
rect 823 10282 934 10285
rect 823 10255 860 10282
rect 889 10258 934 10282
rect 963 10258 966 10285
rect 889 10255 966 10258
rect 823 10253 966 10255
rect 763 10240 966 10253
rect 763 10239 864 10240
rect 656 10094 665 10136
rect 714 10094 728 10136
rect 656 10073 728 10094
rect 656 10031 666 10073
rect 715 10031 728 10073
rect 656 10013 728 10031
rect 1141 10177 1173 10184
rect 1141 10157 1148 10177
rect 1169 10157 1173 10177
rect 1141 10092 1173 10157
rect 1353 10148 1384 10347
rect 1585 10342 1620 10347
rect 1585 10322 1592 10342
rect 1612 10322 1620 10342
rect 1585 10314 1620 10322
rect 1353 10118 1359 10148
rect 1380 10118 1384 10148
rect 1353 10110 1384 10118
rect 1511 10092 1551 10093
rect 1141 10090 1553 10092
rect 1141 10064 1521 10090
rect 1547 10064 1553 10090
rect 1141 10056 1553 10064
rect 1141 10028 1173 10056
rect 1586 10036 1620 10314
rect 1702 10127 1772 10438
rect 3627 10428 3699 10429
rect 3626 10425 3715 10428
rect 2398 10423 3715 10425
rect 2395 10420 3715 10423
rect 2395 10417 3678 10420
rect 2395 10382 3634 10417
rect 3659 10382 3678 10417
rect 3703 10382 3715 10420
rect 2395 10372 3715 10382
rect 3891 10421 3927 10574
rect 3891 10398 3897 10421
rect 3921 10398 3927 10421
rect 3891 10377 3927 10398
rect 2395 10370 3680 10372
rect 2395 10360 2492 10370
rect 2401 10351 2437 10360
rect 3891 10354 3897 10377
rect 3921 10354 3927 10377
rect 1811 10282 2014 10295
rect 1811 10249 1835 10282
rect 1871 10281 2014 10282
rect 1871 10278 1982 10281
rect 1871 10251 1908 10278
rect 1937 10254 1982 10278
rect 2011 10254 2014 10281
rect 1937 10251 2014 10254
rect 1871 10249 2014 10251
rect 1811 10236 2014 10249
rect 1811 10235 1912 10236
rect 1141 10008 1146 10028
rect 1167 10008 1173 10028
rect 1141 10001 1173 10008
rect 1564 10031 1620 10036
rect 1564 10011 1571 10031
rect 1591 10011 1620 10031
rect 1697 10121 1772 10127
rect 1697 10088 1705 10121
rect 1758 10088 1772 10121
rect 1697 10063 1772 10088
rect 1697 10030 1710 10063
rect 1763 10030 1772 10063
rect 1697 10021 1772 10030
rect 2189 10173 2221 10180
rect 2189 10153 2196 10173
rect 2217 10153 2221 10173
rect 2189 10088 2221 10153
rect 2401 10144 2432 10351
rect 2636 10343 2668 10344
rect 3891 10343 3927 10354
rect 2633 10338 2668 10343
rect 2633 10318 2640 10338
rect 2660 10318 2668 10338
rect 2633 10310 2668 10318
rect 2401 10114 2407 10144
rect 2428 10114 2432 10144
rect 2401 10106 2432 10114
rect 2559 10088 2599 10089
rect 2189 10086 2601 10088
rect 2189 10060 2569 10086
rect 2595 10060 2601 10086
rect 2189 10052 2601 10060
rect 2189 10024 2221 10052
rect 2634 10032 2668 10310
rect 1697 10016 1755 10021
rect 1564 10004 1620 10011
rect 2189 10004 2194 10024
rect 2215 10004 2221 10024
rect 1564 10003 1599 10004
rect 2189 9997 2221 10004
rect 2612 10027 2668 10032
rect 2612 10007 2619 10027
rect 2639 10007 2668 10027
rect 2612 10000 2668 10007
rect 2612 9999 2647 10000
rect 855 9948 966 9952
rect 2730 9948 3971 9949
rect 177 9930 3971 9948
rect 177 9910 863 9930
rect 882 9910 940 9930
rect 959 9926 3971 9930
rect 959 9910 1911 9926
rect 177 9906 1911 9910
rect 1930 9906 1988 9926
rect 2007 9906 3971 9926
rect 177 9892 3971 9906
rect 177 9269 284 9892
rect 1903 9889 2014 9892
rect 663 9843 727 9847
rect 659 9837 727 9843
rect 659 9804 676 9837
rect 716 9804 727 9837
rect 659 9792 727 9804
rect 1710 9806 1775 9828
rect 659 9790 716 9792
rect 663 9429 714 9790
rect 1710 9767 1727 9806
rect 1772 9767 1775 9806
rect 1351 9722 1386 9724
rect 1351 9713 1455 9722
rect 1351 9712 1402 9713
rect 1351 9692 1354 9712
rect 1379 9693 1402 9712
rect 1434 9693 1455 9713
rect 1379 9692 1455 9693
rect 1351 9685 1455 9692
rect 1351 9673 1386 9685
rect 763 9607 966 9620
rect 763 9574 787 9607
rect 823 9606 966 9607
rect 823 9603 934 9606
rect 823 9576 860 9603
rect 889 9579 934 9603
rect 963 9579 966 9606
rect 889 9576 966 9579
rect 823 9574 966 9576
rect 763 9561 966 9574
rect 763 9560 864 9561
rect 1141 9498 1173 9505
rect 1141 9478 1148 9498
rect 1169 9478 1173 9498
rect 652 9420 717 9429
rect 652 9383 662 9420
rect 702 9386 717 9420
rect 1141 9413 1173 9478
rect 1353 9469 1384 9673
rect 1588 9668 1620 9669
rect 1585 9663 1620 9668
rect 1585 9643 1592 9663
rect 1612 9643 1620 9663
rect 1585 9635 1620 9643
rect 1353 9439 1359 9469
rect 1380 9439 1384 9469
rect 1353 9431 1384 9439
rect 1511 9413 1551 9414
rect 1141 9411 1553 9413
rect 702 9383 719 9386
rect 652 9364 719 9383
rect 652 9343 666 9364
rect 702 9343 719 9364
rect 652 9336 719 9343
rect 1141 9385 1521 9411
rect 1547 9385 1553 9411
rect 1141 9377 1553 9385
rect 1141 9349 1173 9377
rect 1586 9357 1620 9635
rect 1710 9467 1775 9767
rect 3889 9761 3994 9770
rect 3889 9756 3943 9761
rect 3889 9735 3902 9756
rect 3922 9740 3943 9756
rect 3963 9740 3994 9761
rect 3922 9735 3994 9740
rect 3889 9704 3994 9735
rect 3892 9687 3927 9704
rect 3891 9669 3927 9687
rect 3301 9604 3504 9617
rect 3301 9571 3325 9604
rect 3361 9603 3504 9604
rect 3361 9600 3472 9603
rect 3361 9573 3398 9600
rect 3427 9576 3472 9600
rect 3501 9576 3504 9603
rect 3427 9573 3504 9576
rect 3361 9571 3504 9573
rect 3301 9558 3504 9571
rect 3301 9557 3402 9558
rect 3679 9495 3711 9502
rect 3679 9475 3686 9495
rect 3707 9475 3711 9495
rect 1141 9329 1146 9349
rect 1167 9329 1173 9349
rect 1141 9322 1173 9329
rect 1564 9352 1620 9357
rect 1564 9332 1571 9352
rect 1591 9332 1620 9352
rect 1564 9325 1620 9332
rect 1700 9456 1780 9467
rect 1700 9430 1717 9456
rect 1757 9430 1780 9456
rect 1700 9403 1780 9430
rect 1700 9377 1721 9403
rect 1761 9377 1780 9403
rect 1700 9358 1780 9377
rect 1700 9332 1724 9358
rect 1764 9332 1780 9358
rect 1564 9324 1599 9325
rect 1700 9320 1780 9332
rect 3679 9410 3711 9475
rect 3891 9466 3922 9669
rect 4126 9665 4158 9666
rect 4123 9660 4158 9665
rect 4123 9640 4130 9660
rect 4150 9640 4158 9660
rect 4123 9632 4158 9640
rect 3891 9436 3897 9466
rect 3918 9436 3922 9466
rect 3891 9428 3922 9436
rect 4049 9410 4089 9411
rect 3679 9408 4091 9410
rect 3679 9382 4059 9408
rect 4085 9382 4091 9408
rect 3679 9374 4091 9382
rect 3679 9346 3711 9374
rect 4124 9354 4158 9632
rect 3679 9326 3684 9346
rect 3705 9326 3711 9346
rect 3679 9319 3711 9326
rect 4102 9349 4158 9354
rect 4102 9329 4109 9349
rect 4129 9329 4158 9349
rect 4102 9322 4158 9329
rect 4102 9321 4137 9322
rect 855 9269 966 9273
rect 2610 9269 2817 9270
rect 3393 9269 3504 9270
rect 175 9251 4195 9269
rect 175 9231 863 9251
rect 882 9231 940 9251
rect 959 9248 4195 9251
rect 959 9231 3401 9248
rect 175 9228 3401 9231
rect 3420 9228 3478 9248
rect 3497 9228 4195 9248
rect 175 9213 4195 9228
rect 177 9025 284 9213
rect 2772 9211 4195 9213
rect 645 9174 766 9184
rect 645 9172 714 9174
rect 645 9131 658 9172
rect 695 9133 714 9172
rect 751 9133 766 9174
rect 695 9131 766 9133
rect 645 9113 766 9131
rect 177 9021 285 9025
rect 651 9021 728 9113
rect 1701 9109 1777 9125
rect 1701 9086 1716 9109
rect 178 8428 285 9021
rect 653 8970 728 9021
rect 1694 9072 1716 9086
rect 1760 9072 1777 9109
rect 1694 9052 1777 9072
rect 1694 8986 1711 9052
rect 1765 8986 1777 9052
rect 653 8927 729 8970
rect 657 8616 729 8927
rect 1694 8962 1777 8986
rect 1694 8942 1770 8962
rect 1694 8923 1773 8942
rect 1353 8907 1425 8908
rect 1352 8899 1451 8907
rect 1352 8896 1404 8899
rect 1352 8861 1360 8896
rect 1385 8861 1404 8896
rect 1429 8861 1451 8899
rect 1352 8849 1451 8861
rect 1353 8830 1421 8849
rect 1354 8827 1387 8830
rect 1589 8827 1621 8828
rect 764 8766 967 8779
rect 764 8733 788 8766
rect 824 8765 967 8766
rect 824 8762 935 8765
rect 824 8735 861 8762
rect 890 8738 935 8762
rect 964 8738 967 8765
rect 890 8735 967 8738
rect 824 8733 967 8735
rect 764 8720 967 8733
rect 764 8719 865 8720
rect 657 8574 666 8616
rect 715 8574 729 8616
rect 657 8553 729 8574
rect 657 8511 667 8553
rect 716 8511 729 8553
rect 657 8493 729 8511
rect 1142 8657 1174 8664
rect 1142 8637 1149 8657
rect 1170 8637 1174 8657
rect 1142 8572 1174 8637
rect 1354 8628 1385 8827
rect 1586 8822 1621 8827
rect 1586 8802 1593 8822
rect 1613 8802 1621 8822
rect 1586 8794 1621 8802
rect 1354 8598 1360 8628
rect 1381 8598 1385 8628
rect 1354 8590 1385 8598
rect 1512 8572 1552 8573
rect 1142 8570 1554 8572
rect 1142 8544 1522 8570
rect 1548 8544 1554 8570
rect 1142 8536 1554 8544
rect 1142 8508 1174 8536
rect 1587 8516 1621 8794
rect 1703 8607 1773 8923
rect 3691 8908 3722 8909
rect 3691 8900 3736 8908
rect 2771 8877 2935 8884
rect 3691 8877 3701 8900
rect 2397 8862 3701 8877
rect 3726 8862 3736 8900
rect 2397 8844 3736 8862
rect 2402 8831 2438 8844
rect 2771 8841 2935 8844
rect 1812 8762 2015 8775
rect 1812 8729 1836 8762
rect 1872 8761 2015 8762
rect 1872 8758 1983 8761
rect 1872 8731 1909 8758
rect 1938 8734 1983 8758
rect 2012 8734 2015 8761
rect 1938 8731 2015 8734
rect 1872 8729 2015 8731
rect 1812 8716 2015 8729
rect 1812 8715 1913 8716
rect 1142 8488 1147 8508
rect 1168 8488 1174 8508
rect 1142 8481 1174 8488
rect 1565 8511 1621 8516
rect 1565 8491 1572 8511
rect 1592 8491 1621 8511
rect 1698 8601 1773 8607
rect 1698 8568 1706 8601
rect 1759 8568 1773 8601
rect 1698 8543 1773 8568
rect 1698 8510 1711 8543
rect 1764 8510 1773 8543
rect 1698 8501 1773 8510
rect 2190 8653 2222 8660
rect 2190 8633 2197 8653
rect 2218 8633 2222 8653
rect 2190 8568 2222 8633
rect 2402 8624 2433 8831
rect 2637 8823 2669 8824
rect 2634 8818 2669 8823
rect 2634 8798 2641 8818
rect 2661 8798 2669 8818
rect 2634 8790 2669 8798
rect 2402 8594 2408 8624
rect 2429 8594 2433 8624
rect 2402 8586 2433 8594
rect 2560 8568 2600 8569
rect 2190 8566 2602 8568
rect 2190 8540 2570 8566
rect 2596 8540 2602 8566
rect 2190 8532 2602 8540
rect 2190 8504 2222 8532
rect 2635 8512 2669 8790
rect 1698 8496 1756 8501
rect 1565 8484 1621 8491
rect 2190 8484 2195 8504
rect 2216 8484 2222 8504
rect 1565 8483 1600 8484
rect 2190 8477 2222 8484
rect 2613 8507 2669 8512
rect 2613 8487 2620 8507
rect 2640 8487 2669 8507
rect 2613 8480 2669 8487
rect 2613 8479 2648 8480
rect 856 8428 967 8432
rect 2639 8428 3939 8429
rect 178 8410 3939 8428
rect 178 8390 864 8410
rect 883 8390 941 8410
rect 960 8406 3939 8410
rect 960 8390 1912 8406
rect 178 8386 1912 8390
rect 1931 8386 1989 8406
rect 2008 8386 3939 8406
rect 178 8372 3939 8386
rect 178 7749 285 8372
rect 1904 8369 2015 8372
rect 664 8323 728 8327
rect 660 8317 728 8323
rect 660 8284 677 8317
rect 717 8284 728 8317
rect 660 8272 728 8284
rect 1711 8286 1776 8308
rect 660 8270 717 8272
rect 664 7909 715 8270
rect 1711 8247 1728 8286
rect 1773 8247 1776 8286
rect 1352 8202 1387 8204
rect 1352 8193 1456 8202
rect 1352 8192 1403 8193
rect 1352 8172 1355 8192
rect 1380 8173 1403 8192
rect 1435 8173 1456 8193
rect 1380 8172 1456 8173
rect 1352 8165 1456 8172
rect 1352 8153 1387 8165
rect 764 8087 967 8100
rect 764 8054 788 8087
rect 824 8086 967 8087
rect 824 8083 935 8086
rect 824 8056 861 8083
rect 890 8059 935 8083
rect 964 8059 967 8086
rect 890 8056 967 8059
rect 824 8054 967 8056
rect 764 8041 967 8054
rect 764 8040 865 8041
rect 1142 7978 1174 7985
rect 1142 7958 1149 7978
rect 1170 7958 1174 7978
rect 653 7900 718 7909
rect 653 7863 663 7900
rect 703 7866 718 7900
rect 1142 7893 1174 7958
rect 1354 7949 1385 8153
rect 1589 8148 1621 8149
rect 1586 8143 1621 8148
rect 1586 8123 1593 8143
rect 1613 8123 1621 8143
rect 1586 8115 1621 8123
rect 1354 7919 1360 7949
rect 1381 7919 1385 7949
rect 1354 7911 1385 7919
rect 1512 7893 1552 7894
rect 1142 7891 1554 7893
rect 703 7863 720 7866
rect 653 7844 720 7863
rect 653 7823 667 7844
rect 703 7823 720 7844
rect 653 7816 720 7823
rect 1142 7865 1522 7891
rect 1548 7865 1554 7891
rect 1142 7857 1554 7865
rect 1142 7829 1174 7857
rect 1587 7837 1621 8115
rect 1711 7947 1776 8247
rect 3848 8208 3885 8229
rect 3848 8171 3859 8208
rect 3876 8184 3885 8208
rect 3876 8171 3886 8184
rect 3848 8161 3886 8171
rect 3849 8157 3886 8161
rect 3849 8151 3882 8157
rect 3259 8082 3462 8095
rect 3259 8049 3283 8082
rect 3319 8081 3462 8082
rect 3319 8078 3430 8081
rect 3319 8051 3356 8078
rect 3385 8054 3430 8078
rect 3459 8054 3462 8081
rect 3385 8051 3462 8054
rect 3319 8049 3462 8051
rect 3259 8036 3462 8049
rect 3259 8035 3360 8036
rect 3637 7973 3669 7980
rect 3637 7953 3644 7973
rect 3665 7953 3669 7973
rect 1142 7809 1147 7829
rect 1168 7809 1174 7829
rect 1142 7802 1174 7809
rect 1565 7832 1621 7837
rect 1565 7812 1572 7832
rect 1592 7812 1621 7832
rect 1565 7805 1621 7812
rect 1701 7936 1781 7947
rect 1701 7910 1718 7936
rect 1758 7910 1781 7936
rect 1701 7883 1781 7910
rect 1701 7857 1722 7883
rect 1762 7857 1781 7883
rect 3637 7888 3669 7953
rect 3849 7944 3880 8151
rect 4084 8143 4116 8144
rect 4081 8138 4116 8143
rect 4081 8118 4088 8138
rect 4108 8118 4116 8138
rect 4081 8110 4116 8118
rect 3849 7914 3855 7944
rect 3876 7914 3880 7944
rect 3849 7906 3880 7914
rect 4007 7888 4047 7889
rect 3637 7886 4049 7888
rect 1701 7838 1781 7857
rect 1701 7812 1725 7838
rect 1765 7812 1781 7838
rect 2814 7876 3251 7882
rect 2814 7853 2832 7876
rect 2858 7869 3251 7876
rect 2858 7853 3212 7869
rect 2814 7846 3212 7853
rect 3238 7846 3251 7869
rect 2814 7833 3251 7846
rect 3637 7860 4017 7886
rect 4043 7860 4049 7886
rect 3637 7852 4049 7860
rect 1565 7804 1600 7805
rect 1701 7800 1781 7812
rect 3637 7824 3669 7852
rect 4082 7832 4116 8110
rect 3637 7804 3642 7824
rect 3663 7804 3669 7824
rect 3637 7797 3669 7804
rect 4060 7827 4116 7832
rect 4060 7807 4067 7827
rect 4087 7807 4116 7827
rect 4060 7800 4116 7807
rect 4060 7799 4095 7800
rect 856 7749 967 7753
rect 2598 7749 4148 7752
rect 176 7731 4148 7749
rect 176 7711 864 7731
rect 883 7711 941 7731
rect 960 7726 4148 7731
rect 960 7711 3359 7726
rect 176 7706 3359 7711
rect 3378 7706 3436 7726
rect 3455 7706 4148 7726
rect 176 7696 4148 7706
rect 176 7693 801 7696
rect 988 7693 4148 7696
rect 178 7465 285 7693
rect 2598 7692 4148 7693
rect 3351 7689 3462 7692
rect 646 7654 767 7664
rect 646 7652 715 7654
rect 646 7611 659 7652
rect 696 7613 715 7652
rect 752 7613 767 7654
rect 696 7611 767 7613
rect 646 7593 767 7611
rect 652 7491 731 7593
rect 1704 7553 1771 7572
rect 1704 7533 1724 7553
rect 178 7410 286 7465
rect 653 7410 731 7491
rect 1703 7487 1724 7533
rect 1754 7533 1771 7553
rect 1754 7503 1773 7533
rect 1754 7487 1774 7503
rect 1703 7471 1774 7487
rect 1353 7460 1425 7461
rect 1352 7452 1451 7460
rect 1352 7449 1404 7452
rect 1352 7414 1360 7449
rect 1385 7414 1404 7449
rect 1429 7414 1451 7452
rect 178 6981 285 7410
rect 657 7169 729 7410
rect 1352 7402 1451 7414
rect 1353 7383 1421 7402
rect 1354 7380 1387 7383
rect 1589 7380 1621 7381
rect 764 7319 967 7332
rect 764 7286 788 7319
rect 824 7318 967 7319
rect 824 7315 935 7318
rect 824 7288 861 7315
rect 890 7291 935 7315
rect 964 7291 967 7318
rect 890 7288 967 7291
rect 824 7286 967 7288
rect 764 7273 967 7286
rect 764 7272 865 7273
rect 657 7127 666 7169
rect 715 7127 729 7169
rect 657 7106 729 7127
rect 657 7064 667 7106
rect 716 7064 729 7106
rect 657 7046 729 7064
rect 1142 7210 1174 7217
rect 1142 7190 1149 7210
rect 1170 7190 1174 7210
rect 1142 7125 1174 7190
rect 1354 7181 1385 7380
rect 1586 7375 1621 7380
rect 1586 7355 1593 7375
rect 1613 7355 1621 7375
rect 1586 7347 1621 7355
rect 1354 7151 1360 7181
rect 1381 7151 1385 7181
rect 1354 7143 1385 7151
rect 1512 7125 1552 7126
rect 1142 7123 1554 7125
rect 1142 7097 1522 7123
rect 1548 7097 1554 7123
rect 1142 7089 1554 7097
rect 1142 7061 1174 7089
rect 1587 7069 1621 7347
rect 1703 7160 1773 7471
rect 2400 7462 3742 7467
rect 2400 7460 3699 7462
rect 2397 7434 3699 7460
rect 3727 7434 3742 7462
rect 2397 7426 3742 7434
rect 2397 7401 2436 7426
rect 2397 7384 2438 7401
rect 2397 7377 2436 7384
rect 1812 7315 2015 7328
rect 1812 7282 1836 7315
rect 1872 7314 2015 7315
rect 1872 7311 1983 7314
rect 1872 7284 1909 7311
rect 1938 7287 1983 7311
rect 2012 7287 2015 7314
rect 1938 7284 2015 7287
rect 1872 7282 2015 7284
rect 1812 7269 2015 7282
rect 1812 7268 1913 7269
rect 1142 7041 1147 7061
rect 1168 7041 1174 7061
rect 1142 7034 1174 7041
rect 1565 7064 1621 7069
rect 1565 7044 1572 7064
rect 1592 7044 1621 7064
rect 1698 7154 1773 7160
rect 1698 7121 1706 7154
rect 1759 7121 1773 7154
rect 1698 7096 1773 7121
rect 1698 7063 1711 7096
rect 1764 7063 1773 7096
rect 1698 7054 1773 7063
rect 2190 7206 2222 7213
rect 2190 7186 2197 7206
rect 2218 7186 2222 7206
rect 2190 7121 2222 7186
rect 2402 7177 2433 7377
rect 2637 7376 2669 7377
rect 2634 7371 2669 7376
rect 2634 7351 2641 7371
rect 2661 7351 2669 7371
rect 2634 7343 2669 7351
rect 2402 7147 2408 7177
rect 2429 7147 2433 7177
rect 2402 7139 2433 7147
rect 2560 7121 2600 7122
rect 2190 7119 2602 7121
rect 2190 7093 2570 7119
rect 2596 7093 2602 7119
rect 2190 7085 2602 7093
rect 2190 7057 2222 7085
rect 2635 7065 2669 7343
rect 1698 7049 1756 7054
rect 1565 7037 1621 7044
rect 2190 7037 2195 7057
rect 2216 7037 2222 7057
rect 1565 7036 1600 7037
rect 2190 7030 2222 7037
rect 2613 7060 2669 7065
rect 2613 7040 2620 7060
rect 2640 7040 2669 7060
rect 2613 7033 2669 7040
rect 2613 7032 2648 7033
rect 856 6981 967 6985
rect 2731 6981 3721 6982
rect 178 6963 3721 6981
rect 178 6943 864 6963
rect 883 6943 941 6963
rect 960 6959 3721 6963
rect 960 6943 1912 6959
rect 178 6939 1912 6943
rect 1931 6939 1989 6959
rect 2008 6939 3721 6959
rect 178 6925 3721 6939
rect 178 6302 285 6925
rect 1904 6922 2015 6925
rect 664 6876 728 6880
rect 660 6870 728 6876
rect 660 6837 677 6870
rect 717 6837 728 6870
rect 660 6825 728 6837
rect 1711 6839 1776 6861
rect 660 6823 717 6825
rect 664 6462 715 6823
rect 1711 6800 1728 6839
rect 1773 6800 1776 6839
rect 1352 6755 1387 6757
rect 1352 6746 1456 6755
rect 1352 6745 1403 6746
rect 1352 6725 1355 6745
rect 1380 6726 1403 6745
rect 1435 6726 1456 6746
rect 1380 6725 1456 6726
rect 1352 6718 1456 6725
rect 1352 6706 1387 6718
rect 764 6640 967 6653
rect 764 6607 788 6640
rect 824 6639 967 6640
rect 824 6636 935 6639
rect 824 6609 861 6636
rect 890 6612 935 6636
rect 964 6612 967 6639
rect 890 6609 967 6612
rect 824 6607 967 6609
rect 764 6594 967 6607
rect 764 6593 865 6594
rect 1142 6531 1174 6538
rect 1142 6511 1149 6531
rect 1170 6511 1174 6531
rect 653 6453 718 6462
rect 653 6416 663 6453
rect 703 6419 718 6453
rect 1142 6446 1174 6511
rect 1354 6502 1385 6706
rect 1589 6701 1621 6702
rect 1586 6696 1621 6701
rect 1586 6676 1593 6696
rect 1613 6676 1621 6696
rect 1586 6668 1621 6676
rect 1354 6472 1360 6502
rect 1381 6472 1385 6502
rect 1354 6464 1385 6472
rect 1512 6446 1552 6447
rect 1142 6444 1554 6446
rect 703 6416 720 6419
rect 653 6397 720 6416
rect 653 6376 667 6397
rect 703 6376 720 6397
rect 653 6369 720 6376
rect 1142 6418 1522 6444
rect 1548 6418 1554 6444
rect 1142 6410 1554 6418
rect 1142 6382 1174 6410
rect 1587 6390 1621 6668
rect 1711 6500 1776 6800
rect 1142 6362 1147 6382
rect 1168 6362 1174 6382
rect 1142 6355 1174 6362
rect 1565 6385 1621 6390
rect 1565 6365 1572 6385
rect 1592 6365 1621 6385
rect 1565 6358 1621 6365
rect 1701 6489 1781 6500
rect 1701 6463 1718 6489
rect 1758 6463 1781 6489
rect 1701 6436 1781 6463
rect 4253 6439 4302 11625
rect 5185 11622 5685 11625
rect 5547 11614 5685 11622
rect 8827 11593 8907 11605
rect 9008 11600 9043 11601
rect 8827 11567 8843 11593
rect 8883 11567 8907 11593
rect 8827 11548 8907 11567
rect 8827 11522 8846 11548
rect 8886 11522 8907 11548
rect 8827 11495 8907 11522
rect 8827 11469 8850 11495
rect 8890 11469 8907 11495
rect 8827 11458 8907 11469
rect 8987 11593 9043 11600
rect 8987 11573 9016 11593
rect 9036 11573 9043 11593
rect 8987 11568 9043 11573
rect 9434 11596 9466 11603
rect 9434 11576 9440 11596
rect 9461 11576 9466 11596
rect 5293 11351 5398 11376
rect 5293 11142 5310 11351
rect 5381 11142 5398 11351
rect 4367 6631 4570 6644
rect 4367 6598 4391 6631
rect 4427 6630 4570 6631
rect 4427 6627 4538 6630
rect 4427 6600 4464 6627
rect 4493 6603 4538 6627
rect 4567 6603 4570 6630
rect 4493 6600 4570 6603
rect 4427 6598 4570 6600
rect 4367 6585 4570 6598
rect 4367 6584 4468 6585
rect 4745 6522 4777 6529
rect 4745 6502 4752 6522
rect 4773 6502 4777 6522
rect 1701 6410 1722 6436
rect 1762 6410 1781 6436
rect 1701 6391 1781 6410
rect 4252 6429 4363 6439
rect 4252 6428 4317 6429
rect 4252 6404 4260 6428
rect 4284 6405 4317 6428
rect 4341 6405 4363 6429
rect 4284 6404 4363 6405
rect 4252 6397 4363 6404
rect 4745 6437 4777 6502
rect 4957 6493 4988 6693
rect 5192 6692 5224 6693
rect 5189 6687 5224 6692
rect 5189 6667 5196 6687
rect 5216 6667 5224 6687
rect 5189 6659 5224 6667
rect 4957 6463 4963 6493
rect 4984 6463 4988 6493
rect 4957 6455 4988 6463
rect 5115 6437 5155 6438
rect 4745 6435 5157 6437
rect 4745 6409 5125 6435
rect 5151 6409 5157 6435
rect 4745 6401 5157 6409
rect 1701 6365 1725 6391
rect 1765 6365 1781 6391
rect 1565 6357 1600 6358
rect 1701 6353 1781 6365
rect 4745 6373 4777 6401
rect 5190 6381 5224 6659
rect 4745 6353 4750 6373
rect 4771 6353 4777 6373
rect 4745 6346 4777 6353
rect 4956 6373 4990 6380
rect 4956 6351 4963 6373
rect 4987 6351 4990 6373
rect 856 6302 967 6306
rect 2611 6302 2818 6303
rect 176 6297 4251 6302
rect 176 6284 4570 6297
rect 176 6264 864 6284
rect 883 6264 941 6284
rect 960 6275 4570 6284
rect 960 6264 4467 6275
rect 176 6255 4467 6264
rect 4486 6255 4544 6275
rect 4563 6255 4570 6275
rect 176 6246 4570 6255
rect 178 6073 285 6246
rect 2773 6244 4570 6246
rect 4459 6238 4570 6244
rect 646 6207 767 6217
rect 646 6205 715 6207
rect 646 6164 659 6205
rect 696 6166 715 6205
rect 752 6166 767 6207
rect 696 6164 767 6166
rect 646 6146 767 6164
rect 4794 6196 4846 6227
rect 4794 6162 4803 6196
rect 4832 6162 4846 6196
rect 169 6046 285 6073
rect 652 6054 717 6146
rect 4794 6136 4846 6162
rect 4956 6145 4990 6351
rect 5168 6376 5224 6381
rect 5168 6356 5175 6376
rect 5195 6356 5224 6376
rect 5168 6349 5224 6356
rect 5168 6348 5203 6349
rect 169 5907 280 6046
rect 650 6008 717 6054
rect 1702 6092 1774 6114
rect 1702 6044 1716 6092
rect 1762 6087 1774 6092
rect 4794 6102 4802 6136
rect 4831 6102 4846 6136
rect 1762 6044 1779 6087
rect 650 5907 715 6008
rect 169 5847 282 5907
rect 650 5869 726 5907
rect 175 5387 282 5847
rect 654 5575 726 5869
rect 1350 5866 1422 5867
rect 1349 5858 1448 5866
rect 1702 5861 1779 6044
rect 2990 6045 3074 6056
rect 2990 6017 3018 6045
rect 3062 6017 3074 6045
rect 2804 5966 2878 5994
rect 2804 5918 2827 5966
rect 2864 5918 2878 5966
rect 2990 5988 3074 6017
rect 2990 5960 3015 5988
rect 3059 5960 3074 5988
rect 2990 5927 3074 5960
rect 2804 5909 2878 5918
rect 2400 5867 2472 5868
rect 1349 5855 1401 5858
rect 1349 5820 1357 5855
rect 1382 5820 1401 5855
rect 1426 5820 1448 5858
rect 1349 5808 1448 5820
rect 1700 5832 1779 5861
rect 2399 5859 2488 5867
rect 2399 5856 2451 5859
rect 1350 5789 1418 5808
rect 1351 5786 1384 5789
rect 1586 5786 1618 5787
rect 761 5725 964 5738
rect 761 5692 785 5725
rect 821 5724 964 5725
rect 821 5721 932 5724
rect 821 5694 858 5721
rect 887 5697 932 5721
rect 961 5697 964 5724
rect 887 5694 964 5697
rect 821 5692 964 5694
rect 761 5679 964 5692
rect 761 5678 862 5679
rect 654 5533 663 5575
rect 712 5533 726 5575
rect 654 5512 726 5533
rect 654 5470 664 5512
rect 713 5470 726 5512
rect 654 5452 726 5470
rect 1139 5616 1171 5623
rect 1139 5596 1146 5616
rect 1167 5596 1171 5616
rect 1139 5531 1171 5596
rect 1351 5587 1382 5786
rect 1583 5781 1618 5786
rect 1583 5761 1590 5781
rect 1610 5761 1618 5781
rect 1583 5753 1618 5761
rect 1351 5557 1357 5587
rect 1378 5557 1382 5587
rect 1351 5549 1382 5557
rect 1509 5531 1549 5532
rect 1139 5529 1551 5531
rect 1139 5503 1519 5529
rect 1545 5503 1551 5529
rect 1139 5495 1551 5503
rect 1139 5467 1171 5495
rect 1584 5475 1618 5753
rect 1700 5566 1770 5832
rect 2399 5821 2407 5856
rect 2432 5821 2451 5856
rect 2476 5821 2488 5859
rect 2399 5809 2488 5821
rect 2399 5808 2468 5809
rect 2399 5790 2435 5808
rect 1809 5721 2012 5734
rect 1809 5688 1833 5721
rect 1869 5720 2012 5721
rect 1869 5717 1980 5720
rect 1869 5690 1906 5717
rect 1935 5693 1980 5717
rect 2009 5693 2012 5720
rect 1935 5690 2012 5693
rect 1869 5688 2012 5690
rect 1809 5675 2012 5688
rect 1809 5674 1910 5675
rect 1139 5447 1144 5467
rect 1165 5447 1171 5467
rect 1139 5440 1171 5447
rect 1562 5470 1618 5475
rect 1562 5450 1569 5470
rect 1589 5450 1618 5470
rect 1695 5560 1770 5566
rect 1695 5527 1703 5560
rect 1756 5527 1770 5560
rect 1695 5502 1770 5527
rect 1695 5469 1708 5502
rect 1761 5469 1770 5502
rect 1695 5460 1770 5469
rect 2187 5612 2219 5619
rect 2187 5592 2194 5612
rect 2215 5592 2219 5612
rect 2187 5527 2219 5592
rect 2399 5583 2430 5790
rect 2634 5782 2666 5783
rect 2631 5777 2666 5782
rect 2631 5757 2638 5777
rect 2658 5757 2666 5777
rect 2631 5749 2666 5757
rect 2399 5553 2405 5583
rect 2426 5553 2430 5583
rect 2399 5545 2430 5553
rect 2557 5527 2597 5528
rect 2187 5525 2599 5527
rect 2187 5499 2567 5525
rect 2593 5499 2599 5525
rect 2187 5491 2599 5499
rect 2187 5463 2219 5491
rect 2632 5471 2666 5749
rect 2815 5564 2877 5909
rect 2984 5882 3074 5927
rect 2984 5567 3066 5882
rect 2815 5545 2879 5564
rect 2815 5506 2828 5545
rect 2862 5506 2879 5545
rect 2815 5487 2879 5506
rect 2984 5526 3005 5567
rect 3041 5526 3066 5567
rect 2984 5497 3066 5526
rect 1695 5455 1753 5460
rect 1562 5443 1618 5450
rect 2187 5443 2192 5463
rect 2213 5443 2219 5463
rect 1562 5442 1597 5443
rect 2187 5436 2219 5443
rect 2610 5466 2666 5471
rect 2610 5446 2617 5466
rect 2637 5446 2666 5466
rect 2610 5439 2666 5446
rect 2610 5438 2645 5439
rect 853 5387 964 5391
rect 2636 5387 4206 5388
rect 175 5369 4206 5387
rect 175 5349 861 5369
rect 880 5349 938 5369
rect 957 5365 4206 5369
rect 957 5349 1909 5365
rect 175 5345 1909 5349
rect 1928 5345 1986 5365
rect 2005 5345 4206 5365
rect 175 5331 4206 5345
rect 175 4708 282 5331
rect 1901 5328 2012 5331
rect 661 5282 725 5286
rect 657 5276 725 5282
rect 657 5243 674 5276
rect 714 5243 725 5276
rect 657 5231 725 5243
rect 1708 5245 1773 5267
rect 657 5229 714 5231
rect 661 4868 712 5229
rect 1708 5206 1725 5245
rect 1770 5206 1773 5245
rect 1349 5161 1384 5163
rect 1349 5152 1453 5161
rect 1349 5151 1400 5152
rect 1349 5131 1352 5151
rect 1377 5132 1400 5151
rect 1432 5132 1453 5152
rect 1377 5131 1453 5132
rect 1349 5124 1453 5131
rect 1349 5112 1384 5124
rect 761 5046 964 5059
rect 761 5013 785 5046
rect 821 5045 964 5046
rect 821 5042 932 5045
rect 821 5015 858 5042
rect 887 5018 932 5042
rect 961 5018 964 5045
rect 887 5015 964 5018
rect 821 5013 964 5015
rect 761 5000 964 5013
rect 761 4999 862 5000
rect 1139 4937 1171 4944
rect 1139 4917 1146 4937
rect 1167 4917 1171 4937
rect 650 4859 715 4868
rect 650 4822 660 4859
rect 700 4825 715 4859
rect 1139 4852 1171 4917
rect 1351 4908 1382 5112
rect 1586 5107 1618 5108
rect 1583 5102 1618 5107
rect 1583 5082 1590 5102
rect 1610 5082 1618 5102
rect 1583 5074 1618 5082
rect 1351 4878 1357 4908
rect 1378 4878 1382 4908
rect 1351 4870 1382 4878
rect 1509 4852 1549 4853
rect 1139 4850 1551 4852
rect 700 4822 717 4825
rect 650 4803 717 4822
rect 650 4782 664 4803
rect 700 4782 717 4803
rect 650 4775 717 4782
rect 1139 4824 1519 4850
rect 1545 4824 1551 4850
rect 1139 4816 1551 4824
rect 1139 4788 1171 4816
rect 1584 4796 1618 5074
rect 1708 4906 1773 5206
rect 2979 5230 3072 5245
rect 2979 5186 2994 5230
rect 3054 5186 3072 5230
rect 1139 4768 1144 4788
rect 1165 4768 1171 4788
rect 1139 4761 1171 4768
rect 1562 4791 1618 4796
rect 1562 4771 1569 4791
rect 1589 4771 1618 4791
rect 1562 4764 1618 4771
rect 1698 4895 1778 4906
rect 1698 4869 1715 4895
rect 1755 4869 1778 4895
rect 1698 4842 1778 4869
rect 1698 4816 1719 4842
rect 1759 4816 1778 4842
rect 1698 4797 1778 4816
rect 1698 4771 1722 4797
rect 1762 4771 1778 4797
rect 1562 4763 1597 4764
rect 1698 4759 1778 4771
rect 2979 4813 3072 5186
rect 3256 5041 3459 5054
rect 3256 5008 3280 5041
rect 3316 5040 3459 5041
rect 3316 5037 3427 5040
rect 3316 5010 3353 5037
rect 3382 5013 3427 5037
rect 3456 5013 3459 5040
rect 3382 5010 3459 5013
rect 3316 5008 3459 5010
rect 3256 4995 3459 5008
rect 3256 4994 3357 4995
rect 2979 4772 2994 4813
rect 3048 4772 3072 4813
rect 2979 4765 3072 4772
rect 3634 4932 3666 4939
rect 3634 4912 3641 4932
rect 3662 4912 3666 4932
rect 3634 4847 3666 4912
rect 3846 4903 3877 5104
rect 4081 5102 4113 5103
rect 4078 5097 4113 5102
rect 4078 5077 4085 5097
rect 4105 5077 4113 5097
rect 4078 5069 4113 5077
rect 3846 4873 3852 4903
rect 3873 4873 3877 4903
rect 3846 4865 3877 4873
rect 4004 4847 4044 4848
rect 3634 4845 4046 4847
rect 3634 4819 4014 4845
rect 4040 4819 4046 4845
rect 3634 4811 4046 4819
rect 3634 4783 3666 4811
rect 4079 4791 4113 5069
rect 3634 4763 3639 4783
rect 3660 4763 3666 4783
rect 3634 4756 3666 4763
rect 4057 4786 4113 4791
rect 4057 4766 4064 4786
rect 4084 4766 4113 4786
rect 4057 4759 4113 4766
rect 4057 4758 4092 4759
rect 853 4708 964 4712
rect 2595 4708 4239 4711
rect 173 4690 4239 4708
rect 173 4670 861 4690
rect 880 4670 938 4690
rect 957 4685 4239 4690
rect 957 4670 3356 4685
rect 173 4665 3356 4670
rect 3375 4665 3433 4685
rect 3452 4665 4239 4685
rect 173 4655 4239 4665
rect 173 4652 798 4655
rect 985 4652 4239 4655
rect 175 4424 282 4652
rect 2595 4651 4239 4652
rect 3348 4648 3459 4651
rect 643 4613 764 4623
rect 643 4611 712 4613
rect 643 4570 656 4611
rect 693 4572 712 4611
rect 749 4572 764 4613
rect 693 4570 764 4572
rect 643 4552 764 4570
rect 3848 4593 3934 4597
rect 3848 4575 3863 4593
rect 3915 4575 3934 4593
rect 3848 4566 3934 4575
rect 649 4450 728 4552
rect 1701 4512 1768 4531
rect 1701 4492 1721 4512
rect 175 4369 283 4424
rect 650 4369 728 4450
rect 1700 4446 1721 4492
rect 1751 4492 1768 4512
rect 1751 4462 1770 4492
rect 1751 4446 1771 4462
rect 1700 4430 1771 4446
rect 1350 4419 1422 4420
rect 1349 4411 1448 4419
rect 1349 4408 1401 4411
rect 1349 4373 1357 4408
rect 1382 4373 1401 4408
rect 1426 4373 1448 4411
rect 175 3940 282 4369
rect 654 4128 726 4369
rect 1349 4361 1448 4373
rect 1350 4342 1418 4361
rect 1351 4339 1384 4342
rect 1586 4339 1618 4340
rect 761 4278 964 4291
rect 761 4245 785 4278
rect 821 4277 964 4278
rect 821 4274 932 4277
rect 821 4247 858 4274
rect 887 4250 932 4274
rect 961 4250 964 4277
rect 887 4247 964 4250
rect 821 4245 964 4247
rect 761 4232 964 4245
rect 761 4231 862 4232
rect 654 4086 663 4128
rect 712 4086 726 4128
rect 654 4065 726 4086
rect 654 4023 664 4065
rect 713 4023 726 4065
rect 654 4005 726 4023
rect 1139 4169 1171 4176
rect 1139 4149 1146 4169
rect 1167 4149 1171 4169
rect 1139 4084 1171 4149
rect 1351 4140 1382 4339
rect 1583 4334 1618 4339
rect 1583 4314 1590 4334
rect 1610 4314 1618 4334
rect 1583 4306 1618 4314
rect 1351 4110 1357 4140
rect 1378 4110 1382 4140
rect 1351 4102 1382 4110
rect 1509 4084 1549 4085
rect 1139 4082 1551 4084
rect 1139 4056 1519 4082
rect 1545 4056 1551 4082
rect 1139 4048 1551 4056
rect 1139 4020 1171 4048
rect 1584 4028 1618 4306
rect 1700 4119 1770 4430
rect 3625 4420 3697 4421
rect 3624 4417 3713 4420
rect 2396 4415 3713 4417
rect 2393 4412 3713 4415
rect 2393 4409 3676 4412
rect 2393 4374 3632 4409
rect 3657 4374 3676 4409
rect 3701 4374 3713 4412
rect 2393 4364 3713 4374
rect 3889 4413 3925 4566
rect 3889 4390 3895 4413
rect 3919 4390 3925 4413
rect 3889 4369 3925 4390
rect 2393 4362 3678 4364
rect 2393 4352 2490 4362
rect 2399 4343 2435 4352
rect 3889 4346 3895 4369
rect 3919 4346 3925 4369
rect 1809 4274 2012 4287
rect 1809 4241 1833 4274
rect 1869 4273 2012 4274
rect 1869 4270 1980 4273
rect 1869 4243 1906 4270
rect 1935 4246 1980 4270
rect 2009 4246 2012 4273
rect 1935 4243 2012 4246
rect 1869 4241 2012 4243
rect 1809 4228 2012 4241
rect 1809 4227 1910 4228
rect 1139 4000 1144 4020
rect 1165 4000 1171 4020
rect 1139 3993 1171 4000
rect 1562 4023 1618 4028
rect 1562 4003 1569 4023
rect 1589 4003 1618 4023
rect 1695 4113 1770 4119
rect 1695 4080 1703 4113
rect 1756 4080 1770 4113
rect 1695 4055 1770 4080
rect 1695 4022 1708 4055
rect 1761 4022 1770 4055
rect 1695 4013 1770 4022
rect 2187 4165 2219 4172
rect 2187 4145 2194 4165
rect 2215 4145 2219 4165
rect 2187 4080 2219 4145
rect 2399 4136 2430 4343
rect 2634 4335 2666 4336
rect 3889 4335 3925 4346
rect 2631 4330 2666 4335
rect 2631 4310 2638 4330
rect 2658 4310 2666 4330
rect 2631 4302 2666 4310
rect 2399 4106 2405 4136
rect 2426 4106 2430 4136
rect 2399 4098 2430 4106
rect 2557 4080 2597 4081
rect 2187 4078 2599 4080
rect 2187 4052 2567 4078
rect 2593 4052 2599 4078
rect 2187 4044 2599 4052
rect 2187 4016 2219 4044
rect 2632 4024 2666 4302
rect 1695 4008 1753 4013
rect 1562 3996 1618 4003
rect 2187 3996 2192 4016
rect 2213 3996 2219 4016
rect 1562 3995 1597 3996
rect 2187 3989 2219 3996
rect 2610 4019 2666 4024
rect 2610 3999 2617 4019
rect 2637 3999 2666 4019
rect 2610 3992 2666 3999
rect 2610 3991 2645 3992
rect 853 3940 964 3944
rect 2728 3940 3887 3941
rect 175 3922 3887 3940
rect 175 3902 861 3922
rect 880 3902 938 3922
rect 957 3918 3887 3922
rect 957 3902 1909 3918
rect 175 3898 1909 3902
rect 1928 3898 1986 3918
rect 2005 3898 3887 3918
rect 175 3884 3887 3898
rect 175 3261 282 3884
rect 1901 3881 2012 3884
rect 661 3835 725 3839
rect 657 3829 725 3835
rect 657 3796 674 3829
rect 714 3796 725 3829
rect 657 3784 725 3796
rect 1708 3798 1773 3820
rect 657 3782 714 3784
rect 661 3421 712 3782
rect 1708 3759 1725 3798
rect 1770 3759 1773 3798
rect 4794 3796 4846 6102
rect 4955 6079 4990 6145
rect 4955 4763 4989 6079
rect 5293 5932 5398 11142
rect 8832 11158 8897 11458
rect 8987 11290 9021 11568
rect 9434 11548 9466 11576
rect 9054 11540 9466 11548
rect 9054 11514 9060 11540
rect 9086 11514 9466 11540
rect 9888 11582 9955 11589
rect 9888 11561 9905 11582
rect 9941 11561 9955 11582
rect 9888 11542 9955 11561
rect 9888 11539 9905 11542
rect 9054 11512 9466 11514
rect 9056 11511 9096 11512
rect 9223 11486 9254 11494
rect 9223 11456 9227 11486
rect 9248 11456 9254 11486
rect 8987 11282 9022 11290
rect 8987 11262 8995 11282
rect 9015 11262 9022 11282
rect 8987 11257 9022 11262
rect 8987 11256 9019 11257
rect 9223 11252 9254 11456
rect 9434 11447 9466 11512
rect 9890 11505 9905 11539
rect 9945 11505 9955 11542
rect 9890 11496 9955 11505
rect 9434 11427 9438 11447
rect 9459 11427 9466 11447
rect 9434 11420 9466 11427
rect 9743 11364 9844 11365
rect 9641 11351 9844 11364
rect 9641 11349 9784 11351
rect 9641 11346 9718 11349
rect 9641 11319 9644 11346
rect 9673 11322 9718 11346
rect 9747 11322 9784 11349
rect 9673 11319 9784 11322
rect 9641 11318 9784 11319
rect 9820 11318 9844 11351
rect 9641 11305 9844 11318
rect 9221 11240 9256 11252
rect 9152 11233 9256 11240
rect 9152 11232 9228 11233
rect 9152 11212 9173 11232
rect 9205 11213 9228 11232
rect 9253 11213 9256 11233
rect 9205 11212 9256 11213
rect 9152 11203 9256 11212
rect 9221 11201 9256 11203
rect 8832 11119 8835 11158
rect 8880 11119 8897 11158
rect 9893 11135 9944 11496
rect 9891 11133 9948 11135
rect 8832 11097 8897 11119
rect 9880 11121 9948 11133
rect 9880 11088 9891 11121
rect 9931 11088 9948 11121
rect 9880 11082 9948 11088
rect 9880 11078 9944 11082
rect 8593 11033 8704 11036
rect 10323 11033 10430 11656
rect 6357 11019 10430 11033
rect 6357 10999 8600 11019
rect 8619 10999 8677 11019
rect 8696 11015 10430 11019
rect 8696 10999 9648 11015
rect 6357 10995 9648 10999
rect 9667 10995 9725 11015
rect 9744 10995 10430 11015
rect 6357 10977 10430 10995
rect 6357 10976 7877 10977
rect 9641 10973 9752 10977
rect 7960 10925 7995 10926
rect 7939 10918 7995 10925
rect 7939 10898 7968 10918
rect 7988 10898 7995 10918
rect 7939 10893 7995 10898
rect 8386 10921 8418 10928
rect 9008 10921 9043 10922
rect 8386 10901 8392 10921
rect 8413 10901 8418 10921
rect 8987 10914 9043 10921
rect 8852 10904 8910 10909
rect 7939 10615 7973 10893
rect 8386 10873 8418 10901
rect 8006 10865 8418 10873
rect 8006 10839 8012 10865
rect 8038 10839 8418 10865
rect 8006 10837 8418 10839
rect 8008 10836 8048 10837
rect 8175 10811 8206 10819
rect 8175 10781 8179 10811
rect 8200 10781 8206 10811
rect 7939 10607 7974 10615
rect 7939 10587 7947 10607
rect 7967 10587 7974 10607
rect 7939 10582 7974 10587
rect 7939 10581 7971 10582
rect 8175 10581 8206 10781
rect 8386 10772 8418 10837
rect 8386 10752 8390 10772
rect 8411 10752 8418 10772
rect 8386 10745 8418 10752
rect 8835 10895 8910 10904
rect 8835 10862 8844 10895
rect 8897 10862 8910 10895
rect 8835 10837 8910 10862
rect 8835 10804 8849 10837
rect 8902 10804 8910 10837
rect 8835 10798 8910 10804
rect 8987 10894 9016 10914
rect 9036 10894 9043 10914
rect 8987 10889 9043 10894
rect 9434 10917 9466 10924
rect 9434 10897 9440 10917
rect 9461 10897 9466 10917
rect 8695 10689 8796 10690
rect 8593 10676 8796 10689
rect 8593 10674 8736 10676
rect 8593 10671 8670 10674
rect 8593 10644 8596 10671
rect 8625 10647 8670 10671
rect 8699 10647 8736 10674
rect 8625 10644 8736 10647
rect 8593 10643 8736 10644
rect 8772 10643 8796 10676
rect 8593 10630 8796 10643
rect 8172 10574 8211 10581
rect 8170 10557 8211 10574
rect 8172 10532 8211 10557
rect 6866 10524 8211 10532
rect 6866 10496 6881 10524
rect 6909 10498 8211 10524
rect 6909 10496 8208 10498
rect 6866 10491 8208 10496
rect 8835 10487 8905 10798
rect 8987 10611 9021 10889
rect 9434 10869 9466 10897
rect 9054 10861 9466 10869
rect 9054 10835 9060 10861
rect 9086 10835 9466 10861
rect 9054 10833 9466 10835
rect 9056 10832 9096 10833
rect 9223 10807 9254 10815
rect 9223 10777 9227 10807
rect 9248 10777 9254 10807
rect 8987 10603 9022 10611
rect 8987 10583 8995 10603
rect 9015 10583 9022 10603
rect 8987 10578 9022 10583
rect 9223 10578 9254 10777
rect 9434 10768 9466 10833
rect 9434 10748 9438 10768
rect 9459 10748 9466 10768
rect 9434 10741 9466 10748
rect 9879 10894 9951 10912
rect 9879 10852 9892 10894
rect 9941 10852 9951 10894
rect 9879 10831 9951 10852
rect 9879 10789 9893 10831
rect 9942 10789 9951 10831
rect 9743 10685 9844 10686
rect 9641 10672 9844 10685
rect 9641 10670 9784 10672
rect 9641 10667 9718 10670
rect 9641 10640 9644 10667
rect 9673 10643 9718 10667
rect 9747 10643 9784 10670
rect 9673 10640 9784 10643
rect 9641 10639 9784 10640
rect 9820 10639 9844 10672
rect 9641 10626 9844 10639
rect 8987 10577 9019 10578
rect 9221 10575 9254 10578
rect 9187 10556 9255 10575
rect 9157 10544 9256 10556
rect 9879 10548 9951 10789
rect 10323 10548 10430 10977
rect 9157 10506 9179 10544
rect 9204 10509 9223 10544
rect 9248 10509 9256 10544
rect 9204 10506 9256 10509
rect 9157 10498 9256 10506
rect 9183 10497 9255 10498
rect 8834 10471 8905 10487
rect 8834 10455 8854 10471
rect 8835 10425 8854 10455
rect 8837 10405 8854 10425
rect 8884 10425 8905 10471
rect 9877 10467 9955 10548
rect 10322 10493 10430 10548
rect 8884 10405 8904 10425
rect 8837 10386 8904 10405
rect 9877 10365 9956 10467
rect 9841 10347 9962 10365
rect 9841 10345 9912 10347
rect 9841 10304 9856 10345
rect 9893 10306 9912 10345
rect 9949 10306 9962 10347
rect 9893 10304 9962 10306
rect 9841 10294 9962 10304
rect 7146 10266 7257 10269
rect 6357 10265 8010 10266
rect 10323 10265 10430 10493
rect 6357 10262 9620 10265
rect 9807 10262 10432 10265
rect 6357 10252 10432 10262
rect 6357 10232 7153 10252
rect 7172 10232 7230 10252
rect 7249 10247 10432 10252
rect 7249 10232 9648 10247
rect 6357 10227 9648 10232
rect 9667 10227 9725 10247
rect 9744 10227 10432 10247
rect 6357 10209 10432 10227
rect 6357 10206 8010 10209
rect 9641 10205 9752 10209
rect 6513 10158 6548 10159
rect 6492 10151 6548 10158
rect 6492 10131 6521 10151
rect 6541 10131 6548 10151
rect 6492 10126 6548 10131
rect 6939 10154 6971 10161
rect 6939 10134 6945 10154
rect 6966 10134 6971 10154
rect 6492 9848 6526 10126
rect 6939 10106 6971 10134
rect 8827 10146 8907 10158
rect 9008 10153 9043 10154
rect 6559 10098 6971 10106
rect 6559 10072 6565 10098
rect 6591 10072 6971 10098
rect 7357 10112 7794 10125
rect 7357 10089 7370 10112
rect 7396 10105 7794 10112
rect 7396 10089 7750 10105
rect 7357 10082 7750 10089
rect 7776 10082 7794 10105
rect 7357 10076 7794 10082
rect 8827 10120 8843 10146
rect 8883 10120 8907 10146
rect 8827 10101 8907 10120
rect 6559 10070 6971 10072
rect 6561 10069 6601 10070
rect 6728 10044 6759 10052
rect 6728 10014 6732 10044
rect 6753 10014 6759 10044
rect 6492 9840 6527 9848
rect 6492 9820 6500 9840
rect 6520 9820 6527 9840
rect 6492 9815 6527 9820
rect 6492 9814 6524 9815
rect 6728 9807 6759 10014
rect 6939 10005 6971 10070
rect 8827 10075 8846 10101
rect 8886 10075 8907 10101
rect 8827 10048 8907 10075
rect 8827 10022 8850 10048
rect 8890 10022 8907 10048
rect 8827 10011 8907 10022
rect 8987 10146 9043 10153
rect 8987 10126 9016 10146
rect 9036 10126 9043 10146
rect 8987 10121 9043 10126
rect 9434 10149 9466 10156
rect 9434 10129 9440 10149
rect 9461 10129 9466 10149
rect 6939 9985 6943 10005
rect 6964 9985 6971 10005
rect 6939 9978 6971 9985
rect 7248 9922 7349 9923
rect 7146 9909 7349 9922
rect 7146 9907 7289 9909
rect 7146 9904 7223 9907
rect 7146 9877 7149 9904
rect 7178 9880 7223 9904
rect 7252 9880 7289 9907
rect 7178 9877 7289 9880
rect 7146 9876 7289 9877
rect 7325 9876 7349 9909
rect 7146 9863 7349 9876
rect 6726 9801 6759 9807
rect 6722 9797 6759 9801
rect 6722 9787 6760 9797
rect 6722 9774 6732 9787
rect 6723 9750 6732 9774
rect 6749 9750 6760 9787
rect 6723 9729 6760 9750
rect 8832 9711 8897 10011
rect 8987 9843 9021 10121
rect 9434 10101 9466 10129
rect 9054 10093 9466 10101
rect 9054 10067 9060 10093
rect 9086 10067 9466 10093
rect 9888 10135 9955 10142
rect 9888 10114 9905 10135
rect 9941 10114 9955 10135
rect 9888 10095 9955 10114
rect 9888 10092 9905 10095
rect 9054 10065 9466 10067
rect 9056 10064 9096 10065
rect 9223 10039 9254 10047
rect 9223 10009 9227 10039
rect 9248 10009 9254 10039
rect 8987 9835 9022 9843
rect 8987 9815 8995 9835
rect 9015 9815 9022 9835
rect 8987 9810 9022 9815
rect 8987 9809 9019 9810
rect 9223 9805 9254 10009
rect 9434 10000 9466 10065
rect 9890 10058 9905 10092
rect 9945 10058 9955 10095
rect 9890 10049 9955 10058
rect 9434 9980 9438 10000
rect 9459 9980 9466 10000
rect 9434 9973 9466 9980
rect 9743 9917 9844 9918
rect 9641 9904 9844 9917
rect 9641 9902 9784 9904
rect 9641 9899 9718 9902
rect 9641 9872 9644 9899
rect 9673 9875 9718 9899
rect 9747 9875 9784 9902
rect 9673 9872 9784 9875
rect 9641 9871 9784 9872
rect 9820 9871 9844 9904
rect 9641 9858 9844 9871
rect 9221 9793 9256 9805
rect 9152 9786 9256 9793
rect 9152 9785 9228 9786
rect 9152 9765 9173 9785
rect 9205 9766 9228 9785
rect 9253 9766 9256 9786
rect 9205 9765 9256 9766
rect 9152 9756 9256 9765
rect 9221 9754 9256 9756
rect 8832 9672 8835 9711
rect 8880 9672 8897 9711
rect 9893 9688 9944 10049
rect 9891 9686 9948 9688
rect 8832 9650 8897 9672
rect 9880 9674 9948 9686
rect 9880 9641 9891 9674
rect 9931 9641 9948 9674
rect 9880 9635 9948 9641
rect 9880 9631 9944 9635
rect 8593 9586 8704 9589
rect 10323 9586 10430 10209
rect 5980 9572 10430 9586
rect 5980 9552 8600 9572
rect 8619 9552 8677 9572
rect 8696 9568 10430 9572
rect 8696 9552 9648 9568
rect 5980 9548 9648 9552
rect 9667 9548 9725 9568
rect 9744 9548 10430 9568
rect 5980 9534 10430 9548
rect 6399 9530 10430 9534
rect 6399 9529 7969 9530
rect 9641 9526 9752 9530
rect 7960 9478 7995 9479
rect 7939 9471 7995 9478
rect 7939 9451 7968 9471
rect 7988 9451 7995 9471
rect 7939 9446 7995 9451
rect 8386 9474 8418 9481
rect 9008 9474 9043 9475
rect 8386 9454 8392 9474
rect 8413 9454 8418 9474
rect 8987 9467 9043 9474
rect 8852 9457 8910 9462
rect 7939 9168 7973 9446
rect 8386 9426 8418 9454
rect 8006 9418 8418 9426
rect 8006 9392 8012 9418
rect 8038 9392 8418 9418
rect 8006 9390 8418 9392
rect 8008 9389 8048 9390
rect 8175 9364 8206 9372
rect 8175 9334 8179 9364
rect 8200 9334 8206 9364
rect 7939 9160 7974 9168
rect 7939 9140 7947 9160
rect 7967 9140 7974 9160
rect 7939 9135 7974 9140
rect 7939 9134 7971 9135
rect 8175 9127 8206 9334
rect 8386 9325 8418 9390
rect 8386 9305 8390 9325
rect 8411 9305 8418 9325
rect 8386 9298 8418 9305
rect 8835 9448 8910 9457
rect 8835 9415 8844 9448
rect 8897 9415 8910 9448
rect 8835 9390 8910 9415
rect 8835 9357 8849 9390
rect 8902 9357 8910 9390
rect 8835 9351 8910 9357
rect 8987 9447 9016 9467
rect 9036 9447 9043 9467
rect 8987 9442 9043 9447
rect 9434 9470 9466 9477
rect 9434 9450 9440 9470
rect 9461 9450 9466 9470
rect 8695 9242 8796 9243
rect 8593 9229 8796 9242
rect 8593 9227 8736 9229
rect 8593 9224 8670 9227
rect 8593 9197 8596 9224
rect 8625 9200 8670 9224
rect 8699 9200 8736 9227
rect 8625 9197 8736 9200
rect 8593 9196 8736 9197
rect 8772 9196 8796 9229
rect 8593 9183 8796 9196
rect 7673 9114 7837 9117
rect 8170 9114 8206 9127
rect 6872 9096 8211 9114
rect 6872 9058 6882 9096
rect 6907 9081 8211 9096
rect 6907 9058 6917 9081
rect 7673 9074 7837 9081
rect 6872 9050 6917 9058
rect 6886 9049 6917 9050
rect 8835 9035 8905 9351
rect 8987 9164 9021 9442
rect 9434 9422 9466 9450
rect 9054 9414 9466 9422
rect 9054 9388 9060 9414
rect 9086 9388 9466 9414
rect 9054 9386 9466 9388
rect 9056 9385 9096 9386
rect 9223 9360 9254 9368
rect 9223 9330 9227 9360
rect 9248 9330 9254 9360
rect 8987 9156 9022 9164
rect 8987 9136 8995 9156
rect 9015 9136 9022 9156
rect 8987 9131 9022 9136
rect 9223 9131 9254 9330
rect 9434 9321 9466 9386
rect 9434 9301 9438 9321
rect 9459 9301 9466 9321
rect 9434 9294 9466 9301
rect 9879 9447 9951 9465
rect 9879 9405 9892 9447
rect 9941 9405 9951 9447
rect 9879 9384 9951 9405
rect 9879 9342 9893 9384
rect 9942 9342 9951 9384
rect 9743 9238 9844 9239
rect 9641 9225 9844 9238
rect 9641 9223 9784 9225
rect 9641 9220 9718 9223
rect 9641 9193 9644 9220
rect 9673 9196 9718 9220
rect 9747 9196 9784 9223
rect 9673 9193 9784 9196
rect 9641 9192 9784 9193
rect 9820 9192 9844 9225
rect 9641 9179 9844 9192
rect 8987 9130 9019 9131
rect 9221 9128 9254 9131
rect 9187 9109 9255 9128
rect 9157 9097 9256 9109
rect 9157 9059 9179 9097
rect 9204 9062 9223 9097
rect 9248 9062 9256 9097
rect 9204 9059 9256 9062
rect 9157 9051 9256 9059
rect 9183 9050 9255 9051
rect 8835 9016 8914 9035
rect 8838 8996 8914 9016
rect 8831 8972 8914 8996
rect 9879 9031 9951 9342
rect 9879 8988 9955 9031
rect 8831 8906 8843 8972
rect 8897 8906 8914 8972
rect 8831 8886 8914 8906
rect 8831 8849 8848 8886
rect 8892 8872 8914 8886
rect 9880 8937 9955 8988
rect 10323 8937 10430 9530
rect 8892 8849 8907 8872
rect 8831 8833 8907 8849
rect 9880 8845 9957 8937
rect 10323 8933 10431 8937
rect 9842 8827 9963 8845
rect 9842 8825 9913 8827
rect 9842 8784 9857 8825
rect 9894 8786 9913 8825
rect 9950 8786 9963 8827
rect 9894 8784 9963 8786
rect 9842 8774 9963 8784
rect 6367 8745 7836 8747
rect 10324 8745 10431 8933
rect 6367 8730 10433 8745
rect 6367 8710 7111 8730
rect 7130 8710 7188 8730
rect 7207 8727 10433 8730
rect 7207 8710 9649 8727
rect 6367 8707 9649 8710
rect 9668 8707 9726 8727
rect 9745 8707 10433 8727
rect 6367 8689 10433 8707
rect 7104 8688 7215 8689
rect 7791 8688 7998 8689
rect 9642 8685 9753 8689
rect 6471 8636 6506 8637
rect 6450 8629 6506 8636
rect 6450 8609 6479 8629
rect 6499 8609 6506 8629
rect 6450 8604 6506 8609
rect 6897 8632 6929 8639
rect 6897 8612 6903 8632
rect 6924 8612 6929 8632
rect 6450 8326 6484 8604
rect 6897 8584 6929 8612
rect 6517 8576 6929 8584
rect 6517 8550 6523 8576
rect 6549 8550 6929 8576
rect 6517 8548 6929 8550
rect 6519 8547 6559 8548
rect 6686 8522 6717 8530
rect 6686 8492 6690 8522
rect 6711 8492 6717 8522
rect 6450 8318 6485 8326
rect 6450 8298 6458 8318
rect 6478 8298 6485 8318
rect 6450 8293 6485 8298
rect 6686 8296 6717 8492
rect 6897 8483 6929 8548
rect 8828 8626 8908 8638
rect 9009 8633 9044 8634
rect 8828 8600 8844 8626
rect 8884 8600 8908 8626
rect 8828 8581 8908 8600
rect 8828 8555 8847 8581
rect 8887 8555 8908 8581
rect 8828 8528 8908 8555
rect 8828 8502 8851 8528
rect 8891 8502 8908 8528
rect 8828 8491 8908 8502
rect 8988 8626 9044 8633
rect 8988 8606 9017 8626
rect 9037 8606 9044 8626
rect 8988 8601 9044 8606
rect 9435 8629 9467 8636
rect 9435 8609 9441 8629
rect 9462 8609 9467 8629
rect 6897 8463 6901 8483
rect 6922 8463 6929 8483
rect 6897 8456 6929 8463
rect 7206 8400 7307 8401
rect 7104 8387 7307 8400
rect 7104 8385 7247 8387
rect 7104 8382 7181 8385
rect 7104 8355 7107 8382
rect 7136 8358 7181 8382
rect 7210 8358 7247 8385
rect 7136 8355 7247 8358
rect 7104 8354 7247 8355
rect 7283 8354 7307 8387
rect 7104 8341 7307 8354
rect 6450 8292 6482 8293
rect 6686 8207 6720 8296
rect 6307 8203 6720 8207
rect 5293 5878 5310 5932
rect 5373 5878 5398 5932
rect 5293 5857 5398 5878
rect 5760 8158 6720 8203
rect 8833 8191 8898 8491
rect 8988 8323 9022 8601
rect 9435 8581 9467 8609
rect 9055 8573 9467 8581
rect 9055 8547 9061 8573
rect 9087 8547 9467 8573
rect 9889 8615 9956 8622
rect 9889 8594 9906 8615
rect 9942 8594 9956 8615
rect 9889 8575 9956 8594
rect 9889 8572 9906 8575
rect 9055 8545 9467 8547
rect 9057 8544 9097 8545
rect 9224 8519 9255 8527
rect 9224 8489 9228 8519
rect 9249 8489 9255 8519
rect 8988 8315 9023 8323
rect 8988 8295 8996 8315
rect 9016 8295 9023 8315
rect 8988 8290 9023 8295
rect 8988 8289 9020 8290
rect 9224 8285 9255 8489
rect 9435 8480 9467 8545
rect 9891 8538 9906 8572
rect 9946 8538 9956 8575
rect 9891 8529 9956 8538
rect 9435 8460 9439 8480
rect 9460 8460 9467 8480
rect 9435 8453 9467 8460
rect 9744 8397 9845 8398
rect 9642 8384 9845 8397
rect 9642 8382 9785 8384
rect 9642 8379 9719 8382
rect 9642 8352 9645 8379
rect 9674 8355 9719 8379
rect 9748 8355 9785 8382
rect 9674 8352 9785 8355
rect 9642 8351 9785 8352
rect 9821 8351 9845 8384
rect 9642 8338 9845 8351
rect 9222 8273 9257 8285
rect 9153 8266 9257 8273
rect 9153 8265 9229 8266
rect 9153 8245 9174 8265
rect 9206 8246 9229 8265
rect 9254 8246 9257 8266
rect 9206 8245 9257 8246
rect 9153 8236 9257 8245
rect 9222 8234 9257 8236
rect 5760 8154 6357 8158
rect 5760 5848 5812 8154
rect 8833 8152 8836 8191
rect 8881 8152 8898 8191
rect 9894 8168 9945 8529
rect 9892 8166 9949 8168
rect 8833 8130 8898 8152
rect 9881 8154 9949 8166
rect 9881 8121 9892 8154
rect 9932 8121 9949 8154
rect 9881 8115 9949 8121
rect 9881 8111 9945 8115
rect 8594 8066 8705 8069
rect 10324 8066 10431 8689
rect 6719 8052 10431 8066
rect 6719 8032 8601 8052
rect 8620 8032 8678 8052
rect 8697 8048 10431 8052
rect 8697 8032 9649 8048
rect 6719 8028 9649 8032
rect 9668 8028 9726 8048
rect 9745 8028 10431 8048
rect 6719 8010 10431 8028
rect 6719 8009 7878 8010
rect 9642 8006 9753 8010
rect 7961 7958 7996 7959
rect 7940 7951 7996 7958
rect 7940 7931 7969 7951
rect 7989 7931 7996 7951
rect 7940 7926 7996 7931
rect 8387 7954 8419 7961
rect 9009 7954 9044 7955
rect 8387 7934 8393 7954
rect 8414 7934 8419 7954
rect 8988 7947 9044 7954
rect 8853 7937 8911 7942
rect 7940 7648 7974 7926
rect 8387 7906 8419 7934
rect 8007 7898 8419 7906
rect 8007 7872 8013 7898
rect 8039 7872 8419 7898
rect 8007 7870 8419 7872
rect 8009 7869 8049 7870
rect 8176 7844 8207 7852
rect 8176 7814 8180 7844
rect 8201 7814 8207 7844
rect 7940 7640 7975 7648
rect 7940 7620 7948 7640
rect 7968 7620 7975 7640
rect 7940 7615 7975 7620
rect 6681 7604 6717 7615
rect 7940 7614 7972 7615
rect 8176 7607 8207 7814
rect 8387 7805 8419 7870
rect 8387 7785 8391 7805
rect 8412 7785 8419 7805
rect 8387 7778 8419 7785
rect 8836 7928 8911 7937
rect 8836 7895 8845 7928
rect 8898 7895 8911 7928
rect 8836 7870 8911 7895
rect 8836 7837 8850 7870
rect 8903 7837 8911 7870
rect 8836 7831 8911 7837
rect 8988 7927 9017 7947
rect 9037 7927 9044 7947
rect 8988 7922 9044 7927
rect 9435 7950 9467 7957
rect 9435 7930 9441 7950
rect 9462 7930 9467 7950
rect 8696 7722 8797 7723
rect 8594 7709 8797 7722
rect 8594 7707 8737 7709
rect 8594 7704 8671 7707
rect 8594 7677 8597 7704
rect 8626 7680 8671 7704
rect 8700 7680 8737 7707
rect 8626 7677 8737 7680
rect 8594 7676 8737 7677
rect 8773 7676 8797 7709
rect 8594 7663 8797 7676
rect 6681 7581 6687 7604
rect 6711 7581 6717 7604
rect 8171 7598 8207 7607
rect 8116 7588 8213 7598
rect 6928 7586 8213 7588
rect 6681 7560 6717 7581
rect 6681 7537 6687 7560
rect 6711 7537 6717 7560
rect 6681 7384 6717 7537
rect 6893 7576 8213 7586
rect 6893 7538 6905 7576
rect 6930 7541 6949 7576
rect 6974 7541 8213 7576
rect 6930 7538 8213 7541
rect 6893 7535 8213 7538
rect 6893 7533 8210 7535
rect 6893 7530 6982 7533
rect 6909 7529 6981 7530
rect 8836 7520 8906 7831
rect 8988 7644 9022 7922
rect 9435 7902 9467 7930
rect 9055 7894 9467 7902
rect 9055 7868 9061 7894
rect 9087 7868 9467 7894
rect 9055 7866 9467 7868
rect 9057 7865 9097 7866
rect 9224 7840 9255 7848
rect 9224 7810 9228 7840
rect 9249 7810 9255 7840
rect 8988 7636 9023 7644
rect 8988 7616 8996 7636
rect 9016 7616 9023 7636
rect 8988 7611 9023 7616
rect 9224 7611 9255 7810
rect 9435 7801 9467 7866
rect 9435 7781 9439 7801
rect 9460 7781 9467 7801
rect 9435 7774 9467 7781
rect 9880 7927 9952 7945
rect 9880 7885 9893 7927
rect 9942 7885 9952 7927
rect 9880 7864 9952 7885
rect 9880 7822 9894 7864
rect 9943 7822 9952 7864
rect 9744 7718 9845 7719
rect 9642 7705 9845 7718
rect 9642 7703 9785 7705
rect 9642 7700 9719 7703
rect 9642 7673 9645 7700
rect 9674 7676 9719 7700
rect 9748 7676 9785 7703
rect 9674 7673 9785 7676
rect 9642 7672 9785 7673
rect 9821 7672 9845 7705
rect 9642 7659 9845 7672
rect 8988 7610 9020 7611
rect 9222 7608 9255 7611
rect 9188 7589 9256 7608
rect 9158 7577 9257 7589
rect 9880 7581 9952 7822
rect 10324 7581 10431 8010
rect 9158 7539 9180 7577
rect 9205 7542 9224 7577
rect 9249 7542 9257 7577
rect 9205 7539 9257 7542
rect 9158 7531 9257 7539
rect 9184 7530 9256 7531
rect 8835 7504 8906 7520
rect 8835 7488 8855 7504
rect 8836 7458 8855 7488
rect 8838 7438 8855 7458
rect 8885 7458 8906 7504
rect 9878 7500 9956 7581
rect 10323 7526 10431 7581
rect 8885 7438 8905 7458
rect 8838 7419 8905 7438
rect 9878 7398 9957 7500
rect 6672 7375 6758 7384
rect 6672 7357 6691 7375
rect 6743 7357 6758 7375
rect 6672 7353 6758 7357
rect 9842 7380 9963 7398
rect 9842 7378 9913 7380
rect 9842 7337 9857 7378
rect 9894 7339 9913 7378
rect 9950 7339 9963 7380
rect 9894 7337 9963 7339
rect 9842 7327 9963 7337
rect 7147 7299 7258 7302
rect 6367 7298 8011 7299
rect 10324 7298 10431 7526
rect 6367 7295 9621 7298
rect 9808 7295 10433 7298
rect 6367 7285 10433 7295
rect 6367 7265 7154 7285
rect 7173 7265 7231 7285
rect 7250 7280 10433 7285
rect 7250 7265 9649 7280
rect 6367 7260 9649 7265
rect 9668 7260 9726 7280
rect 9745 7260 10433 7280
rect 6367 7242 10433 7260
rect 6367 7239 8011 7242
rect 9642 7238 9753 7242
rect 6514 7191 6549 7192
rect 6493 7184 6549 7191
rect 6493 7164 6522 7184
rect 6542 7164 6549 7184
rect 6493 7159 6549 7164
rect 6940 7187 6972 7194
rect 6940 7167 6946 7187
rect 6967 7167 6972 7187
rect 6493 6881 6527 7159
rect 6940 7139 6972 7167
rect 6560 7131 6972 7139
rect 6560 7105 6566 7131
rect 6592 7105 6972 7131
rect 6560 7103 6972 7105
rect 6562 7102 6602 7103
rect 6729 7077 6760 7085
rect 6729 7047 6733 7077
rect 6754 7047 6760 7077
rect 6493 6873 6528 6881
rect 6493 6853 6501 6873
rect 6521 6853 6528 6873
rect 6493 6848 6528 6853
rect 6493 6847 6525 6848
rect 6729 6846 6760 7047
rect 6940 7038 6972 7103
rect 6940 7018 6944 7038
rect 6965 7018 6972 7038
rect 6940 7011 6972 7018
rect 7534 7178 7627 7185
rect 7534 7137 7558 7178
rect 7612 7137 7627 7178
rect 7249 6955 7350 6956
rect 7147 6942 7350 6955
rect 7147 6940 7290 6942
rect 7147 6937 7224 6940
rect 7147 6910 7150 6937
rect 7179 6913 7224 6937
rect 7253 6913 7290 6940
rect 7179 6910 7290 6913
rect 7147 6909 7290 6910
rect 7326 6909 7350 6942
rect 7147 6896 7350 6909
rect 7534 6764 7627 7137
rect 8828 7179 8908 7191
rect 9009 7186 9044 7187
rect 8828 7153 8844 7179
rect 8884 7153 8908 7179
rect 8828 7134 8908 7153
rect 8828 7108 8847 7134
rect 8887 7108 8908 7134
rect 8828 7081 8908 7108
rect 8828 7055 8851 7081
rect 8891 7055 8908 7081
rect 8828 7044 8908 7055
rect 8988 7179 9044 7186
rect 8988 7159 9017 7179
rect 9037 7159 9044 7179
rect 8988 7154 9044 7159
rect 9435 7182 9467 7189
rect 9435 7162 9441 7182
rect 9462 7162 9467 7182
rect 7534 6720 7552 6764
rect 7612 6720 7627 6764
rect 7534 6705 7627 6720
rect 8833 6744 8898 7044
rect 8988 6876 9022 7154
rect 9435 7134 9467 7162
rect 9055 7126 9467 7134
rect 9055 7100 9061 7126
rect 9087 7100 9467 7126
rect 9889 7168 9956 7175
rect 9889 7147 9906 7168
rect 9942 7147 9956 7168
rect 9889 7128 9956 7147
rect 9889 7125 9906 7128
rect 9055 7098 9467 7100
rect 9057 7097 9097 7098
rect 9224 7072 9255 7080
rect 9224 7042 9228 7072
rect 9249 7042 9255 7072
rect 8988 6868 9023 6876
rect 8988 6848 8996 6868
rect 9016 6848 9023 6868
rect 8988 6843 9023 6848
rect 8988 6842 9020 6843
rect 9224 6838 9255 7042
rect 9435 7033 9467 7098
rect 9891 7091 9906 7125
rect 9946 7091 9956 7128
rect 9891 7082 9956 7091
rect 9435 7013 9439 7033
rect 9460 7013 9467 7033
rect 9435 7006 9467 7013
rect 9744 6950 9845 6951
rect 9642 6937 9845 6950
rect 9642 6935 9785 6937
rect 9642 6932 9719 6935
rect 9642 6905 9645 6932
rect 9674 6908 9719 6932
rect 9748 6908 9785 6935
rect 9674 6905 9785 6908
rect 9642 6904 9785 6905
rect 9821 6904 9845 6937
rect 9642 6891 9845 6904
rect 9222 6826 9257 6838
rect 9153 6819 9257 6826
rect 9153 6818 9229 6819
rect 9153 6798 9174 6818
rect 9206 6799 9229 6818
rect 9254 6799 9257 6819
rect 9206 6798 9257 6799
rect 9153 6789 9257 6798
rect 9222 6787 9257 6789
rect 8833 6705 8836 6744
rect 8881 6705 8898 6744
rect 9894 6721 9945 7082
rect 9892 6719 9949 6721
rect 8833 6683 8898 6705
rect 9881 6707 9949 6719
rect 9881 6674 9892 6707
rect 9932 6674 9949 6707
rect 9881 6668 9949 6674
rect 9881 6664 9945 6668
rect 8594 6619 8705 6622
rect 10324 6619 10431 7242
rect 6400 6605 10431 6619
rect 6400 6585 8601 6605
rect 8620 6585 8678 6605
rect 8697 6601 10431 6605
rect 8697 6585 9649 6601
rect 6400 6581 9649 6585
rect 9668 6581 9726 6601
rect 9745 6581 10431 6601
rect 6400 6563 10431 6581
rect 6400 6562 7970 6563
rect 9642 6559 9753 6563
rect 7961 6511 7996 6512
rect 7940 6504 7996 6511
rect 7940 6484 7969 6504
rect 7989 6484 7996 6504
rect 7940 6479 7996 6484
rect 8387 6507 8419 6514
rect 9009 6507 9044 6508
rect 8387 6487 8393 6507
rect 8414 6487 8419 6507
rect 8988 6500 9044 6507
rect 8853 6490 8911 6495
rect 7540 6424 7622 6453
rect 7540 6383 7565 6424
rect 7601 6383 7622 6424
rect 7727 6444 7791 6463
rect 7727 6405 7744 6444
rect 7778 6405 7791 6444
rect 7727 6386 7791 6405
rect 7540 6068 7622 6383
rect 7532 6023 7622 6068
rect 7729 6041 7791 6386
rect 7940 6201 7974 6479
rect 8387 6459 8419 6487
rect 8007 6451 8419 6459
rect 8007 6425 8013 6451
rect 8039 6425 8419 6451
rect 8007 6423 8419 6425
rect 8009 6422 8049 6423
rect 8176 6397 8207 6405
rect 8176 6367 8180 6397
rect 8201 6367 8207 6397
rect 7940 6193 7975 6201
rect 7940 6173 7948 6193
rect 7968 6173 7975 6193
rect 7940 6168 7975 6173
rect 7940 6167 7972 6168
rect 8176 6160 8207 6367
rect 8387 6358 8419 6423
rect 8387 6338 8391 6358
rect 8412 6338 8419 6358
rect 8387 6331 8419 6338
rect 8836 6481 8911 6490
rect 8836 6448 8845 6481
rect 8898 6448 8911 6481
rect 8836 6423 8911 6448
rect 8836 6390 8850 6423
rect 8903 6390 8911 6423
rect 8836 6384 8911 6390
rect 8988 6480 9017 6500
rect 9037 6480 9044 6500
rect 8988 6475 9044 6480
rect 9435 6503 9467 6510
rect 9435 6483 9441 6503
rect 9462 6483 9467 6503
rect 8696 6275 8797 6276
rect 8594 6262 8797 6275
rect 8594 6260 8737 6262
rect 8594 6257 8671 6260
rect 8594 6230 8597 6257
rect 8626 6233 8671 6257
rect 8700 6233 8737 6260
rect 8626 6230 8737 6233
rect 8594 6229 8737 6230
rect 8773 6229 8797 6262
rect 8594 6216 8797 6229
rect 8171 6142 8207 6160
rect 8138 6141 8207 6142
rect 8118 6129 8207 6141
rect 8118 6091 8130 6129
rect 8155 6094 8174 6129
rect 8199 6094 8207 6129
rect 8836 6118 8906 6384
rect 8988 6197 9022 6475
rect 9435 6455 9467 6483
rect 9055 6447 9467 6455
rect 9055 6421 9061 6447
rect 9087 6421 9467 6447
rect 9055 6419 9467 6421
rect 9057 6418 9097 6419
rect 9224 6393 9255 6401
rect 9224 6363 9228 6393
rect 9249 6363 9255 6393
rect 8988 6189 9023 6197
rect 8988 6169 8996 6189
rect 9016 6169 9023 6189
rect 8988 6164 9023 6169
rect 9224 6164 9255 6363
rect 9435 6354 9467 6419
rect 9435 6334 9439 6354
rect 9460 6334 9467 6354
rect 9435 6327 9467 6334
rect 9880 6480 9952 6498
rect 9880 6438 9893 6480
rect 9942 6438 9952 6480
rect 9880 6417 9952 6438
rect 9880 6375 9894 6417
rect 9943 6375 9952 6417
rect 9744 6271 9845 6272
rect 9642 6258 9845 6271
rect 9642 6256 9785 6258
rect 9642 6253 9719 6256
rect 9642 6226 9645 6253
rect 9674 6229 9719 6253
rect 9748 6229 9785 6256
rect 9674 6226 9785 6229
rect 9642 6225 9785 6226
rect 9821 6225 9845 6258
rect 9642 6212 9845 6225
rect 8988 6163 9020 6164
rect 9222 6161 9255 6164
rect 9188 6142 9256 6161
rect 8155 6091 8207 6094
rect 8118 6083 8207 6091
rect 8827 6089 8906 6118
rect 9158 6130 9257 6142
rect 9158 6092 9180 6130
rect 9205 6095 9224 6130
rect 9249 6095 9257 6130
rect 9205 6092 9257 6095
rect 8134 6082 8206 6083
rect 7728 6032 7802 6041
rect 7532 5990 7616 6023
rect 7532 5962 7547 5990
rect 7591 5962 7616 5990
rect 7532 5933 7616 5962
rect 7728 5984 7742 6032
rect 7779 5984 7802 6032
rect 7728 5956 7802 5984
rect 7532 5905 7544 5933
rect 7588 5905 7616 5933
rect 7532 5894 7616 5905
rect 8827 5906 8904 6089
rect 9158 6084 9257 6092
rect 9184 6083 9256 6084
rect 9880 6081 9952 6375
rect 10324 6103 10431 6563
rect 9880 6043 9956 6081
rect 10324 6043 10437 6103
rect 9891 5942 9956 6043
rect 8827 5863 8844 5906
rect 5760 5814 5775 5848
rect 5804 5814 5812 5848
rect 8832 5858 8844 5863
rect 8890 5858 8904 5906
rect 8832 5836 8904 5858
rect 9889 5896 9956 5942
rect 10326 5904 10437 6043
rect 5760 5788 5812 5814
rect 9889 5804 9954 5896
rect 10321 5877 10437 5904
rect 5760 5754 5774 5788
rect 5803 5754 5812 5788
rect 5760 5723 5812 5754
rect 9839 5786 9960 5804
rect 9839 5784 9910 5786
rect 9839 5743 9854 5784
rect 9891 5745 9910 5784
rect 9947 5745 9960 5786
rect 9891 5743 9960 5745
rect 9839 5733 9960 5743
rect 6036 5706 6147 5712
rect 6036 5704 7833 5706
rect 10321 5704 10428 5877
rect 6036 5695 10430 5704
rect 6036 5675 6043 5695
rect 6062 5675 6120 5695
rect 6139 5686 10430 5695
rect 6139 5675 9646 5686
rect 6036 5666 9646 5675
rect 9665 5666 9723 5686
rect 9742 5666 10430 5686
rect 6036 5653 10430 5666
rect 6355 5648 10430 5653
rect 7788 5647 7995 5648
rect 9639 5644 9750 5648
rect 5403 5601 5438 5602
rect 5382 5594 5438 5601
rect 5382 5574 5411 5594
rect 5431 5574 5438 5594
rect 5382 5569 5438 5574
rect 5829 5597 5861 5604
rect 5829 5577 5835 5597
rect 5856 5577 5861 5597
rect 5382 5291 5416 5569
rect 5829 5549 5861 5577
rect 8825 5585 8905 5597
rect 9006 5592 9041 5593
rect 8825 5559 8841 5585
rect 8881 5559 8905 5585
rect 5449 5541 5861 5549
rect 5449 5515 5455 5541
rect 5481 5515 5861 5541
rect 5449 5513 5861 5515
rect 5451 5512 5491 5513
rect 5618 5487 5649 5495
rect 5618 5457 5622 5487
rect 5643 5457 5649 5487
rect 5382 5283 5417 5291
rect 5382 5263 5390 5283
rect 5410 5263 5417 5283
rect 5618 5272 5649 5457
rect 5829 5448 5861 5513
rect 6243 5546 6354 5553
rect 6243 5545 6322 5546
rect 6243 5521 6265 5545
rect 6289 5522 6322 5545
rect 6346 5522 6354 5546
rect 6289 5521 6354 5522
rect 6243 5511 6354 5521
rect 8825 5540 8905 5559
rect 8825 5514 8844 5540
rect 8884 5514 8905 5540
rect 6304 5494 6353 5511
rect 8825 5487 8905 5514
rect 8825 5461 8848 5487
rect 8888 5461 8905 5487
rect 8825 5450 8905 5461
rect 8985 5585 9041 5592
rect 8985 5565 9014 5585
rect 9034 5565 9041 5585
rect 8985 5560 9041 5565
rect 9432 5588 9464 5595
rect 9432 5568 9438 5588
rect 9459 5568 9464 5588
rect 5829 5428 5833 5448
rect 5854 5428 5861 5448
rect 5829 5421 5861 5428
rect 6138 5365 6239 5366
rect 6036 5352 6239 5365
rect 6036 5350 6179 5352
rect 6036 5347 6113 5350
rect 6036 5320 6039 5347
rect 6068 5323 6113 5347
rect 6142 5323 6179 5350
rect 6068 5320 6179 5323
rect 6036 5319 6179 5320
rect 6215 5319 6239 5352
rect 6036 5306 6239 5319
rect 5382 5258 5417 5263
rect 5382 5257 5414 5258
rect 5616 5195 5650 5272
rect 4249 3792 4846 3796
rect 1349 3714 1384 3716
rect 1349 3705 1453 3714
rect 1349 3704 1400 3705
rect 1349 3684 1352 3704
rect 1377 3685 1400 3704
rect 1432 3685 1453 3705
rect 1377 3684 1453 3685
rect 1349 3677 1453 3684
rect 1349 3665 1384 3677
rect 761 3599 964 3612
rect 761 3566 785 3599
rect 821 3598 964 3599
rect 821 3595 932 3598
rect 821 3568 858 3595
rect 887 3571 932 3595
rect 961 3571 964 3598
rect 887 3568 964 3571
rect 821 3566 964 3568
rect 761 3553 964 3566
rect 761 3552 862 3553
rect 1139 3490 1171 3497
rect 1139 3470 1146 3490
rect 1167 3470 1171 3490
rect 650 3412 715 3421
rect 650 3375 660 3412
rect 700 3378 715 3412
rect 1139 3405 1171 3470
rect 1351 3461 1382 3665
rect 1586 3660 1618 3661
rect 1583 3655 1618 3660
rect 1583 3635 1590 3655
rect 1610 3635 1618 3655
rect 1583 3627 1618 3635
rect 1351 3431 1357 3461
rect 1378 3431 1382 3461
rect 1351 3423 1382 3431
rect 1509 3405 1549 3406
rect 1139 3403 1551 3405
rect 700 3375 717 3378
rect 650 3356 717 3375
rect 650 3335 664 3356
rect 700 3335 717 3356
rect 650 3328 717 3335
rect 1139 3377 1519 3403
rect 1545 3377 1551 3403
rect 1139 3369 1551 3377
rect 1139 3341 1171 3369
rect 1584 3349 1618 3627
rect 1708 3459 1773 3759
rect 3886 3747 4846 3792
rect 4953 4135 4989 4763
rect 3886 3743 4299 3747
rect 3886 3654 3920 3743
rect 4124 3657 4156 3658
rect 3299 3596 3502 3609
rect 3299 3563 3323 3596
rect 3359 3595 3502 3596
rect 3359 3592 3470 3595
rect 3359 3565 3396 3592
rect 3425 3568 3470 3592
rect 3499 3568 3502 3595
rect 3425 3565 3502 3568
rect 3359 3563 3502 3565
rect 3299 3550 3502 3563
rect 3299 3549 3400 3550
rect 3677 3487 3709 3494
rect 3677 3467 3684 3487
rect 3705 3467 3709 3487
rect 1139 3321 1144 3341
rect 1165 3321 1171 3341
rect 1139 3314 1171 3321
rect 1562 3344 1618 3349
rect 1562 3324 1569 3344
rect 1589 3324 1618 3344
rect 1562 3317 1618 3324
rect 1698 3448 1778 3459
rect 1698 3422 1715 3448
rect 1755 3422 1778 3448
rect 1698 3395 1778 3422
rect 1698 3369 1719 3395
rect 1759 3369 1778 3395
rect 1698 3350 1778 3369
rect 1698 3324 1722 3350
rect 1762 3324 1778 3350
rect 1562 3316 1597 3317
rect 1698 3312 1778 3324
rect 3677 3402 3709 3467
rect 3889 3458 3920 3654
rect 4121 3652 4156 3657
rect 4121 3632 4128 3652
rect 4148 3632 4156 3652
rect 4121 3624 4156 3632
rect 3889 3428 3895 3458
rect 3916 3428 3920 3458
rect 3889 3420 3920 3428
rect 4047 3402 4087 3403
rect 3677 3400 4089 3402
rect 3677 3374 4057 3400
rect 4083 3374 4089 3400
rect 3677 3366 4089 3374
rect 3677 3338 3709 3366
rect 4122 3346 4156 3624
rect 3677 3318 3682 3338
rect 3703 3318 3709 3338
rect 3677 3311 3709 3318
rect 4100 3341 4156 3346
rect 4100 3321 4107 3341
rect 4127 3321 4156 3341
rect 4100 3314 4156 3321
rect 4100 3313 4135 3314
rect 853 3261 964 3265
rect 2608 3261 2815 3262
rect 3391 3261 3502 3262
rect 173 3243 4239 3261
rect 173 3223 861 3243
rect 880 3223 938 3243
rect 957 3240 4239 3243
rect 957 3223 3399 3240
rect 173 3220 3399 3223
rect 3418 3220 3476 3240
rect 3495 3220 4239 3240
rect 173 3205 4239 3220
rect 175 3017 282 3205
rect 2770 3203 4239 3205
rect 643 3166 764 3176
rect 643 3164 712 3166
rect 643 3123 656 3164
rect 693 3125 712 3164
rect 749 3125 764 3166
rect 693 3123 764 3125
rect 643 3105 764 3123
rect 175 3013 283 3017
rect 649 3013 726 3105
rect 1699 3101 1775 3117
rect 1699 3078 1714 3101
rect 176 2420 283 3013
rect 651 2962 726 3013
rect 1692 3064 1714 3078
rect 1758 3064 1775 3101
rect 1692 3044 1775 3064
rect 1692 2978 1709 3044
rect 1763 2978 1775 3044
rect 651 2919 727 2962
rect 655 2608 727 2919
rect 1692 2954 1775 2978
rect 1692 2934 1768 2954
rect 1692 2915 1771 2934
rect 1351 2899 1423 2900
rect 1350 2891 1449 2899
rect 1350 2888 1402 2891
rect 1350 2853 1358 2888
rect 1383 2853 1402 2888
rect 1427 2853 1449 2891
rect 1350 2841 1449 2853
rect 1351 2822 1419 2841
rect 1352 2819 1385 2822
rect 1587 2819 1619 2820
rect 762 2758 965 2771
rect 762 2725 786 2758
rect 822 2757 965 2758
rect 822 2754 933 2757
rect 822 2727 859 2754
rect 888 2730 933 2754
rect 962 2730 965 2757
rect 888 2727 965 2730
rect 822 2725 965 2727
rect 762 2712 965 2725
rect 762 2711 863 2712
rect 655 2566 664 2608
rect 713 2566 727 2608
rect 655 2545 727 2566
rect 655 2503 665 2545
rect 714 2503 727 2545
rect 655 2485 727 2503
rect 1140 2649 1172 2656
rect 1140 2629 1147 2649
rect 1168 2629 1172 2649
rect 1140 2564 1172 2629
rect 1352 2620 1383 2819
rect 1584 2814 1619 2819
rect 1584 2794 1591 2814
rect 1611 2794 1619 2814
rect 1584 2786 1619 2794
rect 1352 2590 1358 2620
rect 1379 2590 1383 2620
rect 1352 2582 1383 2590
rect 1510 2564 1550 2565
rect 1140 2562 1552 2564
rect 1140 2536 1520 2562
rect 1546 2536 1552 2562
rect 1140 2528 1552 2536
rect 1140 2500 1172 2528
rect 1585 2508 1619 2786
rect 1701 2599 1771 2915
rect 3689 2900 3720 2901
rect 3689 2892 3734 2900
rect 2769 2869 2933 2876
rect 3689 2869 3699 2892
rect 2395 2854 3699 2869
rect 3724 2854 3734 2892
rect 4953 2895 4987 4135
rect 4953 2891 5183 2895
rect 4953 2865 5152 2891
rect 5177 2865 5183 2891
rect 4953 2857 5183 2865
rect 2395 2836 3734 2854
rect 2400 2823 2436 2836
rect 2769 2833 2933 2836
rect 1810 2754 2013 2767
rect 1810 2721 1834 2754
rect 1870 2753 2013 2754
rect 1870 2750 1981 2753
rect 1870 2723 1907 2750
rect 1936 2726 1981 2750
rect 2010 2726 2013 2753
rect 1936 2723 2013 2726
rect 1870 2721 2013 2723
rect 1810 2708 2013 2721
rect 1810 2707 1911 2708
rect 1140 2480 1145 2500
rect 1166 2480 1172 2500
rect 1140 2473 1172 2480
rect 1563 2503 1619 2508
rect 1563 2483 1570 2503
rect 1590 2483 1619 2503
rect 1696 2593 1771 2599
rect 1696 2560 1704 2593
rect 1757 2560 1771 2593
rect 1696 2535 1771 2560
rect 1696 2502 1709 2535
rect 1762 2502 1771 2535
rect 1696 2493 1771 2502
rect 2188 2645 2220 2652
rect 2188 2625 2195 2645
rect 2216 2625 2220 2645
rect 2188 2560 2220 2625
rect 2400 2616 2431 2823
rect 2635 2815 2667 2816
rect 2632 2810 2667 2815
rect 2632 2790 2639 2810
rect 2659 2790 2667 2810
rect 2632 2782 2667 2790
rect 2400 2586 2406 2616
rect 2427 2586 2431 2616
rect 2400 2578 2431 2586
rect 2558 2560 2598 2561
rect 2188 2558 2600 2560
rect 2188 2532 2568 2558
rect 2594 2532 2600 2558
rect 2188 2524 2600 2532
rect 2188 2496 2220 2524
rect 2633 2504 2667 2782
rect 4712 2760 4915 2773
rect 4712 2727 4736 2760
rect 4772 2759 4915 2760
rect 4772 2756 4883 2759
rect 4772 2729 4809 2756
rect 4838 2732 4883 2756
rect 4912 2732 4915 2759
rect 4838 2729 4915 2732
rect 4772 2727 4915 2729
rect 4712 2714 4915 2727
rect 4712 2713 4813 2714
rect 1696 2488 1754 2493
rect 1563 2476 1619 2483
rect 2188 2476 2193 2496
rect 2214 2476 2220 2496
rect 1563 2475 1598 2476
rect 2188 2469 2220 2476
rect 2611 2499 2667 2504
rect 2611 2479 2618 2499
rect 2638 2479 2667 2499
rect 2611 2472 2667 2479
rect 5090 2651 5122 2658
rect 5090 2631 5097 2651
rect 5118 2631 5122 2651
rect 5090 2566 5122 2631
rect 5302 2622 5333 2848
rect 5537 2821 5569 2822
rect 5534 2816 5569 2821
rect 5534 2796 5541 2816
rect 5561 2796 5569 2816
rect 5534 2788 5569 2796
rect 5302 2592 5308 2622
rect 5329 2592 5333 2622
rect 5302 2584 5333 2592
rect 5460 2566 5500 2567
rect 5090 2564 5502 2566
rect 5090 2538 5470 2564
rect 5496 2538 5502 2564
rect 5090 2530 5502 2538
rect 5090 2502 5122 2530
rect 5090 2482 5095 2502
rect 5116 2482 5122 2502
rect 5090 2475 5122 2482
rect 5292 2504 5340 2511
rect 5535 2510 5569 2788
rect 5292 2484 5299 2504
rect 5332 2484 5340 2504
rect 2611 2471 2646 2472
rect 854 2420 965 2424
rect 2637 2420 4207 2421
rect 176 2416 4207 2420
rect 4532 2416 4950 2429
rect 176 2404 4950 2416
rect 176 2402 4812 2404
rect 176 2382 862 2402
rect 881 2382 939 2402
rect 958 2398 4812 2402
rect 958 2382 1910 2398
rect 176 2378 1910 2382
rect 1929 2378 1987 2398
rect 2006 2384 4812 2398
rect 4831 2384 4889 2404
rect 4908 2384 4950 2404
rect 2006 2378 4950 2384
rect 176 2364 4950 2378
rect 176 1741 283 2364
rect 1902 2361 2013 2364
rect 4532 2358 4950 2364
rect 662 2315 726 2319
rect 658 2309 726 2315
rect 658 2276 675 2309
rect 715 2276 726 2309
rect 658 2264 726 2276
rect 1709 2278 1774 2300
rect 658 2262 715 2264
rect 662 1901 713 2262
rect 1709 2239 1726 2278
rect 1771 2239 1774 2278
rect 1350 2194 1385 2196
rect 1350 2185 1454 2194
rect 1350 2184 1401 2185
rect 1350 2164 1353 2184
rect 1378 2165 1401 2184
rect 1433 2165 1454 2185
rect 1378 2164 1454 2165
rect 1350 2157 1454 2164
rect 1350 2145 1385 2157
rect 762 2079 965 2092
rect 762 2046 786 2079
rect 822 2078 965 2079
rect 822 2075 933 2078
rect 822 2048 859 2075
rect 888 2051 933 2075
rect 962 2051 965 2078
rect 888 2048 965 2051
rect 822 2046 965 2048
rect 762 2033 965 2046
rect 762 2032 863 2033
rect 1140 1970 1172 1977
rect 1140 1950 1147 1970
rect 1168 1950 1172 1970
rect 651 1892 716 1901
rect 651 1855 661 1892
rect 701 1858 716 1892
rect 1140 1885 1172 1950
rect 1352 1941 1383 2145
rect 1587 2140 1619 2141
rect 1584 2135 1619 2140
rect 1584 2115 1591 2135
rect 1611 2115 1619 2135
rect 1584 2107 1619 2115
rect 1352 1911 1358 1941
rect 1379 1911 1383 1941
rect 1352 1903 1383 1911
rect 1510 1885 1550 1886
rect 1140 1883 1552 1885
rect 701 1855 718 1858
rect 651 1836 718 1855
rect 651 1815 665 1836
rect 701 1815 718 1836
rect 651 1808 718 1815
rect 1140 1857 1520 1883
rect 1546 1857 1552 1883
rect 1140 1849 1552 1857
rect 1140 1821 1172 1849
rect 1585 1829 1619 2107
rect 1709 1939 1774 2239
rect 3846 2200 3883 2221
rect 3846 2163 3857 2200
rect 3874 2176 3883 2200
rect 3874 2163 3884 2176
rect 3846 2153 3884 2163
rect 3847 2149 3884 2153
rect 3847 2143 3880 2149
rect 3257 2074 3460 2087
rect 3257 2041 3281 2074
rect 3317 2073 3460 2074
rect 3317 2070 3428 2073
rect 3317 2043 3354 2070
rect 3383 2046 3428 2070
rect 3457 2046 3460 2073
rect 3383 2043 3460 2046
rect 3317 2041 3460 2043
rect 3257 2028 3460 2041
rect 3257 2027 3358 2028
rect 3635 1965 3667 1972
rect 3635 1945 3642 1965
rect 3663 1945 3667 1965
rect 1140 1801 1145 1821
rect 1166 1801 1172 1821
rect 1140 1794 1172 1801
rect 1563 1824 1619 1829
rect 1563 1804 1570 1824
rect 1590 1804 1619 1824
rect 1563 1797 1619 1804
rect 1699 1928 1779 1939
rect 1699 1902 1716 1928
rect 1756 1902 1779 1928
rect 1699 1875 1779 1902
rect 1699 1849 1720 1875
rect 1760 1849 1779 1875
rect 1699 1830 1779 1849
rect 1699 1804 1723 1830
rect 1763 1804 1779 1830
rect 2773 1874 2878 1895
rect 3635 1880 3667 1945
rect 3847 1936 3878 2143
rect 4082 2135 4114 2136
rect 4079 2130 4114 2135
rect 4079 2110 4086 2130
rect 4106 2110 4114 2130
rect 4079 2102 4114 2110
rect 3847 1906 3853 1936
rect 3874 1906 3878 1936
rect 3847 1898 3878 1906
rect 4005 1880 4045 1881
rect 3635 1878 4047 1880
rect 2773 1868 3249 1874
rect 2773 1866 2830 1868
rect 2773 1835 2785 1866
rect 2810 1845 2830 1866
rect 2856 1861 3249 1868
rect 2856 1845 3210 1861
rect 2810 1838 3210 1845
rect 3236 1838 3249 1861
rect 2810 1835 3249 1838
rect 2773 1825 3249 1835
rect 3635 1852 4015 1878
rect 4041 1852 4047 1878
rect 3635 1844 4047 1852
rect 2773 1823 2878 1825
rect 1563 1796 1598 1797
rect 1699 1792 1779 1804
rect 3635 1816 3667 1844
rect 4080 1824 4114 2102
rect 3635 1796 3640 1816
rect 3661 1796 3667 1816
rect 3635 1789 3667 1796
rect 4058 1819 4114 1824
rect 4058 1799 4065 1819
rect 4085 1799 4114 1819
rect 4058 1792 4114 1799
rect 4058 1791 4093 1792
rect 854 1741 965 1745
rect 2596 1741 4249 1744
rect 174 1723 4249 1741
rect 174 1703 862 1723
rect 881 1703 939 1723
rect 958 1718 4249 1723
rect 958 1703 3357 1718
rect 174 1698 3357 1703
rect 3376 1698 3434 1718
rect 3453 1698 4249 1718
rect 174 1688 4249 1698
rect 174 1685 799 1688
rect 986 1685 4249 1688
rect 176 1457 283 1685
rect 2596 1684 4249 1685
rect 3349 1681 3460 1684
rect 644 1646 765 1656
rect 644 1644 713 1646
rect 644 1603 657 1644
rect 694 1605 713 1644
rect 750 1605 765 1646
rect 694 1603 765 1605
rect 644 1585 765 1603
rect 650 1483 729 1585
rect 1702 1545 1769 1564
rect 1702 1525 1722 1545
rect 176 1402 284 1457
rect 651 1402 729 1483
rect 1701 1479 1722 1525
rect 1752 1525 1769 1545
rect 1752 1495 1771 1525
rect 1752 1479 1772 1495
rect 1701 1463 1772 1479
rect 1351 1452 1423 1453
rect 1350 1444 1449 1452
rect 1350 1441 1402 1444
rect 1350 1406 1358 1441
rect 1383 1406 1402 1441
rect 1427 1406 1449 1444
rect 176 973 283 1402
rect 655 1161 727 1402
rect 1350 1394 1449 1406
rect 1351 1375 1419 1394
rect 1352 1372 1385 1375
rect 1587 1372 1619 1373
rect 762 1311 965 1324
rect 762 1278 786 1311
rect 822 1310 965 1311
rect 822 1307 933 1310
rect 822 1280 859 1307
rect 888 1283 933 1307
rect 962 1283 965 1310
rect 888 1280 965 1283
rect 822 1278 965 1280
rect 762 1265 965 1278
rect 762 1264 863 1265
rect 655 1119 664 1161
rect 713 1119 727 1161
rect 655 1098 727 1119
rect 655 1056 665 1098
rect 714 1056 727 1098
rect 655 1038 727 1056
rect 1140 1202 1172 1209
rect 1140 1182 1147 1202
rect 1168 1182 1172 1202
rect 1140 1117 1172 1182
rect 1352 1173 1383 1372
rect 1584 1367 1619 1372
rect 1584 1347 1591 1367
rect 1611 1347 1619 1367
rect 1584 1339 1619 1347
rect 1352 1143 1358 1173
rect 1379 1143 1383 1173
rect 1352 1135 1383 1143
rect 1510 1117 1550 1118
rect 1140 1115 1552 1117
rect 1140 1089 1520 1115
rect 1546 1089 1552 1115
rect 1140 1081 1552 1089
rect 1140 1053 1172 1081
rect 1585 1061 1619 1339
rect 1701 1152 1771 1463
rect 2398 1454 3740 1459
rect 2398 1452 3697 1454
rect 2395 1426 3697 1452
rect 3725 1426 3740 1454
rect 2395 1418 3740 1426
rect 2395 1393 2434 1418
rect 2395 1376 2436 1393
rect 2395 1369 2434 1376
rect 1810 1307 2013 1320
rect 1810 1274 1834 1307
rect 1870 1306 2013 1307
rect 1870 1303 1981 1306
rect 1870 1276 1907 1303
rect 1936 1279 1981 1303
rect 2010 1279 2013 1306
rect 1936 1276 2013 1279
rect 1870 1274 2013 1276
rect 1810 1261 2013 1274
rect 1810 1260 1911 1261
rect 1140 1033 1145 1053
rect 1166 1033 1172 1053
rect 1140 1026 1172 1033
rect 1563 1056 1619 1061
rect 1563 1036 1570 1056
rect 1590 1036 1619 1056
rect 1696 1146 1771 1152
rect 1696 1113 1704 1146
rect 1757 1113 1771 1146
rect 1696 1088 1771 1113
rect 1696 1055 1709 1088
rect 1762 1055 1771 1088
rect 1696 1046 1771 1055
rect 2188 1198 2220 1205
rect 2188 1178 2195 1198
rect 2216 1178 2220 1198
rect 2188 1113 2220 1178
rect 2400 1169 2431 1369
rect 2635 1368 2667 1369
rect 2632 1363 2667 1368
rect 2632 1343 2639 1363
rect 2659 1343 2667 1363
rect 2632 1335 2667 1343
rect 2400 1139 2406 1169
rect 2427 1139 2431 1169
rect 2400 1131 2431 1139
rect 2558 1113 2598 1114
rect 2188 1111 2600 1113
rect 2188 1085 2568 1111
rect 2594 1085 2600 1111
rect 2188 1077 2600 1085
rect 2188 1049 2220 1077
rect 2633 1057 2667 1335
rect 1696 1041 1754 1046
rect 1563 1029 1619 1036
rect 2188 1029 2193 1049
rect 2214 1029 2220 1049
rect 1563 1028 1598 1029
rect 2188 1022 2220 1029
rect 2611 1052 2667 1057
rect 2611 1032 2618 1052
rect 2638 1032 2667 1052
rect 2611 1025 2667 1032
rect 2611 1024 2646 1025
rect 854 973 965 977
rect 2729 973 4249 974
rect 176 955 4249 973
rect 176 935 862 955
rect 881 935 939 955
rect 958 951 4249 955
rect 958 935 1910 951
rect 176 931 1910 935
rect 1929 931 1987 951
rect 2006 931 4249 951
rect 176 917 4249 931
rect 176 294 283 917
rect 1902 914 2013 917
rect 662 868 726 872
rect 658 862 726 868
rect 658 829 675 862
rect 715 829 726 862
rect 658 817 726 829
rect 1709 831 1774 853
rect 658 815 715 817
rect 662 454 713 815
rect 1709 792 1726 831
rect 1771 792 1774 831
rect 1350 747 1385 749
rect 1350 738 1454 747
rect 1350 737 1401 738
rect 1350 717 1353 737
rect 1378 718 1401 737
rect 1433 718 1454 738
rect 1378 717 1454 718
rect 1350 710 1454 717
rect 1350 698 1385 710
rect 762 632 965 645
rect 762 599 786 632
rect 822 631 965 632
rect 822 628 933 631
rect 822 601 859 628
rect 888 604 933 628
rect 962 604 965 631
rect 888 601 965 604
rect 822 599 965 601
rect 762 586 965 599
rect 762 585 863 586
rect 1140 523 1172 530
rect 1140 503 1147 523
rect 1168 503 1172 523
rect 651 445 716 454
rect 651 408 661 445
rect 701 411 716 445
rect 1140 438 1172 503
rect 1352 494 1383 698
rect 1587 693 1619 694
rect 1584 688 1619 693
rect 1584 668 1591 688
rect 1611 668 1619 688
rect 1584 660 1619 668
rect 1352 464 1358 494
rect 1379 464 1383 494
rect 1352 456 1383 464
rect 1510 438 1550 439
rect 1140 436 1552 438
rect 701 408 718 411
rect 651 389 718 408
rect 651 368 665 389
rect 701 368 718 389
rect 651 361 718 368
rect 1140 410 1520 436
rect 1546 410 1552 436
rect 1140 402 1552 410
rect 1140 374 1172 402
rect 1585 382 1619 660
rect 1709 529 1774 792
rect 1709 525 1770 529
rect 1140 354 1145 374
rect 1166 354 1172 374
rect 1140 347 1172 354
rect 1563 377 1619 382
rect 1563 357 1570 377
rect 1590 357 1619 377
rect 1563 350 1619 357
rect 1563 349 1598 350
rect 854 294 965 298
rect 174 276 1493 294
rect 174 256 862 276
rect 881 256 939 276
rect 958 256 1493 276
rect 174 238 1493 256
rect 176 118 283 238
rect 644 199 765 209
rect 644 197 713 199
rect 644 156 657 197
rect 694 158 713 197
rect 750 158 765 199
rect 694 156 765 158
rect 644 138 765 156
rect -25 45 109 74
rect -25 -67 13 45
rect 92 -67 109 45
rect 176 38 284 118
rect -25 -1020 109 -67
rect 177 -774 284 38
rect 650 66 715 138
rect 650 0 718 66
rect 651 -546 718 0
rect 1705 -362 1770 525
rect 2748 255 2885 259
rect 2735 251 2892 255
rect 2735 144 2772 251
rect 2872 144 2892 251
rect 2735 102 2892 144
rect 2748 -146 2885 102
rect 2738 -188 2904 -146
rect 2738 -263 2767 -188
rect 2884 -263 2904 -188
rect 2738 -279 2904 -263
rect 1694 -383 1831 -362
rect 1694 -458 1719 -383
rect 1789 -458 1831 -383
rect 1694 -489 1831 -458
rect 637 -595 812 -546
rect 637 -674 670 -595
rect 770 -674 812 -595
rect 637 -679 812 -674
rect 177 -816 325 -774
rect 177 -824 217 -816
rect 179 -903 217 -824
rect 287 -903 325 -816
rect 179 -941 325 -903
rect -29 -1056 110 -1020
rect -29 -1151 -15 -1056
rect 75 -1151 110 -1056
rect -29 -1169 110 -1151
rect 5292 -1276 5340 2484
rect 5513 2505 5569 2510
rect 5513 2485 5520 2505
rect 5540 2485 5569 2505
rect 5513 2478 5569 2485
rect 5513 2477 5548 2478
rect 5617 2387 5645 5195
rect 8830 5150 8895 5450
rect 8985 5282 9019 5560
rect 9432 5540 9464 5568
rect 9052 5532 9464 5540
rect 9052 5506 9058 5532
rect 9084 5506 9464 5532
rect 9886 5574 9953 5581
rect 9886 5553 9903 5574
rect 9939 5553 9953 5574
rect 9886 5534 9953 5553
rect 9886 5531 9903 5534
rect 9052 5504 9464 5506
rect 9054 5503 9094 5504
rect 9221 5478 9252 5486
rect 9221 5448 9225 5478
rect 9246 5448 9252 5478
rect 8985 5274 9020 5282
rect 8985 5254 8993 5274
rect 9013 5254 9020 5274
rect 8985 5249 9020 5254
rect 8985 5248 9017 5249
rect 9221 5244 9252 5448
rect 9432 5439 9464 5504
rect 9888 5497 9903 5531
rect 9943 5497 9953 5534
rect 9888 5488 9953 5497
rect 9432 5419 9436 5439
rect 9457 5419 9464 5439
rect 9432 5412 9464 5419
rect 9741 5356 9842 5357
rect 9639 5343 9842 5356
rect 9639 5341 9782 5343
rect 9639 5338 9716 5341
rect 9639 5311 9642 5338
rect 9671 5314 9716 5338
rect 9745 5314 9782 5341
rect 9671 5311 9782 5314
rect 9639 5310 9782 5311
rect 9818 5310 9842 5343
rect 9639 5297 9842 5310
rect 9219 5232 9254 5244
rect 9150 5225 9254 5232
rect 9150 5224 9226 5225
rect 9150 5204 9171 5224
rect 9203 5205 9226 5224
rect 9251 5205 9254 5225
rect 9203 5204 9254 5205
rect 9150 5195 9254 5204
rect 9219 5193 9254 5195
rect 8830 5111 8833 5150
rect 8878 5111 8895 5150
rect 9891 5127 9942 5488
rect 9889 5125 9946 5127
rect 8830 5089 8895 5111
rect 9878 5113 9946 5125
rect 9878 5080 9889 5113
rect 9929 5080 9946 5113
rect 9878 5074 9946 5080
rect 9878 5070 9942 5074
rect 8591 5025 8702 5028
rect 10321 5025 10428 5648
rect 6885 5011 10428 5025
rect 6885 4991 8598 5011
rect 8617 4991 8675 5011
rect 8694 5007 10428 5011
rect 8694 4991 9646 5007
rect 6885 4987 9646 4991
rect 9665 4987 9723 5007
rect 9742 4987 10428 5007
rect 6885 4969 10428 4987
rect 6885 4968 7875 4969
rect 9639 4965 9750 4969
rect 7958 4917 7993 4918
rect 7937 4910 7993 4917
rect 7937 4890 7966 4910
rect 7986 4890 7993 4910
rect 7937 4885 7993 4890
rect 8384 4913 8416 4920
rect 9006 4913 9041 4914
rect 8384 4893 8390 4913
rect 8411 4893 8416 4913
rect 8985 4906 9041 4913
rect 8850 4896 8908 4901
rect 7937 4607 7971 4885
rect 8384 4865 8416 4893
rect 8004 4857 8416 4865
rect 8004 4831 8010 4857
rect 8036 4831 8416 4857
rect 8004 4829 8416 4831
rect 8006 4828 8046 4829
rect 8173 4803 8204 4811
rect 8173 4773 8177 4803
rect 8198 4773 8204 4803
rect 7937 4599 7972 4607
rect 7937 4579 7945 4599
rect 7965 4579 7972 4599
rect 7937 4574 7972 4579
rect 7937 4573 7969 4574
rect 8173 4573 8204 4773
rect 8384 4764 8416 4829
rect 8384 4744 8388 4764
rect 8409 4744 8416 4764
rect 8384 4737 8416 4744
rect 8833 4887 8908 4896
rect 8833 4854 8842 4887
rect 8895 4854 8908 4887
rect 8833 4829 8908 4854
rect 8833 4796 8847 4829
rect 8900 4796 8908 4829
rect 8833 4790 8908 4796
rect 8985 4886 9014 4906
rect 9034 4886 9041 4906
rect 8985 4881 9041 4886
rect 9432 4909 9464 4916
rect 9432 4889 9438 4909
rect 9459 4889 9464 4909
rect 8693 4681 8794 4682
rect 8591 4668 8794 4681
rect 8591 4666 8734 4668
rect 8591 4663 8668 4666
rect 8591 4636 8594 4663
rect 8623 4639 8668 4663
rect 8697 4639 8734 4666
rect 8623 4636 8734 4639
rect 8591 4635 8734 4636
rect 8770 4635 8794 4668
rect 8591 4622 8794 4635
rect 8170 4566 8209 4573
rect 8168 4549 8209 4566
rect 8170 4524 8209 4549
rect 6864 4516 8209 4524
rect 6864 4488 6879 4516
rect 6907 4490 8209 4516
rect 6907 4488 8206 4490
rect 6864 4483 8206 4488
rect 8833 4479 8903 4790
rect 8985 4603 9019 4881
rect 9432 4861 9464 4889
rect 9052 4853 9464 4861
rect 9052 4827 9058 4853
rect 9084 4827 9464 4853
rect 9052 4825 9464 4827
rect 9054 4824 9094 4825
rect 9221 4799 9252 4807
rect 9221 4769 9225 4799
rect 9246 4769 9252 4799
rect 8985 4595 9020 4603
rect 8985 4575 8993 4595
rect 9013 4575 9020 4595
rect 8985 4570 9020 4575
rect 9221 4570 9252 4769
rect 9432 4760 9464 4825
rect 9432 4740 9436 4760
rect 9457 4740 9464 4760
rect 9432 4733 9464 4740
rect 9877 4886 9949 4904
rect 9877 4844 9890 4886
rect 9939 4844 9949 4886
rect 9877 4823 9949 4844
rect 9877 4781 9891 4823
rect 9940 4781 9949 4823
rect 9741 4677 9842 4678
rect 9639 4664 9842 4677
rect 9639 4662 9782 4664
rect 9639 4659 9716 4662
rect 9639 4632 9642 4659
rect 9671 4635 9716 4659
rect 9745 4635 9782 4662
rect 9671 4632 9782 4635
rect 9639 4631 9782 4632
rect 9818 4631 9842 4664
rect 9639 4618 9842 4631
rect 8985 4569 9017 4570
rect 9219 4567 9252 4570
rect 9185 4548 9253 4567
rect 9155 4536 9254 4548
rect 9877 4540 9949 4781
rect 10321 4540 10428 4969
rect 9155 4498 9177 4536
rect 9202 4501 9221 4536
rect 9246 4501 9254 4536
rect 9202 4498 9254 4501
rect 9155 4490 9254 4498
rect 9181 4489 9253 4490
rect 8832 4463 8903 4479
rect 8832 4447 8852 4463
rect 8833 4417 8852 4447
rect 8835 4397 8852 4417
rect 8882 4417 8903 4463
rect 9875 4459 9953 4540
rect 10320 4485 10428 4540
rect 8882 4397 8902 4417
rect 8835 4378 8902 4397
rect 9875 4357 9954 4459
rect 9839 4339 9960 4357
rect 9839 4337 9910 4339
rect 9839 4296 9854 4337
rect 9891 4298 9910 4337
rect 9947 4298 9960 4339
rect 9891 4296 9960 4298
rect 9839 4286 9960 4296
rect 7144 4258 7255 4261
rect 6458 4257 8008 4258
rect 10321 4257 10428 4485
rect 6458 4254 9618 4257
rect 9805 4254 10430 4257
rect 6458 4244 10430 4254
rect 6458 4224 7151 4244
rect 7170 4224 7228 4244
rect 7247 4239 10430 4244
rect 7247 4224 9646 4239
rect 6458 4219 9646 4224
rect 9665 4219 9723 4239
rect 9742 4219 10430 4239
rect 6458 4201 10430 4219
rect 6458 4198 8008 4201
rect 9639 4197 9750 4201
rect 6511 4150 6546 4151
rect 6490 4143 6546 4150
rect 6490 4123 6519 4143
rect 6539 4123 6546 4143
rect 6490 4118 6546 4123
rect 6937 4146 6969 4153
rect 6937 4126 6943 4146
rect 6964 4126 6969 4146
rect 6490 3840 6524 4118
rect 6937 4098 6969 4126
rect 8825 4138 8905 4150
rect 9006 4145 9041 4146
rect 6557 4090 6969 4098
rect 6557 4064 6563 4090
rect 6589 4064 6969 4090
rect 7355 4104 7792 4117
rect 7355 4081 7368 4104
rect 7394 4097 7792 4104
rect 7394 4081 7748 4097
rect 7355 4074 7748 4081
rect 7774 4074 7792 4097
rect 7355 4068 7792 4074
rect 8825 4112 8841 4138
rect 8881 4112 8905 4138
rect 8825 4093 8905 4112
rect 6557 4062 6969 4064
rect 6559 4061 6599 4062
rect 6726 4036 6757 4044
rect 6726 4006 6730 4036
rect 6751 4006 6757 4036
rect 6490 3832 6525 3840
rect 6490 3812 6498 3832
rect 6518 3812 6525 3832
rect 6490 3807 6525 3812
rect 6490 3806 6522 3807
rect 6726 3799 6757 4006
rect 6937 3997 6969 4062
rect 8825 4067 8844 4093
rect 8884 4067 8905 4093
rect 8825 4040 8905 4067
rect 8825 4014 8848 4040
rect 8888 4014 8905 4040
rect 8825 4003 8905 4014
rect 8985 4138 9041 4145
rect 8985 4118 9014 4138
rect 9034 4118 9041 4138
rect 8985 4113 9041 4118
rect 9432 4141 9464 4148
rect 9432 4121 9438 4141
rect 9459 4121 9464 4141
rect 6937 3977 6941 3997
rect 6962 3977 6969 3997
rect 6937 3970 6969 3977
rect 7246 3914 7347 3915
rect 7144 3901 7347 3914
rect 7144 3899 7287 3901
rect 7144 3896 7221 3899
rect 7144 3869 7147 3896
rect 7176 3872 7221 3896
rect 7250 3872 7287 3899
rect 7176 3869 7287 3872
rect 7144 3868 7287 3869
rect 7323 3868 7347 3901
rect 7144 3855 7347 3868
rect 6724 3793 6757 3799
rect 6720 3789 6757 3793
rect 6720 3779 6758 3789
rect 6720 3766 6730 3779
rect 6721 3742 6730 3766
rect 6747 3742 6758 3779
rect 6721 3721 6758 3742
rect 8830 3703 8895 4003
rect 8985 3835 9019 4113
rect 9432 4093 9464 4121
rect 9052 4085 9464 4093
rect 9052 4059 9058 4085
rect 9084 4059 9464 4085
rect 9886 4127 9953 4134
rect 9886 4106 9903 4127
rect 9939 4106 9953 4127
rect 9886 4087 9953 4106
rect 9886 4084 9903 4087
rect 9052 4057 9464 4059
rect 9054 4056 9094 4057
rect 9221 4031 9252 4039
rect 9221 4001 9225 4031
rect 9246 4001 9252 4031
rect 8985 3827 9020 3835
rect 8985 3807 8993 3827
rect 9013 3807 9020 3827
rect 8985 3802 9020 3807
rect 8985 3801 9017 3802
rect 9221 3797 9252 4001
rect 9432 3992 9464 4057
rect 9888 4050 9903 4084
rect 9943 4050 9953 4087
rect 9888 4041 9953 4050
rect 9432 3972 9436 3992
rect 9457 3972 9464 3992
rect 9432 3965 9464 3972
rect 9741 3909 9842 3910
rect 9639 3896 9842 3909
rect 9639 3894 9782 3896
rect 9639 3891 9716 3894
rect 9639 3864 9642 3891
rect 9671 3867 9716 3891
rect 9745 3867 9782 3894
rect 9671 3864 9782 3867
rect 9639 3863 9782 3864
rect 9818 3863 9842 3896
rect 9639 3850 9842 3863
rect 9219 3785 9254 3797
rect 9150 3778 9254 3785
rect 9150 3777 9226 3778
rect 9150 3757 9171 3777
rect 9203 3758 9226 3777
rect 9251 3758 9254 3778
rect 9203 3757 9254 3758
rect 9150 3748 9254 3757
rect 9219 3746 9254 3748
rect 8830 3664 8833 3703
rect 8878 3664 8895 3703
rect 9891 3680 9942 4041
rect 9889 3678 9946 3680
rect 8830 3642 8895 3664
rect 9878 3666 9946 3678
rect 9878 3633 9889 3666
rect 9929 3633 9946 3666
rect 9878 3627 9946 3633
rect 9878 3623 9942 3627
rect 8591 3578 8702 3581
rect 10321 3578 10428 4201
rect 6667 3564 10428 3578
rect 6667 3544 8598 3564
rect 8617 3544 8675 3564
rect 8694 3560 10428 3564
rect 8694 3544 9646 3560
rect 6667 3540 9646 3544
rect 9665 3540 9723 3560
rect 9742 3540 10428 3560
rect 6667 3522 10428 3540
rect 6667 3521 7967 3522
rect 9639 3518 9750 3522
rect 7958 3470 7993 3471
rect 7937 3463 7993 3470
rect 7937 3443 7966 3463
rect 7986 3443 7993 3463
rect 7937 3438 7993 3443
rect 8384 3466 8416 3473
rect 9006 3466 9041 3467
rect 8384 3446 8390 3466
rect 8411 3446 8416 3466
rect 8985 3459 9041 3466
rect 8850 3449 8908 3454
rect 7937 3160 7971 3438
rect 8384 3418 8416 3446
rect 8004 3410 8416 3418
rect 8004 3384 8010 3410
rect 8036 3384 8416 3410
rect 8004 3382 8416 3384
rect 8006 3381 8046 3382
rect 8173 3356 8204 3364
rect 8173 3326 8177 3356
rect 8198 3326 8204 3356
rect 7937 3152 7972 3160
rect 7937 3132 7945 3152
rect 7965 3132 7972 3152
rect 7937 3127 7972 3132
rect 7937 3126 7969 3127
rect 8173 3119 8204 3326
rect 8384 3317 8416 3382
rect 8384 3297 8388 3317
rect 8409 3297 8416 3317
rect 8384 3290 8416 3297
rect 8833 3440 8908 3449
rect 8833 3407 8842 3440
rect 8895 3407 8908 3440
rect 8833 3382 8908 3407
rect 8833 3349 8847 3382
rect 8900 3349 8908 3382
rect 8833 3343 8908 3349
rect 8985 3439 9014 3459
rect 9034 3439 9041 3459
rect 8985 3434 9041 3439
rect 9432 3462 9464 3469
rect 9432 3442 9438 3462
rect 9459 3442 9464 3462
rect 8693 3234 8794 3235
rect 8591 3221 8794 3234
rect 8591 3219 8734 3221
rect 8591 3216 8668 3219
rect 8591 3189 8594 3216
rect 8623 3192 8668 3216
rect 8697 3192 8734 3219
rect 8623 3189 8734 3192
rect 8591 3188 8734 3189
rect 8770 3188 8794 3221
rect 8591 3175 8794 3188
rect 7671 3106 7835 3109
rect 8168 3106 8204 3119
rect 6870 3088 8209 3106
rect 6870 3050 6880 3088
rect 6905 3073 8209 3088
rect 6905 3050 6915 3073
rect 7671 3066 7835 3073
rect 6870 3042 6915 3050
rect 6884 3041 6915 3042
rect 8833 3027 8903 3343
rect 8985 3156 9019 3434
rect 9432 3414 9464 3442
rect 9052 3406 9464 3414
rect 9052 3380 9058 3406
rect 9084 3380 9464 3406
rect 9052 3378 9464 3380
rect 9054 3377 9094 3378
rect 9221 3352 9252 3360
rect 9221 3322 9225 3352
rect 9246 3322 9252 3352
rect 8985 3148 9020 3156
rect 8985 3128 8993 3148
rect 9013 3128 9020 3148
rect 8985 3123 9020 3128
rect 9221 3123 9252 3322
rect 9432 3313 9464 3378
rect 9432 3293 9436 3313
rect 9457 3293 9464 3313
rect 9432 3286 9464 3293
rect 9877 3439 9949 3457
rect 9877 3397 9890 3439
rect 9939 3397 9949 3439
rect 9877 3376 9949 3397
rect 9877 3334 9891 3376
rect 9940 3334 9949 3376
rect 9741 3230 9842 3231
rect 9639 3217 9842 3230
rect 9639 3215 9782 3217
rect 9639 3212 9716 3215
rect 9639 3185 9642 3212
rect 9671 3188 9716 3212
rect 9745 3188 9782 3215
rect 9671 3185 9782 3188
rect 9639 3184 9782 3185
rect 9818 3184 9842 3217
rect 9639 3171 9842 3184
rect 8985 3122 9017 3123
rect 9219 3120 9252 3123
rect 9185 3101 9253 3120
rect 9155 3089 9254 3101
rect 9155 3051 9177 3089
rect 9202 3054 9221 3089
rect 9246 3054 9254 3089
rect 9202 3051 9254 3054
rect 9155 3043 9254 3051
rect 9181 3042 9253 3043
rect 8833 3008 8912 3027
rect 8836 2988 8912 3008
rect 8829 2964 8912 2988
rect 9877 3023 9949 3334
rect 9877 2980 9953 3023
rect 8829 2898 8841 2964
rect 8895 2898 8912 2964
rect 8829 2878 8912 2898
rect 8829 2841 8846 2878
rect 8890 2864 8912 2878
rect 9878 2929 9953 2980
rect 10321 2929 10428 3522
rect 8890 2841 8905 2864
rect 8829 2825 8905 2841
rect 9878 2837 9955 2929
rect 10321 2925 10429 2929
rect 9840 2819 9961 2837
rect 9840 2817 9911 2819
rect 9840 2776 9855 2817
rect 9892 2778 9911 2817
rect 9948 2778 9961 2819
rect 9892 2776 9961 2778
rect 9840 2766 9961 2776
rect 6411 2737 7834 2739
rect 10322 2737 10429 2925
rect 6411 2722 10431 2737
rect 6411 2702 7109 2722
rect 7128 2702 7186 2722
rect 7205 2719 10431 2722
rect 7205 2702 9647 2719
rect 6411 2699 9647 2702
rect 9666 2699 9724 2719
rect 9743 2699 10431 2719
rect 6411 2681 10431 2699
rect 7102 2680 7213 2681
rect 7789 2680 7996 2681
rect 9640 2677 9751 2681
rect 6469 2628 6504 2629
rect 6448 2621 6504 2628
rect 6448 2601 6477 2621
rect 6497 2601 6504 2621
rect 6448 2596 6504 2601
rect 6895 2624 6927 2631
rect 6895 2604 6901 2624
rect 6922 2604 6927 2624
rect 5617 2372 5643 2387
rect 5614 2365 5650 2372
rect 5614 2327 5620 2365
rect 5643 2327 5650 2365
rect 5614 2321 5650 2327
rect 6448 2318 6482 2596
rect 6895 2576 6927 2604
rect 6515 2568 6927 2576
rect 6515 2542 6521 2568
rect 6547 2542 6927 2568
rect 6515 2540 6927 2542
rect 6517 2539 6557 2540
rect 6684 2514 6715 2522
rect 6684 2484 6688 2514
rect 6709 2484 6715 2514
rect 6448 2310 6483 2318
rect 6448 2290 6456 2310
rect 6476 2290 6483 2310
rect 6448 2285 6483 2290
rect 6448 2284 6480 2285
rect 6684 2281 6715 2484
rect 6895 2475 6927 2540
rect 8826 2618 8906 2630
rect 9007 2625 9042 2626
rect 8826 2592 8842 2618
rect 8882 2592 8906 2618
rect 8826 2573 8906 2592
rect 8826 2547 8845 2573
rect 8885 2547 8906 2573
rect 8826 2520 8906 2547
rect 8826 2494 8849 2520
rect 8889 2494 8906 2520
rect 8826 2483 8906 2494
rect 8986 2618 9042 2625
rect 8986 2598 9015 2618
rect 9035 2598 9042 2618
rect 8986 2593 9042 2598
rect 9433 2621 9465 2628
rect 9433 2601 9439 2621
rect 9460 2601 9465 2621
rect 6895 2455 6899 2475
rect 6920 2455 6927 2475
rect 6895 2448 6927 2455
rect 7204 2392 7305 2393
rect 7102 2379 7305 2392
rect 7102 2377 7245 2379
rect 7102 2374 7179 2377
rect 7102 2347 7105 2374
rect 7134 2350 7179 2374
rect 7208 2350 7245 2377
rect 7134 2347 7245 2350
rect 7102 2346 7245 2347
rect 7281 2346 7305 2379
rect 7102 2333 7305 2346
rect 6679 2263 6715 2281
rect 6679 2246 6714 2263
rect 6612 2215 6717 2246
rect 6612 2210 6684 2215
rect 6612 2189 6643 2210
rect 6663 2194 6684 2210
rect 6704 2194 6717 2215
rect 6663 2189 6717 2194
rect 6612 2180 6717 2189
rect 8831 2183 8896 2483
rect 8986 2315 9020 2593
rect 9433 2573 9465 2601
rect 9053 2565 9465 2573
rect 9053 2539 9059 2565
rect 9085 2539 9465 2565
rect 9887 2607 9954 2614
rect 9887 2586 9904 2607
rect 9940 2586 9954 2607
rect 9887 2567 9954 2586
rect 9887 2564 9904 2567
rect 9053 2537 9465 2539
rect 9055 2536 9095 2537
rect 9222 2511 9253 2519
rect 9222 2481 9226 2511
rect 9247 2481 9253 2511
rect 8986 2307 9021 2315
rect 8986 2287 8994 2307
rect 9014 2287 9021 2307
rect 8986 2282 9021 2287
rect 8986 2281 9018 2282
rect 9222 2277 9253 2481
rect 9433 2472 9465 2537
rect 9889 2530 9904 2564
rect 9944 2530 9954 2567
rect 9889 2521 9954 2530
rect 9433 2452 9437 2472
rect 9458 2452 9465 2472
rect 9433 2445 9465 2452
rect 9742 2389 9843 2390
rect 9640 2376 9843 2389
rect 9640 2374 9783 2376
rect 9640 2371 9717 2374
rect 9640 2344 9643 2371
rect 9672 2347 9717 2371
rect 9746 2347 9783 2374
rect 9672 2344 9783 2347
rect 9640 2343 9783 2344
rect 9819 2343 9843 2376
rect 9640 2330 9843 2343
rect 9220 2265 9255 2277
rect 9151 2258 9255 2265
rect 9151 2257 9227 2258
rect 9151 2237 9172 2257
rect 9204 2238 9227 2257
rect 9252 2238 9255 2258
rect 9204 2237 9255 2238
rect 9151 2228 9255 2237
rect 9220 2226 9255 2228
rect 8831 2144 8834 2183
rect 8879 2144 8896 2183
rect 9892 2160 9943 2521
rect 9890 2158 9947 2160
rect 8831 2122 8896 2144
rect 9879 2146 9947 2158
rect 9879 2113 9890 2146
rect 9930 2113 9947 2146
rect 9879 2107 9947 2113
rect 9879 2103 9943 2107
rect 8592 2058 8703 2061
rect 10322 2058 10429 2681
rect 6635 2044 10429 2058
rect 6635 2024 8599 2044
rect 8618 2024 8676 2044
rect 8695 2040 10429 2044
rect 8695 2024 9647 2040
rect 6635 2020 9647 2024
rect 9666 2020 9724 2040
rect 9743 2020 10429 2040
rect 6635 2002 10429 2020
rect 6635 2001 7876 2002
rect 9640 1998 9751 2002
rect 7959 1950 7994 1951
rect 7938 1943 7994 1950
rect 7938 1923 7967 1943
rect 7987 1923 7994 1943
rect 7938 1918 7994 1923
rect 8385 1946 8417 1953
rect 9007 1946 9042 1947
rect 8385 1926 8391 1946
rect 8412 1926 8417 1946
rect 8986 1939 9042 1946
rect 8851 1929 8909 1934
rect 7938 1640 7972 1918
rect 8385 1898 8417 1926
rect 8005 1890 8417 1898
rect 8005 1864 8011 1890
rect 8037 1864 8417 1890
rect 8005 1862 8417 1864
rect 8007 1861 8047 1862
rect 8174 1836 8205 1844
rect 8174 1806 8178 1836
rect 8199 1806 8205 1836
rect 7938 1632 7973 1640
rect 7938 1612 7946 1632
rect 7966 1612 7973 1632
rect 7938 1607 7973 1612
rect 6679 1596 6715 1607
rect 7938 1606 7970 1607
rect 8174 1599 8205 1806
rect 8385 1797 8417 1862
rect 8385 1777 8389 1797
rect 8410 1777 8417 1797
rect 8385 1770 8417 1777
rect 8834 1920 8909 1929
rect 8834 1887 8843 1920
rect 8896 1887 8909 1920
rect 8834 1862 8909 1887
rect 8834 1829 8848 1862
rect 8901 1829 8909 1862
rect 8834 1823 8909 1829
rect 8986 1919 9015 1939
rect 9035 1919 9042 1939
rect 8986 1914 9042 1919
rect 9433 1942 9465 1949
rect 9433 1922 9439 1942
rect 9460 1922 9465 1942
rect 8694 1714 8795 1715
rect 8592 1701 8795 1714
rect 8592 1699 8735 1701
rect 8592 1696 8669 1699
rect 8592 1669 8595 1696
rect 8624 1672 8669 1696
rect 8698 1672 8735 1699
rect 8624 1669 8735 1672
rect 8592 1668 8735 1669
rect 8771 1668 8795 1701
rect 8592 1655 8795 1668
rect 6679 1573 6685 1596
rect 6709 1573 6715 1596
rect 8169 1590 8205 1599
rect 8114 1580 8211 1590
rect 6926 1578 8211 1580
rect 6679 1552 6715 1573
rect 6679 1529 6685 1552
rect 6709 1529 6715 1552
rect 6679 1376 6715 1529
rect 6891 1568 8211 1578
rect 6891 1530 6903 1568
rect 6928 1533 6947 1568
rect 6972 1533 8211 1568
rect 6928 1530 8211 1533
rect 6891 1527 8211 1530
rect 6891 1525 8208 1527
rect 6891 1522 6980 1525
rect 6907 1521 6979 1522
rect 8834 1512 8904 1823
rect 8986 1636 9020 1914
rect 9433 1894 9465 1922
rect 9053 1886 9465 1894
rect 9053 1860 9059 1886
rect 9085 1860 9465 1886
rect 9053 1858 9465 1860
rect 9055 1857 9095 1858
rect 9222 1832 9253 1840
rect 9222 1802 9226 1832
rect 9247 1802 9253 1832
rect 8986 1628 9021 1636
rect 8986 1608 8994 1628
rect 9014 1608 9021 1628
rect 8986 1603 9021 1608
rect 9222 1603 9253 1802
rect 9433 1793 9465 1858
rect 9433 1773 9437 1793
rect 9458 1773 9465 1793
rect 9433 1766 9465 1773
rect 9878 1919 9950 1937
rect 9878 1877 9891 1919
rect 9940 1877 9950 1919
rect 9878 1856 9950 1877
rect 9878 1814 9892 1856
rect 9941 1814 9950 1856
rect 9742 1710 9843 1711
rect 9640 1697 9843 1710
rect 9640 1695 9783 1697
rect 9640 1692 9717 1695
rect 9640 1665 9643 1692
rect 9672 1668 9717 1692
rect 9746 1668 9783 1695
rect 9672 1665 9783 1668
rect 9640 1664 9783 1665
rect 9819 1664 9843 1697
rect 9640 1651 9843 1664
rect 8986 1602 9018 1603
rect 9220 1600 9253 1603
rect 9186 1581 9254 1600
rect 9156 1569 9255 1581
rect 9878 1573 9950 1814
rect 10322 1573 10429 2002
rect 9156 1531 9178 1569
rect 9203 1534 9222 1569
rect 9247 1534 9255 1569
rect 9203 1531 9255 1534
rect 9156 1523 9255 1531
rect 9182 1522 9254 1523
rect 8833 1496 8904 1512
rect 8833 1480 8853 1496
rect 8834 1450 8853 1480
rect 8836 1430 8853 1450
rect 8883 1450 8904 1496
rect 9876 1492 9954 1573
rect 10321 1518 10429 1573
rect 8883 1430 8903 1450
rect 8836 1411 8903 1430
rect 9876 1390 9955 1492
rect 6670 1367 6756 1376
rect 6670 1349 6689 1367
rect 6741 1349 6756 1367
rect 6670 1345 6756 1349
rect 9840 1372 9961 1390
rect 9840 1370 9911 1372
rect 9840 1329 9855 1370
rect 9892 1331 9911 1370
rect 9948 1331 9961 1372
rect 9892 1329 9961 1331
rect 9840 1319 9961 1329
rect 7145 1291 7256 1294
rect 6460 1290 8009 1291
rect 10322 1290 10429 1518
rect 6460 1287 9619 1290
rect 9806 1287 10431 1290
rect 6460 1277 10431 1287
rect 6460 1257 7152 1277
rect 7171 1257 7229 1277
rect 7248 1272 10431 1277
rect 7248 1257 9647 1272
rect 6460 1252 9647 1257
rect 9666 1252 9724 1272
rect 9743 1252 10431 1272
rect 6460 1234 10431 1252
rect 6460 1231 8009 1234
rect 9640 1230 9751 1234
rect 6512 1183 6547 1184
rect 6491 1176 6547 1183
rect 6491 1156 6520 1176
rect 6540 1156 6547 1176
rect 6491 1151 6547 1156
rect 6938 1179 6970 1186
rect 6938 1159 6944 1179
rect 6965 1159 6970 1179
rect 6491 873 6525 1151
rect 6938 1131 6970 1159
rect 6558 1123 6970 1131
rect 6558 1097 6564 1123
rect 6590 1097 6970 1123
rect 6558 1095 6970 1097
rect 6560 1094 6600 1095
rect 6727 1069 6758 1077
rect 6727 1039 6731 1069
rect 6752 1039 6758 1069
rect 6491 865 6526 873
rect 6491 845 6499 865
rect 6519 845 6526 865
rect 6491 840 6526 845
rect 6491 839 6523 840
rect 6727 838 6758 1039
rect 6938 1030 6970 1095
rect 6938 1010 6942 1030
rect 6963 1010 6970 1030
rect 6938 1003 6970 1010
rect 7532 1170 7625 1177
rect 7532 1129 7556 1170
rect 7610 1129 7625 1170
rect 7247 947 7348 948
rect 7145 934 7348 947
rect 7145 932 7288 934
rect 7145 929 7222 932
rect 7145 902 7148 929
rect 7177 905 7222 929
rect 7251 905 7288 932
rect 7177 902 7288 905
rect 7145 901 7288 902
rect 7324 901 7348 934
rect 7145 888 7348 901
rect 7532 756 7625 1129
rect 8826 1171 8906 1183
rect 9007 1178 9042 1179
rect 8826 1145 8842 1171
rect 8882 1145 8906 1171
rect 8826 1126 8906 1145
rect 8826 1100 8845 1126
rect 8885 1100 8906 1126
rect 8826 1073 8906 1100
rect 8826 1047 8849 1073
rect 8889 1047 8906 1073
rect 8826 1036 8906 1047
rect 8986 1171 9042 1178
rect 8986 1151 9015 1171
rect 9035 1151 9042 1171
rect 8986 1146 9042 1151
rect 9433 1174 9465 1181
rect 9433 1154 9439 1174
rect 9460 1154 9465 1174
rect 7532 712 7550 756
rect 7610 712 7625 756
rect 7532 697 7625 712
rect 8831 736 8896 1036
rect 8986 868 9020 1146
rect 9433 1126 9465 1154
rect 9053 1118 9465 1126
rect 9053 1092 9059 1118
rect 9085 1092 9465 1118
rect 9887 1160 9954 1167
rect 9887 1139 9904 1160
rect 9940 1139 9954 1160
rect 9887 1120 9954 1139
rect 9887 1117 9904 1120
rect 9053 1090 9465 1092
rect 9055 1089 9095 1090
rect 9222 1064 9253 1072
rect 9222 1034 9226 1064
rect 9247 1034 9253 1064
rect 8986 860 9021 868
rect 8986 840 8994 860
rect 9014 840 9021 860
rect 8986 835 9021 840
rect 8986 834 9018 835
rect 9222 830 9253 1034
rect 9433 1025 9465 1090
rect 9889 1083 9904 1117
rect 9944 1083 9954 1120
rect 9889 1074 9954 1083
rect 9433 1005 9437 1025
rect 9458 1005 9465 1025
rect 9433 998 9465 1005
rect 9742 942 9843 943
rect 9640 929 9843 942
rect 9640 927 9783 929
rect 9640 924 9717 927
rect 9640 897 9643 924
rect 9672 900 9717 924
rect 9746 900 9783 927
rect 9672 897 9783 900
rect 9640 896 9783 897
rect 9819 896 9843 929
rect 9640 883 9843 896
rect 9220 818 9255 830
rect 9151 811 9255 818
rect 9151 810 9227 811
rect 9151 790 9172 810
rect 9204 791 9227 810
rect 9252 791 9255 811
rect 9204 790 9255 791
rect 9151 781 9255 790
rect 9220 779 9255 781
rect 8831 697 8834 736
rect 8879 697 8896 736
rect 9892 713 9943 1074
rect 9890 711 9947 713
rect 8831 675 8896 697
rect 9879 699 9947 711
rect 9879 666 9890 699
rect 9930 666 9947 699
rect 9879 660 9947 666
rect 9879 656 9943 660
rect 8592 611 8703 614
rect 10322 611 10429 1234
rect 6855 597 10429 611
rect 6855 577 8599 597
rect 8618 577 8676 597
rect 8695 593 10429 597
rect 8695 577 9647 593
rect 6855 573 9647 577
rect 9666 573 9724 593
rect 9743 573 10429 593
rect 6855 555 10429 573
rect 6855 554 7968 555
rect 9640 551 9751 555
rect 7959 503 7994 504
rect 7938 496 7994 503
rect 7938 476 7967 496
rect 7987 476 7994 496
rect 7938 471 7994 476
rect 8385 499 8417 506
rect 9007 499 9042 500
rect 8385 479 8391 499
rect 8412 479 8417 499
rect 8986 492 9042 499
rect 8851 482 8909 487
rect 5774 436 7627 469
rect 5774 371 5839 436
rect 5970 416 7627 436
rect 5970 375 7563 416
rect 7599 375 7627 416
rect 7725 436 7789 455
rect 7725 397 7742 436
rect 7776 397 7789 436
rect 7725 378 7789 397
rect 5970 371 7627 375
rect 5774 346 7627 371
rect 7538 343 7620 346
rect 7727 -134 7789 378
rect 7938 193 7972 471
rect 8385 451 8417 479
rect 8005 443 8417 451
rect 8005 417 8011 443
rect 8037 417 8417 443
rect 8005 415 8417 417
rect 8007 414 8047 415
rect 8174 389 8205 397
rect 8174 359 8178 389
rect 8199 359 8205 389
rect 7938 185 7973 193
rect 7938 165 7946 185
rect 7966 165 7973 185
rect 7938 160 7973 165
rect 7938 159 7970 160
rect 8174 152 8205 359
rect 8385 350 8417 415
rect 8385 330 8389 350
rect 8410 330 8417 350
rect 8385 323 8417 330
rect 8834 473 8909 482
rect 8834 440 8843 473
rect 8896 440 8909 473
rect 8834 415 8909 440
rect 8834 382 8848 415
rect 8901 382 8909 415
rect 8834 376 8909 382
rect 8986 472 9015 492
rect 9035 472 9042 492
rect 8986 467 9042 472
rect 9433 495 9465 502
rect 9433 475 9439 495
rect 9460 475 9465 495
rect 8694 267 8795 268
rect 8592 254 8795 267
rect 8592 252 8735 254
rect 8592 249 8669 252
rect 8592 222 8595 249
rect 8624 225 8669 249
rect 8698 225 8735 252
rect 8624 222 8735 225
rect 8592 221 8735 222
rect 8771 221 8795 254
rect 8592 208 8795 221
rect 8169 134 8205 152
rect 8136 133 8205 134
rect 8116 121 8205 133
rect 8116 83 8128 121
rect 8153 86 8172 121
rect 8197 86 8205 121
rect 8153 83 8205 86
rect 8116 75 8205 83
rect 8132 74 8204 75
rect 7685 -192 7801 -134
rect 8834 -145 8904 376
rect 8986 189 9020 467
rect 9433 447 9465 475
rect 9053 439 9465 447
rect 9053 413 9059 439
rect 9085 413 9465 439
rect 9053 411 9465 413
rect 9055 410 9095 411
rect 9222 385 9253 393
rect 9222 355 9226 385
rect 9247 355 9253 385
rect 8986 181 9021 189
rect 8986 161 8994 181
rect 9014 161 9021 181
rect 8986 156 9021 161
rect 9222 156 9253 355
rect 9433 346 9465 411
rect 9433 326 9437 346
rect 9458 326 9465 346
rect 9433 319 9465 326
rect 9878 472 9950 490
rect 9878 430 9891 472
rect 9940 430 9950 472
rect 9878 409 9950 430
rect 9878 367 9892 409
rect 9941 367 9950 409
rect 9742 263 9843 264
rect 9640 250 9843 263
rect 9640 248 9783 250
rect 9640 245 9717 248
rect 9640 218 9643 245
rect 9672 221 9717 245
rect 9746 221 9783 248
rect 9672 218 9783 221
rect 9640 217 9783 218
rect 9819 217 9843 250
rect 9640 204 9843 217
rect 8986 155 9018 156
rect 9220 153 9253 156
rect 9186 134 9254 153
rect 9156 122 9255 134
rect 9156 84 9178 122
rect 9203 87 9222 122
rect 9247 87 9255 122
rect 9203 84 9255 87
rect 9156 76 9255 84
rect 9182 75 9254 76
rect 7685 -263 7697 -192
rect 7776 -263 7801 -192
rect 7685 -283 7801 -263
rect 8815 -346 8917 -145
rect 9878 -153 9950 367
rect 10322 -57 10429 555
rect 10321 -93 10429 -57
rect 10476 66 10630 91
rect 10476 -46 10489 66
rect 10610 -46 10630 66
rect 8779 -383 8945 -346
rect 8779 -462 8816 -383
rect 8900 -462 8945 -383
rect 8779 -500 8945 -462
rect 9856 -554 9953 -153
rect 10314 -229 10434 -93
rect 10321 -235 10429 -229
rect 9786 -583 9961 -554
rect 9786 -662 9832 -583
rect 9932 -662 9961 -583
rect 9786 -687 9961 -662
rect 10321 -778 10425 -235
rect 10164 -808 10435 -778
rect 10164 -895 10198 -808
rect 10268 -816 10435 -808
rect 10268 -895 10331 -816
rect 10164 -903 10331 -895
rect 10401 -903 10435 -816
rect 10164 -949 10435 -903
rect 10476 -1020 10630 -46
rect 10474 -1036 10630 -1020
rect 10474 -1061 10626 -1036
rect 10474 -1156 10504 -1061
rect 10594 -1156 10626 -1061
rect 10474 -1169 10626 -1156
<< via1 >>
rect 787 11700 823 11733
rect 1835 11696 1871 11729
rect 787 11021 823 11054
rect 3282 11016 3318 11049
rect 787 10253 823 10286
rect 1835 10249 1871 10282
rect 787 9574 823 9607
rect 3325 9571 3361 9604
rect 788 8733 824 8766
rect 1836 8729 1872 8762
rect 788 8054 824 8087
rect 3283 8049 3319 8082
rect 788 7286 824 7319
rect 1836 7282 1872 7315
rect 788 6607 824 6640
rect 5310 11142 5381 11351
rect 4391 6598 4427 6631
rect 785 5692 821 5725
rect 1833 5688 1869 5721
rect 785 5013 821 5046
rect 3280 5008 3316 5041
rect 785 4245 821 4278
rect 1833 4241 1869 4274
rect 9784 11318 9820 11351
rect 8736 10643 8772 10676
rect 9784 10639 9820 10672
rect 7289 9876 7325 9909
rect 9784 9871 9820 9904
rect 8736 9196 8772 9229
rect 9784 9192 9820 9225
rect 7247 8354 7283 8387
rect 9785 8351 9821 8384
rect 8737 7676 8773 7709
rect 9785 7672 9821 7705
rect 7290 6909 7326 6942
rect 9785 6904 9821 6937
rect 8737 6229 8773 6262
rect 9785 6225 9821 6258
rect 6179 5319 6215 5352
rect 785 3566 821 3599
rect 3323 3563 3359 3596
rect 786 2725 822 2758
rect 1834 2721 1870 2754
rect 4736 2727 4772 2760
rect 786 2046 822 2079
rect 3281 2041 3317 2074
rect 786 1278 822 1311
rect 1834 1274 1870 1307
rect 786 599 822 632
rect 13 -67 92 45
rect 2767 -263 2884 -188
rect 1719 -458 1789 -383
rect 670 -674 770 -595
rect 217 -903 287 -816
rect -15 -1151 75 -1056
rect 9782 5310 9818 5343
rect 8734 4635 8770 4668
rect 9782 4631 9818 4664
rect 7287 3868 7323 3901
rect 9782 3863 9818 3896
rect 8734 3188 8770 3221
rect 9782 3184 9818 3217
rect 7245 2346 7281 2379
rect 9783 2343 9819 2376
rect 8735 1668 8771 1701
rect 9783 1664 9819 1697
rect 7288 901 7324 934
rect 9783 896 9819 929
rect 8735 221 8771 254
rect 9783 217 9819 250
rect 7697 -263 7776 -192
rect 10489 -46 10610 66
rect 8816 -462 8900 -383
rect 9832 -662 9932 -583
rect 10198 -895 10268 -808
rect 10331 -903 10401 -816
rect 10504 -1156 10594 -1061
<< metal2 >>
rect 6 11748 113 12182
rect 6 11733 3751 11748
rect 6 11700 787 11733
rect 823 11729 3751 11733
rect 823 11700 1835 11729
rect 6 11696 1835 11700
rect 1871 11696 3751 11729
rect 6 11679 3751 11696
rect 6 11073 113 11679
rect 2613 11677 3751 11679
rect 5293 11351 5398 12246
rect 5293 11142 5310 11351
rect 5381 11142 5398 11351
rect 6357 11368 7862 11369
rect 10494 11368 10601 11914
rect 6357 11351 10601 11368
rect 6357 11318 9784 11351
rect 9820 11318 10601 11351
rect 6357 11299 10601 11318
rect 6357 11297 7862 11299
rect 5293 11100 5398 11142
rect 6 11054 4146 11073
rect 6 11021 787 11054
rect 823 11049 4146 11054
rect 823 11021 3282 11049
rect 6 11016 3282 11021
rect 3318 11016 4146 11049
rect 6 11004 4146 11016
rect 6 10301 113 11004
rect 2534 11003 4146 11004
rect 10494 10693 10601 11299
rect 6357 10676 10601 10693
rect 6357 10643 8736 10676
rect 8772 10672 10601 10676
rect 8772 10643 9784 10672
rect 6357 10639 9784 10643
rect 9820 10639 10601 10672
rect 6357 10624 10601 10639
rect 6357 10621 7896 10624
rect 2763 10304 3006 10309
rect 2711 10301 3971 10304
rect 6 10286 3971 10301
rect 6 10253 787 10286
rect 823 10282 3971 10286
rect 823 10253 1835 10282
rect 6 10249 1835 10253
rect 1871 10249 3971 10282
rect 6 10232 3971 10249
rect 6 9626 113 10232
rect 2763 10223 3006 10232
rect 6358 9921 8073 9922
rect 10494 9921 10601 10624
rect 6358 9909 10601 9921
rect 6358 9876 7289 9909
rect 7325 9904 10601 9909
rect 7325 9876 9784 9904
rect 6358 9871 9784 9876
rect 9820 9871 10601 9904
rect 6358 9852 10601 9871
rect 2745 9626 4195 9628
rect 6 9607 4195 9626
rect 6 9574 787 9607
rect 823 9604 4195 9607
rect 823 9574 3325 9604
rect 6 9571 3325 9574
rect 3361 9571 4195 9604
rect 6 9557 4195 9571
rect 6 9022 113 9557
rect 2745 9556 4195 9557
rect 5980 9246 7994 9248
rect 10494 9246 10601 9852
rect 5980 9229 10601 9246
rect 5980 9196 8736 9229
rect 8772 9225 10601 9229
rect 8772 9196 9784 9225
rect 5980 9192 9784 9196
rect 9820 9192 10601 9225
rect 5980 9177 10601 9192
rect 7665 9175 7853 9177
rect 6 9021 114 9022
rect 7 8998 114 9021
rect 5 8954 114 8998
rect 7 8781 114 8954
rect 10494 9004 10601 9177
rect 10494 8960 10603 9004
rect 10494 8937 10601 8960
rect 10494 8936 10602 8937
rect 2755 8781 2943 8783
rect 7 8766 3939 8781
rect 7 8733 788 8766
rect 824 8762 3939 8766
rect 824 8733 1836 8762
rect 7 8729 1836 8733
rect 1872 8729 3939 8762
rect 7 8712 3939 8729
rect 7 8106 114 8712
rect 2614 8710 3939 8712
rect 6367 8401 7863 8402
rect 10495 8401 10602 8936
rect 6367 8387 10602 8401
rect 6367 8354 7247 8387
rect 7283 8384 10602 8387
rect 7283 8354 9785 8384
rect 6367 8351 9785 8354
rect 9821 8351 10602 8384
rect 6367 8332 10602 8351
rect 6367 8330 7863 8332
rect 7 8087 4148 8106
rect 7 8054 788 8087
rect 824 8082 4148 8087
rect 824 8054 3283 8082
rect 7 8049 3283 8054
rect 3319 8049 4148 8082
rect 7 8037 4148 8049
rect 7 7334 114 8037
rect 2535 8036 4148 8037
rect 7602 7726 7845 7735
rect 10495 7726 10602 8332
rect 6367 7709 10602 7726
rect 6367 7676 8737 7709
rect 8773 7705 10602 7709
rect 8773 7676 9785 7705
rect 6367 7672 9785 7676
rect 9821 7672 10602 7705
rect 6367 7657 10602 7672
rect 6367 7654 7897 7657
rect 7602 7649 7845 7654
rect 2712 7334 3721 7337
rect 7 7319 3721 7334
rect 7 7286 788 7319
rect 824 7315 3721 7319
rect 824 7286 1836 7315
rect 7 7282 1836 7286
rect 1872 7282 3721 7315
rect 7 7265 3721 7282
rect 7 6659 114 7265
rect 6367 6954 8074 6955
rect 10495 6954 10602 7657
rect 6367 6942 10602 6954
rect 6367 6909 7290 6942
rect 7326 6937 10602 6942
rect 7326 6909 9785 6937
rect 6367 6904 9785 6909
rect 9821 6904 10602 6937
rect 6367 6885 10602 6904
rect 2746 6660 4251 6661
rect 2746 6659 4451 6660
rect 7 6644 4451 6659
rect 7 6640 4454 6644
rect 7 6607 788 6640
rect 824 6631 4454 6640
rect 824 6607 4391 6631
rect 7 6598 4391 6607
rect 4427 6598 4454 6631
rect 7 6590 4454 6598
rect 7 6073 114 6590
rect 2746 6589 4454 6590
rect 4216 6586 4454 6589
rect 6423 6279 7995 6281
rect 10495 6279 10602 6885
rect 6423 6262 10602 6279
rect 6423 6229 8737 6262
rect 8773 6258 10602 6262
rect 8773 6229 9785 6258
rect 6423 6225 9785 6229
rect 9821 6225 10602 6258
rect 6423 6210 10602 6225
rect 0 5881 116 6073
rect 10495 6069 10602 6210
rect 4 5740 111 5881
rect 10490 5877 10606 6069
rect 4 5725 4183 5740
rect 4 5692 785 5725
rect 821 5721 4183 5725
rect 821 5692 1833 5721
rect 4 5688 1833 5692
rect 1869 5688 4183 5721
rect 4 5671 4183 5688
rect 4 5065 111 5671
rect 2611 5669 4183 5671
rect 6152 5361 6286 5364
rect 6373 5361 6390 5364
rect 6152 5360 7860 5361
rect 10492 5360 10599 5877
rect 6152 5352 10599 5360
rect 6152 5319 6179 5352
rect 6215 5343 10599 5352
rect 6215 5319 9782 5343
rect 6152 5310 9782 5319
rect 9818 5310 10599 5343
rect 6152 5306 10599 5310
rect 6155 5291 10599 5306
rect 6155 5290 7860 5291
rect 6271 5289 7860 5290
rect 6271 5274 6393 5289
rect 4 5046 4239 5065
rect 4 5013 785 5046
rect 821 5041 4239 5046
rect 821 5013 3280 5041
rect 4 5008 3280 5013
rect 3316 5008 4239 5041
rect 4 4996 4239 5008
rect 4 4293 111 4996
rect 2532 4995 4239 4996
rect 10492 4685 10599 5291
rect 6885 4668 10599 4685
rect 6885 4635 8734 4668
rect 8770 4664 10599 4668
rect 8770 4635 9782 4664
rect 6885 4631 9782 4635
rect 9818 4631 10599 4664
rect 6885 4616 10599 4631
rect 6885 4613 7894 4616
rect 2761 4296 3004 4301
rect 2709 4293 4239 4296
rect 4 4278 4239 4293
rect 4 4245 785 4278
rect 821 4274 4239 4278
rect 821 4245 1833 4274
rect 4 4241 1833 4245
rect 1869 4241 4239 4274
rect 4 4224 4239 4241
rect 4 3618 111 4224
rect 2761 4215 3004 4224
rect 6458 3913 8071 3914
rect 10492 3913 10599 4616
rect 6458 3901 10599 3913
rect 6458 3868 7287 3901
rect 7323 3896 10599 3901
rect 7323 3868 9782 3896
rect 6458 3863 9782 3868
rect 9818 3863 10599 3896
rect 6458 3844 10599 3863
rect 2743 3618 4239 3620
rect 4 3599 4239 3618
rect 4 3566 785 3599
rect 821 3596 4239 3599
rect 821 3566 3323 3596
rect 4 3563 3323 3566
rect 3359 3563 4239 3596
rect 4 3549 4239 3563
rect 4 3014 111 3549
rect 2743 3548 4239 3549
rect 6667 3238 7992 3240
rect 10492 3238 10599 3844
rect 6667 3221 10599 3238
rect 6667 3188 8734 3221
rect 8770 3217 10599 3221
rect 8770 3188 9782 3217
rect 6667 3184 9782 3188
rect 9818 3184 10599 3217
rect 6667 3169 10599 3184
rect 7663 3167 7851 3169
rect 4 3013 112 3014
rect 5 2990 112 3013
rect 3 2946 112 2990
rect 5 2773 112 2946
rect 10492 2996 10599 3169
rect 10492 2952 10601 2996
rect 10492 2929 10599 2952
rect 10492 2928 10600 2929
rect 2753 2773 2941 2775
rect 4532 2773 4950 2780
rect 5 2760 4950 2773
rect 5 2758 4736 2760
rect 5 2725 786 2758
rect 822 2754 4736 2758
rect 822 2725 1834 2754
rect 5 2721 1834 2725
rect 1870 2727 4736 2754
rect 4772 2727 4950 2760
rect 1870 2721 4950 2727
rect 5 2709 4950 2721
rect 5 2704 4626 2709
rect 5 2098 112 2704
rect 2612 2702 4626 2704
rect 6411 2393 7861 2394
rect 10493 2393 10600 2928
rect 6411 2379 10600 2393
rect 6411 2346 7245 2379
rect 7281 2376 10600 2379
rect 7281 2346 9783 2376
rect 6411 2343 9783 2346
rect 9819 2343 10600 2376
rect 6411 2324 10600 2343
rect 6411 2322 7861 2324
rect 5 2079 4248 2098
rect 5 2046 786 2079
rect 822 2074 4248 2079
rect 822 2046 3281 2074
rect 5 2041 3281 2046
rect 3317 2041 4248 2074
rect 5 2029 4248 2041
rect 5 1326 112 2029
rect 2533 2028 4248 2029
rect 7600 1718 7843 1727
rect 10493 1718 10600 2324
rect 6635 1701 10600 1718
rect 6635 1668 8735 1701
rect 8771 1697 10600 1701
rect 8771 1668 9783 1697
rect 6635 1664 9783 1668
rect 9819 1664 10600 1697
rect 6635 1649 10600 1664
rect 6635 1646 7895 1649
rect 7600 1641 7843 1646
rect 2710 1326 4249 1329
rect 5 1311 4249 1326
rect 5 1278 786 1311
rect 822 1307 4249 1311
rect 822 1278 1834 1307
rect 5 1274 1834 1278
rect 1870 1274 4249 1307
rect 5 1257 4249 1274
rect 5 651 112 1257
rect 6460 946 8072 947
rect 10493 946 10600 1649
rect 6460 934 10600 946
rect 6460 901 7288 934
rect 7324 929 10600 934
rect 7324 901 9783 929
rect 6460 896 9783 901
rect 9819 896 10600 929
rect 6460 877 10600 896
rect 2744 651 4249 653
rect 5 632 4249 651
rect 5 599 786 632
rect 822 599 4249 632
rect 5 582 4249 599
rect 5 83 112 582
rect 2744 581 4249 582
rect 7635 271 7993 273
rect 10493 271 10600 877
rect 7635 254 10600 271
rect 7635 221 8735 254
rect 8771 250 10600 254
rect 8771 221 9783 250
rect 7635 217 9783 221
rect 9819 220 10600 250
rect 9819 217 10639 220
rect 7635 202 10639 217
rect -20 45 113 83
rect -20 -67 13 45
rect 92 14 113 45
rect 10468 66 10639 202
rect 92 -30 125 14
rect 92 -67 113 -30
rect -20 -84 113 -67
rect 10468 -46 10489 66
rect 10610 -46 10639 66
rect 10468 -96 10639 -46
rect 2738 -188 7801 -179
rect 2738 -263 2767 -188
rect 2884 -192 7801 -188
rect 2884 -263 7697 -192
rect 7776 -263 7801 -192
rect 2738 -279 7801 -263
rect 1694 -383 8925 -356
rect 1694 -458 1719 -383
rect 1789 -458 8816 -383
rect 1694 -462 8816 -458
rect 8900 -462 8925 -383
rect 1694 -489 8925 -462
rect 645 -583 9952 -566
rect 645 -595 9832 -583
rect 645 -674 670 -595
rect 770 -662 9832 -595
rect 9932 -662 9952 -583
rect 770 -674 9952 -662
rect 645 -683 9952 -674
rect 179 -808 10439 -783
rect 179 -816 10198 -808
rect 179 -903 217 -816
rect 287 -895 10198 -816
rect 10268 -816 10439 -808
rect 10268 -895 10331 -816
rect 287 -903 10331 -895
rect 10401 -903 10439 -816
rect 179 -945 10439 -903
rect -40 -1056 10633 -1027
rect -40 -1151 -15 -1056
rect 75 -1061 10633 -1056
rect 75 -1151 10504 -1061
rect -40 -1156 10504 -1151
rect 10594 -1156 10633 -1061
rect -40 -1181 10633 -1156
<< labels >>
rlabel metal1 4258 12210 4293 12224 1 d4
rlabel metal1 2996 12165 3048 12184 1 d3
rlabel metal1 2820 12182 2870 12195 1 d2
rlabel metal1 1710 12119 1763 12141 1 d1
rlabel metal1 664 12137 726 12164 1 d0
rlabel metal2 9 12122 105 12155 1 vdd
rlabel metal1 185 12122 281 12155 1 gnd
rlabel locali 449 12133 493 12155 1 vref
rlabel metal2 5306 12146 5385 12217 1 d5
rlabel metal1 5307 2826 5330 2839 1 vout
<< end >>
