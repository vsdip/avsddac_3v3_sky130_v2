magic
tech sky130A
timestamp 1620564505
<< nwell >>
rect 282 4310 609 4384
rect 282 4160 1093 4310
rect 1220 4066 1547 4140
rect 1220 3916 2031 4066
rect 281 3756 608 3830
rect 281 3606 1092 3756
rect 1361 3474 1688 3548
rect 1361 3324 2172 3474
rect 283 3207 610 3281
rect 283 3057 1094 3207
rect 1221 2963 1548 3037
rect 1221 2813 2032 2963
rect 282 2653 609 2727
rect 282 2503 1093 2653
rect 1331 2384 1658 2458
rect 1331 2234 2142 2384
rect 283 2104 610 2178
rect 283 1954 1094 2104
rect 1221 1860 1548 1934
rect 1221 1710 2032 1860
rect 282 1550 609 1624
rect 282 1400 1093 1550
rect 1362 1268 1689 1342
rect 1362 1118 2173 1268
rect 284 1001 611 1075
rect 284 851 1095 1001
rect 1222 757 1549 831
rect 1222 607 2033 757
rect 283 447 610 521
rect 283 297 1094 447
rect 1331 184 1658 258
rect 1331 34 2142 184
rect 284 -102 611 -28
rect 284 -252 1095 -102
rect 1222 -346 1549 -272
rect 1222 -496 2033 -346
rect 283 -656 610 -582
rect 283 -806 1094 -656
rect 1363 -938 1690 -864
rect 1363 -1088 2174 -938
rect 285 -1205 612 -1131
rect 285 -1355 1096 -1205
rect 1223 -1449 1550 -1375
rect 1223 -1599 2034 -1449
rect 284 -1759 611 -1685
rect 284 -1909 1095 -1759
rect 1333 -2028 1660 -1954
rect 1333 -2178 2144 -2028
rect 285 -2308 612 -2234
rect 285 -2458 1096 -2308
rect 1223 -2552 1550 -2478
rect 1223 -2702 2034 -2552
rect 284 -2862 611 -2788
rect 284 -3012 1095 -2862
rect 1364 -3144 1691 -3070
rect 1364 -3294 2175 -3144
rect 286 -3411 613 -3337
rect 286 -3561 1097 -3411
rect 1224 -3655 1551 -3581
rect 1224 -3805 2035 -3655
rect 285 -3965 612 -3891
rect 285 -4115 1096 -3965
<< nmos >>
rect 346 4059 396 4101
rect 559 4059 609 4101
rect 767 4059 817 4101
rect 975 4059 1025 4101
rect 1284 3815 1334 3857
rect 1497 3815 1547 3857
rect 1705 3815 1755 3857
rect 1913 3815 1963 3857
rect 345 3505 395 3547
rect 558 3505 608 3547
rect 766 3505 816 3547
rect 974 3505 1024 3547
rect 1425 3223 1475 3265
rect 1638 3223 1688 3265
rect 1846 3223 1896 3265
rect 2054 3223 2104 3265
rect 347 2956 397 2998
rect 560 2956 610 2998
rect 768 2956 818 2998
rect 976 2956 1026 2998
rect 1285 2712 1335 2754
rect 1498 2712 1548 2754
rect 1706 2712 1756 2754
rect 1914 2712 1964 2754
rect 346 2402 396 2444
rect 559 2402 609 2444
rect 767 2402 817 2444
rect 975 2402 1025 2444
rect 1395 2133 1445 2175
rect 1608 2133 1658 2175
rect 1816 2133 1866 2175
rect 2024 2133 2074 2175
rect 347 1853 397 1895
rect 560 1853 610 1895
rect 768 1853 818 1895
rect 976 1853 1026 1895
rect 1285 1609 1335 1651
rect 1498 1609 1548 1651
rect 1706 1609 1756 1651
rect 1914 1609 1964 1651
rect 346 1299 396 1341
rect 559 1299 609 1341
rect 767 1299 817 1341
rect 975 1299 1025 1341
rect 1426 1017 1476 1059
rect 1639 1017 1689 1059
rect 1847 1017 1897 1059
rect 2055 1017 2105 1059
rect 348 750 398 792
rect 561 750 611 792
rect 769 750 819 792
rect 977 750 1027 792
rect 1286 506 1336 548
rect 1499 506 1549 548
rect 1707 506 1757 548
rect 1915 506 1965 548
rect 347 196 397 238
rect 560 196 610 238
rect 768 196 818 238
rect 976 196 1026 238
rect 1395 -67 1445 -25
rect 1608 -67 1658 -25
rect 1816 -67 1866 -25
rect 2024 -67 2074 -25
rect 348 -353 398 -311
rect 561 -353 611 -311
rect 769 -353 819 -311
rect 977 -353 1027 -311
rect 1286 -597 1336 -555
rect 1499 -597 1549 -555
rect 1707 -597 1757 -555
rect 1915 -597 1965 -555
rect 347 -907 397 -865
rect 560 -907 610 -865
rect 768 -907 818 -865
rect 976 -907 1026 -865
rect 1427 -1189 1477 -1147
rect 1640 -1189 1690 -1147
rect 1848 -1189 1898 -1147
rect 2056 -1189 2106 -1147
rect 349 -1456 399 -1414
rect 562 -1456 612 -1414
rect 770 -1456 820 -1414
rect 978 -1456 1028 -1414
rect 1287 -1700 1337 -1658
rect 1500 -1700 1550 -1658
rect 1708 -1700 1758 -1658
rect 1916 -1700 1966 -1658
rect 348 -2010 398 -1968
rect 561 -2010 611 -1968
rect 769 -2010 819 -1968
rect 977 -2010 1027 -1968
rect 1397 -2279 1447 -2237
rect 1610 -2279 1660 -2237
rect 1818 -2279 1868 -2237
rect 2026 -2279 2076 -2237
rect 349 -2559 399 -2517
rect 562 -2559 612 -2517
rect 770 -2559 820 -2517
rect 978 -2559 1028 -2517
rect 1287 -2803 1337 -2761
rect 1500 -2803 1550 -2761
rect 1708 -2803 1758 -2761
rect 1916 -2803 1966 -2761
rect 348 -3113 398 -3071
rect 561 -3113 611 -3071
rect 769 -3113 819 -3071
rect 977 -3113 1027 -3071
rect 1428 -3395 1478 -3353
rect 1641 -3395 1691 -3353
rect 1849 -3395 1899 -3353
rect 2057 -3395 2107 -3353
rect 350 -3662 400 -3620
rect 563 -3662 613 -3620
rect 771 -3662 821 -3620
rect 979 -3662 1029 -3620
rect 1288 -3906 1338 -3864
rect 1501 -3906 1551 -3864
rect 1709 -3906 1759 -3864
rect 1917 -3906 1967 -3864
rect 349 -4216 399 -4174
rect 562 -4216 612 -4174
rect 770 -4216 820 -4174
rect 978 -4216 1028 -4174
<< pmos >>
rect 346 4178 396 4278
rect 559 4178 609 4278
rect 767 4178 817 4278
rect 975 4178 1025 4278
rect 1284 3934 1334 4034
rect 1497 3934 1547 4034
rect 1705 3934 1755 4034
rect 1913 3934 1963 4034
rect 345 3624 395 3724
rect 558 3624 608 3724
rect 766 3624 816 3724
rect 974 3624 1024 3724
rect 1425 3342 1475 3442
rect 1638 3342 1688 3442
rect 1846 3342 1896 3442
rect 2054 3342 2104 3442
rect 347 3075 397 3175
rect 560 3075 610 3175
rect 768 3075 818 3175
rect 976 3075 1026 3175
rect 1285 2831 1335 2931
rect 1498 2831 1548 2931
rect 1706 2831 1756 2931
rect 1914 2831 1964 2931
rect 346 2521 396 2621
rect 559 2521 609 2621
rect 767 2521 817 2621
rect 975 2521 1025 2621
rect 1395 2252 1445 2352
rect 1608 2252 1658 2352
rect 1816 2252 1866 2352
rect 2024 2252 2074 2352
rect 347 1972 397 2072
rect 560 1972 610 2072
rect 768 1972 818 2072
rect 976 1972 1026 2072
rect 1285 1728 1335 1828
rect 1498 1728 1548 1828
rect 1706 1728 1756 1828
rect 1914 1728 1964 1828
rect 346 1418 396 1518
rect 559 1418 609 1518
rect 767 1418 817 1518
rect 975 1418 1025 1518
rect 1426 1136 1476 1236
rect 1639 1136 1689 1236
rect 1847 1136 1897 1236
rect 2055 1136 2105 1236
rect 348 869 398 969
rect 561 869 611 969
rect 769 869 819 969
rect 977 869 1027 969
rect 1286 625 1336 725
rect 1499 625 1549 725
rect 1707 625 1757 725
rect 1915 625 1965 725
rect 347 315 397 415
rect 560 315 610 415
rect 768 315 818 415
rect 976 315 1026 415
rect 1395 52 1445 152
rect 1608 52 1658 152
rect 1816 52 1866 152
rect 2024 52 2074 152
rect 348 -234 398 -134
rect 561 -234 611 -134
rect 769 -234 819 -134
rect 977 -234 1027 -134
rect 1286 -478 1336 -378
rect 1499 -478 1549 -378
rect 1707 -478 1757 -378
rect 1915 -478 1965 -378
rect 347 -788 397 -688
rect 560 -788 610 -688
rect 768 -788 818 -688
rect 976 -788 1026 -688
rect 1427 -1070 1477 -970
rect 1640 -1070 1690 -970
rect 1848 -1070 1898 -970
rect 2056 -1070 2106 -970
rect 349 -1337 399 -1237
rect 562 -1337 612 -1237
rect 770 -1337 820 -1237
rect 978 -1337 1028 -1237
rect 1287 -1581 1337 -1481
rect 1500 -1581 1550 -1481
rect 1708 -1581 1758 -1481
rect 1916 -1581 1966 -1481
rect 348 -1891 398 -1791
rect 561 -1891 611 -1791
rect 769 -1891 819 -1791
rect 977 -1891 1027 -1791
rect 1397 -2160 1447 -2060
rect 1610 -2160 1660 -2060
rect 1818 -2160 1868 -2060
rect 2026 -2160 2076 -2060
rect 349 -2440 399 -2340
rect 562 -2440 612 -2340
rect 770 -2440 820 -2340
rect 978 -2440 1028 -2340
rect 1287 -2684 1337 -2584
rect 1500 -2684 1550 -2584
rect 1708 -2684 1758 -2584
rect 1916 -2684 1966 -2584
rect 348 -2994 398 -2894
rect 561 -2994 611 -2894
rect 769 -2994 819 -2894
rect 977 -2994 1027 -2894
rect 1428 -3276 1478 -3176
rect 1641 -3276 1691 -3176
rect 1849 -3276 1899 -3176
rect 2057 -3276 2107 -3176
rect 350 -3543 400 -3443
rect 563 -3543 613 -3443
rect 771 -3543 821 -3443
rect 979 -3543 1029 -3443
rect 1288 -3787 1338 -3687
rect 1501 -3787 1551 -3687
rect 1709 -3787 1759 -3687
rect 1917 -3787 1967 -3687
rect 349 -4097 399 -3997
rect 562 -4097 612 -3997
rect 770 -4097 820 -3997
rect 978 -4097 1028 -3997
<< ndiff >>
rect 297 4091 346 4101
rect 297 4071 308 4091
rect 328 4071 346 4091
rect 297 4059 346 4071
rect 396 4095 440 4101
rect 396 4075 411 4095
rect 431 4075 440 4095
rect 396 4059 440 4075
rect 510 4091 559 4101
rect 510 4071 521 4091
rect 541 4071 559 4091
rect 510 4059 559 4071
rect 609 4095 653 4101
rect 609 4075 624 4095
rect 644 4075 653 4095
rect 609 4059 653 4075
rect 718 4091 767 4101
rect 718 4071 729 4091
rect 749 4071 767 4091
rect 718 4059 767 4071
rect 817 4095 861 4101
rect 817 4075 832 4095
rect 852 4075 861 4095
rect 817 4059 861 4075
rect 931 4095 975 4101
rect 931 4075 940 4095
rect 960 4075 975 4095
rect 931 4059 975 4075
rect 1025 4091 1074 4101
rect 1025 4071 1043 4091
rect 1063 4071 1074 4091
rect 1025 4059 1074 4071
rect 1235 3847 1284 3857
rect 1235 3827 1246 3847
rect 1266 3827 1284 3847
rect 1235 3815 1284 3827
rect 1334 3851 1378 3857
rect 1334 3831 1349 3851
rect 1369 3831 1378 3851
rect 1334 3815 1378 3831
rect 1448 3847 1497 3857
rect 1448 3827 1459 3847
rect 1479 3827 1497 3847
rect 1448 3815 1497 3827
rect 1547 3851 1591 3857
rect 1547 3831 1562 3851
rect 1582 3831 1591 3851
rect 1547 3815 1591 3831
rect 1656 3847 1705 3857
rect 1656 3827 1667 3847
rect 1687 3827 1705 3847
rect 1656 3815 1705 3827
rect 1755 3851 1799 3857
rect 1755 3831 1770 3851
rect 1790 3831 1799 3851
rect 1755 3815 1799 3831
rect 1869 3851 1913 3857
rect 1869 3831 1878 3851
rect 1898 3831 1913 3851
rect 1869 3815 1913 3831
rect 1963 3847 2012 3857
rect 1963 3827 1981 3847
rect 2001 3827 2012 3847
rect 1963 3815 2012 3827
rect 296 3537 345 3547
rect 296 3517 307 3537
rect 327 3517 345 3537
rect 296 3505 345 3517
rect 395 3541 439 3547
rect 395 3521 410 3541
rect 430 3521 439 3541
rect 395 3505 439 3521
rect 509 3537 558 3547
rect 509 3517 520 3537
rect 540 3517 558 3537
rect 509 3505 558 3517
rect 608 3541 652 3547
rect 608 3521 623 3541
rect 643 3521 652 3541
rect 608 3505 652 3521
rect 717 3537 766 3547
rect 717 3517 728 3537
rect 748 3517 766 3537
rect 717 3505 766 3517
rect 816 3541 860 3547
rect 816 3521 831 3541
rect 851 3521 860 3541
rect 816 3505 860 3521
rect 930 3541 974 3547
rect 930 3521 939 3541
rect 959 3521 974 3541
rect 930 3505 974 3521
rect 1024 3537 1073 3547
rect 1024 3517 1042 3537
rect 1062 3517 1073 3537
rect 1024 3505 1073 3517
rect 1376 3255 1425 3265
rect 1376 3235 1387 3255
rect 1407 3235 1425 3255
rect 1376 3223 1425 3235
rect 1475 3259 1519 3265
rect 1475 3239 1490 3259
rect 1510 3239 1519 3259
rect 1475 3223 1519 3239
rect 1589 3255 1638 3265
rect 1589 3235 1600 3255
rect 1620 3235 1638 3255
rect 1589 3223 1638 3235
rect 1688 3259 1732 3265
rect 1688 3239 1703 3259
rect 1723 3239 1732 3259
rect 1688 3223 1732 3239
rect 1797 3255 1846 3265
rect 1797 3235 1808 3255
rect 1828 3235 1846 3255
rect 1797 3223 1846 3235
rect 1896 3259 1940 3265
rect 1896 3239 1911 3259
rect 1931 3239 1940 3259
rect 1896 3223 1940 3239
rect 2010 3259 2054 3265
rect 2010 3239 2019 3259
rect 2039 3239 2054 3259
rect 2010 3223 2054 3239
rect 2104 3255 2153 3265
rect 2104 3235 2122 3255
rect 2142 3235 2153 3255
rect 2104 3223 2153 3235
rect 298 2988 347 2998
rect 298 2968 309 2988
rect 329 2968 347 2988
rect 298 2956 347 2968
rect 397 2992 441 2998
rect 397 2972 412 2992
rect 432 2972 441 2992
rect 397 2956 441 2972
rect 511 2988 560 2998
rect 511 2968 522 2988
rect 542 2968 560 2988
rect 511 2956 560 2968
rect 610 2992 654 2998
rect 610 2972 625 2992
rect 645 2972 654 2992
rect 610 2956 654 2972
rect 719 2988 768 2998
rect 719 2968 730 2988
rect 750 2968 768 2988
rect 719 2956 768 2968
rect 818 2992 862 2998
rect 818 2972 833 2992
rect 853 2972 862 2992
rect 818 2956 862 2972
rect 932 2992 976 2998
rect 932 2972 941 2992
rect 961 2972 976 2992
rect 932 2956 976 2972
rect 1026 2988 1075 2998
rect 1026 2968 1044 2988
rect 1064 2968 1075 2988
rect 1026 2956 1075 2968
rect 1236 2744 1285 2754
rect 1236 2724 1247 2744
rect 1267 2724 1285 2744
rect 1236 2712 1285 2724
rect 1335 2748 1379 2754
rect 1335 2728 1350 2748
rect 1370 2728 1379 2748
rect 1335 2712 1379 2728
rect 1449 2744 1498 2754
rect 1449 2724 1460 2744
rect 1480 2724 1498 2744
rect 1449 2712 1498 2724
rect 1548 2748 1592 2754
rect 1548 2728 1563 2748
rect 1583 2728 1592 2748
rect 1548 2712 1592 2728
rect 1657 2744 1706 2754
rect 1657 2724 1668 2744
rect 1688 2724 1706 2744
rect 1657 2712 1706 2724
rect 1756 2748 1800 2754
rect 1756 2728 1771 2748
rect 1791 2728 1800 2748
rect 1756 2712 1800 2728
rect 1870 2748 1914 2754
rect 1870 2728 1879 2748
rect 1899 2728 1914 2748
rect 1870 2712 1914 2728
rect 1964 2744 2013 2754
rect 1964 2724 1982 2744
rect 2002 2724 2013 2744
rect 1964 2712 2013 2724
rect 297 2434 346 2444
rect 297 2414 308 2434
rect 328 2414 346 2434
rect 297 2402 346 2414
rect 396 2438 440 2444
rect 396 2418 411 2438
rect 431 2418 440 2438
rect 396 2402 440 2418
rect 510 2434 559 2444
rect 510 2414 521 2434
rect 541 2414 559 2434
rect 510 2402 559 2414
rect 609 2438 653 2444
rect 609 2418 624 2438
rect 644 2418 653 2438
rect 609 2402 653 2418
rect 718 2434 767 2444
rect 718 2414 729 2434
rect 749 2414 767 2434
rect 718 2402 767 2414
rect 817 2438 861 2444
rect 817 2418 832 2438
rect 852 2418 861 2438
rect 817 2402 861 2418
rect 931 2438 975 2444
rect 931 2418 940 2438
rect 960 2418 975 2438
rect 931 2402 975 2418
rect 1025 2434 1074 2444
rect 1025 2414 1043 2434
rect 1063 2414 1074 2434
rect 1025 2402 1074 2414
rect 1346 2165 1395 2175
rect 1346 2145 1357 2165
rect 1377 2145 1395 2165
rect 1346 2133 1395 2145
rect 1445 2169 1489 2175
rect 1445 2149 1460 2169
rect 1480 2149 1489 2169
rect 1445 2133 1489 2149
rect 1559 2165 1608 2175
rect 1559 2145 1570 2165
rect 1590 2145 1608 2165
rect 1559 2133 1608 2145
rect 1658 2169 1702 2175
rect 1658 2149 1673 2169
rect 1693 2149 1702 2169
rect 1658 2133 1702 2149
rect 1767 2165 1816 2175
rect 1767 2145 1778 2165
rect 1798 2145 1816 2165
rect 1767 2133 1816 2145
rect 1866 2169 1910 2175
rect 1866 2149 1881 2169
rect 1901 2149 1910 2169
rect 1866 2133 1910 2149
rect 1980 2169 2024 2175
rect 1980 2149 1989 2169
rect 2009 2149 2024 2169
rect 1980 2133 2024 2149
rect 2074 2165 2123 2175
rect 2074 2145 2092 2165
rect 2112 2145 2123 2165
rect 2074 2133 2123 2145
rect 298 1885 347 1895
rect 298 1865 309 1885
rect 329 1865 347 1885
rect 298 1853 347 1865
rect 397 1889 441 1895
rect 397 1869 412 1889
rect 432 1869 441 1889
rect 397 1853 441 1869
rect 511 1885 560 1895
rect 511 1865 522 1885
rect 542 1865 560 1885
rect 511 1853 560 1865
rect 610 1889 654 1895
rect 610 1869 625 1889
rect 645 1869 654 1889
rect 610 1853 654 1869
rect 719 1885 768 1895
rect 719 1865 730 1885
rect 750 1865 768 1885
rect 719 1853 768 1865
rect 818 1889 862 1895
rect 818 1869 833 1889
rect 853 1869 862 1889
rect 818 1853 862 1869
rect 932 1889 976 1895
rect 932 1869 941 1889
rect 961 1869 976 1889
rect 932 1853 976 1869
rect 1026 1885 1075 1895
rect 1026 1865 1044 1885
rect 1064 1865 1075 1885
rect 1026 1853 1075 1865
rect 1236 1641 1285 1651
rect 1236 1621 1247 1641
rect 1267 1621 1285 1641
rect 1236 1609 1285 1621
rect 1335 1645 1379 1651
rect 1335 1625 1350 1645
rect 1370 1625 1379 1645
rect 1335 1609 1379 1625
rect 1449 1641 1498 1651
rect 1449 1621 1460 1641
rect 1480 1621 1498 1641
rect 1449 1609 1498 1621
rect 1548 1645 1592 1651
rect 1548 1625 1563 1645
rect 1583 1625 1592 1645
rect 1548 1609 1592 1625
rect 1657 1641 1706 1651
rect 1657 1621 1668 1641
rect 1688 1621 1706 1641
rect 1657 1609 1706 1621
rect 1756 1645 1800 1651
rect 1756 1625 1771 1645
rect 1791 1625 1800 1645
rect 1756 1609 1800 1625
rect 1870 1645 1914 1651
rect 1870 1625 1879 1645
rect 1899 1625 1914 1645
rect 1870 1609 1914 1625
rect 1964 1641 2013 1651
rect 1964 1621 1982 1641
rect 2002 1621 2013 1641
rect 1964 1609 2013 1621
rect 297 1331 346 1341
rect 297 1311 308 1331
rect 328 1311 346 1331
rect 297 1299 346 1311
rect 396 1335 440 1341
rect 396 1315 411 1335
rect 431 1315 440 1335
rect 396 1299 440 1315
rect 510 1331 559 1341
rect 510 1311 521 1331
rect 541 1311 559 1331
rect 510 1299 559 1311
rect 609 1335 653 1341
rect 609 1315 624 1335
rect 644 1315 653 1335
rect 609 1299 653 1315
rect 718 1331 767 1341
rect 718 1311 729 1331
rect 749 1311 767 1331
rect 718 1299 767 1311
rect 817 1335 861 1341
rect 817 1315 832 1335
rect 852 1315 861 1335
rect 817 1299 861 1315
rect 931 1335 975 1341
rect 931 1315 940 1335
rect 960 1315 975 1335
rect 931 1299 975 1315
rect 1025 1331 1074 1341
rect 1025 1311 1043 1331
rect 1063 1311 1074 1331
rect 1025 1299 1074 1311
rect 1377 1049 1426 1059
rect 1377 1029 1388 1049
rect 1408 1029 1426 1049
rect 1377 1017 1426 1029
rect 1476 1053 1520 1059
rect 1476 1033 1491 1053
rect 1511 1033 1520 1053
rect 1476 1017 1520 1033
rect 1590 1049 1639 1059
rect 1590 1029 1601 1049
rect 1621 1029 1639 1049
rect 1590 1017 1639 1029
rect 1689 1053 1733 1059
rect 1689 1033 1704 1053
rect 1724 1033 1733 1053
rect 1689 1017 1733 1033
rect 1798 1049 1847 1059
rect 1798 1029 1809 1049
rect 1829 1029 1847 1049
rect 1798 1017 1847 1029
rect 1897 1053 1941 1059
rect 1897 1033 1912 1053
rect 1932 1033 1941 1053
rect 1897 1017 1941 1033
rect 2011 1053 2055 1059
rect 2011 1033 2020 1053
rect 2040 1033 2055 1053
rect 2011 1017 2055 1033
rect 2105 1049 2154 1059
rect 2105 1029 2123 1049
rect 2143 1029 2154 1049
rect 2105 1017 2154 1029
rect 299 782 348 792
rect 299 762 310 782
rect 330 762 348 782
rect 299 750 348 762
rect 398 786 442 792
rect 398 766 413 786
rect 433 766 442 786
rect 398 750 442 766
rect 512 782 561 792
rect 512 762 523 782
rect 543 762 561 782
rect 512 750 561 762
rect 611 786 655 792
rect 611 766 626 786
rect 646 766 655 786
rect 611 750 655 766
rect 720 782 769 792
rect 720 762 731 782
rect 751 762 769 782
rect 720 750 769 762
rect 819 786 863 792
rect 819 766 834 786
rect 854 766 863 786
rect 819 750 863 766
rect 933 786 977 792
rect 933 766 942 786
rect 962 766 977 786
rect 933 750 977 766
rect 1027 782 1076 792
rect 1027 762 1045 782
rect 1065 762 1076 782
rect 1027 750 1076 762
rect 1237 538 1286 548
rect 1237 518 1248 538
rect 1268 518 1286 538
rect 1237 506 1286 518
rect 1336 542 1380 548
rect 1336 522 1351 542
rect 1371 522 1380 542
rect 1336 506 1380 522
rect 1450 538 1499 548
rect 1450 518 1461 538
rect 1481 518 1499 538
rect 1450 506 1499 518
rect 1549 542 1593 548
rect 1549 522 1564 542
rect 1584 522 1593 542
rect 1549 506 1593 522
rect 1658 538 1707 548
rect 1658 518 1669 538
rect 1689 518 1707 538
rect 1658 506 1707 518
rect 1757 542 1801 548
rect 1757 522 1772 542
rect 1792 522 1801 542
rect 1757 506 1801 522
rect 1871 542 1915 548
rect 1871 522 1880 542
rect 1900 522 1915 542
rect 1871 506 1915 522
rect 1965 538 2014 548
rect 1965 518 1983 538
rect 2003 518 2014 538
rect 1965 506 2014 518
rect 298 228 347 238
rect 298 208 309 228
rect 329 208 347 228
rect 298 196 347 208
rect 397 232 441 238
rect 397 212 412 232
rect 432 212 441 232
rect 397 196 441 212
rect 511 228 560 238
rect 511 208 522 228
rect 542 208 560 228
rect 511 196 560 208
rect 610 232 654 238
rect 610 212 625 232
rect 645 212 654 232
rect 610 196 654 212
rect 719 228 768 238
rect 719 208 730 228
rect 750 208 768 228
rect 719 196 768 208
rect 818 232 862 238
rect 818 212 833 232
rect 853 212 862 232
rect 818 196 862 212
rect 932 232 976 238
rect 932 212 941 232
rect 961 212 976 232
rect 932 196 976 212
rect 1026 228 1075 238
rect 1026 208 1044 228
rect 1064 208 1075 228
rect 1026 196 1075 208
rect 1346 -35 1395 -25
rect 1346 -55 1357 -35
rect 1377 -55 1395 -35
rect 1346 -67 1395 -55
rect 1445 -31 1489 -25
rect 1445 -51 1460 -31
rect 1480 -51 1489 -31
rect 1445 -67 1489 -51
rect 1559 -35 1608 -25
rect 1559 -55 1570 -35
rect 1590 -55 1608 -35
rect 1559 -67 1608 -55
rect 1658 -31 1702 -25
rect 1658 -51 1673 -31
rect 1693 -51 1702 -31
rect 1658 -67 1702 -51
rect 1767 -35 1816 -25
rect 1767 -55 1778 -35
rect 1798 -55 1816 -35
rect 1767 -67 1816 -55
rect 1866 -31 1910 -25
rect 1866 -51 1881 -31
rect 1901 -51 1910 -31
rect 1866 -67 1910 -51
rect 1980 -31 2024 -25
rect 1980 -51 1989 -31
rect 2009 -51 2024 -31
rect 1980 -67 2024 -51
rect 2074 -35 2123 -25
rect 2074 -55 2092 -35
rect 2112 -55 2123 -35
rect 2074 -67 2123 -55
rect 299 -321 348 -311
rect 299 -341 310 -321
rect 330 -341 348 -321
rect 299 -353 348 -341
rect 398 -317 442 -311
rect 398 -337 413 -317
rect 433 -337 442 -317
rect 398 -353 442 -337
rect 512 -321 561 -311
rect 512 -341 523 -321
rect 543 -341 561 -321
rect 512 -353 561 -341
rect 611 -317 655 -311
rect 611 -337 626 -317
rect 646 -337 655 -317
rect 611 -353 655 -337
rect 720 -321 769 -311
rect 720 -341 731 -321
rect 751 -341 769 -321
rect 720 -353 769 -341
rect 819 -317 863 -311
rect 819 -337 834 -317
rect 854 -337 863 -317
rect 819 -353 863 -337
rect 933 -317 977 -311
rect 933 -337 942 -317
rect 962 -337 977 -317
rect 933 -353 977 -337
rect 1027 -321 1076 -311
rect 1027 -341 1045 -321
rect 1065 -341 1076 -321
rect 1027 -353 1076 -341
rect 1237 -565 1286 -555
rect 1237 -585 1248 -565
rect 1268 -585 1286 -565
rect 1237 -597 1286 -585
rect 1336 -561 1380 -555
rect 1336 -581 1351 -561
rect 1371 -581 1380 -561
rect 1336 -597 1380 -581
rect 1450 -565 1499 -555
rect 1450 -585 1461 -565
rect 1481 -585 1499 -565
rect 1450 -597 1499 -585
rect 1549 -561 1593 -555
rect 1549 -581 1564 -561
rect 1584 -581 1593 -561
rect 1549 -597 1593 -581
rect 1658 -565 1707 -555
rect 1658 -585 1669 -565
rect 1689 -585 1707 -565
rect 1658 -597 1707 -585
rect 1757 -561 1801 -555
rect 1757 -581 1772 -561
rect 1792 -581 1801 -561
rect 1757 -597 1801 -581
rect 1871 -561 1915 -555
rect 1871 -581 1880 -561
rect 1900 -581 1915 -561
rect 1871 -597 1915 -581
rect 1965 -565 2014 -555
rect 1965 -585 1983 -565
rect 2003 -585 2014 -565
rect 1965 -597 2014 -585
rect 298 -875 347 -865
rect 298 -895 309 -875
rect 329 -895 347 -875
rect 298 -907 347 -895
rect 397 -871 441 -865
rect 397 -891 412 -871
rect 432 -891 441 -871
rect 397 -907 441 -891
rect 511 -875 560 -865
rect 511 -895 522 -875
rect 542 -895 560 -875
rect 511 -907 560 -895
rect 610 -871 654 -865
rect 610 -891 625 -871
rect 645 -891 654 -871
rect 610 -907 654 -891
rect 719 -875 768 -865
rect 719 -895 730 -875
rect 750 -895 768 -875
rect 719 -907 768 -895
rect 818 -871 862 -865
rect 818 -891 833 -871
rect 853 -891 862 -871
rect 818 -907 862 -891
rect 932 -871 976 -865
rect 932 -891 941 -871
rect 961 -891 976 -871
rect 932 -907 976 -891
rect 1026 -875 1075 -865
rect 1026 -895 1044 -875
rect 1064 -895 1075 -875
rect 1026 -907 1075 -895
rect 1378 -1157 1427 -1147
rect 1378 -1177 1389 -1157
rect 1409 -1177 1427 -1157
rect 1378 -1189 1427 -1177
rect 1477 -1153 1521 -1147
rect 1477 -1173 1492 -1153
rect 1512 -1173 1521 -1153
rect 1477 -1189 1521 -1173
rect 1591 -1157 1640 -1147
rect 1591 -1177 1602 -1157
rect 1622 -1177 1640 -1157
rect 1591 -1189 1640 -1177
rect 1690 -1153 1734 -1147
rect 1690 -1173 1705 -1153
rect 1725 -1173 1734 -1153
rect 1690 -1189 1734 -1173
rect 1799 -1157 1848 -1147
rect 1799 -1177 1810 -1157
rect 1830 -1177 1848 -1157
rect 1799 -1189 1848 -1177
rect 1898 -1153 1942 -1147
rect 1898 -1173 1913 -1153
rect 1933 -1173 1942 -1153
rect 1898 -1189 1942 -1173
rect 2012 -1153 2056 -1147
rect 2012 -1173 2021 -1153
rect 2041 -1173 2056 -1153
rect 2012 -1189 2056 -1173
rect 2106 -1157 2155 -1147
rect 2106 -1177 2124 -1157
rect 2144 -1177 2155 -1157
rect 2106 -1189 2155 -1177
rect 300 -1424 349 -1414
rect 300 -1444 311 -1424
rect 331 -1444 349 -1424
rect 300 -1456 349 -1444
rect 399 -1420 443 -1414
rect 399 -1440 414 -1420
rect 434 -1440 443 -1420
rect 399 -1456 443 -1440
rect 513 -1424 562 -1414
rect 513 -1444 524 -1424
rect 544 -1444 562 -1424
rect 513 -1456 562 -1444
rect 612 -1420 656 -1414
rect 612 -1440 627 -1420
rect 647 -1440 656 -1420
rect 612 -1456 656 -1440
rect 721 -1424 770 -1414
rect 721 -1444 732 -1424
rect 752 -1444 770 -1424
rect 721 -1456 770 -1444
rect 820 -1420 864 -1414
rect 820 -1440 835 -1420
rect 855 -1440 864 -1420
rect 820 -1456 864 -1440
rect 934 -1420 978 -1414
rect 934 -1440 943 -1420
rect 963 -1440 978 -1420
rect 934 -1456 978 -1440
rect 1028 -1424 1077 -1414
rect 1028 -1444 1046 -1424
rect 1066 -1444 1077 -1424
rect 1028 -1456 1077 -1444
rect 1238 -1668 1287 -1658
rect 1238 -1688 1249 -1668
rect 1269 -1688 1287 -1668
rect 1238 -1700 1287 -1688
rect 1337 -1664 1381 -1658
rect 1337 -1684 1352 -1664
rect 1372 -1684 1381 -1664
rect 1337 -1700 1381 -1684
rect 1451 -1668 1500 -1658
rect 1451 -1688 1462 -1668
rect 1482 -1688 1500 -1668
rect 1451 -1700 1500 -1688
rect 1550 -1664 1594 -1658
rect 1550 -1684 1565 -1664
rect 1585 -1684 1594 -1664
rect 1550 -1700 1594 -1684
rect 1659 -1668 1708 -1658
rect 1659 -1688 1670 -1668
rect 1690 -1688 1708 -1668
rect 1659 -1700 1708 -1688
rect 1758 -1664 1802 -1658
rect 1758 -1684 1773 -1664
rect 1793 -1684 1802 -1664
rect 1758 -1700 1802 -1684
rect 1872 -1664 1916 -1658
rect 1872 -1684 1881 -1664
rect 1901 -1684 1916 -1664
rect 1872 -1700 1916 -1684
rect 1966 -1668 2015 -1658
rect 1966 -1688 1984 -1668
rect 2004 -1688 2015 -1668
rect 1966 -1700 2015 -1688
rect 299 -1978 348 -1968
rect 299 -1998 310 -1978
rect 330 -1998 348 -1978
rect 299 -2010 348 -1998
rect 398 -1974 442 -1968
rect 398 -1994 413 -1974
rect 433 -1994 442 -1974
rect 398 -2010 442 -1994
rect 512 -1978 561 -1968
rect 512 -1998 523 -1978
rect 543 -1998 561 -1978
rect 512 -2010 561 -1998
rect 611 -1974 655 -1968
rect 611 -1994 626 -1974
rect 646 -1994 655 -1974
rect 611 -2010 655 -1994
rect 720 -1978 769 -1968
rect 720 -1998 731 -1978
rect 751 -1998 769 -1978
rect 720 -2010 769 -1998
rect 819 -1974 863 -1968
rect 819 -1994 834 -1974
rect 854 -1994 863 -1974
rect 819 -2010 863 -1994
rect 933 -1974 977 -1968
rect 933 -1994 942 -1974
rect 962 -1994 977 -1974
rect 933 -2010 977 -1994
rect 1027 -1978 1076 -1968
rect 1027 -1998 1045 -1978
rect 1065 -1998 1076 -1978
rect 1027 -2010 1076 -1998
rect 1348 -2247 1397 -2237
rect 1348 -2267 1359 -2247
rect 1379 -2267 1397 -2247
rect 1348 -2279 1397 -2267
rect 1447 -2243 1491 -2237
rect 1447 -2263 1462 -2243
rect 1482 -2263 1491 -2243
rect 1447 -2279 1491 -2263
rect 1561 -2247 1610 -2237
rect 1561 -2267 1572 -2247
rect 1592 -2267 1610 -2247
rect 1561 -2279 1610 -2267
rect 1660 -2243 1704 -2237
rect 1660 -2263 1675 -2243
rect 1695 -2263 1704 -2243
rect 1660 -2279 1704 -2263
rect 1769 -2247 1818 -2237
rect 1769 -2267 1780 -2247
rect 1800 -2267 1818 -2247
rect 1769 -2279 1818 -2267
rect 1868 -2243 1912 -2237
rect 1868 -2263 1883 -2243
rect 1903 -2263 1912 -2243
rect 1868 -2279 1912 -2263
rect 1982 -2243 2026 -2237
rect 1982 -2263 1991 -2243
rect 2011 -2263 2026 -2243
rect 1982 -2279 2026 -2263
rect 2076 -2247 2125 -2237
rect 2076 -2267 2094 -2247
rect 2114 -2267 2125 -2247
rect 2076 -2279 2125 -2267
rect 300 -2527 349 -2517
rect 300 -2547 311 -2527
rect 331 -2547 349 -2527
rect 300 -2559 349 -2547
rect 399 -2523 443 -2517
rect 399 -2543 414 -2523
rect 434 -2543 443 -2523
rect 399 -2559 443 -2543
rect 513 -2527 562 -2517
rect 513 -2547 524 -2527
rect 544 -2547 562 -2527
rect 513 -2559 562 -2547
rect 612 -2523 656 -2517
rect 612 -2543 627 -2523
rect 647 -2543 656 -2523
rect 612 -2559 656 -2543
rect 721 -2527 770 -2517
rect 721 -2547 732 -2527
rect 752 -2547 770 -2527
rect 721 -2559 770 -2547
rect 820 -2523 864 -2517
rect 820 -2543 835 -2523
rect 855 -2543 864 -2523
rect 820 -2559 864 -2543
rect 934 -2523 978 -2517
rect 934 -2543 943 -2523
rect 963 -2543 978 -2523
rect 934 -2559 978 -2543
rect 1028 -2527 1077 -2517
rect 1028 -2547 1046 -2527
rect 1066 -2547 1077 -2527
rect 1028 -2559 1077 -2547
rect 1238 -2771 1287 -2761
rect 1238 -2791 1249 -2771
rect 1269 -2791 1287 -2771
rect 1238 -2803 1287 -2791
rect 1337 -2767 1381 -2761
rect 1337 -2787 1352 -2767
rect 1372 -2787 1381 -2767
rect 1337 -2803 1381 -2787
rect 1451 -2771 1500 -2761
rect 1451 -2791 1462 -2771
rect 1482 -2791 1500 -2771
rect 1451 -2803 1500 -2791
rect 1550 -2767 1594 -2761
rect 1550 -2787 1565 -2767
rect 1585 -2787 1594 -2767
rect 1550 -2803 1594 -2787
rect 1659 -2771 1708 -2761
rect 1659 -2791 1670 -2771
rect 1690 -2791 1708 -2771
rect 1659 -2803 1708 -2791
rect 1758 -2767 1802 -2761
rect 1758 -2787 1773 -2767
rect 1793 -2787 1802 -2767
rect 1758 -2803 1802 -2787
rect 1872 -2767 1916 -2761
rect 1872 -2787 1881 -2767
rect 1901 -2787 1916 -2767
rect 1872 -2803 1916 -2787
rect 1966 -2771 2015 -2761
rect 1966 -2791 1984 -2771
rect 2004 -2791 2015 -2771
rect 1966 -2803 2015 -2791
rect 299 -3081 348 -3071
rect 299 -3101 310 -3081
rect 330 -3101 348 -3081
rect 299 -3113 348 -3101
rect 398 -3077 442 -3071
rect 398 -3097 413 -3077
rect 433 -3097 442 -3077
rect 398 -3113 442 -3097
rect 512 -3081 561 -3071
rect 512 -3101 523 -3081
rect 543 -3101 561 -3081
rect 512 -3113 561 -3101
rect 611 -3077 655 -3071
rect 611 -3097 626 -3077
rect 646 -3097 655 -3077
rect 611 -3113 655 -3097
rect 720 -3081 769 -3071
rect 720 -3101 731 -3081
rect 751 -3101 769 -3081
rect 720 -3113 769 -3101
rect 819 -3077 863 -3071
rect 819 -3097 834 -3077
rect 854 -3097 863 -3077
rect 819 -3113 863 -3097
rect 933 -3077 977 -3071
rect 933 -3097 942 -3077
rect 962 -3097 977 -3077
rect 933 -3113 977 -3097
rect 1027 -3081 1076 -3071
rect 1027 -3101 1045 -3081
rect 1065 -3101 1076 -3081
rect 1027 -3113 1076 -3101
rect 1379 -3363 1428 -3353
rect 1379 -3383 1390 -3363
rect 1410 -3383 1428 -3363
rect 1379 -3395 1428 -3383
rect 1478 -3359 1522 -3353
rect 1478 -3379 1493 -3359
rect 1513 -3379 1522 -3359
rect 1478 -3395 1522 -3379
rect 1592 -3363 1641 -3353
rect 1592 -3383 1603 -3363
rect 1623 -3383 1641 -3363
rect 1592 -3395 1641 -3383
rect 1691 -3359 1735 -3353
rect 1691 -3379 1706 -3359
rect 1726 -3379 1735 -3359
rect 1691 -3395 1735 -3379
rect 1800 -3363 1849 -3353
rect 1800 -3383 1811 -3363
rect 1831 -3383 1849 -3363
rect 1800 -3395 1849 -3383
rect 1899 -3359 1943 -3353
rect 1899 -3379 1914 -3359
rect 1934 -3379 1943 -3359
rect 1899 -3395 1943 -3379
rect 2013 -3359 2057 -3353
rect 2013 -3379 2022 -3359
rect 2042 -3379 2057 -3359
rect 2013 -3395 2057 -3379
rect 2107 -3363 2156 -3353
rect 2107 -3383 2125 -3363
rect 2145 -3383 2156 -3363
rect 2107 -3395 2156 -3383
rect 301 -3630 350 -3620
rect 301 -3650 312 -3630
rect 332 -3650 350 -3630
rect 301 -3662 350 -3650
rect 400 -3626 444 -3620
rect 400 -3646 415 -3626
rect 435 -3646 444 -3626
rect 400 -3662 444 -3646
rect 514 -3630 563 -3620
rect 514 -3650 525 -3630
rect 545 -3650 563 -3630
rect 514 -3662 563 -3650
rect 613 -3626 657 -3620
rect 613 -3646 628 -3626
rect 648 -3646 657 -3626
rect 613 -3662 657 -3646
rect 722 -3630 771 -3620
rect 722 -3650 733 -3630
rect 753 -3650 771 -3630
rect 722 -3662 771 -3650
rect 821 -3626 865 -3620
rect 821 -3646 836 -3626
rect 856 -3646 865 -3626
rect 821 -3662 865 -3646
rect 935 -3626 979 -3620
rect 935 -3646 944 -3626
rect 964 -3646 979 -3626
rect 935 -3662 979 -3646
rect 1029 -3630 1078 -3620
rect 1029 -3650 1047 -3630
rect 1067 -3650 1078 -3630
rect 1029 -3662 1078 -3650
rect 1239 -3874 1288 -3864
rect 1239 -3894 1250 -3874
rect 1270 -3894 1288 -3874
rect 1239 -3906 1288 -3894
rect 1338 -3870 1382 -3864
rect 1338 -3890 1353 -3870
rect 1373 -3890 1382 -3870
rect 1338 -3906 1382 -3890
rect 1452 -3874 1501 -3864
rect 1452 -3894 1463 -3874
rect 1483 -3894 1501 -3874
rect 1452 -3906 1501 -3894
rect 1551 -3870 1595 -3864
rect 1551 -3890 1566 -3870
rect 1586 -3890 1595 -3870
rect 1551 -3906 1595 -3890
rect 1660 -3874 1709 -3864
rect 1660 -3894 1671 -3874
rect 1691 -3894 1709 -3874
rect 1660 -3906 1709 -3894
rect 1759 -3870 1803 -3864
rect 1759 -3890 1774 -3870
rect 1794 -3890 1803 -3870
rect 1759 -3906 1803 -3890
rect 1873 -3870 1917 -3864
rect 1873 -3890 1882 -3870
rect 1902 -3890 1917 -3870
rect 1873 -3906 1917 -3890
rect 1967 -3874 2016 -3864
rect 1967 -3894 1985 -3874
rect 2005 -3894 2016 -3874
rect 1967 -3906 2016 -3894
rect 300 -4184 349 -4174
rect 300 -4204 311 -4184
rect 331 -4204 349 -4184
rect 300 -4216 349 -4204
rect 399 -4180 443 -4174
rect 399 -4200 414 -4180
rect 434 -4200 443 -4180
rect 399 -4216 443 -4200
rect 513 -4184 562 -4174
rect 513 -4204 524 -4184
rect 544 -4204 562 -4184
rect 513 -4216 562 -4204
rect 612 -4180 656 -4174
rect 612 -4200 627 -4180
rect 647 -4200 656 -4180
rect 612 -4216 656 -4200
rect 721 -4184 770 -4174
rect 721 -4204 732 -4184
rect 752 -4204 770 -4184
rect 721 -4216 770 -4204
rect 820 -4180 864 -4174
rect 820 -4200 835 -4180
rect 855 -4200 864 -4180
rect 820 -4216 864 -4200
rect 934 -4180 978 -4174
rect 934 -4200 943 -4180
rect 963 -4200 978 -4180
rect 934 -4216 978 -4200
rect 1028 -4184 1077 -4174
rect 1028 -4204 1046 -4184
rect 1066 -4204 1077 -4184
rect 1028 -4216 1077 -4204
<< pdiff >>
rect 302 4240 346 4278
rect 302 4220 314 4240
rect 334 4220 346 4240
rect 302 4178 346 4220
rect 396 4240 438 4278
rect 396 4220 410 4240
rect 430 4220 438 4240
rect 396 4178 438 4220
rect 515 4240 559 4278
rect 515 4220 527 4240
rect 547 4220 559 4240
rect 515 4178 559 4220
rect 609 4240 651 4278
rect 609 4220 623 4240
rect 643 4220 651 4240
rect 609 4178 651 4220
rect 723 4240 767 4278
rect 723 4220 735 4240
rect 755 4220 767 4240
rect 723 4178 767 4220
rect 817 4240 859 4278
rect 817 4220 831 4240
rect 851 4220 859 4240
rect 817 4178 859 4220
rect 933 4240 975 4278
rect 933 4220 941 4240
rect 961 4220 975 4240
rect 933 4178 975 4220
rect 1025 4247 1070 4278
rect 1025 4240 1069 4247
rect 1025 4220 1037 4240
rect 1057 4220 1069 4240
rect 1025 4178 1069 4220
rect 1240 3996 1284 4034
rect 1240 3976 1252 3996
rect 1272 3976 1284 3996
rect 1240 3934 1284 3976
rect 1334 3996 1376 4034
rect 1334 3976 1348 3996
rect 1368 3976 1376 3996
rect 1334 3934 1376 3976
rect 1453 3996 1497 4034
rect 1453 3976 1465 3996
rect 1485 3976 1497 3996
rect 1453 3934 1497 3976
rect 1547 3996 1589 4034
rect 1547 3976 1561 3996
rect 1581 3976 1589 3996
rect 1547 3934 1589 3976
rect 1661 3996 1705 4034
rect 1661 3976 1673 3996
rect 1693 3976 1705 3996
rect 1661 3934 1705 3976
rect 1755 3996 1797 4034
rect 1755 3976 1769 3996
rect 1789 3976 1797 3996
rect 1755 3934 1797 3976
rect 1871 3996 1913 4034
rect 1871 3976 1879 3996
rect 1899 3976 1913 3996
rect 1871 3934 1913 3976
rect 1963 4003 2008 4034
rect 1963 3996 2007 4003
rect 1963 3976 1975 3996
rect 1995 3976 2007 3996
rect 1963 3934 2007 3976
rect 301 3686 345 3724
rect 301 3666 313 3686
rect 333 3666 345 3686
rect 301 3624 345 3666
rect 395 3686 437 3724
rect 395 3666 409 3686
rect 429 3666 437 3686
rect 395 3624 437 3666
rect 514 3686 558 3724
rect 514 3666 526 3686
rect 546 3666 558 3686
rect 514 3624 558 3666
rect 608 3686 650 3724
rect 608 3666 622 3686
rect 642 3666 650 3686
rect 608 3624 650 3666
rect 722 3686 766 3724
rect 722 3666 734 3686
rect 754 3666 766 3686
rect 722 3624 766 3666
rect 816 3686 858 3724
rect 816 3666 830 3686
rect 850 3666 858 3686
rect 816 3624 858 3666
rect 932 3686 974 3724
rect 932 3666 940 3686
rect 960 3666 974 3686
rect 932 3624 974 3666
rect 1024 3693 1069 3724
rect 1024 3686 1068 3693
rect 1024 3666 1036 3686
rect 1056 3666 1068 3686
rect 1024 3624 1068 3666
rect 1381 3404 1425 3442
rect 1381 3384 1393 3404
rect 1413 3384 1425 3404
rect 1381 3342 1425 3384
rect 1475 3404 1517 3442
rect 1475 3384 1489 3404
rect 1509 3384 1517 3404
rect 1475 3342 1517 3384
rect 1594 3404 1638 3442
rect 1594 3384 1606 3404
rect 1626 3384 1638 3404
rect 1594 3342 1638 3384
rect 1688 3404 1730 3442
rect 1688 3384 1702 3404
rect 1722 3384 1730 3404
rect 1688 3342 1730 3384
rect 1802 3404 1846 3442
rect 1802 3384 1814 3404
rect 1834 3384 1846 3404
rect 1802 3342 1846 3384
rect 1896 3404 1938 3442
rect 1896 3384 1910 3404
rect 1930 3384 1938 3404
rect 1896 3342 1938 3384
rect 2012 3404 2054 3442
rect 2012 3384 2020 3404
rect 2040 3384 2054 3404
rect 2012 3342 2054 3384
rect 2104 3411 2149 3442
rect 2104 3404 2148 3411
rect 2104 3384 2116 3404
rect 2136 3384 2148 3404
rect 2104 3342 2148 3384
rect 303 3137 347 3175
rect 303 3117 315 3137
rect 335 3117 347 3137
rect 303 3075 347 3117
rect 397 3137 439 3175
rect 397 3117 411 3137
rect 431 3117 439 3137
rect 397 3075 439 3117
rect 516 3137 560 3175
rect 516 3117 528 3137
rect 548 3117 560 3137
rect 516 3075 560 3117
rect 610 3137 652 3175
rect 610 3117 624 3137
rect 644 3117 652 3137
rect 610 3075 652 3117
rect 724 3137 768 3175
rect 724 3117 736 3137
rect 756 3117 768 3137
rect 724 3075 768 3117
rect 818 3137 860 3175
rect 818 3117 832 3137
rect 852 3117 860 3137
rect 818 3075 860 3117
rect 934 3137 976 3175
rect 934 3117 942 3137
rect 962 3117 976 3137
rect 934 3075 976 3117
rect 1026 3144 1071 3175
rect 1026 3137 1070 3144
rect 1026 3117 1038 3137
rect 1058 3117 1070 3137
rect 1026 3075 1070 3117
rect 1241 2893 1285 2931
rect 1241 2873 1253 2893
rect 1273 2873 1285 2893
rect 1241 2831 1285 2873
rect 1335 2893 1377 2931
rect 1335 2873 1349 2893
rect 1369 2873 1377 2893
rect 1335 2831 1377 2873
rect 1454 2893 1498 2931
rect 1454 2873 1466 2893
rect 1486 2873 1498 2893
rect 1454 2831 1498 2873
rect 1548 2893 1590 2931
rect 1548 2873 1562 2893
rect 1582 2873 1590 2893
rect 1548 2831 1590 2873
rect 1662 2893 1706 2931
rect 1662 2873 1674 2893
rect 1694 2873 1706 2893
rect 1662 2831 1706 2873
rect 1756 2893 1798 2931
rect 1756 2873 1770 2893
rect 1790 2873 1798 2893
rect 1756 2831 1798 2873
rect 1872 2893 1914 2931
rect 1872 2873 1880 2893
rect 1900 2873 1914 2893
rect 1872 2831 1914 2873
rect 1964 2900 2009 2931
rect 1964 2893 2008 2900
rect 1964 2873 1976 2893
rect 1996 2873 2008 2893
rect 1964 2831 2008 2873
rect 302 2583 346 2621
rect 302 2563 314 2583
rect 334 2563 346 2583
rect 302 2521 346 2563
rect 396 2583 438 2621
rect 396 2563 410 2583
rect 430 2563 438 2583
rect 396 2521 438 2563
rect 515 2583 559 2621
rect 515 2563 527 2583
rect 547 2563 559 2583
rect 515 2521 559 2563
rect 609 2583 651 2621
rect 609 2563 623 2583
rect 643 2563 651 2583
rect 609 2521 651 2563
rect 723 2583 767 2621
rect 723 2563 735 2583
rect 755 2563 767 2583
rect 723 2521 767 2563
rect 817 2583 859 2621
rect 817 2563 831 2583
rect 851 2563 859 2583
rect 817 2521 859 2563
rect 933 2583 975 2621
rect 933 2563 941 2583
rect 961 2563 975 2583
rect 933 2521 975 2563
rect 1025 2590 1070 2621
rect 1025 2583 1069 2590
rect 1025 2563 1037 2583
rect 1057 2563 1069 2583
rect 1025 2521 1069 2563
rect 1351 2314 1395 2352
rect 1351 2294 1363 2314
rect 1383 2294 1395 2314
rect 1351 2252 1395 2294
rect 1445 2314 1487 2352
rect 1445 2294 1459 2314
rect 1479 2294 1487 2314
rect 1445 2252 1487 2294
rect 1564 2314 1608 2352
rect 1564 2294 1576 2314
rect 1596 2294 1608 2314
rect 1564 2252 1608 2294
rect 1658 2314 1700 2352
rect 1658 2294 1672 2314
rect 1692 2294 1700 2314
rect 1658 2252 1700 2294
rect 1772 2314 1816 2352
rect 1772 2294 1784 2314
rect 1804 2294 1816 2314
rect 1772 2252 1816 2294
rect 1866 2314 1908 2352
rect 1866 2294 1880 2314
rect 1900 2294 1908 2314
rect 1866 2252 1908 2294
rect 1982 2314 2024 2352
rect 1982 2294 1990 2314
rect 2010 2294 2024 2314
rect 1982 2252 2024 2294
rect 2074 2321 2119 2352
rect 2074 2314 2118 2321
rect 2074 2294 2086 2314
rect 2106 2294 2118 2314
rect 2074 2252 2118 2294
rect 303 2034 347 2072
rect 303 2014 315 2034
rect 335 2014 347 2034
rect 303 1972 347 2014
rect 397 2034 439 2072
rect 397 2014 411 2034
rect 431 2014 439 2034
rect 397 1972 439 2014
rect 516 2034 560 2072
rect 516 2014 528 2034
rect 548 2014 560 2034
rect 516 1972 560 2014
rect 610 2034 652 2072
rect 610 2014 624 2034
rect 644 2014 652 2034
rect 610 1972 652 2014
rect 724 2034 768 2072
rect 724 2014 736 2034
rect 756 2014 768 2034
rect 724 1972 768 2014
rect 818 2034 860 2072
rect 818 2014 832 2034
rect 852 2014 860 2034
rect 818 1972 860 2014
rect 934 2034 976 2072
rect 934 2014 942 2034
rect 962 2014 976 2034
rect 934 1972 976 2014
rect 1026 2041 1071 2072
rect 1026 2034 1070 2041
rect 1026 2014 1038 2034
rect 1058 2014 1070 2034
rect 1026 1972 1070 2014
rect 1241 1790 1285 1828
rect 1241 1770 1253 1790
rect 1273 1770 1285 1790
rect 1241 1728 1285 1770
rect 1335 1790 1377 1828
rect 1335 1770 1349 1790
rect 1369 1770 1377 1790
rect 1335 1728 1377 1770
rect 1454 1790 1498 1828
rect 1454 1770 1466 1790
rect 1486 1770 1498 1790
rect 1454 1728 1498 1770
rect 1548 1790 1590 1828
rect 1548 1770 1562 1790
rect 1582 1770 1590 1790
rect 1548 1728 1590 1770
rect 1662 1790 1706 1828
rect 1662 1770 1674 1790
rect 1694 1770 1706 1790
rect 1662 1728 1706 1770
rect 1756 1790 1798 1828
rect 1756 1770 1770 1790
rect 1790 1770 1798 1790
rect 1756 1728 1798 1770
rect 1872 1790 1914 1828
rect 1872 1770 1880 1790
rect 1900 1770 1914 1790
rect 1872 1728 1914 1770
rect 1964 1797 2009 1828
rect 1964 1790 2008 1797
rect 1964 1770 1976 1790
rect 1996 1770 2008 1790
rect 1964 1728 2008 1770
rect 302 1480 346 1518
rect 302 1460 314 1480
rect 334 1460 346 1480
rect 302 1418 346 1460
rect 396 1480 438 1518
rect 396 1460 410 1480
rect 430 1460 438 1480
rect 396 1418 438 1460
rect 515 1480 559 1518
rect 515 1460 527 1480
rect 547 1460 559 1480
rect 515 1418 559 1460
rect 609 1480 651 1518
rect 609 1460 623 1480
rect 643 1460 651 1480
rect 609 1418 651 1460
rect 723 1480 767 1518
rect 723 1460 735 1480
rect 755 1460 767 1480
rect 723 1418 767 1460
rect 817 1480 859 1518
rect 817 1460 831 1480
rect 851 1460 859 1480
rect 817 1418 859 1460
rect 933 1480 975 1518
rect 933 1460 941 1480
rect 961 1460 975 1480
rect 933 1418 975 1460
rect 1025 1487 1070 1518
rect 1025 1480 1069 1487
rect 1025 1460 1037 1480
rect 1057 1460 1069 1480
rect 1025 1418 1069 1460
rect 1382 1198 1426 1236
rect 1382 1178 1394 1198
rect 1414 1178 1426 1198
rect 1382 1136 1426 1178
rect 1476 1198 1518 1236
rect 1476 1178 1490 1198
rect 1510 1178 1518 1198
rect 1476 1136 1518 1178
rect 1595 1198 1639 1236
rect 1595 1178 1607 1198
rect 1627 1178 1639 1198
rect 1595 1136 1639 1178
rect 1689 1198 1731 1236
rect 1689 1178 1703 1198
rect 1723 1178 1731 1198
rect 1689 1136 1731 1178
rect 1803 1198 1847 1236
rect 1803 1178 1815 1198
rect 1835 1178 1847 1198
rect 1803 1136 1847 1178
rect 1897 1198 1939 1236
rect 1897 1178 1911 1198
rect 1931 1178 1939 1198
rect 1897 1136 1939 1178
rect 2013 1198 2055 1236
rect 2013 1178 2021 1198
rect 2041 1178 2055 1198
rect 2013 1136 2055 1178
rect 2105 1205 2150 1236
rect 2105 1198 2149 1205
rect 2105 1178 2117 1198
rect 2137 1178 2149 1198
rect 2105 1136 2149 1178
rect 304 931 348 969
rect 304 911 316 931
rect 336 911 348 931
rect 304 869 348 911
rect 398 931 440 969
rect 398 911 412 931
rect 432 911 440 931
rect 398 869 440 911
rect 517 931 561 969
rect 517 911 529 931
rect 549 911 561 931
rect 517 869 561 911
rect 611 931 653 969
rect 611 911 625 931
rect 645 911 653 931
rect 611 869 653 911
rect 725 931 769 969
rect 725 911 737 931
rect 757 911 769 931
rect 725 869 769 911
rect 819 931 861 969
rect 819 911 833 931
rect 853 911 861 931
rect 819 869 861 911
rect 935 931 977 969
rect 935 911 943 931
rect 963 911 977 931
rect 935 869 977 911
rect 1027 938 1072 969
rect 1027 931 1071 938
rect 1027 911 1039 931
rect 1059 911 1071 931
rect 1027 869 1071 911
rect 1242 687 1286 725
rect 1242 667 1254 687
rect 1274 667 1286 687
rect 1242 625 1286 667
rect 1336 687 1378 725
rect 1336 667 1350 687
rect 1370 667 1378 687
rect 1336 625 1378 667
rect 1455 687 1499 725
rect 1455 667 1467 687
rect 1487 667 1499 687
rect 1455 625 1499 667
rect 1549 687 1591 725
rect 1549 667 1563 687
rect 1583 667 1591 687
rect 1549 625 1591 667
rect 1663 687 1707 725
rect 1663 667 1675 687
rect 1695 667 1707 687
rect 1663 625 1707 667
rect 1757 687 1799 725
rect 1757 667 1771 687
rect 1791 667 1799 687
rect 1757 625 1799 667
rect 1873 687 1915 725
rect 1873 667 1881 687
rect 1901 667 1915 687
rect 1873 625 1915 667
rect 1965 694 2010 725
rect 1965 687 2009 694
rect 1965 667 1977 687
rect 1997 667 2009 687
rect 1965 625 2009 667
rect 303 377 347 415
rect 303 357 315 377
rect 335 357 347 377
rect 303 315 347 357
rect 397 377 439 415
rect 397 357 411 377
rect 431 357 439 377
rect 397 315 439 357
rect 516 377 560 415
rect 516 357 528 377
rect 548 357 560 377
rect 516 315 560 357
rect 610 377 652 415
rect 610 357 624 377
rect 644 357 652 377
rect 610 315 652 357
rect 724 377 768 415
rect 724 357 736 377
rect 756 357 768 377
rect 724 315 768 357
rect 818 377 860 415
rect 818 357 832 377
rect 852 357 860 377
rect 818 315 860 357
rect 934 377 976 415
rect 934 357 942 377
rect 962 357 976 377
rect 934 315 976 357
rect 1026 384 1071 415
rect 1026 377 1070 384
rect 1026 357 1038 377
rect 1058 357 1070 377
rect 1026 315 1070 357
rect 1351 114 1395 152
rect 1351 94 1363 114
rect 1383 94 1395 114
rect 1351 52 1395 94
rect 1445 114 1487 152
rect 1445 94 1459 114
rect 1479 94 1487 114
rect 1445 52 1487 94
rect 1564 114 1608 152
rect 1564 94 1576 114
rect 1596 94 1608 114
rect 1564 52 1608 94
rect 1658 114 1700 152
rect 1658 94 1672 114
rect 1692 94 1700 114
rect 1658 52 1700 94
rect 1772 114 1816 152
rect 1772 94 1784 114
rect 1804 94 1816 114
rect 1772 52 1816 94
rect 1866 114 1908 152
rect 1866 94 1880 114
rect 1900 94 1908 114
rect 1866 52 1908 94
rect 1982 114 2024 152
rect 1982 94 1990 114
rect 2010 94 2024 114
rect 1982 52 2024 94
rect 2074 121 2119 152
rect 2074 114 2118 121
rect 2074 94 2086 114
rect 2106 94 2118 114
rect 2074 52 2118 94
rect 304 -172 348 -134
rect 304 -192 316 -172
rect 336 -192 348 -172
rect 304 -234 348 -192
rect 398 -172 440 -134
rect 398 -192 412 -172
rect 432 -192 440 -172
rect 398 -234 440 -192
rect 517 -172 561 -134
rect 517 -192 529 -172
rect 549 -192 561 -172
rect 517 -234 561 -192
rect 611 -172 653 -134
rect 611 -192 625 -172
rect 645 -192 653 -172
rect 611 -234 653 -192
rect 725 -172 769 -134
rect 725 -192 737 -172
rect 757 -192 769 -172
rect 725 -234 769 -192
rect 819 -172 861 -134
rect 819 -192 833 -172
rect 853 -192 861 -172
rect 819 -234 861 -192
rect 935 -172 977 -134
rect 935 -192 943 -172
rect 963 -192 977 -172
rect 935 -234 977 -192
rect 1027 -165 1072 -134
rect 1027 -172 1071 -165
rect 1027 -192 1039 -172
rect 1059 -192 1071 -172
rect 1027 -234 1071 -192
rect 1242 -416 1286 -378
rect 1242 -436 1254 -416
rect 1274 -436 1286 -416
rect 1242 -478 1286 -436
rect 1336 -416 1378 -378
rect 1336 -436 1350 -416
rect 1370 -436 1378 -416
rect 1336 -478 1378 -436
rect 1455 -416 1499 -378
rect 1455 -436 1467 -416
rect 1487 -436 1499 -416
rect 1455 -478 1499 -436
rect 1549 -416 1591 -378
rect 1549 -436 1563 -416
rect 1583 -436 1591 -416
rect 1549 -478 1591 -436
rect 1663 -416 1707 -378
rect 1663 -436 1675 -416
rect 1695 -436 1707 -416
rect 1663 -478 1707 -436
rect 1757 -416 1799 -378
rect 1757 -436 1771 -416
rect 1791 -436 1799 -416
rect 1757 -478 1799 -436
rect 1873 -416 1915 -378
rect 1873 -436 1881 -416
rect 1901 -436 1915 -416
rect 1873 -478 1915 -436
rect 1965 -409 2010 -378
rect 1965 -416 2009 -409
rect 1965 -436 1977 -416
rect 1997 -436 2009 -416
rect 1965 -478 2009 -436
rect 303 -726 347 -688
rect 303 -746 315 -726
rect 335 -746 347 -726
rect 303 -788 347 -746
rect 397 -726 439 -688
rect 397 -746 411 -726
rect 431 -746 439 -726
rect 397 -788 439 -746
rect 516 -726 560 -688
rect 516 -746 528 -726
rect 548 -746 560 -726
rect 516 -788 560 -746
rect 610 -726 652 -688
rect 610 -746 624 -726
rect 644 -746 652 -726
rect 610 -788 652 -746
rect 724 -726 768 -688
rect 724 -746 736 -726
rect 756 -746 768 -726
rect 724 -788 768 -746
rect 818 -726 860 -688
rect 818 -746 832 -726
rect 852 -746 860 -726
rect 818 -788 860 -746
rect 934 -726 976 -688
rect 934 -746 942 -726
rect 962 -746 976 -726
rect 934 -788 976 -746
rect 1026 -719 1071 -688
rect 1026 -726 1070 -719
rect 1026 -746 1038 -726
rect 1058 -746 1070 -726
rect 1026 -788 1070 -746
rect 1383 -1008 1427 -970
rect 1383 -1028 1395 -1008
rect 1415 -1028 1427 -1008
rect 1383 -1070 1427 -1028
rect 1477 -1008 1519 -970
rect 1477 -1028 1491 -1008
rect 1511 -1028 1519 -1008
rect 1477 -1070 1519 -1028
rect 1596 -1008 1640 -970
rect 1596 -1028 1608 -1008
rect 1628 -1028 1640 -1008
rect 1596 -1070 1640 -1028
rect 1690 -1008 1732 -970
rect 1690 -1028 1704 -1008
rect 1724 -1028 1732 -1008
rect 1690 -1070 1732 -1028
rect 1804 -1008 1848 -970
rect 1804 -1028 1816 -1008
rect 1836 -1028 1848 -1008
rect 1804 -1070 1848 -1028
rect 1898 -1008 1940 -970
rect 1898 -1028 1912 -1008
rect 1932 -1028 1940 -1008
rect 1898 -1070 1940 -1028
rect 2014 -1008 2056 -970
rect 2014 -1028 2022 -1008
rect 2042 -1028 2056 -1008
rect 2014 -1070 2056 -1028
rect 2106 -1001 2151 -970
rect 2106 -1008 2150 -1001
rect 2106 -1028 2118 -1008
rect 2138 -1028 2150 -1008
rect 2106 -1070 2150 -1028
rect 305 -1275 349 -1237
rect 305 -1295 317 -1275
rect 337 -1295 349 -1275
rect 305 -1337 349 -1295
rect 399 -1275 441 -1237
rect 399 -1295 413 -1275
rect 433 -1295 441 -1275
rect 399 -1337 441 -1295
rect 518 -1275 562 -1237
rect 518 -1295 530 -1275
rect 550 -1295 562 -1275
rect 518 -1337 562 -1295
rect 612 -1275 654 -1237
rect 612 -1295 626 -1275
rect 646 -1295 654 -1275
rect 612 -1337 654 -1295
rect 726 -1275 770 -1237
rect 726 -1295 738 -1275
rect 758 -1295 770 -1275
rect 726 -1337 770 -1295
rect 820 -1275 862 -1237
rect 820 -1295 834 -1275
rect 854 -1295 862 -1275
rect 820 -1337 862 -1295
rect 936 -1275 978 -1237
rect 936 -1295 944 -1275
rect 964 -1295 978 -1275
rect 936 -1337 978 -1295
rect 1028 -1268 1073 -1237
rect 1028 -1275 1072 -1268
rect 1028 -1295 1040 -1275
rect 1060 -1295 1072 -1275
rect 1028 -1337 1072 -1295
rect 1243 -1519 1287 -1481
rect 1243 -1539 1255 -1519
rect 1275 -1539 1287 -1519
rect 1243 -1581 1287 -1539
rect 1337 -1519 1379 -1481
rect 1337 -1539 1351 -1519
rect 1371 -1539 1379 -1519
rect 1337 -1581 1379 -1539
rect 1456 -1519 1500 -1481
rect 1456 -1539 1468 -1519
rect 1488 -1539 1500 -1519
rect 1456 -1581 1500 -1539
rect 1550 -1519 1592 -1481
rect 1550 -1539 1564 -1519
rect 1584 -1539 1592 -1519
rect 1550 -1581 1592 -1539
rect 1664 -1519 1708 -1481
rect 1664 -1539 1676 -1519
rect 1696 -1539 1708 -1519
rect 1664 -1581 1708 -1539
rect 1758 -1519 1800 -1481
rect 1758 -1539 1772 -1519
rect 1792 -1539 1800 -1519
rect 1758 -1581 1800 -1539
rect 1874 -1519 1916 -1481
rect 1874 -1539 1882 -1519
rect 1902 -1539 1916 -1519
rect 1874 -1581 1916 -1539
rect 1966 -1512 2011 -1481
rect 1966 -1519 2010 -1512
rect 1966 -1539 1978 -1519
rect 1998 -1539 2010 -1519
rect 1966 -1581 2010 -1539
rect 304 -1829 348 -1791
rect 304 -1849 316 -1829
rect 336 -1849 348 -1829
rect 304 -1891 348 -1849
rect 398 -1829 440 -1791
rect 398 -1849 412 -1829
rect 432 -1849 440 -1829
rect 398 -1891 440 -1849
rect 517 -1829 561 -1791
rect 517 -1849 529 -1829
rect 549 -1849 561 -1829
rect 517 -1891 561 -1849
rect 611 -1829 653 -1791
rect 611 -1849 625 -1829
rect 645 -1849 653 -1829
rect 611 -1891 653 -1849
rect 725 -1829 769 -1791
rect 725 -1849 737 -1829
rect 757 -1849 769 -1829
rect 725 -1891 769 -1849
rect 819 -1829 861 -1791
rect 819 -1849 833 -1829
rect 853 -1849 861 -1829
rect 819 -1891 861 -1849
rect 935 -1829 977 -1791
rect 935 -1849 943 -1829
rect 963 -1849 977 -1829
rect 935 -1891 977 -1849
rect 1027 -1822 1072 -1791
rect 1027 -1829 1071 -1822
rect 1027 -1849 1039 -1829
rect 1059 -1849 1071 -1829
rect 1027 -1891 1071 -1849
rect 1353 -2098 1397 -2060
rect 1353 -2118 1365 -2098
rect 1385 -2118 1397 -2098
rect 1353 -2160 1397 -2118
rect 1447 -2098 1489 -2060
rect 1447 -2118 1461 -2098
rect 1481 -2118 1489 -2098
rect 1447 -2160 1489 -2118
rect 1566 -2098 1610 -2060
rect 1566 -2118 1578 -2098
rect 1598 -2118 1610 -2098
rect 1566 -2160 1610 -2118
rect 1660 -2098 1702 -2060
rect 1660 -2118 1674 -2098
rect 1694 -2118 1702 -2098
rect 1660 -2160 1702 -2118
rect 1774 -2098 1818 -2060
rect 1774 -2118 1786 -2098
rect 1806 -2118 1818 -2098
rect 1774 -2160 1818 -2118
rect 1868 -2098 1910 -2060
rect 1868 -2118 1882 -2098
rect 1902 -2118 1910 -2098
rect 1868 -2160 1910 -2118
rect 1984 -2098 2026 -2060
rect 1984 -2118 1992 -2098
rect 2012 -2118 2026 -2098
rect 1984 -2160 2026 -2118
rect 2076 -2091 2121 -2060
rect 2076 -2098 2120 -2091
rect 2076 -2118 2088 -2098
rect 2108 -2118 2120 -2098
rect 2076 -2160 2120 -2118
rect 305 -2378 349 -2340
rect 305 -2398 317 -2378
rect 337 -2398 349 -2378
rect 305 -2440 349 -2398
rect 399 -2378 441 -2340
rect 399 -2398 413 -2378
rect 433 -2398 441 -2378
rect 399 -2440 441 -2398
rect 518 -2378 562 -2340
rect 518 -2398 530 -2378
rect 550 -2398 562 -2378
rect 518 -2440 562 -2398
rect 612 -2378 654 -2340
rect 612 -2398 626 -2378
rect 646 -2398 654 -2378
rect 612 -2440 654 -2398
rect 726 -2378 770 -2340
rect 726 -2398 738 -2378
rect 758 -2398 770 -2378
rect 726 -2440 770 -2398
rect 820 -2378 862 -2340
rect 820 -2398 834 -2378
rect 854 -2398 862 -2378
rect 820 -2440 862 -2398
rect 936 -2378 978 -2340
rect 936 -2398 944 -2378
rect 964 -2398 978 -2378
rect 936 -2440 978 -2398
rect 1028 -2371 1073 -2340
rect 1028 -2378 1072 -2371
rect 1028 -2398 1040 -2378
rect 1060 -2398 1072 -2378
rect 1028 -2440 1072 -2398
rect 1243 -2622 1287 -2584
rect 1243 -2642 1255 -2622
rect 1275 -2642 1287 -2622
rect 1243 -2684 1287 -2642
rect 1337 -2622 1379 -2584
rect 1337 -2642 1351 -2622
rect 1371 -2642 1379 -2622
rect 1337 -2684 1379 -2642
rect 1456 -2622 1500 -2584
rect 1456 -2642 1468 -2622
rect 1488 -2642 1500 -2622
rect 1456 -2684 1500 -2642
rect 1550 -2622 1592 -2584
rect 1550 -2642 1564 -2622
rect 1584 -2642 1592 -2622
rect 1550 -2684 1592 -2642
rect 1664 -2622 1708 -2584
rect 1664 -2642 1676 -2622
rect 1696 -2642 1708 -2622
rect 1664 -2684 1708 -2642
rect 1758 -2622 1800 -2584
rect 1758 -2642 1772 -2622
rect 1792 -2642 1800 -2622
rect 1758 -2684 1800 -2642
rect 1874 -2622 1916 -2584
rect 1874 -2642 1882 -2622
rect 1902 -2642 1916 -2622
rect 1874 -2684 1916 -2642
rect 1966 -2615 2011 -2584
rect 1966 -2622 2010 -2615
rect 1966 -2642 1978 -2622
rect 1998 -2642 2010 -2622
rect 1966 -2684 2010 -2642
rect 304 -2932 348 -2894
rect 304 -2952 316 -2932
rect 336 -2952 348 -2932
rect 304 -2994 348 -2952
rect 398 -2932 440 -2894
rect 398 -2952 412 -2932
rect 432 -2952 440 -2932
rect 398 -2994 440 -2952
rect 517 -2932 561 -2894
rect 517 -2952 529 -2932
rect 549 -2952 561 -2932
rect 517 -2994 561 -2952
rect 611 -2932 653 -2894
rect 611 -2952 625 -2932
rect 645 -2952 653 -2932
rect 611 -2994 653 -2952
rect 725 -2932 769 -2894
rect 725 -2952 737 -2932
rect 757 -2952 769 -2932
rect 725 -2994 769 -2952
rect 819 -2932 861 -2894
rect 819 -2952 833 -2932
rect 853 -2952 861 -2932
rect 819 -2994 861 -2952
rect 935 -2932 977 -2894
rect 935 -2952 943 -2932
rect 963 -2952 977 -2932
rect 935 -2994 977 -2952
rect 1027 -2925 1072 -2894
rect 1027 -2932 1071 -2925
rect 1027 -2952 1039 -2932
rect 1059 -2952 1071 -2932
rect 1027 -2994 1071 -2952
rect 1384 -3214 1428 -3176
rect 1384 -3234 1396 -3214
rect 1416 -3234 1428 -3214
rect 1384 -3276 1428 -3234
rect 1478 -3214 1520 -3176
rect 1478 -3234 1492 -3214
rect 1512 -3234 1520 -3214
rect 1478 -3276 1520 -3234
rect 1597 -3214 1641 -3176
rect 1597 -3234 1609 -3214
rect 1629 -3234 1641 -3214
rect 1597 -3276 1641 -3234
rect 1691 -3214 1733 -3176
rect 1691 -3234 1705 -3214
rect 1725 -3234 1733 -3214
rect 1691 -3276 1733 -3234
rect 1805 -3214 1849 -3176
rect 1805 -3234 1817 -3214
rect 1837 -3234 1849 -3214
rect 1805 -3276 1849 -3234
rect 1899 -3214 1941 -3176
rect 1899 -3234 1913 -3214
rect 1933 -3234 1941 -3214
rect 1899 -3276 1941 -3234
rect 2015 -3214 2057 -3176
rect 2015 -3234 2023 -3214
rect 2043 -3234 2057 -3214
rect 2015 -3276 2057 -3234
rect 2107 -3207 2152 -3176
rect 2107 -3214 2151 -3207
rect 2107 -3234 2119 -3214
rect 2139 -3234 2151 -3214
rect 2107 -3276 2151 -3234
rect 306 -3481 350 -3443
rect 306 -3501 318 -3481
rect 338 -3501 350 -3481
rect 306 -3543 350 -3501
rect 400 -3481 442 -3443
rect 400 -3501 414 -3481
rect 434 -3501 442 -3481
rect 400 -3543 442 -3501
rect 519 -3481 563 -3443
rect 519 -3501 531 -3481
rect 551 -3501 563 -3481
rect 519 -3543 563 -3501
rect 613 -3481 655 -3443
rect 613 -3501 627 -3481
rect 647 -3501 655 -3481
rect 613 -3543 655 -3501
rect 727 -3481 771 -3443
rect 727 -3501 739 -3481
rect 759 -3501 771 -3481
rect 727 -3543 771 -3501
rect 821 -3481 863 -3443
rect 821 -3501 835 -3481
rect 855 -3501 863 -3481
rect 821 -3543 863 -3501
rect 937 -3481 979 -3443
rect 937 -3501 945 -3481
rect 965 -3501 979 -3481
rect 937 -3543 979 -3501
rect 1029 -3474 1074 -3443
rect 1029 -3481 1073 -3474
rect 1029 -3501 1041 -3481
rect 1061 -3501 1073 -3481
rect 1029 -3543 1073 -3501
rect 1244 -3725 1288 -3687
rect 1244 -3745 1256 -3725
rect 1276 -3745 1288 -3725
rect 1244 -3787 1288 -3745
rect 1338 -3725 1380 -3687
rect 1338 -3745 1352 -3725
rect 1372 -3745 1380 -3725
rect 1338 -3787 1380 -3745
rect 1457 -3725 1501 -3687
rect 1457 -3745 1469 -3725
rect 1489 -3745 1501 -3725
rect 1457 -3787 1501 -3745
rect 1551 -3725 1593 -3687
rect 1551 -3745 1565 -3725
rect 1585 -3745 1593 -3725
rect 1551 -3787 1593 -3745
rect 1665 -3725 1709 -3687
rect 1665 -3745 1677 -3725
rect 1697 -3745 1709 -3725
rect 1665 -3787 1709 -3745
rect 1759 -3725 1801 -3687
rect 1759 -3745 1773 -3725
rect 1793 -3745 1801 -3725
rect 1759 -3787 1801 -3745
rect 1875 -3725 1917 -3687
rect 1875 -3745 1883 -3725
rect 1903 -3745 1917 -3725
rect 1875 -3787 1917 -3745
rect 1967 -3718 2012 -3687
rect 1967 -3725 2011 -3718
rect 1967 -3745 1979 -3725
rect 1999 -3745 2011 -3725
rect 1967 -3787 2011 -3745
rect 305 -4035 349 -3997
rect 305 -4055 317 -4035
rect 337 -4055 349 -4035
rect 305 -4097 349 -4055
rect 399 -4035 441 -3997
rect 399 -4055 413 -4035
rect 433 -4055 441 -4035
rect 399 -4097 441 -4055
rect 518 -4035 562 -3997
rect 518 -4055 530 -4035
rect 550 -4055 562 -4035
rect 518 -4097 562 -4055
rect 612 -4035 654 -3997
rect 612 -4055 626 -4035
rect 646 -4055 654 -4035
rect 612 -4097 654 -4055
rect 726 -4035 770 -3997
rect 726 -4055 738 -4035
rect 758 -4055 770 -4035
rect 726 -4097 770 -4055
rect 820 -4035 862 -3997
rect 820 -4055 834 -4035
rect 854 -4055 862 -4035
rect 820 -4097 862 -4055
rect 936 -4035 978 -3997
rect 936 -4055 944 -4035
rect 964 -4055 978 -4035
rect 936 -4097 978 -4055
rect 1028 -4028 1073 -3997
rect 1028 -4035 1072 -4028
rect 1028 -4055 1040 -4035
rect 1060 -4055 1072 -4035
rect 1028 -4097 1072 -4055
<< ndiffc >>
rect 80 4356 98 4374
rect 82 4257 100 4275
rect 80 4169 98 4187
rect 82 4070 100 4088
rect 308 4071 328 4091
rect 411 4075 431 4095
rect 521 4071 541 4091
rect 624 4075 644 4095
rect 729 4071 749 4091
rect 832 4075 852 4095
rect 940 4075 960 4095
rect 1043 4071 1063 4091
rect 80 3940 98 3958
rect 82 3841 100 3859
rect 1246 3827 1266 3847
rect 1349 3831 1369 3851
rect 1459 3827 1479 3847
rect 1562 3831 1582 3851
rect 1667 3827 1687 3847
rect 1770 3831 1790 3851
rect 1878 3831 1898 3851
rect 1981 3827 2001 3847
rect 80 3710 98 3728
rect 82 3611 100 3629
rect 307 3517 327 3537
rect 410 3521 430 3541
rect 520 3517 540 3537
rect 623 3521 643 3541
rect 728 3517 748 3537
rect 831 3521 851 3541
rect 939 3521 959 3541
rect 1042 3517 1062 3537
rect 81 3253 99 3271
rect 1387 3235 1407 3255
rect 1490 3239 1510 3259
rect 1600 3235 1620 3255
rect 1703 3239 1723 3259
rect 1808 3235 1828 3255
rect 1911 3239 1931 3259
rect 2019 3239 2039 3259
rect 2122 3235 2142 3255
rect 83 3154 101 3172
rect 81 3066 99 3084
rect 83 2967 101 2985
rect 309 2968 329 2988
rect 412 2972 432 2992
rect 522 2968 542 2988
rect 625 2972 645 2992
rect 730 2968 750 2988
rect 833 2972 853 2992
rect 941 2972 961 2992
rect 1044 2968 1064 2988
rect 81 2837 99 2855
rect 83 2738 101 2756
rect 1247 2724 1267 2744
rect 1350 2728 1370 2748
rect 1460 2724 1480 2744
rect 1563 2728 1583 2748
rect 1668 2724 1688 2744
rect 1771 2728 1791 2748
rect 1879 2728 1899 2748
rect 1982 2724 2002 2744
rect 81 2607 99 2625
rect 83 2508 101 2526
rect 308 2414 328 2434
rect 411 2418 431 2438
rect 521 2414 541 2434
rect 624 2418 644 2438
rect 729 2414 749 2434
rect 832 2418 852 2438
rect 940 2418 960 2438
rect 1043 2414 1063 2434
rect 81 2150 99 2168
rect 1357 2145 1377 2165
rect 1460 2149 1480 2169
rect 1570 2145 1590 2165
rect 1673 2149 1693 2169
rect 1778 2145 1798 2165
rect 1881 2149 1901 2169
rect 1989 2149 2009 2169
rect 2092 2145 2112 2165
rect 83 2051 101 2069
rect 81 1963 99 1981
rect 83 1864 101 1882
rect 309 1865 329 1885
rect 412 1869 432 1889
rect 522 1865 542 1885
rect 625 1869 645 1889
rect 730 1865 750 1885
rect 833 1869 853 1889
rect 941 1869 961 1889
rect 1044 1865 1064 1885
rect 81 1734 99 1752
rect 83 1635 101 1653
rect 1247 1621 1267 1641
rect 1350 1625 1370 1645
rect 1460 1621 1480 1641
rect 1563 1625 1583 1645
rect 1668 1621 1688 1641
rect 1771 1625 1791 1645
rect 1879 1625 1899 1645
rect 1982 1621 2002 1641
rect 81 1504 99 1522
rect 83 1405 101 1423
rect 308 1311 328 1331
rect 411 1315 431 1335
rect 521 1311 541 1331
rect 624 1315 644 1335
rect 729 1311 749 1331
rect 832 1315 852 1335
rect 940 1315 960 1335
rect 1043 1311 1063 1331
rect 82 1047 100 1065
rect 1388 1029 1408 1049
rect 1491 1033 1511 1053
rect 1601 1029 1621 1049
rect 1704 1033 1724 1053
rect 1809 1029 1829 1049
rect 1912 1033 1932 1053
rect 2020 1033 2040 1053
rect 2123 1029 2143 1049
rect 84 948 102 966
rect 82 860 100 878
rect 84 761 102 779
rect 310 762 330 782
rect 413 766 433 786
rect 523 762 543 782
rect 626 766 646 786
rect 731 762 751 782
rect 834 766 854 786
rect 942 766 962 786
rect 1045 762 1065 782
rect 82 631 100 649
rect 84 532 102 550
rect 1248 518 1268 538
rect 1351 522 1371 542
rect 1461 518 1481 538
rect 1564 522 1584 542
rect 1669 518 1689 538
rect 1772 522 1792 542
rect 1880 522 1900 542
rect 1983 518 2003 538
rect 82 401 100 419
rect 84 302 102 320
rect 309 208 329 228
rect 412 212 432 232
rect 522 208 542 228
rect 625 212 645 232
rect 730 208 750 228
rect 833 212 853 232
rect 941 212 961 232
rect 1044 208 1064 228
rect 82 -56 100 -38
rect 1357 -55 1377 -35
rect 1460 -51 1480 -31
rect 1570 -55 1590 -35
rect 1673 -51 1693 -31
rect 1778 -55 1798 -35
rect 1881 -51 1901 -31
rect 1989 -51 2009 -31
rect 2092 -55 2112 -35
rect 84 -155 102 -137
rect 82 -243 100 -225
rect 84 -342 102 -324
rect 310 -341 330 -321
rect 413 -337 433 -317
rect 523 -341 543 -321
rect 626 -337 646 -317
rect 731 -341 751 -321
rect 834 -337 854 -317
rect 942 -337 962 -317
rect 1045 -341 1065 -321
rect 82 -472 100 -454
rect 84 -571 102 -553
rect 1248 -585 1268 -565
rect 1351 -581 1371 -561
rect 1461 -585 1481 -565
rect 1564 -581 1584 -561
rect 1669 -585 1689 -565
rect 1772 -581 1792 -561
rect 1880 -581 1900 -561
rect 1983 -585 2003 -565
rect 82 -702 100 -684
rect 84 -801 102 -783
rect 309 -895 329 -875
rect 412 -891 432 -871
rect 522 -895 542 -875
rect 625 -891 645 -871
rect 730 -895 750 -875
rect 833 -891 853 -871
rect 941 -891 961 -871
rect 1044 -895 1064 -875
rect 83 -1159 101 -1141
rect 1389 -1177 1409 -1157
rect 1492 -1173 1512 -1153
rect 1602 -1177 1622 -1157
rect 1705 -1173 1725 -1153
rect 1810 -1177 1830 -1157
rect 1913 -1173 1933 -1153
rect 2021 -1173 2041 -1153
rect 2124 -1177 2144 -1157
rect 85 -1258 103 -1240
rect 83 -1346 101 -1328
rect 85 -1445 103 -1427
rect 311 -1444 331 -1424
rect 414 -1440 434 -1420
rect 524 -1444 544 -1424
rect 627 -1440 647 -1420
rect 732 -1444 752 -1424
rect 835 -1440 855 -1420
rect 943 -1440 963 -1420
rect 1046 -1444 1066 -1424
rect 83 -1575 101 -1557
rect 85 -1674 103 -1656
rect 1249 -1688 1269 -1668
rect 1352 -1684 1372 -1664
rect 1462 -1688 1482 -1668
rect 1565 -1684 1585 -1664
rect 1670 -1688 1690 -1668
rect 1773 -1684 1793 -1664
rect 1881 -1684 1901 -1664
rect 1984 -1688 2004 -1668
rect 83 -1805 101 -1787
rect 85 -1904 103 -1886
rect 310 -1998 330 -1978
rect 413 -1994 433 -1974
rect 523 -1998 543 -1978
rect 626 -1994 646 -1974
rect 731 -1998 751 -1978
rect 834 -1994 854 -1974
rect 942 -1994 962 -1974
rect 1045 -1998 1065 -1978
rect 83 -2262 101 -2244
rect 1359 -2267 1379 -2247
rect 1462 -2263 1482 -2243
rect 1572 -2267 1592 -2247
rect 1675 -2263 1695 -2243
rect 1780 -2267 1800 -2247
rect 1883 -2263 1903 -2243
rect 1991 -2263 2011 -2243
rect 2094 -2267 2114 -2247
rect 85 -2361 103 -2343
rect 83 -2449 101 -2431
rect 85 -2548 103 -2530
rect 311 -2547 331 -2527
rect 414 -2543 434 -2523
rect 524 -2547 544 -2527
rect 627 -2543 647 -2523
rect 732 -2547 752 -2527
rect 835 -2543 855 -2523
rect 943 -2543 963 -2523
rect 1046 -2547 1066 -2527
rect 83 -2678 101 -2660
rect 85 -2777 103 -2759
rect 1249 -2791 1269 -2771
rect 1352 -2787 1372 -2767
rect 1462 -2791 1482 -2771
rect 1565 -2787 1585 -2767
rect 1670 -2791 1690 -2771
rect 1773 -2787 1793 -2767
rect 1881 -2787 1901 -2767
rect 1984 -2791 2004 -2771
rect 83 -2908 101 -2890
rect 85 -3007 103 -2989
rect 310 -3101 330 -3081
rect 413 -3097 433 -3077
rect 523 -3101 543 -3081
rect 626 -3097 646 -3077
rect 731 -3101 751 -3081
rect 834 -3097 854 -3077
rect 942 -3097 962 -3077
rect 1045 -3101 1065 -3081
rect 84 -3365 102 -3347
rect 1390 -3383 1410 -3363
rect 1493 -3379 1513 -3359
rect 1603 -3383 1623 -3363
rect 1706 -3379 1726 -3359
rect 1811 -3383 1831 -3363
rect 1914 -3379 1934 -3359
rect 2022 -3379 2042 -3359
rect 2125 -3383 2145 -3363
rect 86 -3464 104 -3446
rect 84 -3552 102 -3534
rect 86 -3651 104 -3633
rect 312 -3650 332 -3630
rect 415 -3646 435 -3626
rect 525 -3650 545 -3630
rect 628 -3646 648 -3626
rect 733 -3650 753 -3630
rect 836 -3646 856 -3626
rect 944 -3646 964 -3626
rect 1047 -3650 1067 -3630
rect 84 -3781 102 -3763
rect 86 -3880 104 -3862
rect 1250 -3894 1270 -3874
rect 1353 -3890 1373 -3870
rect 1463 -3894 1483 -3874
rect 1566 -3890 1586 -3870
rect 1671 -3894 1691 -3874
rect 1774 -3890 1794 -3870
rect 1882 -3890 1902 -3870
rect 1985 -3894 2005 -3874
rect 84 -4011 102 -3993
rect 86 -4110 104 -4092
rect 311 -4204 331 -4184
rect 414 -4200 434 -4180
rect 524 -4204 544 -4184
rect 627 -4200 647 -4180
rect 732 -4204 752 -4184
rect 835 -4200 855 -4180
rect 943 -4200 963 -4180
rect 1046 -4204 1066 -4184
<< pdiffc >>
rect 314 4220 334 4240
rect 410 4220 430 4240
rect 527 4220 547 4240
rect 623 4220 643 4240
rect 735 4220 755 4240
rect 831 4220 851 4240
rect 941 4220 961 4240
rect 1037 4220 1057 4240
rect 1252 3976 1272 3996
rect 1348 3976 1368 3996
rect 1465 3976 1485 3996
rect 1561 3976 1581 3996
rect 1673 3976 1693 3996
rect 1769 3976 1789 3996
rect 1879 3976 1899 3996
rect 1975 3976 1995 3996
rect 313 3666 333 3686
rect 409 3666 429 3686
rect 526 3666 546 3686
rect 622 3666 642 3686
rect 734 3666 754 3686
rect 830 3666 850 3686
rect 940 3666 960 3686
rect 1036 3666 1056 3686
rect 1393 3384 1413 3404
rect 1489 3384 1509 3404
rect 1606 3384 1626 3404
rect 1702 3384 1722 3404
rect 1814 3384 1834 3404
rect 1910 3384 1930 3404
rect 2020 3384 2040 3404
rect 2116 3384 2136 3404
rect 315 3117 335 3137
rect 411 3117 431 3137
rect 528 3117 548 3137
rect 624 3117 644 3137
rect 736 3117 756 3137
rect 832 3117 852 3137
rect 942 3117 962 3137
rect 1038 3117 1058 3137
rect 1253 2873 1273 2893
rect 1349 2873 1369 2893
rect 1466 2873 1486 2893
rect 1562 2873 1582 2893
rect 1674 2873 1694 2893
rect 1770 2873 1790 2893
rect 1880 2873 1900 2893
rect 1976 2873 1996 2893
rect 314 2563 334 2583
rect 410 2563 430 2583
rect 527 2563 547 2583
rect 623 2563 643 2583
rect 735 2563 755 2583
rect 831 2563 851 2583
rect 941 2563 961 2583
rect 1037 2563 1057 2583
rect 1363 2294 1383 2314
rect 1459 2294 1479 2314
rect 1576 2294 1596 2314
rect 1672 2294 1692 2314
rect 1784 2294 1804 2314
rect 1880 2294 1900 2314
rect 1990 2294 2010 2314
rect 2086 2294 2106 2314
rect 315 2014 335 2034
rect 411 2014 431 2034
rect 528 2014 548 2034
rect 624 2014 644 2034
rect 736 2014 756 2034
rect 832 2014 852 2034
rect 942 2014 962 2034
rect 1038 2014 1058 2034
rect 1253 1770 1273 1790
rect 1349 1770 1369 1790
rect 1466 1770 1486 1790
rect 1562 1770 1582 1790
rect 1674 1770 1694 1790
rect 1770 1770 1790 1790
rect 1880 1770 1900 1790
rect 1976 1770 1996 1790
rect 314 1460 334 1480
rect 410 1460 430 1480
rect 527 1460 547 1480
rect 623 1460 643 1480
rect 735 1460 755 1480
rect 831 1460 851 1480
rect 941 1460 961 1480
rect 1037 1460 1057 1480
rect 1394 1178 1414 1198
rect 1490 1178 1510 1198
rect 1607 1178 1627 1198
rect 1703 1178 1723 1198
rect 1815 1178 1835 1198
rect 1911 1178 1931 1198
rect 2021 1178 2041 1198
rect 2117 1178 2137 1198
rect 316 911 336 931
rect 412 911 432 931
rect 529 911 549 931
rect 625 911 645 931
rect 737 911 757 931
rect 833 911 853 931
rect 943 911 963 931
rect 1039 911 1059 931
rect 1254 667 1274 687
rect 1350 667 1370 687
rect 1467 667 1487 687
rect 1563 667 1583 687
rect 1675 667 1695 687
rect 1771 667 1791 687
rect 1881 667 1901 687
rect 1977 667 1997 687
rect 315 357 335 377
rect 411 357 431 377
rect 528 357 548 377
rect 624 357 644 377
rect 736 357 756 377
rect 832 357 852 377
rect 942 357 962 377
rect 1038 357 1058 377
rect 1363 94 1383 114
rect 1459 94 1479 114
rect 1576 94 1596 114
rect 1672 94 1692 114
rect 1784 94 1804 114
rect 1880 94 1900 114
rect 1990 94 2010 114
rect 2086 94 2106 114
rect 316 -192 336 -172
rect 412 -192 432 -172
rect 529 -192 549 -172
rect 625 -192 645 -172
rect 737 -192 757 -172
rect 833 -192 853 -172
rect 943 -192 963 -172
rect 1039 -192 1059 -172
rect 1254 -436 1274 -416
rect 1350 -436 1370 -416
rect 1467 -436 1487 -416
rect 1563 -436 1583 -416
rect 1675 -436 1695 -416
rect 1771 -436 1791 -416
rect 1881 -436 1901 -416
rect 1977 -436 1997 -416
rect 315 -746 335 -726
rect 411 -746 431 -726
rect 528 -746 548 -726
rect 624 -746 644 -726
rect 736 -746 756 -726
rect 832 -746 852 -726
rect 942 -746 962 -726
rect 1038 -746 1058 -726
rect 1395 -1028 1415 -1008
rect 1491 -1028 1511 -1008
rect 1608 -1028 1628 -1008
rect 1704 -1028 1724 -1008
rect 1816 -1028 1836 -1008
rect 1912 -1028 1932 -1008
rect 2022 -1028 2042 -1008
rect 2118 -1028 2138 -1008
rect 317 -1295 337 -1275
rect 413 -1295 433 -1275
rect 530 -1295 550 -1275
rect 626 -1295 646 -1275
rect 738 -1295 758 -1275
rect 834 -1295 854 -1275
rect 944 -1295 964 -1275
rect 1040 -1295 1060 -1275
rect 1255 -1539 1275 -1519
rect 1351 -1539 1371 -1519
rect 1468 -1539 1488 -1519
rect 1564 -1539 1584 -1519
rect 1676 -1539 1696 -1519
rect 1772 -1539 1792 -1519
rect 1882 -1539 1902 -1519
rect 1978 -1539 1998 -1519
rect 316 -1849 336 -1829
rect 412 -1849 432 -1829
rect 529 -1849 549 -1829
rect 625 -1849 645 -1829
rect 737 -1849 757 -1829
rect 833 -1849 853 -1829
rect 943 -1849 963 -1829
rect 1039 -1849 1059 -1829
rect 1365 -2118 1385 -2098
rect 1461 -2118 1481 -2098
rect 1578 -2118 1598 -2098
rect 1674 -2118 1694 -2098
rect 1786 -2118 1806 -2098
rect 1882 -2118 1902 -2098
rect 1992 -2118 2012 -2098
rect 2088 -2118 2108 -2098
rect 317 -2398 337 -2378
rect 413 -2398 433 -2378
rect 530 -2398 550 -2378
rect 626 -2398 646 -2378
rect 738 -2398 758 -2378
rect 834 -2398 854 -2378
rect 944 -2398 964 -2378
rect 1040 -2398 1060 -2378
rect 1255 -2642 1275 -2622
rect 1351 -2642 1371 -2622
rect 1468 -2642 1488 -2622
rect 1564 -2642 1584 -2622
rect 1676 -2642 1696 -2622
rect 1772 -2642 1792 -2622
rect 1882 -2642 1902 -2622
rect 1978 -2642 1998 -2622
rect 316 -2952 336 -2932
rect 412 -2952 432 -2932
rect 529 -2952 549 -2932
rect 625 -2952 645 -2932
rect 737 -2952 757 -2932
rect 833 -2952 853 -2932
rect 943 -2952 963 -2932
rect 1039 -2952 1059 -2932
rect 1396 -3234 1416 -3214
rect 1492 -3234 1512 -3214
rect 1609 -3234 1629 -3214
rect 1705 -3234 1725 -3214
rect 1817 -3234 1837 -3214
rect 1913 -3234 1933 -3214
rect 2023 -3234 2043 -3214
rect 2119 -3234 2139 -3214
rect 318 -3501 338 -3481
rect 414 -3501 434 -3481
rect 531 -3501 551 -3481
rect 627 -3501 647 -3481
rect 739 -3501 759 -3481
rect 835 -3501 855 -3481
rect 945 -3501 965 -3481
rect 1041 -3501 1061 -3481
rect 1256 -3745 1276 -3725
rect 1352 -3745 1372 -3725
rect 1469 -3745 1489 -3725
rect 1565 -3745 1585 -3725
rect 1677 -3745 1697 -3725
rect 1773 -3745 1793 -3725
rect 1883 -3745 1903 -3725
rect 1979 -3745 1999 -3725
rect 317 -4055 337 -4035
rect 413 -4055 433 -4035
rect 530 -4055 550 -4035
rect 626 -4055 646 -4035
rect 738 -4055 758 -4035
rect 834 -4055 854 -4035
rect 944 -4055 964 -4035
rect 1040 -4055 1060 -4035
<< psubdiff >>
rect 382 4004 493 4018
rect 382 3974 423 4004
rect 451 3974 493 4004
rect 382 3959 493 3974
rect 1320 3760 1431 3774
rect 1320 3730 1361 3760
rect 1389 3730 1431 3760
rect 1320 3715 1431 3730
rect 381 3450 492 3464
rect 381 3420 422 3450
rect 450 3420 492 3450
rect 381 3405 492 3420
rect 1461 3168 1572 3182
rect 1461 3138 1502 3168
rect 1530 3138 1572 3168
rect 1461 3123 1572 3138
rect 383 2901 494 2915
rect 383 2871 424 2901
rect 452 2871 494 2901
rect 383 2856 494 2871
rect 1321 2657 1432 2671
rect 1321 2627 1362 2657
rect 1390 2627 1432 2657
rect 1321 2612 1432 2627
rect 382 2347 493 2361
rect 382 2317 423 2347
rect 451 2317 493 2347
rect 382 2303 493 2317
rect 1431 2078 1542 2092
rect 1431 2048 1472 2078
rect 1500 2048 1542 2078
rect 1431 2033 1542 2048
rect 383 1798 494 1812
rect 383 1768 424 1798
rect 452 1768 494 1798
rect 383 1753 494 1768
rect 1321 1554 1432 1568
rect 1321 1524 1362 1554
rect 1390 1524 1432 1554
rect 1321 1509 1432 1524
rect 382 1244 493 1258
rect 382 1214 423 1244
rect 451 1214 493 1244
rect 382 1199 493 1214
rect 1462 962 1573 976
rect 1462 932 1503 962
rect 1531 932 1573 962
rect 1462 917 1573 932
rect 384 695 495 709
rect 384 665 425 695
rect 453 665 495 695
rect 384 650 495 665
rect 1322 451 1433 465
rect 1322 421 1363 451
rect 1391 421 1433 451
rect 1322 406 1433 421
rect 383 141 494 155
rect 383 111 424 141
rect 452 111 494 141
rect 383 96 494 111
rect 1431 -122 1542 -108
rect 1431 -152 1472 -122
rect 1500 -152 1542 -122
rect 1431 -167 1542 -152
rect 384 -408 495 -394
rect 384 -438 425 -408
rect 453 -438 495 -408
rect 384 -453 495 -438
rect 1322 -652 1433 -638
rect 1322 -682 1363 -652
rect 1391 -682 1433 -652
rect 1322 -697 1433 -682
rect 383 -962 494 -948
rect 383 -992 424 -962
rect 452 -992 494 -962
rect 383 -1007 494 -992
rect 1463 -1244 1574 -1230
rect 1463 -1274 1504 -1244
rect 1532 -1274 1574 -1244
rect 1463 -1289 1574 -1274
rect 385 -1511 496 -1497
rect 385 -1541 426 -1511
rect 454 -1541 496 -1511
rect 385 -1556 496 -1541
rect 1323 -1755 1434 -1741
rect 1323 -1785 1364 -1755
rect 1392 -1785 1434 -1755
rect 1323 -1800 1434 -1785
rect 384 -2065 495 -2051
rect 384 -2095 425 -2065
rect 453 -2095 495 -2065
rect 384 -2109 495 -2095
rect 1433 -2334 1544 -2320
rect 1433 -2364 1474 -2334
rect 1502 -2364 1544 -2334
rect 1433 -2379 1544 -2364
rect 385 -2614 496 -2600
rect 385 -2644 426 -2614
rect 454 -2644 496 -2614
rect 385 -2659 496 -2644
rect 1323 -2858 1434 -2844
rect 1323 -2888 1364 -2858
rect 1392 -2888 1434 -2858
rect 1323 -2903 1434 -2888
rect 384 -3168 495 -3154
rect 384 -3198 425 -3168
rect 453 -3198 495 -3168
rect 384 -3213 495 -3198
rect 1464 -3450 1575 -3436
rect 1464 -3480 1505 -3450
rect 1533 -3480 1575 -3450
rect 1464 -3495 1575 -3480
rect 386 -3717 497 -3703
rect 386 -3747 427 -3717
rect 455 -3747 497 -3717
rect 386 -3762 497 -3747
rect 1324 -3961 1435 -3947
rect 1324 -3991 1365 -3961
rect 1393 -3991 1435 -3961
rect 1324 -4006 1435 -3991
rect 385 -4271 496 -4257
rect 385 -4301 426 -4271
rect 454 -4301 496 -4271
rect 385 -4316 496 -4301
<< nsubdiff >>
rect 383 4351 493 4365
rect 383 4321 426 4351
rect 454 4321 493 4351
rect 383 4306 493 4321
rect 1321 4107 1431 4121
rect 1321 4077 1364 4107
rect 1392 4077 1431 4107
rect 1321 4062 1431 4077
rect 382 3797 492 3811
rect 382 3767 425 3797
rect 453 3767 492 3797
rect 382 3752 492 3767
rect 1462 3515 1572 3529
rect 1462 3485 1505 3515
rect 1533 3485 1572 3515
rect 1462 3470 1572 3485
rect 384 3248 494 3262
rect 384 3218 427 3248
rect 455 3218 494 3248
rect 384 3203 494 3218
rect 1322 3004 1432 3018
rect 1322 2974 1365 3004
rect 1393 2974 1432 3004
rect 1322 2959 1432 2974
rect 383 2694 493 2708
rect 383 2664 426 2694
rect 454 2664 493 2694
rect 383 2649 493 2664
rect 1432 2425 1542 2439
rect 1432 2395 1475 2425
rect 1503 2395 1542 2425
rect 1432 2380 1542 2395
rect 384 2145 494 2159
rect 384 2115 427 2145
rect 455 2115 494 2145
rect 384 2100 494 2115
rect 1322 1901 1432 1915
rect 1322 1871 1365 1901
rect 1393 1871 1432 1901
rect 1322 1856 1432 1871
rect 383 1591 493 1605
rect 383 1561 426 1591
rect 454 1561 493 1591
rect 383 1546 493 1561
rect 1463 1309 1573 1323
rect 1463 1279 1506 1309
rect 1534 1279 1573 1309
rect 1463 1264 1573 1279
rect 385 1042 495 1056
rect 385 1012 428 1042
rect 456 1012 495 1042
rect 385 997 495 1012
rect 1323 798 1433 812
rect 1323 768 1366 798
rect 1394 768 1433 798
rect 1323 753 1433 768
rect 384 488 494 502
rect 384 458 427 488
rect 455 458 494 488
rect 384 443 494 458
rect 1432 225 1542 239
rect 1432 195 1475 225
rect 1503 195 1542 225
rect 1432 180 1542 195
rect 385 -61 495 -47
rect 385 -91 428 -61
rect 456 -91 495 -61
rect 385 -106 495 -91
rect 1323 -305 1433 -291
rect 1323 -335 1366 -305
rect 1394 -335 1433 -305
rect 1323 -350 1433 -335
rect 384 -615 494 -601
rect 384 -645 427 -615
rect 455 -645 494 -615
rect 384 -660 494 -645
rect 1464 -897 1574 -883
rect 1464 -927 1507 -897
rect 1535 -927 1574 -897
rect 1464 -942 1574 -927
rect 386 -1164 496 -1150
rect 386 -1194 429 -1164
rect 457 -1194 496 -1164
rect 386 -1209 496 -1194
rect 1324 -1408 1434 -1394
rect 1324 -1438 1367 -1408
rect 1395 -1438 1434 -1408
rect 1324 -1453 1434 -1438
rect 385 -1718 495 -1704
rect 385 -1748 428 -1718
rect 456 -1748 495 -1718
rect 385 -1763 495 -1748
rect 1434 -1987 1544 -1973
rect 1434 -2017 1477 -1987
rect 1505 -2017 1544 -1987
rect 1434 -2032 1544 -2017
rect 386 -2267 496 -2253
rect 386 -2297 429 -2267
rect 457 -2297 496 -2267
rect 386 -2312 496 -2297
rect 1324 -2511 1434 -2497
rect 1324 -2541 1367 -2511
rect 1395 -2541 1434 -2511
rect 1324 -2556 1434 -2541
rect 385 -2821 495 -2807
rect 385 -2851 428 -2821
rect 456 -2851 495 -2821
rect 385 -2866 495 -2851
rect 1465 -3103 1575 -3089
rect 1465 -3133 1508 -3103
rect 1536 -3133 1575 -3103
rect 1465 -3148 1575 -3133
rect 387 -3370 497 -3356
rect 387 -3400 430 -3370
rect 458 -3400 497 -3370
rect 387 -3415 497 -3400
rect 1325 -3614 1435 -3600
rect 1325 -3644 1368 -3614
rect 1396 -3644 1435 -3614
rect 1325 -3659 1435 -3644
rect 386 -3924 496 -3910
rect 386 -3954 429 -3924
rect 457 -3954 496 -3924
rect 386 -3969 496 -3954
<< psubdiffcont >>
rect 423 3974 451 4004
rect 1361 3730 1389 3760
rect 422 3420 450 3450
rect 1502 3138 1530 3168
rect 424 2871 452 2901
rect 1362 2627 1390 2657
rect 423 2317 451 2347
rect 1472 2048 1500 2078
rect 424 1768 452 1798
rect 1362 1524 1390 1554
rect 423 1214 451 1244
rect 1503 932 1531 962
rect 425 665 453 695
rect 1363 421 1391 451
rect 424 111 452 141
rect 1472 -152 1500 -122
rect 425 -438 453 -408
rect 1363 -682 1391 -652
rect 424 -992 452 -962
rect 1504 -1274 1532 -1244
rect 426 -1541 454 -1511
rect 1364 -1785 1392 -1755
rect 425 -2095 453 -2065
rect 1474 -2364 1502 -2334
rect 426 -2644 454 -2614
rect 1364 -2888 1392 -2858
rect 425 -3198 453 -3168
rect 1505 -3480 1533 -3450
rect 427 -3747 455 -3717
rect 1365 -3991 1393 -3961
rect 426 -4301 454 -4271
<< nsubdiffcont >>
rect 426 4321 454 4351
rect 1364 4077 1392 4107
rect 425 3767 453 3797
rect 1505 3485 1533 3515
rect 427 3218 455 3248
rect 1365 2974 1393 3004
rect 426 2664 454 2694
rect 1475 2395 1503 2425
rect 427 2115 455 2145
rect 1365 1871 1393 1901
rect 426 1561 454 1591
rect 1506 1279 1534 1309
rect 428 1012 456 1042
rect 1366 768 1394 798
rect 427 458 455 488
rect 1475 195 1503 225
rect 428 -91 456 -61
rect 1366 -335 1394 -305
rect 427 -645 455 -615
rect 1507 -927 1535 -897
rect 429 -1194 457 -1164
rect 1367 -1438 1395 -1408
rect 428 -1748 456 -1718
rect 1477 -2017 1505 -1987
rect 429 -2297 457 -2267
rect 1367 -2541 1395 -2511
rect 428 -2851 456 -2821
rect 1508 -3133 1536 -3103
rect 430 -3400 458 -3370
rect 1368 -3644 1396 -3614
rect 429 -3954 457 -3924
<< poly >>
rect 346 4278 396 4291
rect 559 4278 609 4291
rect 767 4278 817 4291
rect 975 4278 1025 4291
rect 346 4150 396 4178
rect 346 4130 359 4150
rect 379 4130 396 4150
rect 346 4101 396 4130
rect 559 4149 609 4178
rect 559 4125 570 4149
rect 594 4125 609 4149
rect 559 4101 609 4125
rect 767 4154 817 4178
rect 767 4130 779 4154
rect 803 4130 817 4154
rect 767 4101 817 4130
rect 975 4152 1025 4178
rect 975 4126 993 4152
rect 1019 4126 1025 4152
rect 975 4101 1025 4126
rect 346 4043 396 4059
rect 559 4043 609 4059
rect 767 4043 817 4059
rect 975 4043 1025 4059
rect 1284 4034 1334 4047
rect 1497 4034 1547 4047
rect 1705 4034 1755 4047
rect 1913 4034 1963 4047
rect 1284 3906 1334 3934
rect 1284 3886 1297 3906
rect 1317 3886 1334 3906
rect 1284 3857 1334 3886
rect 1497 3905 1547 3934
rect 1497 3881 1508 3905
rect 1532 3881 1547 3905
rect 1497 3857 1547 3881
rect 1705 3910 1755 3934
rect 1705 3886 1717 3910
rect 1741 3886 1755 3910
rect 1705 3857 1755 3886
rect 1913 3908 1963 3934
rect 1913 3882 1931 3908
rect 1957 3882 1963 3908
rect 1913 3857 1963 3882
rect 1284 3799 1334 3815
rect 1497 3799 1547 3815
rect 1705 3799 1755 3815
rect 1913 3799 1963 3815
rect 345 3724 395 3737
rect 558 3724 608 3737
rect 766 3724 816 3737
rect 974 3724 1024 3737
rect 345 3596 395 3624
rect 345 3576 358 3596
rect 378 3576 395 3596
rect 345 3547 395 3576
rect 558 3595 608 3624
rect 558 3571 569 3595
rect 593 3571 608 3595
rect 558 3547 608 3571
rect 766 3600 816 3624
rect 766 3576 778 3600
rect 802 3576 816 3600
rect 766 3547 816 3576
rect 974 3598 1024 3624
rect 974 3572 992 3598
rect 1018 3572 1024 3598
rect 974 3547 1024 3572
rect 345 3489 395 3505
rect 558 3489 608 3505
rect 766 3489 816 3505
rect 974 3489 1024 3505
rect 1425 3442 1475 3455
rect 1638 3442 1688 3455
rect 1846 3442 1896 3455
rect 2054 3442 2104 3455
rect 1425 3314 1475 3342
rect 1425 3294 1438 3314
rect 1458 3294 1475 3314
rect 1425 3265 1475 3294
rect 1638 3313 1688 3342
rect 1638 3289 1649 3313
rect 1673 3289 1688 3313
rect 1638 3265 1688 3289
rect 1846 3318 1896 3342
rect 1846 3294 1858 3318
rect 1882 3294 1896 3318
rect 1846 3265 1896 3294
rect 2054 3316 2104 3342
rect 2054 3290 2072 3316
rect 2098 3290 2104 3316
rect 2054 3265 2104 3290
rect 1425 3207 1475 3223
rect 1638 3207 1688 3223
rect 1846 3207 1896 3223
rect 2054 3207 2104 3223
rect 347 3175 397 3188
rect 560 3175 610 3188
rect 768 3175 818 3188
rect 976 3175 1026 3188
rect 347 3047 397 3075
rect 347 3027 360 3047
rect 380 3027 397 3047
rect 347 2998 397 3027
rect 560 3046 610 3075
rect 560 3022 571 3046
rect 595 3022 610 3046
rect 560 2998 610 3022
rect 768 3051 818 3075
rect 768 3027 780 3051
rect 804 3027 818 3051
rect 768 2998 818 3027
rect 976 3049 1026 3075
rect 976 3023 994 3049
rect 1020 3023 1026 3049
rect 976 2998 1026 3023
rect 347 2940 397 2956
rect 560 2940 610 2956
rect 768 2940 818 2956
rect 976 2940 1026 2956
rect 1285 2931 1335 2944
rect 1498 2931 1548 2944
rect 1706 2931 1756 2944
rect 1914 2931 1964 2944
rect 1285 2803 1335 2831
rect 1285 2783 1298 2803
rect 1318 2783 1335 2803
rect 1285 2754 1335 2783
rect 1498 2802 1548 2831
rect 1498 2778 1509 2802
rect 1533 2778 1548 2802
rect 1498 2754 1548 2778
rect 1706 2807 1756 2831
rect 1706 2783 1718 2807
rect 1742 2783 1756 2807
rect 1706 2754 1756 2783
rect 1914 2805 1964 2831
rect 1914 2779 1932 2805
rect 1958 2779 1964 2805
rect 1914 2754 1964 2779
rect 1285 2696 1335 2712
rect 1498 2696 1548 2712
rect 1706 2696 1756 2712
rect 1914 2696 1964 2712
rect 346 2621 396 2634
rect 559 2621 609 2634
rect 767 2621 817 2634
rect 975 2621 1025 2634
rect 346 2493 396 2521
rect 346 2473 359 2493
rect 379 2473 396 2493
rect 346 2444 396 2473
rect 559 2492 609 2521
rect 559 2468 570 2492
rect 594 2468 609 2492
rect 559 2444 609 2468
rect 767 2497 817 2521
rect 767 2473 779 2497
rect 803 2473 817 2497
rect 767 2444 817 2473
rect 975 2495 1025 2521
rect 975 2469 993 2495
rect 1019 2469 1025 2495
rect 975 2444 1025 2469
rect 346 2386 396 2402
rect 559 2386 609 2402
rect 767 2386 817 2402
rect 975 2386 1025 2402
rect 1395 2352 1445 2365
rect 1608 2352 1658 2365
rect 1816 2352 1866 2365
rect 2024 2352 2074 2365
rect 1395 2224 1445 2252
rect 1395 2204 1408 2224
rect 1428 2204 1445 2224
rect 1395 2175 1445 2204
rect 1608 2223 1658 2252
rect 1608 2199 1619 2223
rect 1643 2199 1658 2223
rect 1608 2175 1658 2199
rect 1816 2228 1866 2252
rect 1816 2204 1828 2228
rect 1852 2204 1866 2228
rect 1816 2175 1866 2204
rect 2024 2226 2074 2252
rect 2024 2200 2042 2226
rect 2068 2200 2074 2226
rect 2024 2175 2074 2200
rect 1395 2117 1445 2133
rect 1608 2117 1658 2133
rect 1816 2117 1866 2133
rect 2024 2117 2074 2133
rect 347 2072 397 2085
rect 560 2072 610 2085
rect 768 2072 818 2085
rect 976 2072 1026 2085
rect 347 1944 397 1972
rect 347 1924 360 1944
rect 380 1924 397 1944
rect 347 1895 397 1924
rect 560 1943 610 1972
rect 560 1919 571 1943
rect 595 1919 610 1943
rect 560 1895 610 1919
rect 768 1948 818 1972
rect 768 1924 780 1948
rect 804 1924 818 1948
rect 768 1895 818 1924
rect 976 1946 1026 1972
rect 976 1920 994 1946
rect 1020 1920 1026 1946
rect 976 1895 1026 1920
rect 347 1837 397 1853
rect 560 1837 610 1853
rect 768 1837 818 1853
rect 976 1837 1026 1853
rect 1285 1828 1335 1841
rect 1498 1828 1548 1841
rect 1706 1828 1756 1841
rect 1914 1828 1964 1841
rect 1285 1700 1335 1728
rect 1285 1680 1298 1700
rect 1318 1680 1335 1700
rect 1285 1651 1335 1680
rect 1498 1699 1548 1728
rect 1498 1675 1509 1699
rect 1533 1675 1548 1699
rect 1498 1651 1548 1675
rect 1706 1704 1756 1728
rect 1706 1680 1718 1704
rect 1742 1680 1756 1704
rect 1706 1651 1756 1680
rect 1914 1702 1964 1728
rect 1914 1676 1932 1702
rect 1958 1676 1964 1702
rect 1914 1651 1964 1676
rect 1285 1593 1335 1609
rect 1498 1593 1548 1609
rect 1706 1593 1756 1609
rect 1914 1593 1964 1609
rect 346 1518 396 1531
rect 559 1518 609 1531
rect 767 1518 817 1531
rect 975 1518 1025 1531
rect 346 1390 396 1418
rect 346 1370 359 1390
rect 379 1370 396 1390
rect 346 1341 396 1370
rect 559 1389 609 1418
rect 559 1365 570 1389
rect 594 1365 609 1389
rect 559 1341 609 1365
rect 767 1394 817 1418
rect 767 1370 779 1394
rect 803 1370 817 1394
rect 767 1341 817 1370
rect 975 1392 1025 1418
rect 975 1366 993 1392
rect 1019 1366 1025 1392
rect 975 1341 1025 1366
rect 346 1283 396 1299
rect 559 1283 609 1299
rect 767 1283 817 1299
rect 975 1283 1025 1299
rect 1426 1236 1476 1249
rect 1639 1236 1689 1249
rect 1847 1236 1897 1249
rect 2055 1236 2105 1249
rect 1426 1108 1476 1136
rect 1426 1088 1439 1108
rect 1459 1088 1476 1108
rect 1426 1059 1476 1088
rect 1639 1107 1689 1136
rect 1639 1083 1650 1107
rect 1674 1083 1689 1107
rect 1639 1059 1689 1083
rect 1847 1112 1897 1136
rect 1847 1088 1859 1112
rect 1883 1088 1897 1112
rect 1847 1059 1897 1088
rect 2055 1110 2105 1136
rect 2055 1084 2073 1110
rect 2099 1084 2105 1110
rect 2055 1059 2105 1084
rect 1426 1001 1476 1017
rect 1639 1001 1689 1017
rect 1847 1001 1897 1017
rect 2055 1001 2105 1017
rect 348 969 398 982
rect 561 969 611 982
rect 769 969 819 982
rect 977 969 1027 982
rect 348 841 398 869
rect 348 821 361 841
rect 381 821 398 841
rect 348 792 398 821
rect 561 840 611 869
rect 561 816 572 840
rect 596 816 611 840
rect 561 792 611 816
rect 769 845 819 869
rect 769 821 781 845
rect 805 821 819 845
rect 769 792 819 821
rect 977 843 1027 869
rect 977 817 995 843
rect 1021 817 1027 843
rect 977 792 1027 817
rect 348 734 398 750
rect 561 734 611 750
rect 769 734 819 750
rect 977 734 1027 750
rect 1286 725 1336 738
rect 1499 725 1549 738
rect 1707 725 1757 738
rect 1915 725 1965 738
rect 1286 597 1336 625
rect 1286 577 1299 597
rect 1319 577 1336 597
rect 1286 548 1336 577
rect 1499 596 1549 625
rect 1499 572 1510 596
rect 1534 572 1549 596
rect 1499 548 1549 572
rect 1707 601 1757 625
rect 1707 577 1719 601
rect 1743 577 1757 601
rect 1707 548 1757 577
rect 1915 599 1965 625
rect 1915 573 1933 599
rect 1959 573 1965 599
rect 1915 548 1965 573
rect 1286 490 1336 506
rect 1499 490 1549 506
rect 1707 490 1757 506
rect 1915 490 1965 506
rect 347 415 397 428
rect 560 415 610 428
rect 768 415 818 428
rect 976 415 1026 428
rect 347 287 397 315
rect 347 267 360 287
rect 380 267 397 287
rect 347 238 397 267
rect 560 286 610 315
rect 560 262 571 286
rect 595 262 610 286
rect 560 238 610 262
rect 768 291 818 315
rect 768 267 780 291
rect 804 267 818 291
rect 768 238 818 267
rect 976 289 1026 315
rect 976 263 994 289
rect 1020 263 1026 289
rect 976 238 1026 263
rect 347 180 397 196
rect 560 180 610 196
rect 768 180 818 196
rect 976 180 1026 196
rect 1395 152 1445 165
rect 1608 152 1658 165
rect 1816 152 1866 165
rect 2024 152 2074 165
rect 1395 24 1445 52
rect 1395 4 1408 24
rect 1428 4 1445 24
rect 1395 -25 1445 4
rect 1608 23 1658 52
rect 1608 -1 1619 23
rect 1643 -1 1658 23
rect 1608 -25 1658 -1
rect 1816 28 1866 52
rect 1816 4 1828 28
rect 1852 4 1866 28
rect 1816 -25 1866 4
rect 2024 26 2074 52
rect 2024 0 2042 26
rect 2068 0 2074 26
rect 2024 -25 2074 0
rect 1395 -83 1445 -67
rect 1608 -83 1658 -67
rect 1816 -83 1866 -67
rect 2024 -83 2074 -67
rect 348 -134 398 -121
rect 561 -134 611 -121
rect 769 -134 819 -121
rect 977 -134 1027 -121
rect 348 -262 398 -234
rect 348 -282 361 -262
rect 381 -282 398 -262
rect 348 -311 398 -282
rect 561 -263 611 -234
rect 561 -287 572 -263
rect 596 -287 611 -263
rect 561 -311 611 -287
rect 769 -258 819 -234
rect 769 -282 781 -258
rect 805 -282 819 -258
rect 769 -311 819 -282
rect 977 -260 1027 -234
rect 977 -286 995 -260
rect 1021 -286 1027 -260
rect 977 -311 1027 -286
rect 348 -369 398 -353
rect 561 -369 611 -353
rect 769 -369 819 -353
rect 977 -369 1027 -353
rect 1286 -378 1336 -365
rect 1499 -378 1549 -365
rect 1707 -378 1757 -365
rect 1915 -378 1965 -365
rect 1286 -506 1336 -478
rect 1286 -526 1299 -506
rect 1319 -526 1336 -506
rect 1286 -555 1336 -526
rect 1499 -507 1549 -478
rect 1499 -531 1510 -507
rect 1534 -531 1549 -507
rect 1499 -555 1549 -531
rect 1707 -502 1757 -478
rect 1707 -526 1719 -502
rect 1743 -526 1757 -502
rect 1707 -555 1757 -526
rect 1915 -504 1965 -478
rect 1915 -530 1933 -504
rect 1959 -530 1965 -504
rect 1915 -555 1965 -530
rect 1286 -613 1336 -597
rect 1499 -613 1549 -597
rect 1707 -613 1757 -597
rect 1915 -613 1965 -597
rect 347 -688 397 -675
rect 560 -688 610 -675
rect 768 -688 818 -675
rect 976 -688 1026 -675
rect 347 -816 397 -788
rect 347 -836 360 -816
rect 380 -836 397 -816
rect 347 -865 397 -836
rect 560 -817 610 -788
rect 560 -841 571 -817
rect 595 -841 610 -817
rect 560 -865 610 -841
rect 768 -812 818 -788
rect 768 -836 780 -812
rect 804 -836 818 -812
rect 768 -865 818 -836
rect 976 -814 1026 -788
rect 976 -840 994 -814
rect 1020 -840 1026 -814
rect 976 -865 1026 -840
rect 347 -923 397 -907
rect 560 -923 610 -907
rect 768 -923 818 -907
rect 976 -923 1026 -907
rect 1427 -970 1477 -957
rect 1640 -970 1690 -957
rect 1848 -970 1898 -957
rect 2056 -970 2106 -957
rect 1427 -1098 1477 -1070
rect 1427 -1118 1440 -1098
rect 1460 -1118 1477 -1098
rect 1427 -1147 1477 -1118
rect 1640 -1099 1690 -1070
rect 1640 -1123 1651 -1099
rect 1675 -1123 1690 -1099
rect 1640 -1147 1690 -1123
rect 1848 -1094 1898 -1070
rect 1848 -1118 1860 -1094
rect 1884 -1118 1898 -1094
rect 1848 -1147 1898 -1118
rect 2056 -1096 2106 -1070
rect 2056 -1122 2074 -1096
rect 2100 -1122 2106 -1096
rect 2056 -1147 2106 -1122
rect 1427 -1205 1477 -1189
rect 1640 -1205 1690 -1189
rect 1848 -1205 1898 -1189
rect 2056 -1205 2106 -1189
rect 349 -1237 399 -1224
rect 562 -1237 612 -1224
rect 770 -1237 820 -1224
rect 978 -1237 1028 -1224
rect 349 -1365 399 -1337
rect 349 -1385 362 -1365
rect 382 -1385 399 -1365
rect 349 -1414 399 -1385
rect 562 -1366 612 -1337
rect 562 -1390 573 -1366
rect 597 -1390 612 -1366
rect 562 -1414 612 -1390
rect 770 -1361 820 -1337
rect 770 -1385 782 -1361
rect 806 -1385 820 -1361
rect 770 -1414 820 -1385
rect 978 -1363 1028 -1337
rect 978 -1389 996 -1363
rect 1022 -1389 1028 -1363
rect 978 -1414 1028 -1389
rect 349 -1472 399 -1456
rect 562 -1472 612 -1456
rect 770 -1472 820 -1456
rect 978 -1472 1028 -1456
rect 1287 -1481 1337 -1468
rect 1500 -1481 1550 -1468
rect 1708 -1481 1758 -1468
rect 1916 -1481 1966 -1468
rect 1287 -1609 1337 -1581
rect 1287 -1629 1300 -1609
rect 1320 -1629 1337 -1609
rect 1287 -1658 1337 -1629
rect 1500 -1610 1550 -1581
rect 1500 -1634 1511 -1610
rect 1535 -1634 1550 -1610
rect 1500 -1658 1550 -1634
rect 1708 -1605 1758 -1581
rect 1708 -1629 1720 -1605
rect 1744 -1629 1758 -1605
rect 1708 -1658 1758 -1629
rect 1916 -1607 1966 -1581
rect 1916 -1633 1934 -1607
rect 1960 -1633 1966 -1607
rect 1916 -1658 1966 -1633
rect 1287 -1716 1337 -1700
rect 1500 -1716 1550 -1700
rect 1708 -1716 1758 -1700
rect 1916 -1716 1966 -1700
rect 348 -1791 398 -1778
rect 561 -1791 611 -1778
rect 769 -1791 819 -1778
rect 977 -1791 1027 -1778
rect 348 -1919 398 -1891
rect 348 -1939 361 -1919
rect 381 -1939 398 -1919
rect 348 -1968 398 -1939
rect 561 -1920 611 -1891
rect 561 -1944 572 -1920
rect 596 -1944 611 -1920
rect 561 -1968 611 -1944
rect 769 -1915 819 -1891
rect 769 -1939 781 -1915
rect 805 -1939 819 -1915
rect 769 -1968 819 -1939
rect 977 -1917 1027 -1891
rect 977 -1943 995 -1917
rect 1021 -1943 1027 -1917
rect 977 -1968 1027 -1943
rect 348 -2026 398 -2010
rect 561 -2026 611 -2010
rect 769 -2026 819 -2010
rect 977 -2026 1027 -2010
rect 1397 -2060 1447 -2047
rect 1610 -2060 1660 -2047
rect 1818 -2060 1868 -2047
rect 2026 -2060 2076 -2047
rect 1397 -2188 1447 -2160
rect 1397 -2208 1410 -2188
rect 1430 -2208 1447 -2188
rect 1397 -2237 1447 -2208
rect 1610 -2189 1660 -2160
rect 1610 -2213 1621 -2189
rect 1645 -2213 1660 -2189
rect 1610 -2237 1660 -2213
rect 1818 -2184 1868 -2160
rect 1818 -2208 1830 -2184
rect 1854 -2208 1868 -2184
rect 1818 -2237 1868 -2208
rect 2026 -2186 2076 -2160
rect 2026 -2212 2044 -2186
rect 2070 -2212 2076 -2186
rect 2026 -2237 2076 -2212
rect 1397 -2295 1447 -2279
rect 1610 -2295 1660 -2279
rect 1818 -2295 1868 -2279
rect 2026 -2295 2076 -2279
rect 349 -2340 399 -2327
rect 562 -2340 612 -2327
rect 770 -2340 820 -2327
rect 978 -2340 1028 -2327
rect 349 -2468 399 -2440
rect 349 -2488 362 -2468
rect 382 -2488 399 -2468
rect 349 -2517 399 -2488
rect 562 -2469 612 -2440
rect 562 -2493 573 -2469
rect 597 -2493 612 -2469
rect 562 -2517 612 -2493
rect 770 -2464 820 -2440
rect 770 -2488 782 -2464
rect 806 -2488 820 -2464
rect 770 -2517 820 -2488
rect 978 -2466 1028 -2440
rect 978 -2492 996 -2466
rect 1022 -2492 1028 -2466
rect 978 -2517 1028 -2492
rect 349 -2575 399 -2559
rect 562 -2575 612 -2559
rect 770 -2575 820 -2559
rect 978 -2575 1028 -2559
rect 1287 -2584 1337 -2571
rect 1500 -2584 1550 -2571
rect 1708 -2584 1758 -2571
rect 1916 -2584 1966 -2571
rect 1287 -2712 1337 -2684
rect 1287 -2732 1300 -2712
rect 1320 -2732 1337 -2712
rect 1287 -2761 1337 -2732
rect 1500 -2713 1550 -2684
rect 1500 -2737 1511 -2713
rect 1535 -2737 1550 -2713
rect 1500 -2761 1550 -2737
rect 1708 -2708 1758 -2684
rect 1708 -2732 1720 -2708
rect 1744 -2732 1758 -2708
rect 1708 -2761 1758 -2732
rect 1916 -2710 1966 -2684
rect 1916 -2736 1934 -2710
rect 1960 -2736 1966 -2710
rect 1916 -2761 1966 -2736
rect 1287 -2819 1337 -2803
rect 1500 -2819 1550 -2803
rect 1708 -2819 1758 -2803
rect 1916 -2819 1966 -2803
rect 348 -2894 398 -2881
rect 561 -2894 611 -2881
rect 769 -2894 819 -2881
rect 977 -2894 1027 -2881
rect 348 -3022 398 -2994
rect 348 -3042 361 -3022
rect 381 -3042 398 -3022
rect 348 -3071 398 -3042
rect 561 -3023 611 -2994
rect 561 -3047 572 -3023
rect 596 -3047 611 -3023
rect 561 -3071 611 -3047
rect 769 -3018 819 -2994
rect 769 -3042 781 -3018
rect 805 -3042 819 -3018
rect 769 -3071 819 -3042
rect 977 -3020 1027 -2994
rect 977 -3046 995 -3020
rect 1021 -3046 1027 -3020
rect 977 -3071 1027 -3046
rect 348 -3129 398 -3113
rect 561 -3129 611 -3113
rect 769 -3129 819 -3113
rect 977 -3129 1027 -3113
rect 1428 -3176 1478 -3163
rect 1641 -3176 1691 -3163
rect 1849 -3176 1899 -3163
rect 2057 -3176 2107 -3163
rect 1428 -3304 1478 -3276
rect 1428 -3324 1441 -3304
rect 1461 -3324 1478 -3304
rect 1428 -3353 1478 -3324
rect 1641 -3305 1691 -3276
rect 1641 -3329 1652 -3305
rect 1676 -3329 1691 -3305
rect 1641 -3353 1691 -3329
rect 1849 -3300 1899 -3276
rect 1849 -3324 1861 -3300
rect 1885 -3324 1899 -3300
rect 1849 -3353 1899 -3324
rect 2057 -3302 2107 -3276
rect 2057 -3328 2075 -3302
rect 2101 -3328 2107 -3302
rect 2057 -3353 2107 -3328
rect 1428 -3411 1478 -3395
rect 1641 -3411 1691 -3395
rect 1849 -3411 1899 -3395
rect 2057 -3411 2107 -3395
rect 350 -3443 400 -3430
rect 563 -3443 613 -3430
rect 771 -3443 821 -3430
rect 979 -3443 1029 -3430
rect 350 -3571 400 -3543
rect 350 -3591 363 -3571
rect 383 -3591 400 -3571
rect 350 -3620 400 -3591
rect 563 -3572 613 -3543
rect 563 -3596 574 -3572
rect 598 -3596 613 -3572
rect 563 -3620 613 -3596
rect 771 -3567 821 -3543
rect 771 -3591 783 -3567
rect 807 -3591 821 -3567
rect 771 -3620 821 -3591
rect 979 -3569 1029 -3543
rect 979 -3595 997 -3569
rect 1023 -3595 1029 -3569
rect 979 -3620 1029 -3595
rect 350 -3678 400 -3662
rect 563 -3678 613 -3662
rect 771 -3678 821 -3662
rect 979 -3678 1029 -3662
rect 1288 -3687 1338 -3674
rect 1501 -3687 1551 -3674
rect 1709 -3687 1759 -3674
rect 1917 -3687 1967 -3674
rect 1288 -3815 1338 -3787
rect 1288 -3835 1301 -3815
rect 1321 -3835 1338 -3815
rect 1288 -3864 1338 -3835
rect 1501 -3816 1551 -3787
rect 1501 -3840 1512 -3816
rect 1536 -3840 1551 -3816
rect 1501 -3864 1551 -3840
rect 1709 -3811 1759 -3787
rect 1709 -3835 1721 -3811
rect 1745 -3835 1759 -3811
rect 1709 -3864 1759 -3835
rect 1917 -3813 1967 -3787
rect 1917 -3839 1935 -3813
rect 1961 -3839 1967 -3813
rect 1917 -3864 1967 -3839
rect 1288 -3922 1338 -3906
rect 1501 -3922 1551 -3906
rect 1709 -3922 1759 -3906
rect 1917 -3922 1967 -3906
rect 349 -3997 399 -3984
rect 562 -3997 612 -3984
rect 770 -3997 820 -3984
rect 978 -3997 1028 -3984
rect 349 -4125 399 -4097
rect 349 -4145 362 -4125
rect 382 -4145 399 -4125
rect 349 -4174 399 -4145
rect 562 -4126 612 -4097
rect 562 -4150 573 -4126
rect 597 -4150 612 -4126
rect 562 -4174 612 -4150
rect 770 -4121 820 -4097
rect 770 -4145 782 -4121
rect 806 -4145 820 -4121
rect 770 -4174 820 -4145
rect 978 -4123 1028 -4097
rect 978 -4149 996 -4123
rect 1022 -4149 1028 -4123
rect 978 -4174 1028 -4149
rect 349 -4232 399 -4216
rect 562 -4232 612 -4216
rect 770 -4232 820 -4216
rect 978 -4232 1028 -4216
<< polycont >>
rect 359 4130 379 4150
rect 570 4125 594 4149
rect 779 4130 803 4154
rect 993 4126 1019 4152
rect 1297 3886 1317 3906
rect 1508 3881 1532 3905
rect 1717 3886 1741 3910
rect 1931 3882 1957 3908
rect 358 3576 378 3596
rect 569 3571 593 3595
rect 778 3576 802 3600
rect 992 3572 1018 3598
rect 1438 3294 1458 3314
rect 1649 3289 1673 3313
rect 1858 3294 1882 3318
rect 2072 3290 2098 3316
rect 360 3027 380 3047
rect 571 3022 595 3046
rect 780 3027 804 3051
rect 994 3023 1020 3049
rect 1298 2783 1318 2803
rect 1509 2778 1533 2802
rect 1718 2783 1742 2807
rect 1932 2779 1958 2805
rect 359 2473 379 2493
rect 570 2468 594 2492
rect 779 2473 803 2497
rect 993 2469 1019 2495
rect 1408 2204 1428 2224
rect 1619 2199 1643 2223
rect 1828 2204 1852 2228
rect 2042 2200 2068 2226
rect 360 1924 380 1944
rect 571 1919 595 1943
rect 780 1924 804 1948
rect 994 1920 1020 1946
rect 1298 1680 1318 1700
rect 1509 1675 1533 1699
rect 1718 1680 1742 1704
rect 1932 1676 1958 1702
rect 359 1370 379 1390
rect 570 1365 594 1389
rect 779 1370 803 1394
rect 993 1366 1019 1392
rect 1439 1088 1459 1108
rect 1650 1083 1674 1107
rect 1859 1088 1883 1112
rect 2073 1084 2099 1110
rect 361 821 381 841
rect 572 816 596 840
rect 781 821 805 845
rect 995 817 1021 843
rect 1299 577 1319 597
rect 1510 572 1534 596
rect 1719 577 1743 601
rect 1933 573 1959 599
rect 360 267 380 287
rect 571 262 595 286
rect 780 267 804 291
rect 994 263 1020 289
rect 1408 4 1428 24
rect 1619 -1 1643 23
rect 1828 4 1852 28
rect 2042 0 2068 26
rect 361 -282 381 -262
rect 572 -287 596 -263
rect 781 -282 805 -258
rect 995 -286 1021 -260
rect 1299 -526 1319 -506
rect 1510 -531 1534 -507
rect 1719 -526 1743 -502
rect 1933 -530 1959 -504
rect 360 -836 380 -816
rect 571 -841 595 -817
rect 780 -836 804 -812
rect 994 -840 1020 -814
rect 1440 -1118 1460 -1098
rect 1651 -1123 1675 -1099
rect 1860 -1118 1884 -1094
rect 2074 -1122 2100 -1096
rect 362 -1385 382 -1365
rect 573 -1390 597 -1366
rect 782 -1385 806 -1361
rect 996 -1389 1022 -1363
rect 1300 -1629 1320 -1609
rect 1511 -1634 1535 -1610
rect 1720 -1629 1744 -1605
rect 1934 -1633 1960 -1607
rect 361 -1939 381 -1919
rect 572 -1944 596 -1920
rect 781 -1939 805 -1915
rect 995 -1943 1021 -1917
rect 1410 -2208 1430 -2188
rect 1621 -2213 1645 -2189
rect 1830 -2208 1854 -2184
rect 2044 -2212 2070 -2186
rect 362 -2488 382 -2468
rect 573 -2493 597 -2469
rect 782 -2488 806 -2464
rect 996 -2492 1022 -2466
rect 1300 -2732 1320 -2712
rect 1511 -2737 1535 -2713
rect 1720 -2732 1744 -2708
rect 1934 -2736 1960 -2710
rect 361 -3042 381 -3022
rect 572 -3047 596 -3023
rect 781 -3042 805 -3018
rect 995 -3046 1021 -3020
rect 1441 -3324 1461 -3304
rect 1652 -3329 1676 -3305
rect 1861 -3324 1885 -3300
rect 2075 -3328 2101 -3302
rect 363 -3591 383 -3571
rect 574 -3596 598 -3572
rect 783 -3591 807 -3567
rect 997 -3595 1023 -3569
rect 1301 -3835 1321 -3815
rect 1512 -3840 1536 -3816
rect 1721 -3835 1745 -3811
rect 1935 -3839 1961 -3813
rect 362 -4145 382 -4125
rect 573 -4150 597 -4126
rect 782 -4145 806 -4121
rect 996 -4149 1022 -4123
<< ndiffres >>
rect 59 4374 116 4393
rect 59 4371 80 4374
rect -35 4356 80 4371
rect 98 4356 116 4374
rect -35 4333 116 4356
rect -35 4297 7 4333
rect -36 4296 64 4297
rect -36 4275 120 4296
rect -36 4257 82 4275
rect 100 4257 120 4275
rect -36 4253 120 4257
rect 59 4237 120 4253
rect 59 4187 116 4206
rect 59 4184 80 4187
rect -35 4169 80 4184
rect 98 4169 116 4187
rect -35 4146 116 4169
rect -35 4110 7 4146
rect -36 4109 64 4110
rect -36 4088 120 4109
rect -36 4070 82 4088
rect 100 4070 120 4088
rect -36 4066 120 4070
rect 59 4050 120 4066
rect 59 3958 116 3977
rect 59 3955 80 3958
rect -35 3940 80 3955
rect 98 3940 116 3958
rect -35 3917 116 3940
rect -35 3881 7 3917
rect -36 3880 64 3881
rect -36 3859 120 3880
rect -36 3841 82 3859
rect 100 3841 120 3859
rect -36 3837 120 3841
rect 59 3821 120 3837
rect 59 3728 116 3747
rect 59 3725 80 3728
rect -35 3710 80 3725
rect 98 3710 116 3728
rect -35 3687 116 3710
rect -35 3651 7 3687
rect -36 3650 64 3651
rect -36 3629 120 3650
rect -36 3611 82 3629
rect 100 3611 120 3629
rect -36 3607 120 3611
rect 59 3591 120 3607
rect 60 3271 117 3290
rect 60 3268 81 3271
rect -34 3253 81 3268
rect 99 3253 117 3271
rect -34 3230 117 3253
rect -34 3194 8 3230
rect -35 3193 65 3194
rect -35 3172 121 3193
rect -35 3154 83 3172
rect 101 3154 121 3172
rect -35 3150 121 3154
rect 60 3134 121 3150
rect 60 3084 117 3103
rect 60 3081 81 3084
rect -34 3066 81 3081
rect 99 3066 117 3084
rect -34 3043 117 3066
rect -34 3007 8 3043
rect -35 3006 65 3007
rect -35 2985 121 3006
rect -35 2967 83 2985
rect 101 2967 121 2985
rect -35 2963 121 2967
rect 60 2947 121 2963
rect 60 2855 117 2874
rect 60 2852 81 2855
rect -34 2837 81 2852
rect 99 2837 117 2855
rect -34 2814 117 2837
rect -34 2778 8 2814
rect -35 2777 65 2778
rect -35 2756 121 2777
rect -35 2738 83 2756
rect 101 2738 121 2756
rect -35 2734 121 2738
rect 60 2718 121 2734
rect 60 2625 117 2644
rect 60 2622 81 2625
rect -34 2607 81 2622
rect 99 2607 117 2625
rect -34 2584 117 2607
rect -34 2548 8 2584
rect -35 2547 65 2548
rect -35 2526 121 2547
rect -35 2508 83 2526
rect 101 2508 121 2526
rect -35 2504 121 2508
rect 60 2488 121 2504
rect 60 2168 117 2187
rect 60 2165 81 2168
rect -34 2150 81 2165
rect 99 2150 117 2168
rect -34 2127 117 2150
rect -34 2091 8 2127
rect -35 2090 65 2091
rect -35 2069 121 2090
rect -35 2051 83 2069
rect 101 2051 121 2069
rect -35 2047 121 2051
rect 60 2031 121 2047
rect 60 1981 117 2000
rect 60 1978 81 1981
rect -34 1963 81 1978
rect 99 1963 117 1981
rect -34 1940 117 1963
rect -34 1904 8 1940
rect -35 1903 65 1904
rect -35 1882 121 1903
rect -35 1864 83 1882
rect 101 1864 121 1882
rect -35 1860 121 1864
rect 60 1844 121 1860
rect 60 1752 117 1771
rect 60 1749 81 1752
rect -34 1734 81 1749
rect 99 1734 117 1752
rect -34 1711 117 1734
rect -34 1675 8 1711
rect -35 1674 65 1675
rect -35 1653 121 1674
rect -35 1635 83 1653
rect 101 1635 121 1653
rect -35 1631 121 1635
rect 60 1615 121 1631
rect 60 1522 117 1541
rect 60 1519 81 1522
rect -34 1504 81 1519
rect 99 1504 117 1522
rect -34 1481 117 1504
rect -34 1445 8 1481
rect -35 1444 65 1445
rect -35 1423 121 1444
rect -35 1405 83 1423
rect 101 1405 121 1423
rect -35 1401 121 1405
rect 60 1385 121 1401
rect 61 1065 118 1084
rect 61 1062 82 1065
rect -33 1047 82 1062
rect 100 1047 118 1065
rect -33 1024 118 1047
rect -33 988 9 1024
rect -34 987 66 988
rect -34 966 122 987
rect -34 948 84 966
rect 102 948 122 966
rect -34 944 122 948
rect 61 928 122 944
rect 61 878 118 897
rect 61 875 82 878
rect -33 860 82 875
rect 100 860 118 878
rect -33 837 118 860
rect -33 801 9 837
rect -34 800 66 801
rect -34 779 122 800
rect -34 761 84 779
rect 102 761 122 779
rect -34 757 122 761
rect 61 741 122 757
rect 61 649 118 668
rect 61 646 82 649
rect -33 631 82 646
rect 100 631 118 649
rect -33 608 118 631
rect -33 572 9 608
rect -34 571 66 572
rect -34 550 122 571
rect -34 532 84 550
rect 102 532 122 550
rect -34 528 122 532
rect 61 512 122 528
rect 61 419 118 438
rect 61 416 82 419
rect -33 401 82 416
rect 100 401 118 419
rect -33 378 118 401
rect -33 342 9 378
rect -34 341 66 342
rect -34 320 122 341
rect -34 302 84 320
rect 102 302 122 320
rect -34 298 122 302
rect 61 282 122 298
rect 61 -38 118 -19
rect 61 -41 82 -38
rect -33 -56 82 -41
rect 100 -56 118 -38
rect -33 -79 118 -56
rect -33 -115 9 -79
rect -34 -116 66 -115
rect -34 -137 122 -116
rect -34 -155 84 -137
rect 102 -155 122 -137
rect -34 -159 122 -155
rect 61 -175 122 -159
rect 61 -225 118 -206
rect 61 -228 82 -225
rect -33 -243 82 -228
rect 100 -243 118 -225
rect -33 -266 118 -243
rect -33 -302 9 -266
rect -34 -303 66 -302
rect -34 -324 122 -303
rect -34 -342 84 -324
rect 102 -342 122 -324
rect -34 -346 122 -342
rect 61 -362 122 -346
rect 61 -454 118 -435
rect 61 -457 82 -454
rect -33 -472 82 -457
rect 100 -472 118 -454
rect -33 -495 118 -472
rect -33 -531 9 -495
rect -34 -532 66 -531
rect -34 -553 122 -532
rect -34 -571 84 -553
rect 102 -571 122 -553
rect -34 -575 122 -571
rect 61 -591 122 -575
rect 61 -684 118 -665
rect 61 -687 82 -684
rect -33 -702 82 -687
rect 100 -702 118 -684
rect -33 -725 118 -702
rect -33 -761 9 -725
rect -34 -762 66 -761
rect -34 -783 122 -762
rect -34 -801 84 -783
rect 102 -801 122 -783
rect -34 -805 122 -801
rect 61 -821 122 -805
rect 62 -1141 119 -1122
rect 62 -1144 83 -1141
rect -32 -1159 83 -1144
rect 101 -1159 119 -1141
rect -32 -1182 119 -1159
rect -32 -1218 10 -1182
rect -33 -1219 67 -1218
rect -33 -1240 123 -1219
rect -33 -1258 85 -1240
rect 103 -1258 123 -1240
rect -33 -1262 123 -1258
rect 62 -1278 123 -1262
rect 62 -1328 119 -1309
rect 62 -1331 83 -1328
rect -32 -1346 83 -1331
rect 101 -1346 119 -1328
rect -32 -1369 119 -1346
rect -32 -1405 10 -1369
rect -33 -1406 67 -1405
rect -33 -1427 123 -1406
rect -33 -1445 85 -1427
rect 103 -1445 123 -1427
rect -33 -1449 123 -1445
rect 62 -1465 123 -1449
rect 62 -1557 119 -1538
rect 62 -1560 83 -1557
rect -32 -1575 83 -1560
rect 101 -1575 119 -1557
rect -32 -1598 119 -1575
rect -32 -1634 10 -1598
rect -33 -1635 67 -1634
rect -33 -1656 123 -1635
rect -33 -1674 85 -1656
rect 103 -1674 123 -1656
rect -33 -1678 123 -1674
rect 62 -1694 123 -1678
rect 62 -1787 119 -1768
rect 62 -1790 83 -1787
rect -32 -1805 83 -1790
rect 101 -1805 119 -1787
rect -32 -1828 119 -1805
rect -32 -1864 10 -1828
rect -33 -1865 67 -1864
rect -33 -1886 123 -1865
rect -33 -1904 85 -1886
rect 103 -1904 123 -1886
rect -33 -1908 123 -1904
rect 62 -1924 123 -1908
rect 62 -2244 119 -2225
rect 62 -2247 83 -2244
rect -32 -2262 83 -2247
rect 101 -2262 119 -2244
rect -32 -2285 119 -2262
rect -32 -2321 10 -2285
rect -33 -2322 67 -2321
rect -33 -2343 123 -2322
rect -33 -2361 85 -2343
rect 103 -2361 123 -2343
rect -33 -2365 123 -2361
rect 62 -2381 123 -2365
rect 62 -2431 119 -2412
rect 62 -2434 83 -2431
rect -32 -2449 83 -2434
rect 101 -2449 119 -2431
rect -32 -2472 119 -2449
rect -32 -2508 10 -2472
rect -33 -2509 67 -2508
rect -33 -2530 123 -2509
rect -33 -2548 85 -2530
rect 103 -2548 123 -2530
rect -33 -2552 123 -2548
rect 62 -2568 123 -2552
rect 62 -2660 119 -2641
rect 62 -2663 83 -2660
rect -32 -2678 83 -2663
rect 101 -2678 119 -2660
rect -32 -2701 119 -2678
rect -32 -2737 10 -2701
rect -33 -2738 67 -2737
rect -33 -2759 123 -2738
rect -33 -2777 85 -2759
rect 103 -2777 123 -2759
rect -33 -2781 123 -2777
rect 62 -2797 123 -2781
rect 62 -2890 119 -2871
rect 62 -2893 83 -2890
rect -32 -2908 83 -2893
rect 101 -2908 119 -2890
rect -32 -2931 119 -2908
rect -32 -2967 10 -2931
rect -33 -2968 67 -2967
rect -33 -2989 123 -2968
rect -33 -3007 85 -2989
rect 103 -3007 123 -2989
rect -33 -3011 123 -3007
rect 62 -3027 123 -3011
rect 63 -3347 120 -3328
rect 63 -3350 84 -3347
rect -31 -3365 84 -3350
rect 102 -3365 120 -3347
rect -31 -3388 120 -3365
rect -31 -3424 11 -3388
rect -32 -3425 68 -3424
rect -32 -3446 124 -3425
rect -32 -3464 86 -3446
rect 104 -3464 124 -3446
rect -32 -3468 124 -3464
rect 63 -3484 124 -3468
rect 63 -3534 120 -3515
rect 63 -3537 84 -3534
rect -31 -3552 84 -3537
rect 102 -3552 120 -3534
rect -31 -3575 120 -3552
rect -31 -3611 11 -3575
rect -32 -3612 68 -3611
rect -32 -3633 124 -3612
rect -32 -3651 86 -3633
rect 104 -3651 124 -3633
rect -32 -3655 124 -3651
rect 63 -3671 124 -3655
rect 63 -3763 120 -3744
rect 63 -3766 84 -3763
rect -31 -3781 84 -3766
rect 102 -3781 120 -3763
rect -31 -3804 120 -3781
rect -31 -3840 11 -3804
rect -32 -3841 68 -3840
rect -32 -3862 124 -3841
rect -32 -3880 86 -3862
rect 104 -3880 124 -3862
rect -32 -3884 124 -3880
rect 63 -3900 124 -3884
rect 63 -3993 120 -3974
rect 63 -3996 84 -3993
rect -31 -4011 84 -3996
rect 102 -4011 120 -3993
rect -31 -4034 120 -4011
rect -31 -4070 11 -4034
rect -32 -4071 68 -4070
rect -32 -4092 124 -4071
rect -32 -4110 86 -4092
rect 104 -4110 124 -4092
rect -32 -4114 124 -4110
rect 63 -4130 124 -4114
<< locali >>
rect 69 4376 108 4433
rect 69 4374 117 4376
rect 69 4356 80 4374
rect 98 4356 117 4374
rect 69 4347 117 4356
rect 70 4346 117 4347
rect 383 4351 493 4365
rect 383 4348 426 4351
rect 383 4343 387 4348
rect 305 4321 387 4343
rect 416 4321 426 4348
rect 454 4324 461 4351
rect 490 4343 493 4351
rect 490 4324 555 4343
rect 454 4321 555 4324
rect 305 4319 555 4321
rect 73 4283 110 4284
rect 69 4280 110 4283
rect 69 4275 111 4280
rect 69 4257 82 4275
rect 100 4257 111 4275
rect 69 4243 111 4257
rect 149 4243 196 4247
rect 69 4237 196 4243
rect 69 4208 157 4237
rect 186 4208 196 4237
rect 305 4240 342 4319
rect 383 4306 493 4319
rect 457 4250 488 4251
rect 305 4220 314 4240
rect 334 4220 342 4240
rect 305 4210 342 4220
rect 401 4240 488 4250
rect 401 4220 410 4240
rect 430 4220 488 4240
rect 401 4211 488 4220
rect 401 4210 438 4211
rect 69 4204 196 4208
rect 69 4187 108 4204
rect 149 4203 196 4204
rect 69 4169 80 4187
rect 98 4169 108 4187
rect 69 4160 108 4169
rect 70 4159 107 4160
rect 457 4158 488 4211
rect 518 4240 555 4319
rect 726 4316 1119 4336
rect 1139 4316 1142 4336
rect 726 4311 1142 4316
rect 726 4310 1067 4311
rect 670 4250 701 4251
rect 518 4220 527 4240
rect 547 4220 555 4240
rect 518 4210 555 4220
rect 614 4243 701 4250
rect 614 4240 675 4243
rect 614 4220 623 4240
rect 643 4223 675 4240
rect 696 4223 701 4243
rect 643 4220 701 4223
rect 614 4213 701 4220
rect 726 4240 763 4310
rect 1029 4309 1066 4310
rect 878 4250 914 4251
rect 726 4220 735 4240
rect 755 4220 763 4240
rect 614 4211 670 4213
rect 614 4210 651 4211
rect 726 4210 763 4220
rect 822 4240 970 4250
rect 1070 4247 1166 4249
rect 822 4220 831 4240
rect 851 4220 941 4240
rect 961 4220 970 4240
rect 822 4211 970 4220
rect 1028 4240 1166 4247
rect 1028 4220 1037 4240
rect 1057 4220 1166 4240
rect 1028 4211 1166 4220
rect 822 4210 859 4211
rect 878 4159 914 4211
rect 933 4210 970 4211
rect 1029 4210 1066 4211
rect 349 4157 390 4158
rect 241 4150 390 4157
rect 241 4130 359 4150
rect 379 4130 390 4150
rect 241 4122 390 4130
rect 457 4154 816 4158
rect 457 4149 779 4154
rect 457 4125 570 4149
rect 594 4130 779 4149
rect 803 4130 816 4154
rect 594 4125 816 4130
rect 457 4122 816 4125
rect 878 4122 913 4159
rect 981 4156 1081 4159
rect 981 4152 1048 4156
rect 981 4126 993 4152
rect 1019 4130 1048 4152
rect 1074 4130 1081 4156
rect 1019 4126 1081 4130
rect 981 4122 1081 4126
rect 457 4101 488 4122
rect 878 4101 914 4122
rect 300 4100 337 4101
rect 74 4097 108 4098
rect 73 4088 110 4097
rect 73 4070 82 4088
rect 100 4070 110 4088
rect 73 4060 110 4070
rect 299 4091 337 4100
rect 299 4071 308 4091
rect 328 4071 337 4091
rect 299 4063 337 4071
rect 403 4095 488 4101
rect 513 4100 550 4101
rect 403 4075 411 4095
rect 431 4075 488 4095
rect 403 4067 488 4075
rect 512 4091 550 4100
rect 512 4071 521 4091
rect 541 4071 550 4091
rect 403 4066 439 4067
rect 512 4063 550 4071
rect 616 4095 701 4101
rect 721 4100 758 4101
rect 616 4075 624 4095
rect 644 4094 701 4095
rect 644 4075 673 4094
rect 616 4074 673 4075
rect 694 4074 701 4094
rect 616 4067 701 4074
rect 720 4091 758 4100
rect 720 4071 729 4091
rect 749 4071 758 4091
rect 616 4066 652 4067
rect 720 4063 758 4071
rect 824 4095 968 4101
rect 824 4075 832 4095
rect 852 4094 940 4095
rect 852 4075 883 4094
rect 824 4074 883 4075
rect 908 4075 940 4094
rect 960 4075 968 4095
rect 908 4074 968 4075
rect 824 4067 968 4074
rect 824 4066 860 4067
rect 932 4066 968 4067
rect 1034 4100 1071 4101
rect 1034 4099 1072 4100
rect 1034 4091 1098 4099
rect 1034 4071 1043 4091
rect 1063 4077 1098 4091
rect 1118 4077 1121 4097
rect 1063 4072 1121 4077
rect 1063 4071 1098 4072
rect 74 4032 108 4060
rect 300 4034 337 4063
rect 301 4032 337 4034
rect 513 4032 550 4063
rect 74 4031 246 4032
rect 74 3999 260 4031
rect 301 4010 550 4032
rect 721 4031 758 4063
rect 1034 4059 1098 4071
rect 1138 4033 1165 4211
rect 1321 4107 1431 4121
rect 1321 4104 1364 4107
rect 1321 4099 1325 4104
rect 997 4031 1165 4033
rect 721 4025 1165 4031
rect 74 3967 108 3999
rect 70 3958 108 3967
rect 70 3940 80 3958
rect 98 3940 108 3958
rect 70 3934 108 3940
rect 226 3936 260 3999
rect 382 4004 493 4010
rect 382 3996 423 4004
rect 382 3976 390 3996
rect 409 3976 423 3996
rect 382 3974 423 3976
rect 451 3996 493 4004
rect 451 3976 467 3996
rect 486 3976 493 3996
rect 451 3974 493 3976
rect 382 3959 493 3974
rect 720 4005 1165 4025
rect 720 3936 758 4005
rect 997 4004 1165 4005
rect 1243 4077 1325 4099
rect 1354 4077 1364 4104
rect 1392 4080 1399 4107
rect 1428 4099 1431 4107
rect 1428 4080 1493 4099
rect 1392 4077 1493 4080
rect 1243 4075 1493 4077
rect 1243 3996 1280 4075
rect 1321 4062 1431 4075
rect 1395 4006 1426 4007
rect 1243 3976 1252 3996
rect 1272 3976 1280 3996
rect 1243 3966 1280 3976
rect 1339 3996 1426 4006
rect 1339 3976 1348 3996
rect 1368 3976 1426 3996
rect 1339 3967 1426 3976
rect 1339 3966 1376 3967
rect 70 3930 107 3934
rect 226 3925 758 3936
rect 225 3909 758 3925
rect 1395 3914 1426 3967
rect 1456 3996 1493 4075
rect 1664 4072 2057 4092
rect 2077 4072 2080 4092
rect 1664 4067 2080 4072
rect 1664 4066 2005 4067
rect 1608 4006 1639 4007
rect 1456 3976 1465 3996
rect 1485 3976 1493 3996
rect 1456 3966 1493 3976
rect 1552 3999 1639 4006
rect 1552 3996 1613 3999
rect 1552 3976 1561 3996
rect 1581 3979 1613 3996
rect 1634 3979 1639 3999
rect 1581 3976 1639 3979
rect 1552 3969 1639 3976
rect 1664 3996 1701 4066
rect 1967 4065 2004 4066
rect 1816 4006 1852 4007
rect 1664 3976 1673 3996
rect 1693 3976 1701 3996
rect 1552 3967 1608 3969
rect 1552 3966 1589 3967
rect 1664 3966 1701 3976
rect 1760 3996 1908 4006
rect 2008 4003 2104 4005
rect 1760 3976 1769 3996
rect 1789 3976 1879 3996
rect 1899 3976 1908 3996
rect 1760 3967 1908 3976
rect 1966 3996 2104 4003
rect 1966 3976 1975 3996
rect 1995 3976 2104 3996
rect 1966 3967 2104 3976
rect 1760 3966 1797 3967
rect 1816 3915 1852 3967
rect 1871 3966 1908 3967
rect 1967 3966 2004 3967
rect 1287 3913 1328 3914
rect 225 3908 739 3909
rect 1179 3906 1328 3913
rect 1179 3886 1297 3906
rect 1317 3886 1328 3906
rect 1179 3878 1328 3886
rect 1395 3910 1754 3914
rect 1395 3905 1717 3910
rect 1395 3881 1508 3905
rect 1532 3886 1717 3905
rect 1741 3886 1754 3910
rect 1532 3881 1754 3886
rect 1395 3878 1754 3881
rect 1816 3878 1851 3915
rect 1919 3912 2019 3915
rect 1919 3908 1986 3912
rect 1919 3882 1931 3908
rect 1957 3886 1986 3908
rect 2012 3886 2019 3912
rect 1957 3882 2019 3886
rect 1919 3878 2019 3882
rect 73 3867 110 3868
rect 71 3859 111 3867
rect 71 3841 82 3859
rect 100 3841 111 3859
rect 1395 3857 1426 3878
rect 1816 3857 1852 3878
rect 1238 3856 1275 3857
rect 71 3793 111 3841
rect 1237 3847 1275 3856
rect 1237 3827 1246 3847
rect 1266 3827 1275 3847
rect 1237 3819 1275 3827
rect 1341 3851 1426 3857
rect 1451 3856 1488 3857
rect 1341 3831 1349 3851
rect 1369 3831 1426 3851
rect 1341 3823 1426 3831
rect 1450 3847 1488 3856
rect 1450 3827 1459 3847
rect 1479 3827 1488 3847
rect 1341 3822 1377 3823
rect 1450 3819 1488 3827
rect 1554 3851 1639 3857
rect 1659 3856 1696 3857
rect 1554 3831 1562 3851
rect 1582 3850 1639 3851
rect 1582 3831 1611 3850
rect 1554 3830 1611 3831
rect 1632 3830 1639 3850
rect 1554 3823 1639 3830
rect 1658 3847 1696 3856
rect 1658 3827 1667 3847
rect 1687 3827 1696 3847
rect 1554 3822 1590 3823
rect 1658 3819 1696 3827
rect 1762 3851 1906 3857
rect 1762 3831 1770 3851
rect 1790 3834 1826 3851
rect 1846 3834 1878 3851
rect 1790 3831 1878 3834
rect 1898 3831 1906 3851
rect 1762 3823 1906 3831
rect 1762 3822 1798 3823
rect 1870 3822 1906 3823
rect 1972 3856 2009 3857
rect 1972 3855 2010 3856
rect 1972 3847 2036 3855
rect 1972 3827 1981 3847
rect 2001 3833 2036 3847
rect 2056 3833 2059 3853
rect 2001 3828 2059 3833
rect 2001 3827 2036 3828
rect 382 3797 492 3811
rect 382 3794 425 3797
rect 71 3786 196 3793
rect 382 3789 386 3794
rect 71 3767 163 3786
rect 188 3767 196 3786
rect 71 3757 196 3767
rect 304 3767 386 3789
rect 415 3767 425 3794
rect 453 3770 460 3797
rect 489 3789 492 3797
rect 1238 3790 1275 3819
rect 489 3770 554 3789
rect 1239 3788 1275 3790
rect 1451 3788 1488 3819
rect 1659 3792 1696 3819
rect 1972 3815 2036 3827
rect 453 3767 554 3770
rect 304 3765 554 3767
rect 71 3737 111 3757
rect 70 3728 111 3737
rect 70 3710 80 3728
rect 98 3710 111 3728
rect 70 3701 111 3710
rect 70 3700 107 3701
rect 304 3686 341 3765
rect 382 3752 492 3765
rect 456 3696 487 3697
rect 304 3666 313 3686
rect 333 3666 341 3686
rect 304 3656 341 3666
rect 400 3686 487 3696
rect 400 3666 409 3686
rect 429 3666 487 3686
rect 400 3657 487 3666
rect 400 3656 437 3657
rect 73 3634 110 3638
rect 70 3629 110 3634
rect 70 3611 82 3629
rect 100 3611 110 3629
rect 70 3431 110 3611
rect 456 3604 487 3657
rect 517 3686 554 3765
rect 725 3762 1118 3782
rect 1138 3762 1141 3782
rect 1239 3766 1488 3788
rect 1657 3787 1698 3792
rect 2076 3789 2103 3967
rect 1935 3787 2103 3789
rect 1657 3781 2103 3787
rect 725 3757 1141 3762
rect 1320 3760 1431 3766
rect 725 3756 1066 3757
rect 669 3696 700 3697
rect 517 3666 526 3686
rect 546 3666 554 3686
rect 517 3656 554 3666
rect 613 3689 700 3696
rect 613 3686 674 3689
rect 613 3666 622 3686
rect 642 3669 674 3686
rect 695 3669 700 3689
rect 642 3666 700 3669
rect 613 3659 700 3666
rect 725 3686 762 3756
rect 1028 3755 1065 3756
rect 1320 3752 1361 3760
rect 1320 3732 1328 3752
rect 1347 3732 1361 3752
rect 1320 3730 1361 3732
rect 1389 3752 1431 3760
rect 1389 3732 1405 3752
rect 1424 3732 1431 3752
rect 1657 3759 1663 3781
rect 1689 3761 2103 3781
rect 1689 3759 1698 3761
rect 1935 3760 2103 3761
rect 1657 3750 1698 3759
rect 1389 3730 1431 3732
rect 1320 3715 1431 3730
rect 877 3696 913 3697
rect 725 3666 734 3686
rect 754 3666 762 3686
rect 613 3657 669 3659
rect 613 3656 650 3657
rect 725 3656 762 3666
rect 821 3686 969 3696
rect 1069 3693 1165 3695
rect 821 3666 830 3686
rect 850 3666 940 3686
rect 960 3666 969 3686
rect 821 3657 969 3666
rect 1027 3686 1165 3693
rect 1027 3666 1036 3686
rect 1056 3666 1165 3686
rect 1027 3657 1165 3666
rect 821 3656 858 3657
rect 877 3605 913 3657
rect 932 3656 969 3657
rect 1028 3656 1065 3657
rect 348 3603 389 3604
rect 240 3596 389 3603
rect 240 3576 358 3596
rect 378 3576 389 3596
rect 240 3568 389 3576
rect 456 3600 815 3604
rect 456 3595 778 3600
rect 456 3571 569 3595
rect 593 3576 778 3595
rect 802 3576 815 3600
rect 593 3571 815 3576
rect 456 3568 815 3571
rect 877 3568 912 3605
rect 980 3602 1080 3605
rect 980 3598 1047 3602
rect 980 3572 992 3598
rect 1018 3576 1047 3598
rect 1073 3576 1080 3602
rect 1018 3572 1080 3576
rect 980 3568 1080 3572
rect 456 3547 487 3568
rect 877 3547 913 3568
rect 299 3546 336 3547
rect 298 3537 336 3546
rect 298 3517 307 3537
rect 327 3517 336 3537
rect 298 3509 336 3517
rect 402 3541 487 3547
rect 512 3546 549 3547
rect 402 3521 410 3541
rect 430 3521 487 3541
rect 402 3513 487 3521
rect 511 3537 549 3546
rect 511 3517 520 3537
rect 540 3517 549 3537
rect 402 3512 438 3513
rect 511 3509 549 3517
rect 615 3541 700 3547
rect 720 3546 757 3547
rect 615 3521 623 3541
rect 643 3540 700 3541
rect 643 3521 672 3540
rect 615 3520 672 3521
rect 693 3520 700 3540
rect 615 3513 700 3520
rect 719 3537 757 3546
rect 719 3517 728 3537
rect 748 3517 757 3537
rect 615 3512 651 3513
rect 719 3509 757 3517
rect 823 3541 967 3547
rect 823 3521 831 3541
rect 851 3538 939 3541
rect 851 3521 882 3538
rect 823 3518 882 3521
rect 905 3521 939 3538
rect 959 3521 967 3541
rect 905 3518 967 3521
rect 823 3513 967 3518
rect 823 3512 859 3513
rect 931 3512 967 3513
rect 1033 3546 1070 3547
rect 1033 3545 1071 3546
rect 1033 3537 1097 3545
rect 1033 3517 1042 3537
rect 1062 3523 1097 3537
rect 1117 3523 1120 3543
rect 1062 3518 1120 3523
rect 1062 3517 1097 3518
rect 299 3480 336 3509
rect 300 3478 336 3480
rect 512 3478 549 3509
rect 300 3456 549 3478
rect 720 3477 757 3509
rect 1033 3505 1097 3517
rect 1137 3479 1164 3657
rect 1462 3515 1572 3529
rect 1462 3512 1505 3515
rect 1462 3507 1466 3512
rect 996 3477 1164 3479
rect 720 3474 1164 3477
rect 381 3450 492 3456
rect 381 3442 422 3450
rect 70 3387 109 3431
rect 381 3422 389 3442
rect 408 3422 422 3442
rect 381 3420 422 3422
rect 450 3442 492 3450
rect 450 3422 466 3442
rect 485 3422 492 3442
rect 450 3420 492 3422
rect 381 3405 492 3420
rect 718 3451 1164 3474
rect 70 3363 110 3387
rect 410 3363 457 3365
rect 718 3363 756 3451
rect 996 3450 1164 3451
rect 1384 3485 1466 3507
rect 1495 3485 1505 3512
rect 1533 3488 1540 3515
rect 1569 3507 1572 3515
rect 1569 3488 1634 3507
rect 1533 3485 1634 3488
rect 1384 3483 1634 3485
rect 1384 3404 1421 3483
rect 1462 3470 1572 3483
rect 1536 3414 1567 3415
rect 1384 3384 1393 3404
rect 1413 3384 1421 3404
rect 1384 3374 1421 3384
rect 1480 3404 1567 3414
rect 1480 3384 1489 3404
rect 1509 3384 1567 3404
rect 1480 3375 1567 3384
rect 1480 3374 1517 3375
rect 70 3330 756 3363
rect 70 3273 109 3330
rect 718 3328 756 3330
rect 1536 3322 1567 3375
rect 1597 3404 1634 3483
rect 1805 3496 2198 3500
rect 1805 3479 1824 3496
rect 1844 3480 2198 3496
rect 2218 3480 2221 3500
rect 1844 3479 2221 3480
rect 1805 3475 2221 3479
rect 1805 3474 2146 3475
rect 1749 3414 1780 3415
rect 1597 3384 1606 3404
rect 1626 3384 1634 3404
rect 1597 3374 1634 3384
rect 1693 3407 1780 3414
rect 1693 3404 1754 3407
rect 1693 3384 1702 3404
rect 1722 3387 1754 3404
rect 1775 3387 1780 3407
rect 1722 3384 1780 3387
rect 1693 3377 1780 3384
rect 1805 3404 1842 3474
rect 2108 3473 2145 3474
rect 1957 3414 1993 3415
rect 1805 3384 1814 3404
rect 1834 3384 1842 3404
rect 1693 3375 1749 3377
rect 1693 3374 1730 3375
rect 1805 3374 1842 3384
rect 1901 3404 2049 3414
rect 2149 3411 2245 3413
rect 1901 3384 1910 3404
rect 1930 3384 2020 3404
rect 2040 3384 2049 3404
rect 1901 3375 2049 3384
rect 2107 3404 2245 3411
rect 2107 3384 2116 3404
rect 2136 3384 2245 3404
rect 2107 3375 2245 3384
rect 1901 3374 1938 3375
rect 1957 3323 1993 3375
rect 2012 3374 2049 3375
rect 2108 3374 2145 3375
rect 1428 3321 1469 3322
rect 1320 3314 1469 3321
rect 1320 3294 1438 3314
rect 1458 3294 1469 3314
rect 1320 3286 1469 3294
rect 1536 3318 1895 3322
rect 1536 3313 1858 3318
rect 1536 3289 1649 3313
rect 1673 3294 1858 3313
rect 1882 3294 1895 3318
rect 1673 3289 1895 3294
rect 1536 3286 1895 3289
rect 1957 3286 1992 3323
rect 2060 3320 2160 3323
rect 2060 3316 2127 3320
rect 2060 3290 2072 3316
rect 2098 3294 2127 3316
rect 2153 3294 2160 3320
rect 2098 3290 2160 3294
rect 2060 3286 2160 3290
rect 70 3271 118 3273
rect 70 3253 81 3271
rect 99 3253 118 3271
rect 1536 3265 1567 3286
rect 1957 3265 1993 3286
rect 1379 3264 1416 3265
rect 70 3244 118 3253
rect 71 3243 118 3244
rect 384 3248 494 3262
rect 384 3245 427 3248
rect 384 3240 388 3245
rect 306 3218 388 3240
rect 417 3218 427 3245
rect 455 3221 462 3248
rect 491 3240 494 3248
rect 1378 3255 1416 3264
rect 491 3221 556 3240
rect 1378 3235 1387 3255
rect 1407 3235 1416 3255
rect 455 3218 556 3221
rect 306 3216 556 3218
rect 74 3180 111 3181
rect 70 3177 111 3180
rect 70 3172 112 3177
rect 70 3154 83 3172
rect 101 3154 112 3172
rect 70 3140 112 3154
rect 150 3140 197 3144
rect 70 3134 197 3140
rect 70 3105 158 3134
rect 187 3105 197 3134
rect 306 3137 343 3216
rect 384 3203 494 3216
rect 458 3147 489 3148
rect 306 3117 315 3137
rect 335 3117 343 3137
rect 306 3107 343 3117
rect 402 3137 489 3147
rect 402 3117 411 3137
rect 431 3117 489 3137
rect 402 3108 489 3117
rect 402 3107 439 3108
rect 70 3101 197 3105
rect 70 3084 109 3101
rect 150 3100 197 3101
rect 70 3066 81 3084
rect 99 3066 109 3084
rect 70 3057 109 3066
rect 71 3056 108 3057
rect 458 3055 489 3108
rect 519 3137 556 3216
rect 727 3213 1120 3233
rect 1140 3213 1143 3233
rect 1378 3227 1416 3235
rect 1482 3259 1567 3265
rect 1592 3264 1629 3265
rect 1482 3239 1490 3259
rect 1510 3239 1567 3259
rect 1482 3231 1567 3239
rect 1591 3255 1629 3264
rect 1591 3235 1600 3255
rect 1620 3235 1629 3255
rect 1482 3230 1518 3231
rect 1591 3227 1629 3235
rect 1695 3259 1780 3265
rect 1800 3264 1837 3265
rect 1695 3239 1703 3259
rect 1723 3258 1780 3259
rect 1723 3239 1752 3258
rect 1695 3238 1752 3239
rect 1773 3238 1780 3258
rect 1695 3231 1780 3238
rect 1799 3255 1837 3264
rect 1799 3235 1808 3255
rect 1828 3235 1837 3255
rect 1695 3230 1731 3231
rect 1799 3227 1837 3235
rect 1903 3259 2047 3265
rect 1903 3239 1911 3259
rect 1931 3257 2019 3259
rect 1931 3239 1960 3257
rect 1903 3236 1960 3239
rect 1987 3239 2019 3257
rect 2039 3239 2047 3259
rect 1987 3236 2047 3239
rect 1903 3231 2047 3236
rect 1903 3230 1939 3231
rect 2011 3230 2047 3231
rect 2113 3264 2150 3265
rect 2113 3263 2151 3264
rect 2113 3255 2177 3263
rect 2113 3235 2122 3255
rect 2142 3241 2177 3255
rect 2197 3241 2200 3261
rect 2142 3236 2200 3241
rect 2142 3235 2177 3236
rect 727 3208 1143 3213
rect 727 3207 1068 3208
rect 671 3147 702 3148
rect 519 3117 528 3137
rect 548 3117 556 3137
rect 519 3107 556 3117
rect 615 3140 702 3147
rect 615 3137 676 3140
rect 615 3117 624 3137
rect 644 3120 676 3137
rect 697 3120 702 3140
rect 644 3117 702 3120
rect 615 3110 702 3117
rect 727 3137 764 3207
rect 1030 3206 1067 3207
rect 1379 3198 1416 3227
rect 1380 3196 1416 3198
rect 1592 3196 1629 3227
rect 1380 3174 1629 3196
rect 1800 3195 1837 3227
rect 2113 3223 2177 3235
rect 2217 3197 2244 3375
rect 2076 3195 2244 3197
rect 1797 3188 2244 3195
rect 1461 3168 1572 3174
rect 1461 3160 1502 3168
rect 879 3147 915 3148
rect 727 3117 736 3137
rect 756 3117 764 3137
rect 615 3108 671 3110
rect 615 3107 652 3108
rect 727 3107 764 3117
rect 823 3137 971 3147
rect 1071 3144 1167 3146
rect 823 3117 832 3137
rect 852 3117 942 3137
rect 962 3117 971 3137
rect 823 3108 971 3117
rect 1029 3137 1167 3144
rect 1029 3117 1038 3137
rect 1058 3117 1167 3137
rect 1461 3140 1469 3160
rect 1488 3140 1502 3160
rect 1461 3138 1502 3140
rect 1530 3160 1572 3168
rect 1530 3140 1546 3160
rect 1565 3140 1572 3160
rect 1797 3161 1822 3188
rect 1853 3169 2244 3188
rect 1853 3161 1902 3169
rect 2076 3168 2244 3169
rect 1797 3159 1902 3161
rect 1530 3138 1572 3140
rect 1461 3123 1572 3138
rect 1029 3108 1167 3117
rect 823 3107 860 3108
rect 879 3056 915 3108
rect 934 3107 971 3108
rect 1030 3107 1067 3108
rect 350 3054 391 3055
rect 242 3047 391 3054
rect 242 3027 360 3047
rect 380 3027 391 3047
rect 242 3019 391 3027
rect 458 3051 817 3055
rect 458 3046 780 3051
rect 458 3022 571 3046
rect 595 3027 780 3046
rect 804 3027 817 3051
rect 595 3022 817 3027
rect 458 3019 817 3022
rect 879 3019 914 3056
rect 982 3053 1082 3056
rect 982 3049 1049 3053
rect 982 3023 994 3049
rect 1020 3027 1049 3049
rect 1075 3027 1082 3053
rect 1020 3023 1082 3027
rect 982 3019 1082 3023
rect 458 2998 489 3019
rect 879 2998 915 3019
rect 301 2997 338 2998
rect 75 2994 109 2995
rect 74 2985 111 2994
rect 74 2967 83 2985
rect 101 2967 111 2985
rect 74 2957 111 2967
rect 300 2988 338 2997
rect 300 2968 309 2988
rect 329 2968 338 2988
rect 300 2960 338 2968
rect 404 2992 489 2998
rect 514 2997 551 2998
rect 404 2972 412 2992
rect 432 2972 489 2992
rect 404 2964 489 2972
rect 513 2988 551 2997
rect 513 2968 522 2988
rect 542 2968 551 2988
rect 404 2963 440 2964
rect 513 2960 551 2968
rect 617 2992 702 2998
rect 722 2997 759 2998
rect 617 2972 625 2992
rect 645 2991 702 2992
rect 645 2972 674 2991
rect 617 2971 674 2972
rect 695 2971 702 2991
rect 617 2964 702 2971
rect 721 2988 759 2997
rect 721 2968 730 2988
rect 750 2968 759 2988
rect 617 2963 653 2964
rect 721 2960 759 2968
rect 825 2992 969 2998
rect 825 2972 833 2992
rect 853 2991 941 2992
rect 853 2972 884 2991
rect 825 2971 884 2972
rect 909 2972 941 2991
rect 961 2972 969 2992
rect 909 2971 969 2972
rect 825 2964 969 2971
rect 825 2963 861 2964
rect 933 2963 969 2964
rect 1035 2997 1072 2998
rect 1035 2996 1073 2997
rect 1035 2988 1099 2996
rect 1035 2968 1044 2988
rect 1064 2974 1099 2988
rect 1119 2974 1122 2994
rect 1064 2969 1122 2974
rect 1064 2968 1099 2969
rect 75 2929 109 2957
rect 301 2931 338 2960
rect 302 2929 338 2931
rect 514 2929 551 2960
rect 75 2928 247 2929
rect 75 2896 261 2928
rect 302 2907 551 2929
rect 722 2928 759 2960
rect 1035 2956 1099 2968
rect 1139 2930 1166 3108
rect 1322 3004 1432 3018
rect 1322 3001 1365 3004
rect 1322 2996 1326 3001
rect 998 2928 1166 2930
rect 722 2922 1166 2928
rect 75 2864 109 2896
rect 71 2855 109 2864
rect 71 2837 81 2855
rect 99 2837 109 2855
rect 71 2831 109 2837
rect 227 2833 261 2896
rect 383 2901 494 2907
rect 383 2893 424 2901
rect 383 2873 391 2893
rect 410 2873 424 2893
rect 383 2871 424 2873
rect 452 2893 494 2901
rect 452 2873 468 2893
rect 487 2873 494 2893
rect 452 2871 494 2873
rect 383 2856 494 2871
rect 721 2902 1166 2922
rect 721 2833 759 2902
rect 998 2901 1166 2902
rect 1244 2974 1326 2996
rect 1355 2974 1365 3001
rect 1393 2977 1400 3004
rect 1429 2996 1432 3004
rect 1429 2977 1494 2996
rect 1393 2974 1494 2977
rect 1244 2972 1494 2974
rect 1244 2893 1281 2972
rect 1322 2959 1432 2972
rect 1396 2903 1427 2904
rect 1244 2873 1253 2893
rect 1273 2873 1281 2893
rect 1244 2863 1281 2873
rect 1340 2893 1427 2903
rect 1340 2873 1349 2893
rect 1369 2873 1427 2893
rect 1340 2864 1427 2873
rect 1340 2863 1377 2864
rect 71 2827 108 2831
rect 227 2822 759 2833
rect 226 2806 759 2822
rect 1396 2811 1427 2864
rect 1457 2893 1494 2972
rect 1665 2982 2058 2989
rect 1665 2965 1673 2982
rect 1705 2969 2058 2982
rect 2078 2969 2081 2989
rect 1705 2965 2081 2969
rect 1665 2964 2081 2965
rect 1665 2963 2006 2964
rect 1609 2903 1640 2904
rect 1457 2873 1466 2893
rect 1486 2873 1494 2893
rect 1457 2863 1494 2873
rect 1553 2896 1640 2903
rect 1553 2893 1614 2896
rect 1553 2873 1562 2893
rect 1582 2876 1614 2893
rect 1635 2876 1640 2896
rect 1582 2873 1640 2876
rect 1553 2866 1640 2873
rect 1665 2893 1702 2963
rect 1968 2962 2005 2963
rect 1817 2903 1853 2904
rect 1665 2873 1674 2893
rect 1694 2873 1702 2893
rect 1553 2864 1609 2866
rect 1553 2863 1590 2864
rect 1665 2863 1702 2873
rect 1761 2893 1909 2903
rect 2009 2900 2105 2902
rect 1761 2873 1770 2893
rect 1790 2888 1880 2893
rect 1790 2873 1825 2888
rect 1761 2864 1825 2873
rect 1761 2863 1798 2864
rect 1817 2847 1825 2864
rect 1846 2873 1880 2888
rect 1900 2873 1909 2893
rect 1846 2864 1909 2873
rect 1967 2893 2105 2900
rect 1967 2873 1976 2893
rect 1996 2873 2105 2893
rect 1967 2864 2105 2873
rect 1846 2847 1853 2864
rect 1872 2863 1909 2864
rect 1968 2863 2005 2864
rect 1817 2812 1853 2847
rect 1288 2810 1329 2811
rect 226 2805 740 2806
rect 1180 2803 1329 2810
rect 1180 2783 1298 2803
rect 1318 2783 1329 2803
rect 1180 2775 1329 2783
rect 1396 2807 1755 2811
rect 1396 2802 1718 2807
rect 1396 2778 1509 2802
rect 1533 2783 1718 2802
rect 1742 2783 1755 2807
rect 1533 2778 1755 2783
rect 1396 2775 1755 2778
rect 1817 2775 1852 2812
rect 1920 2809 2020 2812
rect 1920 2805 1987 2809
rect 1920 2779 1932 2805
rect 1958 2783 1987 2805
rect 2013 2783 2020 2809
rect 1958 2779 2020 2783
rect 1920 2775 2020 2779
rect 74 2764 111 2765
rect 72 2756 112 2764
rect 72 2738 83 2756
rect 101 2738 112 2756
rect 1396 2754 1427 2775
rect 1817 2754 1853 2775
rect 1239 2753 1276 2754
rect 72 2690 112 2738
rect 1238 2744 1276 2753
rect 1238 2724 1247 2744
rect 1267 2724 1276 2744
rect 1238 2716 1276 2724
rect 1342 2748 1427 2754
rect 1452 2753 1489 2754
rect 1342 2728 1350 2748
rect 1370 2728 1427 2748
rect 1342 2720 1427 2728
rect 1451 2744 1489 2753
rect 1451 2724 1460 2744
rect 1480 2724 1489 2744
rect 1342 2719 1378 2720
rect 1451 2716 1489 2724
rect 1555 2748 1640 2754
rect 1660 2753 1697 2754
rect 1555 2728 1563 2748
rect 1583 2747 1640 2748
rect 1583 2728 1612 2747
rect 1555 2727 1612 2728
rect 1633 2727 1640 2747
rect 1555 2720 1640 2727
rect 1659 2744 1697 2753
rect 1659 2724 1668 2744
rect 1688 2724 1697 2744
rect 1555 2719 1591 2720
rect 1659 2716 1697 2724
rect 1763 2748 1907 2754
rect 1763 2728 1771 2748
rect 1791 2728 1879 2748
rect 1899 2728 1907 2748
rect 1763 2720 1907 2728
rect 1763 2719 1799 2720
rect 1871 2719 1907 2720
rect 1973 2753 2010 2754
rect 1973 2752 2011 2753
rect 1973 2744 2037 2752
rect 1973 2724 1982 2744
rect 2002 2730 2037 2744
rect 2057 2730 2060 2750
rect 2002 2725 2060 2730
rect 2002 2724 2037 2725
rect 383 2694 493 2708
rect 383 2691 426 2694
rect 72 2683 197 2690
rect 383 2686 387 2691
rect 72 2664 164 2683
rect 189 2664 197 2683
rect 72 2654 197 2664
rect 305 2664 387 2686
rect 416 2664 426 2691
rect 454 2667 461 2694
rect 490 2686 493 2694
rect 1239 2687 1276 2716
rect 490 2667 555 2686
rect 1240 2685 1276 2687
rect 1452 2685 1489 2716
rect 1660 2689 1697 2716
rect 1973 2712 2037 2724
rect 454 2664 555 2667
rect 305 2662 555 2664
rect 72 2634 112 2654
rect 71 2625 112 2634
rect 71 2607 81 2625
rect 99 2607 112 2625
rect 71 2598 112 2607
rect 71 2597 108 2598
rect 305 2583 342 2662
rect 383 2649 493 2662
rect 457 2593 488 2594
rect 305 2563 314 2583
rect 334 2563 342 2583
rect 305 2553 342 2563
rect 401 2583 488 2593
rect 401 2563 410 2583
rect 430 2563 488 2583
rect 401 2554 488 2563
rect 401 2553 438 2554
rect 74 2531 111 2535
rect 71 2526 111 2531
rect 71 2508 83 2526
rect 101 2508 111 2526
rect 71 2328 111 2508
rect 457 2501 488 2554
rect 518 2583 555 2662
rect 726 2659 1119 2679
rect 1139 2659 1142 2679
rect 1240 2663 1489 2685
rect 1658 2684 1699 2689
rect 2077 2686 2104 2864
rect 1936 2684 2104 2686
rect 1658 2678 2104 2684
rect 726 2654 1142 2659
rect 1321 2657 1432 2663
rect 726 2653 1067 2654
rect 670 2593 701 2594
rect 518 2563 527 2583
rect 547 2563 555 2583
rect 518 2553 555 2563
rect 614 2586 701 2593
rect 614 2583 675 2586
rect 614 2563 623 2583
rect 643 2566 675 2583
rect 696 2566 701 2586
rect 643 2563 701 2566
rect 614 2556 701 2563
rect 726 2583 763 2653
rect 1029 2652 1066 2653
rect 1321 2649 1362 2657
rect 1321 2629 1329 2649
rect 1348 2629 1362 2649
rect 1321 2627 1362 2629
rect 1390 2649 1432 2657
rect 1390 2629 1406 2649
rect 1425 2629 1432 2649
rect 1658 2656 1664 2678
rect 1690 2658 2104 2678
rect 1690 2656 1699 2658
rect 1936 2657 2104 2658
rect 1658 2647 1699 2656
rect 1390 2627 1432 2629
rect 1321 2612 1432 2627
rect 878 2593 914 2594
rect 726 2563 735 2583
rect 755 2563 763 2583
rect 614 2554 670 2556
rect 614 2553 651 2554
rect 726 2553 763 2563
rect 822 2583 970 2593
rect 1070 2590 1166 2592
rect 822 2563 831 2583
rect 851 2563 941 2583
rect 961 2563 970 2583
rect 822 2554 970 2563
rect 1028 2583 1166 2590
rect 1028 2563 1037 2583
rect 1057 2563 1166 2583
rect 1028 2554 1166 2563
rect 822 2553 859 2554
rect 878 2502 914 2554
rect 933 2553 970 2554
rect 1029 2553 1066 2554
rect 349 2500 390 2501
rect 241 2493 390 2500
rect 241 2473 359 2493
rect 379 2473 390 2493
rect 241 2465 390 2473
rect 457 2497 816 2501
rect 457 2492 779 2497
rect 457 2468 570 2492
rect 594 2473 779 2492
rect 803 2473 816 2497
rect 594 2468 816 2473
rect 457 2465 816 2468
rect 878 2465 913 2502
rect 981 2499 1081 2502
rect 981 2495 1048 2499
rect 981 2469 993 2495
rect 1019 2473 1048 2495
rect 1074 2473 1081 2499
rect 1019 2469 1081 2473
rect 981 2465 1081 2469
rect 457 2444 488 2465
rect 878 2444 914 2465
rect 300 2443 337 2444
rect 299 2434 337 2443
rect 299 2414 308 2434
rect 328 2414 337 2434
rect 299 2406 337 2414
rect 403 2438 488 2444
rect 513 2443 550 2444
rect 403 2418 411 2438
rect 431 2418 488 2438
rect 403 2410 488 2418
rect 512 2434 550 2443
rect 512 2414 521 2434
rect 541 2414 550 2434
rect 403 2409 439 2410
rect 512 2406 550 2414
rect 616 2438 701 2444
rect 721 2443 758 2444
rect 616 2418 624 2438
rect 644 2437 701 2438
rect 644 2418 673 2437
rect 616 2417 673 2418
rect 694 2417 701 2437
rect 616 2410 701 2417
rect 720 2434 758 2443
rect 720 2414 729 2434
rect 749 2414 758 2434
rect 616 2409 652 2410
rect 720 2406 758 2414
rect 824 2438 968 2444
rect 824 2418 832 2438
rect 852 2435 940 2438
rect 852 2418 883 2435
rect 824 2415 883 2418
rect 906 2418 940 2435
rect 960 2418 968 2438
rect 906 2415 968 2418
rect 824 2410 968 2415
rect 824 2409 860 2410
rect 932 2409 968 2410
rect 1034 2443 1071 2444
rect 1034 2442 1072 2443
rect 1034 2434 1098 2442
rect 1034 2414 1043 2434
rect 1063 2420 1098 2434
rect 1118 2420 1121 2440
rect 1063 2415 1121 2420
rect 1063 2414 1098 2415
rect 300 2377 337 2406
rect 301 2375 337 2377
rect 513 2375 550 2406
rect 301 2353 550 2375
rect 721 2374 758 2406
rect 1034 2402 1098 2414
rect 1138 2376 1165 2554
rect 1432 2425 1542 2439
rect 1432 2422 1475 2425
rect 1432 2417 1436 2422
rect 997 2374 1165 2376
rect 721 2371 1165 2374
rect 382 2347 493 2353
rect 382 2339 423 2347
rect 71 2284 110 2328
rect 382 2319 390 2339
rect 409 2319 423 2339
rect 382 2317 423 2319
rect 451 2339 493 2347
rect 451 2319 467 2339
rect 486 2319 493 2339
rect 451 2317 493 2319
rect 382 2303 493 2317
rect 719 2348 1165 2371
rect 71 2260 111 2284
rect 411 2260 458 2262
rect 719 2260 757 2348
rect 997 2347 1165 2348
rect 1354 2395 1436 2417
rect 1465 2395 1475 2422
rect 1503 2398 1510 2425
rect 1539 2417 1542 2425
rect 1539 2398 1604 2417
rect 1503 2395 1604 2398
rect 1354 2393 1604 2395
rect 1354 2314 1391 2393
rect 1432 2380 1542 2393
rect 1506 2324 1537 2325
rect 1354 2294 1363 2314
rect 1383 2294 1391 2314
rect 1354 2284 1391 2294
rect 1450 2314 1537 2324
rect 1450 2294 1459 2314
rect 1479 2294 1537 2314
rect 1450 2285 1537 2294
rect 1450 2284 1487 2285
rect 71 2227 757 2260
rect 1506 2232 1537 2285
rect 1567 2314 1604 2393
rect 1775 2390 2168 2410
rect 2188 2390 2191 2410
rect 1775 2385 2191 2390
rect 1775 2384 2116 2385
rect 1719 2324 1750 2325
rect 1567 2294 1576 2314
rect 1596 2294 1604 2314
rect 1567 2284 1604 2294
rect 1663 2317 1750 2324
rect 1663 2314 1724 2317
rect 1663 2294 1672 2314
rect 1692 2297 1724 2314
rect 1745 2297 1750 2317
rect 1692 2294 1750 2297
rect 1663 2287 1750 2294
rect 1775 2314 1812 2384
rect 2078 2383 2115 2384
rect 1927 2324 1963 2325
rect 1775 2294 1784 2314
rect 1804 2294 1812 2314
rect 1663 2285 1719 2287
rect 1663 2284 1700 2285
rect 1775 2284 1812 2294
rect 1871 2314 2019 2324
rect 2119 2321 2215 2323
rect 1871 2294 1880 2314
rect 1900 2294 1990 2314
rect 2010 2294 2019 2314
rect 1871 2285 2019 2294
rect 2077 2314 2215 2321
rect 2077 2294 2086 2314
rect 2106 2294 2215 2314
rect 2077 2285 2215 2294
rect 1871 2284 1908 2285
rect 1927 2233 1963 2285
rect 1982 2284 2019 2285
rect 2078 2284 2115 2285
rect 1398 2231 1439 2232
rect 70 2170 109 2227
rect 719 2225 757 2227
rect 1290 2224 1439 2231
rect 1290 2204 1408 2224
rect 1428 2204 1439 2224
rect 1290 2196 1439 2204
rect 1506 2228 1865 2232
rect 1506 2223 1828 2228
rect 1506 2199 1619 2223
rect 1643 2204 1828 2223
rect 1852 2204 1865 2228
rect 1643 2199 1865 2204
rect 1506 2196 1865 2199
rect 1927 2196 1962 2233
rect 2030 2230 2130 2233
rect 2030 2226 2097 2230
rect 2030 2200 2042 2226
rect 2068 2204 2097 2226
rect 2123 2204 2130 2230
rect 2068 2200 2130 2204
rect 2030 2196 2130 2200
rect 1506 2175 1537 2196
rect 1927 2175 1963 2196
rect 1349 2174 1386 2175
rect 70 2168 118 2170
rect 70 2150 81 2168
rect 99 2150 118 2168
rect 1348 2165 1386 2174
rect 70 2141 118 2150
rect 71 2140 118 2141
rect 384 2145 494 2159
rect 384 2142 427 2145
rect 384 2137 388 2142
rect 306 2115 388 2137
rect 417 2115 427 2142
rect 455 2118 462 2145
rect 491 2137 494 2145
rect 1348 2145 1357 2165
rect 1377 2145 1386 2165
rect 1348 2137 1386 2145
rect 1452 2169 1537 2175
rect 1562 2174 1599 2175
rect 1452 2149 1460 2169
rect 1480 2149 1537 2169
rect 1452 2141 1537 2149
rect 1561 2165 1599 2174
rect 1561 2145 1570 2165
rect 1590 2145 1599 2165
rect 1452 2140 1488 2141
rect 1561 2137 1599 2145
rect 1665 2169 1750 2175
rect 1770 2174 1807 2175
rect 1665 2149 1673 2169
rect 1693 2168 1750 2169
rect 1693 2149 1722 2168
rect 1665 2148 1722 2149
rect 1743 2148 1750 2168
rect 1665 2141 1750 2148
rect 1769 2165 1807 2174
rect 1769 2145 1778 2165
rect 1798 2145 1807 2165
rect 1665 2140 1701 2141
rect 1769 2137 1807 2145
rect 1873 2169 2017 2175
rect 1873 2149 1881 2169
rect 1901 2167 1989 2169
rect 1901 2149 1930 2167
rect 1873 2148 1930 2149
rect 1959 2149 1989 2167
rect 2009 2149 2017 2169
rect 1959 2148 2017 2149
rect 1873 2141 2017 2148
rect 1873 2140 1909 2141
rect 1981 2140 2017 2141
rect 2083 2174 2120 2175
rect 2083 2173 2121 2174
rect 2083 2165 2147 2173
rect 2083 2145 2092 2165
rect 2112 2151 2147 2165
rect 2167 2151 2170 2171
rect 2112 2146 2170 2151
rect 2112 2145 2147 2146
rect 491 2118 556 2137
rect 455 2115 556 2118
rect 306 2113 556 2115
rect 74 2077 111 2078
rect 70 2074 111 2077
rect 70 2069 112 2074
rect 70 2051 83 2069
rect 101 2051 112 2069
rect 70 2037 112 2051
rect 150 2037 197 2041
rect 70 2031 197 2037
rect 70 2002 158 2031
rect 187 2002 197 2031
rect 306 2034 343 2113
rect 384 2100 494 2113
rect 458 2044 489 2045
rect 306 2014 315 2034
rect 335 2014 343 2034
rect 306 2004 343 2014
rect 402 2034 489 2044
rect 402 2014 411 2034
rect 431 2014 489 2034
rect 402 2005 489 2014
rect 402 2004 439 2005
rect 70 1998 197 2002
rect 70 1981 109 1998
rect 150 1997 197 1998
rect 70 1963 81 1981
rect 99 1963 109 1981
rect 70 1954 109 1963
rect 71 1953 108 1954
rect 458 1952 489 2005
rect 519 2034 556 2113
rect 727 2110 1120 2130
rect 1140 2110 1143 2130
rect 727 2105 1143 2110
rect 1349 2108 1386 2137
rect 1350 2106 1386 2108
rect 1562 2106 1599 2137
rect 727 2104 1068 2105
rect 671 2044 702 2045
rect 519 2014 528 2034
rect 548 2014 556 2034
rect 519 2004 556 2014
rect 615 2037 702 2044
rect 615 2034 676 2037
rect 615 2014 624 2034
rect 644 2017 676 2034
rect 697 2017 702 2037
rect 644 2014 702 2017
rect 615 2007 702 2014
rect 727 2034 764 2104
rect 1030 2103 1067 2104
rect 1350 2084 1599 2106
rect 1770 2105 1807 2137
rect 2083 2133 2147 2145
rect 2187 2109 2214 2285
rect 2095 2107 2214 2109
rect 2046 2105 2214 2107
rect 1431 2078 1542 2084
rect 1770 2079 2214 2105
rect 2046 2078 2214 2079
rect 1431 2070 1472 2078
rect 1431 2050 1439 2070
rect 1458 2050 1472 2070
rect 1431 2048 1472 2050
rect 1500 2070 1542 2078
rect 2095 2077 2203 2078
rect 1500 2050 1516 2070
rect 1535 2050 1542 2070
rect 1500 2048 1542 2050
rect 879 2044 915 2045
rect 727 2014 736 2034
rect 756 2014 764 2034
rect 615 2005 671 2007
rect 615 2004 652 2005
rect 727 2004 764 2014
rect 823 2034 971 2044
rect 1071 2041 1167 2043
rect 823 2014 832 2034
rect 852 2014 942 2034
rect 962 2014 971 2034
rect 823 2005 971 2014
rect 1029 2034 1167 2041
rect 1029 2014 1038 2034
rect 1058 2014 1167 2034
rect 1431 2033 1542 2048
rect 2133 2076 2203 2077
rect 1029 2005 1167 2014
rect 823 2004 860 2005
rect 879 1953 915 2005
rect 934 2004 971 2005
rect 1030 2004 1067 2005
rect 350 1951 391 1952
rect 242 1944 391 1951
rect 242 1924 360 1944
rect 380 1924 391 1944
rect 242 1916 391 1924
rect 458 1948 817 1952
rect 458 1943 780 1948
rect 458 1919 571 1943
rect 595 1924 780 1943
rect 804 1924 817 1948
rect 595 1919 817 1924
rect 458 1916 817 1919
rect 879 1916 914 1953
rect 982 1950 1082 1953
rect 982 1946 1049 1950
rect 982 1920 994 1946
rect 1020 1924 1049 1946
rect 1075 1924 1082 1950
rect 1020 1920 1082 1924
rect 982 1916 1082 1920
rect 458 1895 489 1916
rect 879 1895 915 1916
rect 301 1894 338 1895
rect 75 1891 109 1892
rect 74 1882 111 1891
rect 74 1864 83 1882
rect 101 1864 111 1882
rect 74 1854 111 1864
rect 300 1885 338 1894
rect 300 1865 309 1885
rect 329 1865 338 1885
rect 300 1857 338 1865
rect 404 1889 489 1895
rect 514 1894 551 1895
rect 404 1869 412 1889
rect 432 1869 489 1889
rect 404 1861 489 1869
rect 513 1885 551 1894
rect 513 1865 522 1885
rect 542 1865 551 1885
rect 404 1860 440 1861
rect 513 1857 551 1865
rect 617 1889 702 1895
rect 722 1894 759 1895
rect 617 1869 625 1889
rect 645 1888 702 1889
rect 645 1869 674 1888
rect 617 1868 674 1869
rect 695 1868 702 1888
rect 617 1861 702 1868
rect 721 1885 759 1894
rect 721 1865 730 1885
rect 750 1865 759 1885
rect 617 1860 653 1861
rect 721 1857 759 1865
rect 825 1889 969 1895
rect 825 1869 833 1889
rect 853 1888 941 1889
rect 853 1869 884 1888
rect 825 1868 884 1869
rect 909 1869 941 1888
rect 961 1869 969 1889
rect 909 1868 969 1869
rect 825 1861 969 1868
rect 825 1860 861 1861
rect 933 1860 969 1861
rect 1035 1894 1072 1895
rect 1035 1893 1073 1894
rect 1035 1885 1099 1893
rect 1035 1865 1044 1885
rect 1064 1871 1099 1885
rect 1119 1871 1122 1891
rect 1064 1866 1122 1871
rect 1064 1865 1099 1866
rect 75 1826 109 1854
rect 301 1828 338 1857
rect 302 1826 338 1828
rect 514 1826 551 1857
rect 75 1825 247 1826
rect 75 1793 261 1825
rect 302 1804 551 1826
rect 722 1825 759 1857
rect 1035 1853 1099 1865
rect 1139 1827 1166 2005
rect 2133 1969 2194 2076
rect 2133 1958 2203 1969
rect 2133 1949 2140 1958
rect 2135 1929 2140 1949
rect 2188 1929 2203 1958
rect 2135 1920 2203 1929
rect 1322 1901 1432 1915
rect 1322 1898 1365 1901
rect 1322 1893 1326 1898
rect 998 1825 1166 1827
rect 722 1819 1166 1825
rect 75 1761 109 1793
rect 71 1752 109 1761
rect 71 1734 81 1752
rect 99 1734 109 1752
rect 71 1728 109 1734
rect 227 1730 261 1793
rect 383 1798 494 1804
rect 383 1790 424 1798
rect 383 1770 391 1790
rect 410 1770 424 1790
rect 383 1768 424 1770
rect 452 1790 494 1798
rect 452 1770 468 1790
rect 487 1770 494 1790
rect 452 1768 494 1770
rect 383 1753 494 1768
rect 721 1799 1166 1819
rect 721 1730 759 1799
rect 998 1798 1166 1799
rect 1244 1871 1326 1893
rect 1355 1871 1365 1898
rect 1393 1874 1400 1901
rect 1429 1893 1432 1901
rect 1429 1874 1494 1893
rect 1393 1871 1494 1874
rect 1244 1869 1494 1871
rect 1244 1790 1281 1869
rect 1322 1856 1432 1869
rect 1396 1800 1427 1801
rect 1244 1770 1253 1790
rect 1273 1770 1281 1790
rect 1244 1760 1281 1770
rect 1340 1790 1427 1800
rect 1340 1770 1349 1790
rect 1369 1770 1427 1790
rect 1340 1761 1427 1770
rect 1340 1760 1377 1761
rect 71 1724 108 1728
rect 227 1719 759 1730
rect 226 1703 759 1719
rect 1396 1708 1427 1761
rect 1457 1790 1494 1869
rect 1665 1866 2058 1886
rect 2078 1866 2081 1886
rect 1665 1861 2081 1866
rect 1665 1860 2006 1861
rect 1609 1800 1640 1801
rect 1457 1770 1466 1790
rect 1486 1770 1494 1790
rect 1457 1760 1494 1770
rect 1553 1793 1640 1800
rect 1553 1790 1614 1793
rect 1553 1770 1562 1790
rect 1582 1773 1614 1790
rect 1635 1773 1640 1793
rect 1582 1770 1640 1773
rect 1553 1763 1640 1770
rect 1665 1790 1702 1860
rect 1968 1859 2005 1860
rect 1817 1800 1853 1801
rect 1665 1770 1674 1790
rect 1694 1770 1702 1790
rect 1553 1761 1609 1763
rect 1553 1760 1590 1761
rect 1665 1760 1702 1770
rect 1761 1790 1909 1800
rect 2009 1797 2105 1799
rect 1761 1770 1770 1790
rect 1790 1770 1880 1790
rect 1900 1770 1909 1790
rect 1761 1761 1909 1770
rect 1967 1790 2105 1797
rect 1967 1770 1976 1790
rect 1996 1770 2105 1790
rect 1967 1761 2105 1770
rect 1761 1760 1798 1761
rect 1817 1709 1853 1761
rect 1872 1760 1909 1761
rect 1968 1760 2005 1761
rect 1288 1707 1329 1708
rect 226 1702 740 1703
rect 1180 1700 1329 1707
rect 1180 1680 1298 1700
rect 1318 1680 1329 1700
rect 1180 1672 1329 1680
rect 1396 1704 1755 1708
rect 1396 1699 1718 1704
rect 1396 1675 1509 1699
rect 1533 1680 1718 1699
rect 1742 1680 1755 1704
rect 1533 1675 1755 1680
rect 1396 1672 1755 1675
rect 1817 1672 1852 1709
rect 1920 1706 2020 1709
rect 1920 1702 1987 1706
rect 1920 1676 1932 1702
rect 1958 1680 1987 1702
rect 2013 1680 2020 1706
rect 1958 1676 2020 1680
rect 1920 1672 2020 1676
rect 74 1661 111 1662
rect 72 1653 112 1661
rect 72 1635 83 1653
rect 101 1635 112 1653
rect 1396 1651 1427 1672
rect 1817 1651 1853 1672
rect 1239 1650 1276 1651
rect 72 1587 112 1635
rect 1238 1641 1276 1650
rect 1238 1621 1247 1641
rect 1267 1621 1276 1641
rect 1238 1613 1276 1621
rect 1342 1645 1427 1651
rect 1452 1650 1489 1651
rect 1342 1625 1350 1645
rect 1370 1625 1427 1645
rect 1342 1617 1427 1625
rect 1451 1641 1489 1650
rect 1451 1621 1460 1641
rect 1480 1621 1489 1641
rect 1342 1616 1378 1617
rect 1451 1613 1489 1621
rect 1555 1645 1640 1651
rect 1660 1650 1697 1651
rect 1555 1625 1563 1645
rect 1583 1644 1640 1645
rect 1583 1625 1612 1644
rect 1555 1624 1612 1625
rect 1633 1624 1640 1644
rect 1555 1617 1640 1624
rect 1659 1641 1697 1650
rect 1659 1621 1668 1641
rect 1688 1621 1697 1641
rect 1555 1616 1591 1617
rect 1659 1613 1697 1621
rect 1763 1645 1907 1651
rect 1763 1625 1771 1645
rect 1791 1628 1827 1645
rect 1847 1628 1879 1645
rect 1791 1625 1879 1628
rect 1899 1625 1907 1645
rect 1763 1617 1907 1625
rect 1763 1616 1799 1617
rect 1871 1616 1907 1617
rect 1973 1650 2010 1651
rect 1973 1649 2011 1650
rect 1973 1641 2037 1649
rect 1973 1621 1982 1641
rect 2002 1627 2037 1641
rect 2057 1627 2060 1647
rect 2002 1622 2060 1627
rect 2002 1621 2037 1622
rect 383 1591 493 1605
rect 383 1588 426 1591
rect 72 1580 197 1587
rect 383 1583 387 1588
rect 72 1561 164 1580
rect 189 1561 197 1580
rect 72 1551 197 1561
rect 305 1561 387 1583
rect 416 1561 426 1588
rect 454 1564 461 1591
rect 490 1583 493 1591
rect 1239 1584 1276 1613
rect 490 1564 555 1583
rect 1240 1582 1276 1584
rect 1452 1582 1489 1613
rect 1660 1586 1697 1613
rect 1973 1609 2037 1621
rect 454 1561 555 1564
rect 305 1559 555 1561
rect 72 1531 112 1551
rect 71 1522 112 1531
rect 71 1504 81 1522
rect 99 1504 112 1522
rect 71 1495 112 1504
rect 71 1494 108 1495
rect 305 1480 342 1559
rect 383 1546 493 1559
rect 457 1490 488 1491
rect 305 1460 314 1480
rect 334 1460 342 1480
rect 305 1450 342 1460
rect 401 1480 488 1490
rect 401 1460 410 1480
rect 430 1460 488 1480
rect 401 1451 488 1460
rect 401 1450 438 1451
rect 74 1428 111 1432
rect 71 1423 111 1428
rect 71 1405 83 1423
rect 101 1405 111 1423
rect 71 1225 111 1405
rect 457 1398 488 1451
rect 518 1480 555 1559
rect 726 1556 1119 1576
rect 1139 1556 1142 1576
rect 1240 1560 1489 1582
rect 1658 1581 1699 1586
rect 2077 1583 2104 1761
rect 1936 1581 2104 1583
rect 1658 1575 2104 1581
rect 726 1551 1142 1556
rect 1321 1554 1432 1560
rect 726 1550 1067 1551
rect 670 1490 701 1491
rect 518 1460 527 1480
rect 547 1460 555 1480
rect 518 1450 555 1460
rect 614 1483 701 1490
rect 614 1480 675 1483
rect 614 1460 623 1480
rect 643 1463 675 1480
rect 696 1463 701 1483
rect 643 1460 701 1463
rect 614 1453 701 1460
rect 726 1480 763 1550
rect 1029 1549 1066 1550
rect 1321 1546 1362 1554
rect 1321 1526 1329 1546
rect 1348 1526 1362 1546
rect 1321 1524 1362 1526
rect 1390 1546 1432 1554
rect 1390 1526 1406 1546
rect 1425 1526 1432 1546
rect 1658 1553 1664 1575
rect 1690 1555 2104 1575
rect 1690 1553 1699 1555
rect 1936 1554 2104 1555
rect 1658 1544 1699 1553
rect 1390 1524 1432 1526
rect 1321 1509 1432 1524
rect 878 1490 914 1491
rect 726 1460 735 1480
rect 755 1460 763 1480
rect 614 1451 670 1453
rect 614 1450 651 1451
rect 726 1450 763 1460
rect 822 1480 970 1490
rect 1070 1487 1166 1489
rect 822 1460 831 1480
rect 851 1460 941 1480
rect 961 1460 970 1480
rect 822 1451 970 1460
rect 1028 1480 1166 1487
rect 1028 1460 1037 1480
rect 1057 1460 1166 1480
rect 1028 1451 1166 1460
rect 822 1450 859 1451
rect 878 1399 914 1451
rect 933 1450 970 1451
rect 1029 1450 1066 1451
rect 349 1397 390 1398
rect 241 1390 390 1397
rect 241 1370 359 1390
rect 379 1370 390 1390
rect 241 1362 390 1370
rect 457 1394 816 1398
rect 457 1389 779 1394
rect 457 1365 570 1389
rect 594 1370 779 1389
rect 803 1370 816 1394
rect 594 1365 816 1370
rect 457 1362 816 1365
rect 878 1362 913 1399
rect 981 1396 1081 1399
rect 981 1392 1048 1396
rect 981 1366 993 1392
rect 1019 1370 1048 1392
rect 1074 1370 1081 1396
rect 1019 1366 1081 1370
rect 981 1362 1081 1366
rect 457 1341 488 1362
rect 878 1341 914 1362
rect 300 1340 337 1341
rect 299 1331 337 1340
rect 299 1311 308 1331
rect 328 1311 337 1331
rect 299 1303 337 1311
rect 403 1335 488 1341
rect 513 1340 550 1341
rect 403 1315 411 1335
rect 431 1315 488 1335
rect 403 1307 488 1315
rect 512 1331 550 1340
rect 512 1311 521 1331
rect 541 1311 550 1331
rect 403 1306 439 1307
rect 512 1303 550 1311
rect 616 1335 701 1341
rect 721 1340 758 1341
rect 616 1315 624 1335
rect 644 1334 701 1335
rect 644 1315 673 1334
rect 616 1314 673 1315
rect 694 1314 701 1334
rect 616 1307 701 1314
rect 720 1331 758 1340
rect 720 1311 729 1331
rect 749 1311 758 1331
rect 616 1306 652 1307
rect 720 1303 758 1311
rect 824 1335 968 1341
rect 824 1315 832 1335
rect 852 1332 940 1335
rect 852 1315 883 1332
rect 824 1312 883 1315
rect 906 1315 940 1332
rect 960 1315 968 1335
rect 906 1312 968 1315
rect 824 1307 968 1312
rect 824 1306 860 1307
rect 932 1306 968 1307
rect 1034 1340 1071 1341
rect 1034 1339 1072 1340
rect 1034 1331 1098 1339
rect 1034 1311 1043 1331
rect 1063 1317 1098 1331
rect 1118 1317 1121 1337
rect 1063 1312 1121 1317
rect 1063 1311 1098 1312
rect 300 1274 337 1303
rect 301 1272 337 1274
rect 513 1272 550 1303
rect 301 1250 550 1272
rect 721 1271 758 1303
rect 1034 1299 1098 1311
rect 1138 1273 1165 1451
rect 1463 1309 1573 1323
rect 1463 1306 1506 1309
rect 1463 1301 1467 1306
rect 997 1271 1165 1273
rect 721 1268 1165 1271
rect 382 1244 493 1250
rect 382 1236 423 1244
rect 71 1181 110 1225
rect 382 1216 390 1236
rect 409 1216 423 1236
rect 382 1214 423 1216
rect 451 1236 493 1244
rect 451 1216 467 1236
rect 486 1216 493 1236
rect 451 1214 493 1216
rect 382 1199 493 1214
rect 719 1245 1165 1268
rect 71 1157 111 1181
rect 411 1157 458 1159
rect 719 1157 757 1245
rect 997 1244 1165 1245
rect 1385 1279 1467 1301
rect 1496 1279 1506 1306
rect 1534 1282 1541 1309
rect 1570 1301 1573 1309
rect 1570 1282 1635 1301
rect 1534 1279 1635 1282
rect 1385 1277 1635 1279
rect 1385 1198 1422 1277
rect 1463 1264 1573 1277
rect 1537 1208 1568 1209
rect 1385 1178 1394 1198
rect 1414 1178 1422 1198
rect 1385 1168 1422 1178
rect 1481 1198 1568 1208
rect 1481 1178 1490 1198
rect 1510 1178 1568 1198
rect 1481 1169 1568 1178
rect 1481 1168 1518 1169
rect 71 1124 757 1157
rect 71 1067 110 1124
rect 719 1122 757 1124
rect 1537 1116 1568 1169
rect 1598 1198 1635 1277
rect 1806 1290 2199 1294
rect 1806 1273 1825 1290
rect 1845 1274 2199 1290
rect 2219 1274 2222 1294
rect 1845 1273 2222 1274
rect 1806 1269 2222 1273
rect 1806 1268 2147 1269
rect 1750 1208 1781 1209
rect 1598 1178 1607 1198
rect 1627 1178 1635 1198
rect 1598 1168 1635 1178
rect 1694 1201 1781 1208
rect 1694 1198 1755 1201
rect 1694 1178 1703 1198
rect 1723 1181 1755 1198
rect 1776 1181 1781 1201
rect 1723 1178 1781 1181
rect 1694 1171 1781 1178
rect 1806 1198 1843 1268
rect 2109 1267 2146 1268
rect 1958 1208 1994 1209
rect 1806 1178 1815 1198
rect 1835 1178 1843 1198
rect 1694 1169 1750 1171
rect 1694 1168 1731 1169
rect 1806 1168 1843 1178
rect 1902 1198 2050 1208
rect 2218 1207 2247 1208
rect 2150 1205 2247 1207
rect 1902 1178 1911 1198
rect 1931 1194 2021 1198
rect 1931 1178 1964 1194
rect 1902 1169 1964 1178
rect 1902 1168 1939 1169
rect 1958 1156 1964 1169
rect 1987 1178 2021 1194
rect 2041 1178 2050 1198
rect 1987 1169 2050 1178
rect 2108 1198 2247 1205
rect 2108 1178 2117 1198
rect 2137 1178 2247 1198
rect 2108 1169 2247 1178
rect 1987 1156 1994 1169
rect 2013 1168 2050 1169
rect 2109 1168 2146 1169
rect 1958 1117 1994 1156
rect 1429 1115 1470 1116
rect 1321 1108 1470 1115
rect 1321 1088 1439 1108
rect 1459 1088 1470 1108
rect 1321 1080 1470 1088
rect 1537 1112 1896 1116
rect 1537 1107 1859 1112
rect 1537 1083 1650 1107
rect 1674 1088 1859 1107
rect 1883 1088 1896 1112
rect 1674 1083 1896 1088
rect 1537 1080 1896 1083
rect 1958 1080 1993 1117
rect 2061 1114 2161 1117
rect 2061 1110 2128 1114
rect 2061 1084 2073 1110
rect 2099 1088 2128 1110
rect 2154 1088 2161 1114
rect 2099 1084 2161 1088
rect 2061 1080 2161 1084
rect 71 1065 119 1067
rect 71 1047 82 1065
rect 100 1047 119 1065
rect 1537 1059 1568 1080
rect 1958 1059 1994 1080
rect 1380 1058 1417 1059
rect 71 1038 119 1047
rect 72 1037 119 1038
rect 385 1042 495 1056
rect 385 1039 428 1042
rect 385 1034 389 1039
rect 307 1012 389 1034
rect 418 1012 428 1039
rect 456 1015 463 1042
rect 492 1034 495 1042
rect 1379 1049 1417 1058
rect 492 1015 557 1034
rect 1379 1029 1388 1049
rect 1408 1029 1417 1049
rect 456 1012 557 1015
rect 307 1010 557 1012
rect 75 974 112 975
rect 71 971 112 974
rect 71 966 113 971
rect 71 948 84 966
rect 102 948 113 966
rect 71 934 113 948
rect 151 934 198 938
rect 71 928 198 934
rect 71 899 159 928
rect 188 899 198 928
rect 307 931 344 1010
rect 385 997 495 1010
rect 459 941 490 942
rect 307 911 316 931
rect 336 911 344 931
rect 307 901 344 911
rect 403 931 490 941
rect 403 911 412 931
rect 432 911 490 931
rect 403 902 490 911
rect 403 901 440 902
rect 71 895 198 899
rect 71 878 110 895
rect 151 894 198 895
rect 71 860 82 878
rect 100 860 110 878
rect 71 851 110 860
rect 72 850 109 851
rect 459 849 490 902
rect 520 931 557 1010
rect 728 1007 1121 1027
rect 1141 1007 1144 1027
rect 1379 1021 1417 1029
rect 1483 1053 1568 1059
rect 1593 1058 1630 1059
rect 1483 1033 1491 1053
rect 1511 1033 1568 1053
rect 1483 1025 1568 1033
rect 1592 1049 1630 1058
rect 1592 1029 1601 1049
rect 1621 1029 1630 1049
rect 1483 1024 1519 1025
rect 1592 1021 1630 1029
rect 1696 1053 1781 1059
rect 1801 1058 1838 1059
rect 1696 1033 1704 1053
rect 1724 1052 1781 1053
rect 1724 1033 1753 1052
rect 1696 1032 1753 1033
rect 1774 1032 1781 1052
rect 1696 1025 1781 1032
rect 1800 1049 1838 1058
rect 1800 1029 1809 1049
rect 1829 1029 1838 1049
rect 1696 1024 1732 1025
rect 1800 1021 1838 1029
rect 1904 1053 2048 1059
rect 1904 1033 1912 1053
rect 1932 1033 2020 1053
rect 2040 1033 2048 1053
rect 1904 1025 2048 1033
rect 1904 1024 1940 1025
rect 2012 1024 2048 1025
rect 2114 1058 2151 1059
rect 2114 1057 2152 1058
rect 2114 1049 2178 1057
rect 2114 1029 2123 1049
rect 2143 1035 2178 1049
rect 2198 1035 2201 1055
rect 2143 1030 2201 1035
rect 2143 1029 2178 1030
rect 728 1002 1144 1007
rect 728 1001 1069 1002
rect 672 941 703 942
rect 520 911 529 931
rect 549 911 557 931
rect 520 901 557 911
rect 616 934 703 941
rect 616 931 677 934
rect 616 911 625 931
rect 645 914 677 931
rect 698 914 703 934
rect 645 911 703 914
rect 616 904 703 911
rect 728 931 765 1001
rect 1031 1000 1068 1001
rect 1380 992 1417 1021
rect 1381 990 1417 992
rect 1593 990 1630 1021
rect 1381 968 1630 990
rect 1801 989 1838 1021
rect 2114 1017 2178 1029
rect 2218 991 2247 1169
rect 2077 989 2247 991
rect 1798 982 2247 989
rect 1462 962 1573 968
rect 1462 954 1503 962
rect 880 941 916 942
rect 728 911 737 931
rect 757 911 765 931
rect 616 902 672 904
rect 616 901 653 902
rect 728 901 765 911
rect 824 931 972 941
rect 1072 938 1168 940
rect 824 911 833 931
rect 853 911 943 931
rect 963 911 972 931
rect 824 902 972 911
rect 1030 931 1168 938
rect 1030 911 1039 931
rect 1059 911 1168 931
rect 1462 934 1470 954
rect 1489 934 1503 954
rect 1462 932 1503 934
rect 1531 954 1573 962
rect 1531 934 1547 954
rect 1566 934 1573 954
rect 1798 955 1823 982
rect 1854 963 2247 982
rect 1854 955 1903 963
rect 2077 962 2247 963
rect 1798 953 1903 955
rect 1531 932 1573 934
rect 1462 917 1573 932
rect 1030 902 1168 911
rect 824 901 861 902
rect 880 850 916 902
rect 935 901 972 902
rect 1031 901 1068 902
rect 351 848 392 849
rect 243 841 392 848
rect 243 821 361 841
rect 381 821 392 841
rect 243 813 392 821
rect 459 845 818 849
rect 459 840 781 845
rect 459 816 572 840
rect 596 821 781 840
rect 805 821 818 845
rect 596 816 818 821
rect 459 813 818 816
rect 880 813 915 850
rect 983 847 1083 850
rect 983 843 1050 847
rect 983 817 995 843
rect 1021 821 1050 843
rect 1076 821 1083 847
rect 1021 817 1083 821
rect 983 813 1083 817
rect 459 792 490 813
rect 880 792 916 813
rect 302 791 339 792
rect 76 788 110 789
rect 75 779 112 788
rect 75 761 84 779
rect 102 761 112 779
rect 75 751 112 761
rect 301 782 339 791
rect 301 762 310 782
rect 330 762 339 782
rect 301 754 339 762
rect 405 786 490 792
rect 515 791 552 792
rect 405 766 413 786
rect 433 766 490 786
rect 405 758 490 766
rect 514 782 552 791
rect 514 762 523 782
rect 543 762 552 782
rect 405 757 441 758
rect 514 754 552 762
rect 618 786 703 792
rect 723 791 760 792
rect 618 766 626 786
rect 646 785 703 786
rect 646 766 675 785
rect 618 765 675 766
rect 696 765 703 785
rect 618 758 703 765
rect 722 782 760 791
rect 722 762 731 782
rect 751 762 760 782
rect 618 757 654 758
rect 722 754 760 762
rect 826 786 970 792
rect 826 766 834 786
rect 854 785 942 786
rect 854 766 885 785
rect 826 765 885 766
rect 910 766 942 785
rect 962 766 970 786
rect 910 765 970 766
rect 826 758 970 765
rect 826 757 862 758
rect 934 757 970 758
rect 1036 791 1073 792
rect 1036 790 1074 791
rect 1036 782 1100 790
rect 1036 762 1045 782
rect 1065 768 1100 782
rect 1120 768 1123 788
rect 1065 763 1123 768
rect 1065 762 1100 763
rect 76 723 110 751
rect 302 725 339 754
rect 303 723 339 725
rect 515 723 552 754
rect 76 722 248 723
rect 76 690 262 722
rect 303 701 552 723
rect 723 722 760 754
rect 1036 750 1100 762
rect 1140 724 1167 902
rect 1323 798 1433 812
rect 1323 795 1366 798
rect 1323 790 1327 795
rect 999 722 1167 724
rect 723 716 1167 722
rect 76 658 110 690
rect 72 649 110 658
rect 72 631 82 649
rect 100 631 110 649
rect 72 625 110 631
rect 228 627 262 690
rect 384 695 495 701
rect 384 687 425 695
rect 384 667 392 687
rect 411 667 425 687
rect 384 665 425 667
rect 453 687 495 695
rect 453 667 469 687
rect 488 667 495 687
rect 453 665 495 667
rect 384 650 495 665
rect 722 696 1167 716
rect 722 627 760 696
rect 999 695 1167 696
rect 1245 768 1327 790
rect 1356 768 1366 795
rect 1394 771 1401 798
rect 1430 790 1433 798
rect 1430 771 1495 790
rect 1394 768 1495 771
rect 1245 766 1495 768
rect 1245 687 1282 766
rect 1323 753 1433 766
rect 1397 697 1428 698
rect 1245 667 1254 687
rect 1274 667 1282 687
rect 1245 657 1282 667
rect 1341 687 1428 697
rect 1341 667 1350 687
rect 1370 667 1428 687
rect 1341 658 1428 667
rect 1341 657 1378 658
rect 72 621 109 625
rect 228 616 760 627
rect 227 600 760 616
rect 1397 605 1428 658
rect 1458 687 1495 766
rect 1666 776 2059 783
rect 1666 759 1674 776
rect 1706 763 2059 776
rect 2079 763 2082 783
rect 1706 759 2082 763
rect 1666 758 2082 759
rect 1666 757 2007 758
rect 1610 697 1641 698
rect 1458 667 1467 687
rect 1487 667 1495 687
rect 1458 657 1495 667
rect 1554 690 1641 697
rect 1554 687 1615 690
rect 1554 667 1563 687
rect 1583 670 1615 687
rect 1636 670 1641 690
rect 1583 667 1641 670
rect 1554 660 1641 667
rect 1666 687 1703 757
rect 1969 756 2006 757
rect 1818 697 1854 698
rect 1666 667 1675 687
rect 1695 667 1703 687
rect 1554 658 1610 660
rect 1554 657 1591 658
rect 1666 657 1703 667
rect 1762 687 1910 697
rect 2010 694 2106 696
rect 1762 667 1771 687
rect 1791 682 1881 687
rect 1791 667 1826 682
rect 1762 658 1826 667
rect 1762 657 1799 658
rect 1818 641 1826 658
rect 1847 667 1881 682
rect 1901 667 1910 687
rect 1847 658 1910 667
rect 1968 687 2106 694
rect 1968 667 1977 687
rect 1997 667 2106 687
rect 1968 658 2106 667
rect 1847 641 1854 658
rect 1873 657 1910 658
rect 1969 657 2006 658
rect 1818 606 1854 641
rect 1289 604 1330 605
rect 227 599 741 600
rect 1181 597 1330 604
rect 1181 577 1299 597
rect 1319 577 1330 597
rect 1181 569 1330 577
rect 1397 601 1756 605
rect 1397 596 1719 601
rect 1397 572 1510 596
rect 1534 577 1719 596
rect 1743 577 1756 601
rect 1534 572 1756 577
rect 1397 569 1756 572
rect 1818 569 1853 606
rect 1921 603 2021 606
rect 1921 599 1988 603
rect 1921 573 1933 599
rect 1959 577 1988 599
rect 2014 577 2021 603
rect 1959 573 2021 577
rect 1921 569 2021 573
rect 75 558 112 559
rect 73 550 113 558
rect 73 532 84 550
rect 102 532 113 550
rect 1397 548 1428 569
rect 1818 548 1854 569
rect 1240 547 1277 548
rect 73 484 113 532
rect 1239 538 1277 547
rect 1239 518 1248 538
rect 1268 518 1277 538
rect 1239 510 1277 518
rect 1343 542 1428 548
rect 1453 547 1490 548
rect 1343 522 1351 542
rect 1371 522 1428 542
rect 1343 514 1428 522
rect 1452 538 1490 547
rect 1452 518 1461 538
rect 1481 518 1490 538
rect 1343 513 1379 514
rect 1452 510 1490 518
rect 1556 542 1641 548
rect 1661 547 1698 548
rect 1556 522 1564 542
rect 1584 541 1641 542
rect 1584 522 1613 541
rect 1556 521 1613 522
rect 1634 521 1641 541
rect 1556 514 1641 521
rect 1660 538 1698 547
rect 1660 518 1669 538
rect 1689 518 1698 538
rect 1556 513 1592 514
rect 1660 510 1698 518
rect 1764 542 1908 548
rect 1764 522 1772 542
rect 1792 522 1880 542
rect 1900 522 1908 542
rect 1764 514 1908 522
rect 1764 513 1800 514
rect 1872 513 1908 514
rect 1974 547 2011 548
rect 1974 546 2012 547
rect 1974 538 2038 546
rect 1974 518 1983 538
rect 2003 524 2038 538
rect 2058 524 2061 544
rect 2003 519 2061 524
rect 2003 518 2038 519
rect 384 488 494 502
rect 384 485 427 488
rect 73 477 198 484
rect 384 480 388 485
rect 73 458 165 477
rect 190 458 198 477
rect 73 448 198 458
rect 306 458 388 480
rect 417 458 427 485
rect 455 461 462 488
rect 491 480 494 488
rect 1240 481 1277 510
rect 491 461 556 480
rect 1241 479 1277 481
rect 1453 479 1490 510
rect 1661 483 1698 510
rect 1974 506 2038 518
rect 455 458 556 461
rect 306 456 556 458
rect 73 428 113 448
rect 72 419 113 428
rect 72 401 82 419
rect 100 401 113 419
rect 72 392 113 401
rect 72 391 109 392
rect 306 377 343 456
rect 384 443 494 456
rect 458 387 489 388
rect 306 357 315 377
rect 335 357 343 377
rect 306 347 343 357
rect 402 377 489 387
rect 402 357 411 377
rect 431 357 489 377
rect 402 348 489 357
rect 402 347 439 348
rect 75 325 112 329
rect 72 320 112 325
rect 72 302 84 320
rect 102 302 112 320
rect 72 122 112 302
rect 458 295 489 348
rect 519 377 556 456
rect 727 453 1120 473
rect 1140 453 1143 473
rect 1241 457 1490 479
rect 1659 478 1700 483
rect 2078 480 2105 658
rect 1937 478 2105 480
rect 1659 472 2105 478
rect 727 448 1143 453
rect 1322 451 1433 457
rect 727 447 1068 448
rect 671 387 702 388
rect 519 357 528 377
rect 548 357 556 377
rect 519 347 556 357
rect 615 380 702 387
rect 615 377 676 380
rect 615 357 624 377
rect 644 360 676 377
rect 697 360 702 380
rect 644 357 702 360
rect 615 350 702 357
rect 727 377 764 447
rect 1030 446 1067 447
rect 1322 443 1363 451
rect 1322 423 1330 443
rect 1349 423 1363 443
rect 1322 421 1363 423
rect 1391 443 1433 451
rect 1391 423 1407 443
rect 1426 423 1433 443
rect 1659 450 1665 472
rect 1691 452 2105 472
rect 1691 450 1700 452
rect 1937 451 2105 452
rect 1659 441 1700 450
rect 1391 421 1433 423
rect 1322 406 1433 421
rect 879 387 915 388
rect 727 357 736 377
rect 756 357 764 377
rect 615 348 671 350
rect 615 347 652 348
rect 727 347 764 357
rect 823 377 971 387
rect 1071 384 1167 386
rect 823 357 832 377
rect 852 357 942 377
rect 962 357 971 377
rect 823 348 971 357
rect 1029 377 1167 384
rect 1029 357 1038 377
rect 1058 357 1167 377
rect 1029 348 1167 357
rect 823 347 860 348
rect 879 296 915 348
rect 934 347 971 348
rect 1030 347 1067 348
rect 350 294 391 295
rect 242 287 391 294
rect 242 267 360 287
rect 380 267 391 287
rect 242 259 391 267
rect 458 291 817 295
rect 458 286 780 291
rect 458 262 571 286
rect 595 267 780 286
rect 804 267 817 291
rect 595 262 817 267
rect 458 259 817 262
rect 879 259 914 296
rect 982 293 1082 296
rect 982 289 1049 293
rect 982 263 994 289
rect 1020 267 1049 289
rect 1075 267 1082 293
rect 1020 263 1082 267
rect 982 259 1082 263
rect 458 238 489 259
rect 879 238 915 259
rect 301 237 338 238
rect 300 228 338 237
rect 300 208 309 228
rect 329 208 338 228
rect 300 200 338 208
rect 404 232 489 238
rect 514 237 551 238
rect 404 212 412 232
rect 432 212 489 232
rect 404 204 489 212
rect 513 228 551 237
rect 513 208 522 228
rect 542 208 551 228
rect 404 203 440 204
rect 513 200 551 208
rect 617 232 702 238
rect 722 237 759 238
rect 617 212 625 232
rect 645 231 702 232
rect 645 212 674 231
rect 617 211 674 212
rect 695 211 702 231
rect 617 204 702 211
rect 721 228 759 237
rect 721 208 730 228
rect 750 208 759 228
rect 617 203 653 204
rect 721 200 759 208
rect 825 232 969 238
rect 825 212 833 232
rect 853 229 941 232
rect 853 212 884 229
rect 825 209 884 212
rect 907 212 941 229
rect 961 212 969 232
rect 907 209 969 212
rect 825 204 969 209
rect 825 203 861 204
rect 933 203 969 204
rect 1035 237 1072 238
rect 1035 236 1073 237
rect 1035 228 1099 236
rect 1035 208 1044 228
rect 1064 214 1099 228
rect 1119 214 1122 234
rect 1064 209 1122 214
rect 1064 208 1099 209
rect 301 171 338 200
rect 302 169 338 171
rect 514 169 551 200
rect 302 147 551 169
rect 722 168 759 200
rect 1035 196 1099 208
rect 1139 170 1166 348
rect 1432 225 1542 239
rect 1432 222 1475 225
rect 1432 217 1436 222
rect 998 168 1166 170
rect 722 165 1166 168
rect 383 141 494 147
rect 383 133 424 141
rect 72 78 111 122
rect 383 113 391 133
rect 410 113 424 133
rect 383 111 424 113
rect 452 133 494 141
rect 452 113 468 133
rect 487 113 494 133
rect 452 112 494 113
rect 720 142 1166 165
rect 452 111 495 112
rect 383 92 495 111
rect 72 54 112 78
rect 412 54 459 55
rect 720 54 758 142
rect 998 141 1166 142
rect 1354 195 1436 217
rect 1465 195 1475 222
rect 1503 198 1510 225
rect 1539 217 1542 225
rect 1539 198 1604 217
rect 1503 195 1604 198
rect 1354 193 1604 195
rect 1354 114 1391 193
rect 1432 180 1542 193
rect 1506 124 1537 125
rect 1354 94 1363 114
rect 1383 94 1391 114
rect 1354 84 1391 94
rect 1450 114 1537 124
rect 1450 94 1459 114
rect 1479 94 1537 114
rect 1450 85 1537 94
rect 1450 84 1487 85
rect 72 44 758 54
rect 68 21 758 44
rect 1506 32 1537 85
rect 1567 114 1604 193
rect 1775 190 2168 210
rect 2188 190 2191 210
rect 1775 185 2191 190
rect 1775 184 2116 185
rect 1719 124 1750 125
rect 1567 94 1576 114
rect 1596 94 1604 114
rect 1567 84 1604 94
rect 1663 117 1750 124
rect 1663 114 1724 117
rect 1663 94 1672 114
rect 1692 97 1724 114
rect 1745 97 1750 117
rect 1692 94 1750 97
rect 1663 87 1750 94
rect 1775 114 1812 184
rect 2078 183 2115 184
rect 1927 124 1963 125
rect 1775 94 1784 114
rect 1804 94 1812 114
rect 1663 85 1719 87
rect 1663 84 1700 85
rect 1775 84 1812 94
rect 1871 114 2019 124
rect 2119 121 2215 123
rect 1871 94 1880 114
rect 1900 94 1990 114
rect 2010 94 2019 114
rect 1871 85 2019 94
rect 2077 114 2215 121
rect 2077 94 2086 114
rect 2106 94 2215 114
rect 2077 85 2215 94
rect 1871 84 1908 85
rect 1927 33 1963 85
rect 1982 84 2019 85
rect 2078 84 2115 85
rect 1398 31 1439 32
rect 68 2 110 21
rect 720 19 758 21
rect 1290 24 1439 31
rect 71 -36 110 2
rect 1290 4 1408 24
rect 1428 4 1439 24
rect 1290 -4 1439 4
rect 1506 28 1865 32
rect 1506 23 1828 28
rect 1506 -1 1619 23
rect 1643 4 1828 23
rect 1852 4 1865 28
rect 1643 -1 1865 4
rect 1506 -4 1865 -1
rect 1927 -4 1962 33
rect 2030 30 2130 33
rect 2030 26 2097 30
rect 2030 0 2042 26
rect 2068 4 2097 26
rect 2123 4 2130 30
rect 2068 0 2130 4
rect 2030 -4 2130 0
rect 1506 -25 1537 -4
rect 1927 -25 1963 -4
rect 1349 -26 1386 -25
rect 1348 -35 1386 -26
rect 71 -38 119 -36
rect 71 -56 82 -38
rect 100 -56 119 -38
rect 71 -65 119 -56
rect 72 -66 119 -65
rect 385 -61 495 -47
rect 385 -64 428 -61
rect 385 -69 389 -64
rect 307 -91 389 -69
rect 418 -91 428 -64
rect 456 -88 463 -61
rect 492 -69 495 -61
rect 1348 -55 1357 -35
rect 1377 -55 1386 -35
rect 1348 -63 1386 -55
rect 1452 -31 1537 -25
rect 1562 -26 1599 -25
rect 1452 -51 1460 -31
rect 1480 -51 1537 -31
rect 1452 -59 1537 -51
rect 1561 -35 1599 -26
rect 1561 -55 1570 -35
rect 1590 -55 1599 -35
rect 1452 -60 1488 -59
rect 1561 -63 1599 -55
rect 1665 -31 1750 -25
rect 1770 -26 1807 -25
rect 1665 -51 1673 -31
rect 1693 -32 1750 -31
rect 1693 -51 1722 -32
rect 1665 -52 1722 -51
rect 1743 -52 1750 -32
rect 1665 -59 1750 -52
rect 1769 -35 1807 -26
rect 1769 -55 1778 -35
rect 1798 -55 1807 -35
rect 1665 -60 1701 -59
rect 1769 -63 1807 -55
rect 1873 -31 2017 -25
rect 1873 -51 1881 -31
rect 1901 -51 1989 -31
rect 2009 -51 2017 -31
rect 1873 -59 2017 -51
rect 1873 -60 1909 -59
rect 1981 -60 2017 -59
rect 2083 -26 2120 -25
rect 2083 -27 2121 -26
rect 2083 -35 2147 -27
rect 2083 -55 2092 -35
rect 2112 -49 2147 -35
rect 2167 -49 2170 -29
rect 2112 -54 2170 -49
rect 2112 -55 2147 -54
rect 492 -88 557 -69
rect 456 -91 557 -88
rect 307 -93 557 -91
rect 75 -129 112 -128
rect 71 -132 112 -129
rect 71 -137 113 -132
rect 71 -155 84 -137
rect 102 -155 113 -137
rect 71 -169 113 -155
rect 151 -169 198 -165
rect 71 -175 198 -169
rect 71 -204 159 -175
rect 188 -204 198 -175
rect 307 -172 344 -93
rect 385 -106 495 -93
rect 459 -162 490 -161
rect 307 -192 316 -172
rect 336 -192 344 -172
rect 307 -202 344 -192
rect 403 -172 490 -162
rect 403 -192 412 -172
rect 432 -192 490 -172
rect 403 -201 490 -192
rect 403 -202 440 -201
rect 71 -208 198 -204
rect 71 -225 110 -208
rect 151 -209 198 -208
rect 71 -243 82 -225
rect 100 -243 110 -225
rect 71 -252 110 -243
rect 72 -253 109 -252
rect 459 -254 490 -201
rect 520 -172 557 -93
rect 728 -96 1121 -76
rect 1141 -96 1144 -76
rect 1349 -92 1386 -63
rect 728 -101 1144 -96
rect 1350 -94 1386 -92
rect 1562 -94 1599 -63
rect 728 -102 1069 -101
rect 672 -162 703 -161
rect 520 -192 529 -172
rect 549 -192 557 -172
rect 520 -202 557 -192
rect 616 -169 703 -162
rect 616 -172 677 -169
rect 616 -192 625 -172
rect 645 -189 677 -172
rect 698 -189 703 -169
rect 645 -192 703 -189
rect 616 -199 703 -192
rect 728 -172 765 -102
rect 1031 -103 1068 -102
rect 1350 -116 1599 -94
rect 1770 -95 1807 -63
rect 2083 -67 2147 -55
rect 2187 -92 2214 85
rect 2295 -92 2348 -84
rect 2162 -93 2348 -92
rect 2046 -95 2348 -93
rect 1431 -122 1542 -116
rect 1770 -121 2348 -95
rect 2046 -122 2348 -121
rect 1431 -130 1472 -122
rect 1431 -150 1439 -130
rect 1458 -150 1472 -130
rect 1431 -152 1472 -150
rect 1500 -130 1542 -122
rect 1500 -150 1516 -130
rect 1535 -150 1542 -130
rect 1500 -152 1542 -150
rect 880 -162 916 -161
rect 728 -192 737 -172
rect 757 -192 765 -172
rect 616 -201 672 -199
rect 616 -202 653 -201
rect 728 -202 765 -192
rect 824 -172 972 -162
rect 1072 -165 1168 -163
rect 824 -192 833 -172
rect 853 -192 943 -172
rect 963 -192 972 -172
rect 824 -201 972 -192
rect 1030 -172 1168 -165
rect 1431 -167 1542 -152
rect 1030 -192 1039 -172
rect 1059 -192 1168 -172
rect 1030 -201 1168 -192
rect 824 -202 861 -201
rect 880 -253 916 -201
rect 935 -202 972 -201
rect 1031 -202 1068 -201
rect 351 -255 392 -254
rect 243 -262 392 -255
rect 243 -282 361 -262
rect 381 -282 392 -262
rect 243 -290 392 -282
rect 459 -258 818 -254
rect 459 -263 781 -258
rect 459 -287 572 -263
rect 596 -282 781 -263
rect 805 -282 818 -258
rect 596 -287 818 -282
rect 459 -290 818 -287
rect 880 -290 915 -253
rect 983 -256 1083 -253
rect 983 -260 1050 -256
rect 983 -286 995 -260
rect 1021 -282 1050 -260
rect 1076 -282 1083 -256
rect 1021 -286 1083 -282
rect 983 -290 1083 -286
rect 459 -311 490 -290
rect 880 -311 916 -290
rect 302 -312 339 -311
rect 76 -315 110 -314
rect 75 -324 112 -315
rect 75 -342 84 -324
rect 102 -342 112 -324
rect 75 -352 112 -342
rect 301 -321 339 -312
rect 301 -341 310 -321
rect 330 -341 339 -321
rect 301 -349 339 -341
rect 405 -317 490 -311
rect 515 -312 552 -311
rect 405 -337 413 -317
rect 433 -337 490 -317
rect 405 -345 490 -337
rect 514 -321 552 -312
rect 514 -341 523 -321
rect 543 -341 552 -321
rect 405 -346 441 -345
rect 514 -349 552 -341
rect 618 -317 703 -311
rect 723 -312 760 -311
rect 618 -337 626 -317
rect 646 -318 703 -317
rect 646 -337 675 -318
rect 618 -338 675 -337
rect 696 -338 703 -318
rect 618 -345 703 -338
rect 722 -321 760 -312
rect 722 -341 731 -321
rect 751 -341 760 -321
rect 618 -346 654 -345
rect 722 -349 760 -341
rect 826 -317 970 -311
rect 826 -337 834 -317
rect 854 -318 942 -317
rect 854 -337 885 -318
rect 826 -338 885 -337
rect 910 -337 942 -318
rect 962 -337 970 -317
rect 910 -338 970 -337
rect 826 -345 970 -338
rect 826 -346 862 -345
rect 934 -346 970 -345
rect 1036 -312 1073 -311
rect 1036 -313 1074 -312
rect 1036 -321 1100 -313
rect 1036 -341 1045 -321
rect 1065 -335 1100 -321
rect 1120 -335 1123 -315
rect 1065 -340 1123 -335
rect 1065 -341 1100 -340
rect 76 -380 110 -352
rect 302 -378 339 -349
rect 303 -380 339 -378
rect 515 -380 552 -349
rect 76 -381 248 -380
rect 76 -413 262 -381
rect 303 -402 552 -380
rect 723 -381 760 -349
rect 1036 -353 1100 -341
rect 1140 -379 1167 -201
rect 2295 -229 2348 -122
rect 2295 -247 2343 -229
rect 2295 -287 2303 -247
rect 2330 -287 2343 -247
rect 1323 -305 1433 -291
rect 2295 -301 2343 -287
rect 1323 -308 1366 -305
rect 1323 -313 1327 -308
rect 999 -381 1167 -379
rect 723 -387 1167 -381
rect 76 -445 110 -413
rect 72 -454 110 -445
rect 72 -472 82 -454
rect 100 -472 110 -454
rect 72 -478 110 -472
rect 228 -476 262 -413
rect 384 -408 495 -402
rect 384 -416 425 -408
rect 384 -436 392 -416
rect 411 -436 425 -416
rect 384 -438 425 -436
rect 453 -416 495 -408
rect 453 -436 469 -416
rect 488 -436 495 -416
rect 453 -438 495 -436
rect 384 -453 495 -438
rect 722 -407 1167 -387
rect 722 -476 760 -407
rect 999 -408 1167 -407
rect 1245 -335 1327 -313
rect 1356 -335 1366 -308
rect 1394 -332 1401 -305
rect 1430 -313 1433 -305
rect 1430 -332 1495 -313
rect 1394 -335 1495 -332
rect 1245 -337 1495 -335
rect 1245 -416 1282 -337
rect 1323 -350 1433 -337
rect 1397 -406 1428 -405
rect 1245 -436 1254 -416
rect 1274 -436 1282 -416
rect 1245 -446 1282 -436
rect 1341 -416 1428 -406
rect 1341 -436 1350 -416
rect 1370 -436 1428 -416
rect 1341 -445 1428 -436
rect 1341 -446 1378 -445
rect 72 -482 109 -478
rect 228 -487 760 -476
rect 227 -503 760 -487
rect 1397 -498 1428 -445
rect 1458 -416 1495 -337
rect 1666 -340 2059 -320
rect 2079 -340 2082 -320
rect 1666 -345 2082 -340
rect 1666 -346 2007 -345
rect 1610 -406 1641 -405
rect 1458 -436 1467 -416
rect 1487 -436 1495 -416
rect 1458 -446 1495 -436
rect 1554 -413 1641 -406
rect 1554 -416 1615 -413
rect 1554 -436 1563 -416
rect 1583 -433 1615 -416
rect 1636 -433 1641 -413
rect 1583 -436 1641 -433
rect 1554 -443 1641 -436
rect 1666 -416 1703 -346
rect 1969 -347 2006 -346
rect 1818 -406 1854 -405
rect 1666 -436 1675 -416
rect 1695 -436 1703 -416
rect 1554 -445 1610 -443
rect 1554 -446 1591 -445
rect 1666 -446 1703 -436
rect 1762 -416 1910 -406
rect 2010 -409 2106 -407
rect 1762 -436 1771 -416
rect 1791 -436 1881 -416
rect 1901 -436 1910 -416
rect 1762 -445 1910 -436
rect 1968 -416 2106 -409
rect 1968 -436 1977 -416
rect 1997 -436 2106 -416
rect 1968 -445 2106 -436
rect 1762 -446 1799 -445
rect 1818 -497 1854 -445
rect 1873 -446 1910 -445
rect 1969 -446 2006 -445
rect 1289 -499 1330 -498
rect 227 -504 741 -503
rect 1181 -506 1330 -499
rect 1181 -526 1299 -506
rect 1319 -526 1330 -506
rect 1181 -534 1330 -526
rect 1397 -502 1756 -498
rect 1397 -507 1719 -502
rect 1397 -531 1510 -507
rect 1534 -526 1719 -507
rect 1743 -526 1756 -502
rect 1534 -531 1756 -526
rect 1397 -534 1756 -531
rect 1818 -534 1853 -497
rect 1921 -500 2021 -497
rect 1921 -504 1988 -500
rect 1921 -530 1933 -504
rect 1959 -526 1988 -504
rect 2014 -526 2021 -500
rect 1959 -530 2021 -526
rect 1921 -534 2021 -530
rect 75 -545 112 -544
rect 73 -553 113 -545
rect 73 -571 84 -553
rect 102 -571 113 -553
rect 1397 -555 1428 -534
rect 1818 -555 1854 -534
rect 1240 -556 1277 -555
rect 73 -619 113 -571
rect 1239 -565 1277 -556
rect 1239 -585 1248 -565
rect 1268 -585 1277 -565
rect 1239 -593 1277 -585
rect 1343 -561 1428 -555
rect 1453 -556 1490 -555
rect 1343 -581 1351 -561
rect 1371 -581 1428 -561
rect 1343 -589 1428 -581
rect 1452 -565 1490 -556
rect 1452 -585 1461 -565
rect 1481 -585 1490 -565
rect 1343 -590 1379 -589
rect 1452 -593 1490 -585
rect 1556 -561 1641 -555
rect 1661 -556 1698 -555
rect 1556 -581 1564 -561
rect 1584 -562 1641 -561
rect 1584 -581 1613 -562
rect 1556 -582 1613 -581
rect 1634 -582 1641 -562
rect 1556 -589 1641 -582
rect 1660 -565 1698 -556
rect 1660 -585 1669 -565
rect 1689 -585 1698 -565
rect 1556 -590 1592 -589
rect 1660 -593 1698 -585
rect 1764 -561 1908 -555
rect 1764 -581 1772 -561
rect 1792 -578 1828 -561
rect 1848 -578 1880 -561
rect 1792 -581 1880 -578
rect 1900 -581 1908 -561
rect 1764 -589 1908 -581
rect 1764 -590 1800 -589
rect 1872 -590 1908 -589
rect 1974 -556 2011 -555
rect 1974 -557 2012 -556
rect 1974 -565 2038 -557
rect 1974 -585 1983 -565
rect 2003 -579 2038 -565
rect 2058 -579 2061 -559
rect 2003 -584 2061 -579
rect 2003 -585 2038 -584
rect 384 -615 494 -601
rect 384 -618 427 -615
rect 73 -626 198 -619
rect 384 -623 388 -618
rect 73 -645 165 -626
rect 190 -645 198 -626
rect 73 -655 198 -645
rect 306 -645 388 -623
rect 417 -645 427 -618
rect 455 -642 462 -615
rect 491 -623 494 -615
rect 1240 -622 1277 -593
rect 491 -642 556 -623
rect 1241 -624 1277 -622
rect 1453 -624 1490 -593
rect 1661 -620 1698 -593
rect 1974 -597 2038 -585
rect 455 -645 556 -642
rect 306 -647 556 -645
rect 73 -675 113 -655
rect 72 -684 113 -675
rect 72 -702 82 -684
rect 100 -702 113 -684
rect 72 -711 113 -702
rect 72 -712 109 -711
rect 306 -726 343 -647
rect 384 -660 494 -647
rect 458 -716 489 -715
rect 306 -746 315 -726
rect 335 -746 343 -726
rect 306 -756 343 -746
rect 402 -726 489 -716
rect 402 -746 411 -726
rect 431 -746 489 -726
rect 402 -755 489 -746
rect 402 -756 439 -755
rect 75 -778 112 -774
rect 72 -783 112 -778
rect 72 -801 84 -783
rect 102 -801 112 -783
rect 72 -981 112 -801
rect 458 -808 489 -755
rect 519 -726 556 -647
rect 727 -650 1120 -630
rect 1140 -650 1143 -630
rect 1241 -646 1490 -624
rect 1659 -625 1700 -620
rect 2078 -623 2105 -445
rect 1937 -625 2105 -623
rect 1659 -631 2105 -625
rect 727 -655 1143 -650
rect 1322 -652 1433 -646
rect 727 -656 1068 -655
rect 671 -716 702 -715
rect 519 -746 528 -726
rect 548 -746 556 -726
rect 519 -756 556 -746
rect 615 -723 702 -716
rect 615 -726 676 -723
rect 615 -746 624 -726
rect 644 -743 676 -726
rect 697 -743 702 -723
rect 644 -746 702 -743
rect 615 -753 702 -746
rect 727 -726 764 -656
rect 1030 -657 1067 -656
rect 1322 -660 1363 -652
rect 1322 -680 1330 -660
rect 1349 -680 1363 -660
rect 1322 -682 1363 -680
rect 1391 -660 1433 -652
rect 1391 -680 1407 -660
rect 1426 -680 1433 -660
rect 1659 -653 1665 -631
rect 1691 -651 2105 -631
rect 1691 -653 1700 -651
rect 1937 -652 2105 -651
rect 1659 -662 1700 -653
rect 1391 -682 1433 -680
rect 1322 -697 1433 -682
rect 879 -716 915 -715
rect 727 -746 736 -726
rect 756 -746 764 -726
rect 615 -755 671 -753
rect 615 -756 652 -755
rect 727 -756 764 -746
rect 823 -726 971 -716
rect 1071 -719 1167 -717
rect 823 -746 832 -726
rect 852 -746 942 -726
rect 962 -746 971 -726
rect 823 -755 971 -746
rect 1029 -726 1167 -719
rect 1029 -746 1038 -726
rect 1058 -746 1167 -726
rect 1029 -755 1167 -746
rect 823 -756 860 -755
rect 879 -807 915 -755
rect 934 -756 971 -755
rect 1030 -756 1067 -755
rect 350 -809 391 -808
rect 242 -816 391 -809
rect 242 -836 360 -816
rect 380 -836 391 -816
rect 242 -844 391 -836
rect 458 -812 817 -808
rect 458 -817 780 -812
rect 458 -841 571 -817
rect 595 -836 780 -817
rect 804 -836 817 -812
rect 595 -841 817 -836
rect 458 -844 817 -841
rect 879 -844 914 -807
rect 982 -810 1082 -807
rect 982 -814 1049 -810
rect 982 -840 994 -814
rect 1020 -836 1049 -814
rect 1075 -836 1082 -810
rect 1020 -840 1082 -836
rect 982 -844 1082 -840
rect 458 -865 489 -844
rect 879 -865 915 -844
rect 301 -866 338 -865
rect 300 -875 338 -866
rect 300 -895 309 -875
rect 329 -895 338 -875
rect 300 -903 338 -895
rect 404 -871 489 -865
rect 514 -866 551 -865
rect 404 -891 412 -871
rect 432 -891 489 -871
rect 404 -899 489 -891
rect 513 -875 551 -866
rect 513 -895 522 -875
rect 542 -895 551 -875
rect 404 -900 440 -899
rect 513 -903 551 -895
rect 617 -871 702 -865
rect 722 -866 759 -865
rect 617 -891 625 -871
rect 645 -872 702 -871
rect 645 -891 674 -872
rect 617 -892 674 -891
rect 695 -892 702 -872
rect 617 -899 702 -892
rect 721 -875 759 -866
rect 721 -895 730 -875
rect 750 -895 759 -875
rect 617 -900 653 -899
rect 721 -903 759 -895
rect 825 -871 969 -865
rect 825 -891 833 -871
rect 853 -874 941 -871
rect 853 -891 884 -874
rect 825 -894 884 -891
rect 907 -891 941 -874
rect 961 -891 969 -871
rect 907 -894 969 -891
rect 825 -899 969 -894
rect 825 -900 861 -899
rect 933 -900 969 -899
rect 1035 -866 1072 -865
rect 1035 -867 1073 -866
rect 1035 -875 1099 -867
rect 1035 -895 1044 -875
rect 1064 -889 1099 -875
rect 1119 -889 1122 -869
rect 1064 -894 1122 -889
rect 1064 -895 1099 -894
rect 301 -932 338 -903
rect 302 -934 338 -932
rect 514 -934 551 -903
rect 302 -956 551 -934
rect 722 -935 759 -903
rect 1035 -907 1099 -895
rect 1139 -933 1166 -755
rect 1464 -897 1574 -883
rect 1464 -900 1507 -897
rect 1464 -905 1468 -900
rect 998 -935 1166 -933
rect 722 -938 1166 -935
rect 383 -962 494 -956
rect 383 -970 424 -962
rect 72 -1025 111 -981
rect 383 -990 391 -970
rect 410 -990 424 -970
rect 383 -992 424 -990
rect 452 -970 494 -962
rect 452 -990 468 -970
rect 487 -990 494 -970
rect 452 -992 494 -990
rect 383 -1007 494 -992
rect 720 -961 1166 -938
rect 72 -1049 112 -1025
rect 412 -1049 459 -1047
rect 720 -1049 758 -961
rect 998 -962 1166 -961
rect 1386 -927 1468 -905
rect 1497 -927 1507 -900
rect 1535 -924 1542 -897
rect 1571 -905 1574 -897
rect 1571 -924 1636 -905
rect 1535 -927 1636 -924
rect 1386 -929 1636 -927
rect 1386 -1008 1423 -929
rect 1464 -942 1574 -929
rect 1538 -998 1569 -997
rect 1386 -1028 1395 -1008
rect 1415 -1028 1423 -1008
rect 1386 -1038 1423 -1028
rect 1482 -1008 1569 -998
rect 1482 -1028 1491 -1008
rect 1511 -1028 1569 -1008
rect 1482 -1037 1569 -1028
rect 1482 -1038 1519 -1037
rect 72 -1082 758 -1049
rect 72 -1139 111 -1082
rect 720 -1084 758 -1082
rect 1538 -1090 1569 -1037
rect 1599 -1008 1636 -929
rect 1807 -916 2200 -912
rect 1807 -933 1826 -916
rect 1846 -932 2200 -916
rect 2220 -932 2223 -912
rect 1846 -933 2223 -932
rect 1807 -937 2223 -933
rect 1807 -938 2148 -937
rect 1751 -998 1782 -997
rect 1599 -1028 1608 -1008
rect 1628 -1028 1636 -1008
rect 1599 -1038 1636 -1028
rect 1695 -1005 1782 -998
rect 1695 -1008 1756 -1005
rect 1695 -1028 1704 -1008
rect 1724 -1025 1756 -1008
rect 1777 -1025 1782 -1005
rect 1724 -1028 1782 -1025
rect 1695 -1035 1782 -1028
rect 1807 -1008 1844 -938
rect 2110 -939 2147 -938
rect 1959 -998 1995 -997
rect 1807 -1028 1816 -1008
rect 1836 -1028 1844 -1008
rect 1695 -1037 1751 -1035
rect 1695 -1038 1732 -1037
rect 1807 -1038 1844 -1028
rect 1903 -1008 2051 -998
rect 2151 -1001 2247 -999
rect 1903 -1028 1912 -1008
rect 1932 -1028 2022 -1008
rect 2042 -1028 2051 -1008
rect 1903 -1037 2051 -1028
rect 2109 -1008 2247 -1001
rect 2109 -1028 2118 -1008
rect 2138 -1028 2247 -1008
rect 2109 -1037 2247 -1028
rect 1903 -1038 1940 -1037
rect 1959 -1089 1995 -1037
rect 2014 -1038 2051 -1037
rect 2110 -1038 2147 -1037
rect 1430 -1091 1471 -1090
rect 1322 -1098 1471 -1091
rect 1322 -1118 1440 -1098
rect 1460 -1118 1471 -1098
rect 1322 -1126 1471 -1118
rect 1538 -1094 1897 -1090
rect 1538 -1099 1860 -1094
rect 1538 -1123 1651 -1099
rect 1675 -1118 1860 -1099
rect 1884 -1118 1897 -1094
rect 1675 -1123 1897 -1118
rect 1538 -1126 1897 -1123
rect 1959 -1126 1994 -1089
rect 2062 -1092 2162 -1089
rect 2062 -1096 2129 -1092
rect 2062 -1122 2074 -1096
rect 2100 -1118 2129 -1096
rect 2155 -1118 2162 -1092
rect 2100 -1122 2162 -1118
rect 2062 -1126 2162 -1122
rect 72 -1141 120 -1139
rect 72 -1159 83 -1141
rect 101 -1159 120 -1141
rect 1538 -1147 1569 -1126
rect 1959 -1147 1995 -1126
rect 1381 -1148 1418 -1147
rect 72 -1168 120 -1159
rect 73 -1169 120 -1168
rect 386 -1164 496 -1150
rect 386 -1167 429 -1164
rect 386 -1172 390 -1167
rect 308 -1194 390 -1172
rect 419 -1194 429 -1167
rect 457 -1191 464 -1164
rect 493 -1172 496 -1164
rect 1380 -1157 1418 -1148
rect 493 -1191 558 -1172
rect 1380 -1177 1389 -1157
rect 1409 -1177 1418 -1157
rect 457 -1194 558 -1191
rect 308 -1196 558 -1194
rect 76 -1232 113 -1231
rect 72 -1235 113 -1232
rect 72 -1240 114 -1235
rect 72 -1258 85 -1240
rect 103 -1258 114 -1240
rect 72 -1272 114 -1258
rect 152 -1272 199 -1268
rect 72 -1278 199 -1272
rect 72 -1307 160 -1278
rect 189 -1307 199 -1278
rect 308 -1275 345 -1196
rect 386 -1209 496 -1196
rect 460 -1265 491 -1264
rect 308 -1295 317 -1275
rect 337 -1295 345 -1275
rect 308 -1305 345 -1295
rect 404 -1275 491 -1265
rect 404 -1295 413 -1275
rect 433 -1295 491 -1275
rect 404 -1304 491 -1295
rect 404 -1305 441 -1304
rect 72 -1311 199 -1307
rect 72 -1328 111 -1311
rect 152 -1312 199 -1311
rect 72 -1346 83 -1328
rect 101 -1346 111 -1328
rect 72 -1355 111 -1346
rect 73 -1356 110 -1355
rect 460 -1357 491 -1304
rect 521 -1275 558 -1196
rect 729 -1199 1122 -1179
rect 1142 -1199 1145 -1179
rect 1380 -1185 1418 -1177
rect 1484 -1153 1569 -1147
rect 1594 -1148 1631 -1147
rect 1484 -1173 1492 -1153
rect 1512 -1173 1569 -1153
rect 1484 -1181 1569 -1173
rect 1593 -1157 1631 -1148
rect 1593 -1177 1602 -1157
rect 1622 -1177 1631 -1157
rect 1484 -1182 1520 -1181
rect 1593 -1185 1631 -1177
rect 1697 -1153 1782 -1147
rect 1802 -1148 1839 -1147
rect 1697 -1173 1705 -1153
rect 1725 -1154 1782 -1153
rect 1725 -1173 1754 -1154
rect 1697 -1174 1754 -1173
rect 1775 -1174 1782 -1154
rect 1697 -1181 1782 -1174
rect 1801 -1157 1839 -1148
rect 1801 -1177 1810 -1157
rect 1830 -1177 1839 -1157
rect 1697 -1182 1733 -1181
rect 1801 -1185 1839 -1177
rect 1905 -1153 2049 -1147
rect 1905 -1173 1913 -1153
rect 1933 -1155 2021 -1153
rect 1933 -1173 1962 -1155
rect 1905 -1176 1962 -1173
rect 1989 -1173 2021 -1155
rect 2041 -1173 2049 -1153
rect 1989 -1176 2049 -1173
rect 1905 -1181 2049 -1176
rect 1905 -1182 1941 -1181
rect 2013 -1182 2049 -1181
rect 2115 -1148 2152 -1147
rect 2115 -1149 2153 -1148
rect 2115 -1157 2179 -1149
rect 2115 -1177 2124 -1157
rect 2144 -1171 2179 -1157
rect 2199 -1171 2202 -1151
rect 2144 -1176 2202 -1171
rect 2144 -1177 2179 -1176
rect 729 -1204 1145 -1199
rect 729 -1205 1070 -1204
rect 673 -1265 704 -1264
rect 521 -1295 530 -1275
rect 550 -1295 558 -1275
rect 521 -1305 558 -1295
rect 617 -1272 704 -1265
rect 617 -1275 678 -1272
rect 617 -1295 626 -1275
rect 646 -1292 678 -1275
rect 699 -1292 704 -1272
rect 646 -1295 704 -1292
rect 617 -1302 704 -1295
rect 729 -1275 766 -1205
rect 1032 -1206 1069 -1205
rect 1381 -1214 1418 -1185
rect 1382 -1216 1418 -1214
rect 1594 -1216 1631 -1185
rect 1382 -1238 1631 -1216
rect 1802 -1217 1839 -1185
rect 2115 -1189 2179 -1177
rect 2219 -1215 2246 -1037
rect 2078 -1217 2246 -1215
rect 1799 -1224 2246 -1217
rect 1463 -1244 1574 -1238
rect 1463 -1252 1504 -1244
rect 881 -1265 917 -1264
rect 729 -1295 738 -1275
rect 758 -1295 766 -1275
rect 617 -1304 673 -1302
rect 617 -1305 654 -1304
rect 729 -1305 766 -1295
rect 825 -1275 973 -1265
rect 1073 -1268 1169 -1266
rect 825 -1295 834 -1275
rect 854 -1295 944 -1275
rect 964 -1295 973 -1275
rect 825 -1304 973 -1295
rect 1031 -1275 1169 -1268
rect 1031 -1295 1040 -1275
rect 1060 -1295 1169 -1275
rect 1463 -1272 1471 -1252
rect 1490 -1272 1504 -1252
rect 1463 -1274 1504 -1272
rect 1532 -1252 1574 -1244
rect 1532 -1272 1548 -1252
rect 1567 -1272 1574 -1252
rect 1799 -1251 1824 -1224
rect 1855 -1243 2246 -1224
rect 1855 -1251 1904 -1243
rect 2078 -1244 2246 -1243
rect 1799 -1253 1904 -1251
rect 1532 -1274 1574 -1272
rect 1463 -1289 1574 -1274
rect 1031 -1304 1169 -1295
rect 825 -1305 862 -1304
rect 881 -1356 917 -1304
rect 936 -1305 973 -1304
rect 1032 -1305 1069 -1304
rect 352 -1358 393 -1357
rect 244 -1365 393 -1358
rect 244 -1385 362 -1365
rect 382 -1385 393 -1365
rect 244 -1393 393 -1385
rect 460 -1361 819 -1357
rect 460 -1366 782 -1361
rect 460 -1390 573 -1366
rect 597 -1385 782 -1366
rect 806 -1385 819 -1361
rect 597 -1390 819 -1385
rect 460 -1393 819 -1390
rect 881 -1393 916 -1356
rect 984 -1359 1084 -1356
rect 984 -1363 1051 -1359
rect 984 -1389 996 -1363
rect 1022 -1385 1051 -1363
rect 1077 -1385 1084 -1359
rect 1022 -1389 1084 -1385
rect 984 -1393 1084 -1389
rect 460 -1414 491 -1393
rect 881 -1414 917 -1393
rect 303 -1415 340 -1414
rect 77 -1418 111 -1417
rect 76 -1427 113 -1418
rect 76 -1445 85 -1427
rect 103 -1445 113 -1427
rect 76 -1455 113 -1445
rect 302 -1424 340 -1415
rect 302 -1444 311 -1424
rect 331 -1444 340 -1424
rect 302 -1452 340 -1444
rect 406 -1420 491 -1414
rect 516 -1415 553 -1414
rect 406 -1440 414 -1420
rect 434 -1440 491 -1420
rect 406 -1448 491 -1440
rect 515 -1424 553 -1415
rect 515 -1444 524 -1424
rect 544 -1444 553 -1424
rect 406 -1449 442 -1448
rect 515 -1452 553 -1444
rect 619 -1420 704 -1414
rect 724 -1415 761 -1414
rect 619 -1440 627 -1420
rect 647 -1421 704 -1420
rect 647 -1440 676 -1421
rect 619 -1441 676 -1440
rect 697 -1441 704 -1421
rect 619 -1448 704 -1441
rect 723 -1424 761 -1415
rect 723 -1444 732 -1424
rect 752 -1444 761 -1424
rect 619 -1449 655 -1448
rect 723 -1452 761 -1444
rect 827 -1420 971 -1414
rect 827 -1440 835 -1420
rect 855 -1421 943 -1420
rect 855 -1440 886 -1421
rect 827 -1441 886 -1440
rect 911 -1440 943 -1421
rect 963 -1440 971 -1420
rect 911 -1441 971 -1440
rect 827 -1448 971 -1441
rect 827 -1449 863 -1448
rect 935 -1449 971 -1448
rect 1037 -1415 1074 -1414
rect 1037 -1416 1075 -1415
rect 1037 -1424 1101 -1416
rect 1037 -1444 1046 -1424
rect 1066 -1438 1101 -1424
rect 1121 -1438 1124 -1418
rect 1066 -1443 1124 -1438
rect 1066 -1444 1101 -1443
rect 77 -1483 111 -1455
rect 303 -1481 340 -1452
rect 304 -1483 340 -1481
rect 516 -1483 553 -1452
rect 77 -1484 249 -1483
rect 77 -1516 263 -1484
rect 304 -1505 553 -1483
rect 724 -1484 761 -1452
rect 1037 -1456 1101 -1444
rect 1141 -1482 1168 -1304
rect 1324 -1408 1434 -1394
rect 1324 -1411 1367 -1408
rect 1324 -1416 1328 -1411
rect 1000 -1484 1168 -1482
rect 724 -1490 1168 -1484
rect 77 -1548 111 -1516
rect 73 -1557 111 -1548
rect 73 -1575 83 -1557
rect 101 -1575 111 -1557
rect 73 -1581 111 -1575
rect 229 -1579 263 -1516
rect 385 -1511 496 -1505
rect 385 -1519 426 -1511
rect 385 -1539 393 -1519
rect 412 -1539 426 -1519
rect 385 -1541 426 -1539
rect 454 -1519 496 -1511
rect 454 -1539 470 -1519
rect 489 -1539 496 -1519
rect 454 -1541 496 -1539
rect 385 -1556 496 -1541
rect 723 -1510 1168 -1490
rect 723 -1579 761 -1510
rect 1000 -1511 1168 -1510
rect 1246 -1438 1328 -1416
rect 1357 -1438 1367 -1411
rect 1395 -1435 1402 -1408
rect 1431 -1416 1434 -1408
rect 1431 -1435 1496 -1416
rect 1395 -1438 1496 -1435
rect 1246 -1440 1496 -1438
rect 1246 -1519 1283 -1440
rect 1324 -1453 1434 -1440
rect 1398 -1509 1429 -1508
rect 1246 -1539 1255 -1519
rect 1275 -1539 1283 -1519
rect 1246 -1549 1283 -1539
rect 1342 -1519 1429 -1509
rect 1342 -1539 1351 -1519
rect 1371 -1539 1429 -1519
rect 1342 -1548 1429 -1539
rect 1342 -1549 1379 -1548
rect 73 -1585 110 -1581
rect 229 -1590 761 -1579
rect 228 -1606 761 -1590
rect 1398 -1601 1429 -1548
rect 1459 -1519 1496 -1440
rect 1667 -1430 2060 -1423
rect 1667 -1447 1675 -1430
rect 1707 -1443 2060 -1430
rect 2080 -1443 2083 -1423
rect 1707 -1447 2083 -1443
rect 1667 -1448 2083 -1447
rect 1667 -1449 2008 -1448
rect 1611 -1509 1642 -1508
rect 1459 -1539 1468 -1519
rect 1488 -1539 1496 -1519
rect 1459 -1549 1496 -1539
rect 1555 -1516 1642 -1509
rect 1555 -1519 1616 -1516
rect 1555 -1539 1564 -1519
rect 1584 -1536 1616 -1519
rect 1637 -1536 1642 -1516
rect 1584 -1539 1642 -1536
rect 1555 -1546 1642 -1539
rect 1667 -1519 1704 -1449
rect 1970 -1450 2007 -1449
rect 1819 -1509 1855 -1508
rect 1667 -1539 1676 -1519
rect 1696 -1539 1704 -1519
rect 1555 -1548 1611 -1546
rect 1555 -1549 1592 -1548
rect 1667 -1549 1704 -1539
rect 1763 -1519 1911 -1509
rect 2011 -1512 2107 -1510
rect 1763 -1539 1772 -1519
rect 1792 -1524 1882 -1519
rect 1792 -1539 1827 -1524
rect 1763 -1548 1827 -1539
rect 1763 -1549 1800 -1548
rect 1819 -1565 1827 -1548
rect 1848 -1539 1882 -1524
rect 1902 -1539 1911 -1519
rect 1848 -1548 1911 -1539
rect 1969 -1519 2107 -1512
rect 1969 -1539 1978 -1519
rect 1998 -1539 2107 -1519
rect 1969 -1548 2107 -1539
rect 1848 -1565 1855 -1548
rect 1874 -1549 1911 -1548
rect 1970 -1549 2007 -1548
rect 1819 -1600 1855 -1565
rect 1290 -1602 1331 -1601
rect 228 -1607 742 -1606
rect 1182 -1609 1331 -1602
rect 1182 -1629 1300 -1609
rect 1320 -1629 1331 -1609
rect 1182 -1637 1331 -1629
rect 1398 -1605 1757 -1601
rect 1398 -1610 1720 -1605
rect 1398 -1634 1511 -1610
rect 1535 -1629 1720 -1610
rect 1744 -1629 1757 -1605
rect 1535 -1634 1757 -1629
rect 1398 -1637 1757 -1634
rect 1819 -1637 1854 -1600
rect 1922 -1603 2022 -1600
rect 1922 -1607 1989 -1603
rect 1922 -1633 1934 -1607
rect 1960 -1629 1989 -1607
rect 2015 -1629 2022 -1603
rect 1960 -1633 2022 -1629
rect 1922 -1637 2022 -1633
rect 76 -1648 113 -1647
rect 74 -1656 114 -1648
rect 74 -1674 85 -1656
rect 103 -1674 114 -1656
rect 1398 -1658 1429 -1637
rect 1819 -1658 1855 -1637
rect 1241 -1659 1278 -1658
rect 74 -1722 114 -1674
rect 1240 -1668 1278 -1659
rect 1240 -1688 1249 -1668
rect 1269 -1688 1278 -1668
rect 1240 -1696 1278 -1688
rect 1344 -1664 1429 -1658
rect 1454 -1659 1491 -1658
rect 1344 -1684 1352 -1664
rect 1372 -1684 1429 -1664
rect 1344 -1692 1429 -1684
rect 1453 -1668 1491 -1659
rect 1453 -1688 1462 -1668
rect 1482 -1688 1491 -1668
rect 1344 -1693 1380 -1692
rect 1453 -1696 1491 -1688
rect 1557 -1664 1642 -1658
rect 1662 -1659 1699 -1658
rect 1557 -1684 1565 -1664
rect 1585 -1665 1642 -1664
rect 1585 -1684 1614 -1665
rect 1557 -1685 1614 -1684
rect 1635 -1685 1642 -1665
rect 1557 -1692 1642 -1685
rect 1661 -1668 1699 -1659
rect 1661 -1688 1670 -1668
rect 1690 -1688 1699 -1668
rect 1557 -1693 1593 -1692
rect 1661 -1696 1699 -1688
rect 1765 -1664 1909 -1658
rect 1765 -1684 1773 -1664
rect 1793 -1684 1881 -1664
rect 1901 -1684 1909 -1664
rect 1765 -1692 1909 -1684
rect 1765 -1693 1801 -1692
rect 1873 -1693 1909 -1692
rect 1975 -1659 2012 -1658
rect 1975 -1660 2013 -1659
rect 1975 -1668 2039 -1660
rect 1975 -1688 1984 -1668
rect 2004 -1682 2039 -1668
rect 2059 -1682 2062 -1662
rect 2004 -1687 2062 -1682
rect 2004 -1688 2039 -1687
rect 385 -1718 495 -1704
rect 385 -1721 428 -1718
rect 74 -1729 199 -1722
rect 385 -1726 389 -1721
rect 74 -1748 166 -1729
rect 191 -1748 199 -1729
rect 74 -1758 199 -1748
rect 307 -1748 389 -1726
rect 418 -1748 428 -1721
rect 456 -1745 463 -1718
rect 492 -1726 495 -1718
rect 1241 -1725 1278 -1696
rect 492 -1745 557 -1726
rect 1242 -1727 1278 -1725
rect 1454 -1727 1491 -1696
rect 1662 -1723 1699 -1696
rect 1975 -1700 2039 -1688
rect 456 -1748 557 -1745
rect 307 -1750 557 -1748
rect 74 -1778 114 -1758
rect 73 -1787 114 -1778
rect 73 -1805 83 -1787
rect 101 -1805 114 -1787
rect 73 -1814 114 -1805
rect 73 -1815 110 -1814
rect 307 -1829 344 -1750
rect 385 -1763 495 -1750
rect 459 -1819 490 -1818
rect 307 -1849 316 -1829
rect 336 -1849 344 -1829
rect 307 -1859 344 -1849
rect 403 -1829 490 -1819
rect 403 -1849 412 -1829
rect 432 -1849 490 -1829
rect 403 -1858 490 -1849
rect 403 -1859 440 -1858
rect 76 -1881 113 -1877
rect 73 -1886 113 -1881
rect 73 -1904 85 -1886
rect 103 -1904 113 -1886
rect 73 -2084 113 -1904
rect 459 -1911 490 -1858
rect 520 -1829 557 -1750
rect 728 -1753 1121 -1733
rect 1141 -1753 1144 -1733
rect 1242 -1749 1491 -1727
rect 1660 -1728 1701 -1723
rect 2079 -1726 2106 -1548
rect 1938 -1728 2106 -1726
rect 1660 -1734 2106 -1728
rect 728 -1758 1144 -1753
rect 1323 -1755 1434 -1749
rect 728 -1759 1069 -1758
rect 672 -1819 703 -1818
rect 520 -1849 529 -1829
rect 549 -1849 557 -1829
rect 520 -1859 557 -1849
rect 616 -1826 703 -1819
rect 616 -1829 677 -1826
rect 616 -1849 625 -1829
rect 645 -1846 677 -1829
rect 698 -1846 703 -1826
rect 645 -1849 703 -1846
rect 616 -1856 703 -1849
rect 728 -1829 765 -1759
rect 1031 -1760 1068 -1759
rect 1323 -1763 1364 -1755
rect 1323 -1783 1331 -1763
rect 1350 -1783 1364 -1763
rect 1323 -1785 1364 -1783
rect 1392 -1763 1434 -1755
rect 1392 -1783 1408 -1763
rect 1427 -1783 1434 -1763
rect 1660 -1756 1666 -1734
rect 1692 -1754 2106 -1734
rect 1692 -1756 1701 -1754
rect 1938 -1755 2106 -1754
rect 1660 -1765 1701 -1756
rect 1392 -1785 1434 -1783
rect 1323 -1800 1434 -1785
rect 880 -1819 916 -1818
rect 728 -1849 737 -1829
rect 757 -1849 765 -1829
rect 616 -1858 672 -1856
rect 616 -1859 653 -1858
rect 728 -1859 765 -1849
rect 824 -1829 972 -1819
rect 1072 -1822 1168 -1820
rect 824 -1849 833 -1829
rect 853 -1849 943 -1829
rect 963 -1849 972 -1829
rect 824 -1858 972 -1849
rect 1030 -1829 1168 -1822
rect 1030 -1849 1039 -1829
rect 1059 -1849 1168 -1829
rect 1030 -1858 1168 -1849
rect 824 -1859 861 -1858
rect 880 -1910 916 -1858
rect 935 -1859 972 -1858
rect 1031 -1859 1068 -1858
rect 351 -1912 392 -1911
rect 243 -1919 392 -1912
rect 243 -1939 361 -1919
rect 381 -1939 392 -1919
rect 243 -1947 392 -1939
rect 459 -1915 818 -1911
rect 459 -1920 781 -1915
rect 459 -1944 572 -1920
rect 596 -1939 781 -1920
rect 805 -1939 818 -1915
rect 596 -1944 818 -1939
rect 459 -1947 818 -1944
rect 880 -1947 915 -1910
rect 983 -1913 1083 -1910
rect 983 -1917 1050 -1913
rect 983 -1943 995 -1917
rect 1021 -1939 1050 -1917
rect 1076 -1939 1083 -1913
rect 1021 -1943 1083 -1939
rect 983 -1947 1083 -1943
rect 459 -1968 490 -1947
rect 880 -1968 916 -1947
rect 302 -1969 339 -1968
rect 301 -1978 339 -1969
rect 301 -1998 310 -1978
rect 330 -1998 339 -1978
rect 301 -2006 339 -1998
rect 405 -1974 490 -1968
rect 515 -1969 552 -1968
rect 405 -1994 413 -1974
rect 433 -1994 490 -1974
rect 405 -2002 490 -1994
rect 514 -1978 552 -1969
rect 514 -1998 523 -1978
rect 543 -1998 552 -1978
rect 405 -2003 441 -2002
rect 514 -2006 552 -1998
rect 618 -1974 703 -1968
rect 723 -1969 760 -1968
rect 618 -1994 626 -1974
rect 646 -1975 703 -1974
rect 646 -1994 675 -1975
rect 618 -1995 675 -1994
rect 696 -1995 703 -1975
rect 618 -2002 703 -1995
rect 722 -1978 760 -1969
rect 722 -1998 731 -1978
rect 751 -1998 760 -1978
rect 618 -2003 654 -2002
rect 722 -2006 760 -1998
rect 826 -1974 970 -1968
rect 826 -1994 834 -1974
rect 854 -1977 942 -1974
rect 854 -1994 885 -1977
rect 826 -1997 885 -1994
rect 908 -1994 942 -1977
rect 962 -1994 970 -1974
rect 908 -1997 970 -1994
rect 826 -2002 970 -1997
rect 826 -2003 862 -2002
rect 934 -2003 970 -2002
rect 1036 -1969 1073 -1968
rect 1036 -1970 1074 -1969
rect 1036 -1978 1100 -1970
rect 1036 -1998 1045 -1978
rect 1065 -1992 1100 -1978
rect 1120 -1992 1123 -1972
rect 1065 -1997 1123 -1992
rect 1065 -1998 1100 -1997
rect 302 -2035 339 -2006
rect 303 -2037 339 -2035
rect 515 -2037 552 -2006
rect 303 -2059 552 -2037
rect 723 -2038 760 -2006
rect 1036 -2010 1100 -1998
rect 1140 -2036 1167 -1858
rect 1434 -1987 1544 -1973
rect 1434 -1990 1477 -1987
rect 1434 -1995 1438 -1990
rect 999 -2038 1167 -2036
rect 723 -2041 1167 -2038
rect 384 -2065 495 -2059
rect 384 -2073 425 -2065
rect 73 -2128 112 -2084
rect 384 -2093 392 -2073
rect 411 -2093 425 -2073
rect 384 -2095 425 -2093
rect 453 -2073 495 -2065
rect 453 -2093 469 -2073
rect 488 -2093 495 -2073
rect 453 -2095 495 -2093
rect 384 -2109 495 -2095
rect 721 -2064 1167 -2041
rect 73 -2152 113 -2128
rect 413 -2152 460 -2150
rect 721 -2152 759 -2064
rect 999 -2065 1167 -2064
rect 1356 -2017 1438 -1995
rect 1467 -2017 1477 -1990
rect 1505 -2014 1512 -1987
rect 1541 -1995 1544 -1987
rect 1541 -2014 1606 -1995
rect 1505 -2017 1606 -2014
rect 1356 -2019 1606 -2017
rect 1356 -2098 1393 -2019
rect 1434 -2032 1544 -2019
rect 1508 -2088 1539 -2087
rect 1356 -2118 1365 -2098
rect 1385 -2118 1393 -2098
rect 1356 -2128 1393 -2118
rect 1452 -2098 1539 -2088
rect 1452 -2118 1461 -2098
rect 1481 -2118 1539 -2098
rect 1452 -2127 1539 -2118
rect 1452 -2128 1489 -2127
rect 73 -2185 759 -2152
rect 1508 -2180 1539 -2127
rect 1569 -2098 1606 -2019
rect 1777 -2000 1809 -1988
rect 1777 -2020 1779 -2000
rect 1800 -2002 1809 -2000
rect 1800 -2004 2152 -2002
rect 1800 -2020 2170 -2004
rect 1777 -2022 2170 -2020
rect 2190 -2022 2193 -2004
rect 1777 -2027 2193 -2022
rect 1777 -2028 2118 -2027
rect 1721 -2088 1752 -2087
rect 1569 -2118 1578 -2098
rect 1598 -2118 1606 -2098
rect 1569 -2128 1606 -2118
rect 1665 -2095 1752 -2088
rect 1665 -2098 1726 -2095
rect 1665 -2118 1674 -2098
rect 1694 -2115 1726 -2098
rect 1747 -2115 1752 -2095
rect 1694 -2118 1752 -2115
rect 1665 -2125 1752 -2118
rect 1777 -2098 1814 -2028
rect 2080 -2029 2117 -2028
rect 1929 -2088 1965 -2087
rect 1777 -2118 1786 -2098
rect 1806 -2118 1814 -2098
rect 1665 -2127 1721 -2125
rect 1665 -2128 1702 -2127
rect 1777 -2128 1814 -2118
rect 1873 -2098 2021 -2088
rect 2121 -2091 2217 -2089
rect 1873 -2118 1882 -2098
rect 1902 -2107 1992 -2098
rect 1902 -2118 1933 -2107
rect 1873 -2127 1933 -2118
rect 1873 -2128 1910 -2127
rect 1929 -2139 1933 -2127
rect 1960 -2118 1992 -2107
rect 2012 -2118 2021 -2098
rect 1960 -2127 2021 -2118
rect 2079 -2098 2217 -2091
rect 2079 -2118 2088 -2098
rect 2108 -2118 2217 -2098
rect 2079 -2127 2217 -2118
rect 1960 -2139 1965 -2127
rect 1984 -2128 2021 -2127
rect 2080 -2128 2117 -2127
rect 1929 -2179 1965 -2139
rect 1400 -2181 1441 -2180
rect 72 -2242 111 -2185
rect 721 -2187 759 -2185
rect 1292 -2188 1441 -2181
rect 1292 -2208 1410 -2188
rect 1430 -2208 1441 -2188
rect 1292 -2216 1441 -2208
rect 1508 -2184 1867 -2180
rect 1508 -2189 1830 -2184
rect 1508 -2213 1621 -2189
rect 1645 -2208 1830 -2189
rect 1854 -2208 1867 -2184
rect 1645 -2213 1867 -2208
rect 1508 -2216 1867 -2213
rect 1929 -2216 1964 -2179
rect 2032 -2182 2132 -2179
rect 2032 -2186 2099 -2182
rect 2032 -2212 2044 -2186
rect 2070 -2208 2099 -2186
rect 2125 -2208 2132 -2182
rect 2070 -2212 2132 -2208
rect 2032 -2216 2132 -2212
rect 1508 -2237 1539 -2216
rect 1929 -2237 1965 -2216
rect 1351 -2238 1388 -2237
rect 72 -2244 120 -2242
rect 72 -2262 83 -2244
rect 101 -2262 120 -2244
rect 1350 -2247 1388 -2238
rect 72 -2271 120 -2262
rect 73 -2272 120 -2271
rect 386 -2267 496 -2253
rect 386 -2270 429 -2267
rect 386 -2275 390 -2270
rect 308 -2297 390 -2275
rect 419 -2297 429 -2270
rect 457 -2294 464 -2267
rect 493 -2275 496 -2267
rect 1350 -2267 1359 -2247
rect 1379 -2267 1388 -2247
rect 1350 -2275 1388 -2267
rect 1454 -2243 1539 -2237
rect 1564 -2238 1601 -2237
rect 1454 -2263 1462 -2243
rect 1482 -2263 1539 -2243
rect 1454 -2271 1539 -2263
rect 1563 -2247 1601 -2238
rect 1563 -2267 1572 -2247
rect 1592 -2267 1601 -2247
rect 1454 -2272 1490 -2271
rect 1563 -2275 1601 -2267
rect 1667 -2243 1752 -2237
rect 1772 -2238 1809 -2237
rect 1667 -2263 1675 -2243
rect 1695 -2244 1752 -2243
rect 1695 -2263 1724 -2244
rect 1667 -2264 1724 -2263
rect 1745 -2264 1752 -2244
rect 1667 -2271 1752 -2264
rect 1771 -2247 1809 -2238
rect 1771 -2267 1780 -2247
rect 1800 -2267 1809 -2247
rect 1667 -2272 1703 -2271
rect 1771 -2275 1809 -2267
rect 1875 -2243 2019 -2237
rect 1875 -2263 1883 -2243
rect 1903 -2263 1991 -2243
rect 2011 -2263 2019 -2243
rect 1875 -2271 2019 -2263
rect 1875 -2272 1911 -2271
rect 1983 -2272 2019 -2271
rect 2085 -2238 2122 -2237
rect 2085 -2239 2123 -2238
rect 2085 -2247 2149 -2239
rect 2085 -2267 2094 -2247
rect 2114 -2261 2149 -2247
rect 2169 -2261 2172 -2241
rect 2114 -2266 2172 -2261
rect 2114 -2267 2149 -2266
rect 493 -2294 558 -2275
rect 457 -2297 558 -2294
rect 308 -2299 558 -2297
rect 76 -2335 113 -2334
rect 72 -2338 113 -2335
rect 72 -2343 114 -2338
rect 72 -2361 85 -2343
rect 103 -2361 114 -2343
rect 72 -2375 114 -2361
rect 152 -2375 199 -2371
rect 72 -2381 199 -2375
rect 72 -2410 160 -2381
rect 189 -2410 199 -2381
rect 308 -2378 345 -2299
rect 386 -2312 496 -2299
rect 460 -2368 491 -2367
rect 308 -2398 317 -2378
rect 337 -2398 345 -2378
rect 308 -2408 345 -2398
rect 404 -2378 491 -2368
rect 404 -2398 413 -2378
rect 433 -2398 491 -2378
rect 404 -2407 491 -2398
rect 404 -2408 441 -2407
rect 72 -2414 199 -2410
rect 72 -2431 111 -2414
rect 152 -2415 199 -2414
rect 72 -2449 83 -2431
rect 101 -2449 111 -2431
rect 72 -2458 111 -2449
rect 73 -2459 110 -2458
rect 460 -2460 491 -2407
rect 521 -2378 558 -2299
rect 729 -2302 1122 -2282
rect 1142 -2302 1145 -2282
rect 729 -2307 1145 -2302
rect 1351 -2304 1388 -2275
rect 1352 -2306 1388 -2304
rect 1564 -2306 1601 -2275
rect 729 -2308 1070 -2307
rect 673 -2368 704 -2367
rect 521 -2398 530 -2378
rect 550 -2398 558 -2378
rect 521 -2408 558 -2398
rect 617 -2375 704 -2368
rect 617 -2378 678 -2375
rect 617 -2398 626 -2378
rect 646 -2395 678 -2378
rect 699 -2395 704 -2375
rect 646 -2398 704 -2395
rect 617 -2405 704 -2398
rect 729 -2378 766 -2308
rect 1032 -2309 1069 -2308
rect 1352 -2328 1601 -2306
rect 1772 -2307 1809 -2275
rect 2085 -2279 2149 -2267
rect 2189 -2297 2216 -2127
rect 2137 -2305 2216 -2297
rect 2048 -2307 2216 -2305
rect 1772 -2314 2216 -2307
rect 1433 -2334 1544 -2328
rect 1772 -2333 2142 -2314
rect 2048 -2334 2142 -2333
rect 1433 -2342 1474 -2334
rect 1433 -2362 1441 -2342
rect 1460 -2362 1474 -2342
rect 1433 -2364 1474 -2362
rect 1502 -2342 1544 -2334
rect 1502 -2362 1518 -2342
rect 1537 -2362 1544 -2342
rect 2137 -2343 2142 -2334
rect 2190 -2334 2216 -2314
rect 2190 -2343 2207 -2334
rect 2137 -2352 2207 -2343
rect 1502 -2364 1544 -2362
rect 881 -2368 917 -2367
rect 729 -2398 738 -2378
rect 758 -2398 766 -2378
rect 617 -2407 673 -2405
rect 617 -2408 654 -2407
rect 729 -2408 766 -2398
rect 825 -2378 973 -2368
rect 1073 -2371 1169 -2369
rect 825 -2398 834 -2378
rect 854 -2398 944 -2378
rect 964 -2398 973 -2378
rect 825 -2407 973 -2398
rect 1031 -2378 1169 -2371
rect 1031 -2398 1040 -2378
rect 1060 -2398 1169 -2378
rect 1433 -2379 1544 -2364
rect 1031 -2407 1169 -2398
rect 825 -2408 862 -2407
rect 881 -2459 917 -2407
rect 936 -2408 973 -2407
rect 1032 -2408 1069 -2407
rect 352 -2461 393 -2460
rect 244 -2468 393 -2461
rect 244 -2488 362 -2468
rect 382 -2488 393 -2468
rect 244 -2496 393 -2488
rect 460 -2464 819 -2460
rect 460 -2469 782 -2464
rect 460 -2493 573 -2469
rect 597 -2488 782 -2469
rect 806 -2488 819 -2464
rect 597 -2493 819 -2488
rect 460 -2496 819 -2493
rect 881 -2496 916 -2459
rect 984 -2462 1084 -2459
rect 984 -2466 1051 -2462
rect 984 -2492 996 -2466
rect 1022 -2488 1051 -2466
rect 1077 -2488 1084 -2462
rect 1022 -2492 1084 -2488
rect 984 -2496 1084 -2492
rect 460 -2517 491 -2496
rect 881 -2517 917 -2496
rect 303 -2518 340 -2517
rect 77 -2521 111 -2520
rect 76 -2530 113 -2521
rect 76 -2548 85 -2530
rect 103 -2548 113 -2530
rect 76 -2558 113 -2548
rect 302 -2527 340 -2518
rect 302 -2547 311 -2527
rect 331 -2547 340 -2527
rect 302 -2555 340 -2547
rect 406 -2523 491 -2517
rect 516 -2518 553 -2517
rect 406 -2543 414 -2523
rect 434 -2543 491 -2523
rect 406 -2551 491 -2543
rect 515 -2527 553 -2518
rect 515 -2547 524 -2527
rect 544 -2547 553 -2527
rect 406 -2552 442 -2551
rect 515 -2555 553 -2547
rect 619 -2523 704 -2517
rect 724 -2518 761 -2517
rect 619 -2543 627 -2523
rect 647 -2524 704 -2523
rect 647 -2543 676 -2524
rect 619 -2544 676 -2543
rect 697 -2544 704 -2524
rect 619 -2551 704 -2544
rect 723 -2527 761 -2518
rect 723 -2547 732 -2527
rect 752 -2547 761 -2527
rect 619 -2552 655 -2551
rect 723 -2555 761 -2547
rect 827 -2523 971 -2517
rect 827 -2543 835 -2523
rect 855 -2524 943 -2523
rect 855 -2543 886 -2524
rect 827 -2544 886 -2543
rect 911 -2543 943 -2524
rect 963 -2543 971 -2523
rect 911 -2544 971 -2543
rect 827 -2551 971 -2544
rect 827 -2552 863 -2551
rect 935 -2552 971 -2551
rect 1037 -2518 1074 -2517
rect 1037 -2519 1075 -2518
rect 1037 -2527 1101 -2519
rect 1037 -2547 1046 -2527
rect 1066 -2541 1101 -2527
rect 1121 -2541 1124 -2521
rect 1066 -2546 1124 -2541
rect 1066 -2547 1101 -2546
rect 77 -2586 111 -2558
rect 303 -2584 340 -2555
rect 304 -2586 340 -2584
rect 516 -2586 553 -2555
rect 77 -2587 249 -2586
rect 77 -2619 263 -2587
rect 304 -2608 553 -2586
rect 724 -2587 761 -2555
rect 1037 -2559 1101 -2547
rect 1141 -2585 1168 -2407
rect 1324 -2511 1434 -2497
rect 1324 -2514 1367 -2511
rect 1324 -2519 1328 -2514
rect 1000 -2587 1168 -2585
rect 724 -2593 1168 -2587
rect 77 -2651 111 -2619
rect 73 -2660 111 -2651
rect 73 -2678 83 -2660
rect 101 -2678 111 -2660
rect 73 -2684 111 -2678
rect 229 -2682 263 -2619
rect 385 -2614 496 -2608
rect 385 -2622 426 -2614
rect 385 -2642 393 -2622
rect 412 -2642 426 -2622
rect 385 -2644 426 -2642
rect 454 -2622 496 -2614
rect 454 -2642 470 -2622
rect 489 -2642 496 -2622
rect 454 -2644 496 -2642
rect 385 -2659 496 -2644
rect 723 -2613 1168 -2593
rect 723 -2682 761 -2613
rect 1000 -2614 1168 -2613
rect 1246 -2541 1328 -2519
rect 1357 -2541 1367 -2514
rect 1395 -2538 1402 -2511
rect 1431 -2519 1434 -2511
rect 1431 -2538 1496 -2519
rect 1395 -2541 1496 -2538
rect 1246 -2543 1496 -2541
rect 1246 -2622 1283 -2543
rect 1324 -2556 1434 -2543
rect 1398 -2612 1429 -2611
rect 1246 -2642 1255 -2622
rect 1275 -2642 1283 -2622
rect 1246 -2652 1283 -2642
rect 1342 -2622 1429 -2612
rect 1342 -2642 1351 -2622
rect 1371 -2642 1429 -2622
rect 1342 -2651 1429 -2642
rect 1342 -2652 1379 -2651
rect 73 -2688 110 -2684
rect 229 -2693 761 -2682
rect 228 -2709 761 -2693
rect 1398 -2704 1429 -2651
rect 1459 -2622 1496 -2543
rect 1667 -2546 2060 -2526
rect 2080 -2546 2083 -2526
rect 1667 -2551 2083 -2546
rect 1667 -2552 2008 -2551
rect 1611 -2612 1642 -2611
rect 1459 -2642 1468 -2622
rect 1488 -2642 1496 -2622
rect 1459 -2652 1496 -2642
rect 1555 -2619 1642 -2612
rect 1555 -2622 1616 -2619
rect 1555 -2642 1564 -2622
rect 1584 -2639 1616 -2622
rect 1637 -2639 1642 -2619
rect 1584 -2642 1642 -2639
rect 1555 -2649 1642 -2642
rect 1667 -2622 1704 -2552
rect 1970 -2553 2007 -2552
rect 1819 -2612 1855 -2611
rect 1667 -2642 1676 -2622
rect 1696 -2642 1704 -2622
rect 1555 -2651 1611 -2649
rect 1555 -2652 1592 -2651
rect 1667 -2652 1704 -2642
rect 1763 -2622 1911 -2612
rect 2011 -2615 2107 -2613
rect 1763 -2642 1772 -2622
rect 1792 -2642 1882 -2622
rect 1902 -2642 1911 -2622
rect 1763 -2651 1911 -2642
rect 1969 -2622 2107 -2615
rect 1969 -2642 1978 -2622
rect 1998 -2642 2107 -2622
rect 1969 -2651 2107 -2642
rect 1763 -2652 1800 -2651
rect 1819 -2703 1855 -2651
rect 1874 -2652 1911 -2651
rect 1970 -2652 2007 -2651
rect 1290 -2705 1331 -2704
rect 228 -2710 742 -2709
rect 1182 -2712 1331 -2705
rect 1182 -2732 1300 -2712
rect 1320 -2732 1331 -2712
rect 1182 -2740 1331 -2732
rect 1398 -2708 1757 -2704
rect 1398 -2713 1720 -2708
rect 1398 -2737 1511 -2713
rect 1535 -2732 1720 -2713
rect 1744 -2732 1757 -2708
rect 1535 -2737 1757 -2732
rect 1398 -2740 1757 -2737
rect 1819 -2740 1854 -2703
rect 1922 -2706 2022 -2703
rect 1922 -2710 1989 -2706
rect 1922 -2736 1934 -2710
rect 1960 -2732 1989 -2710
rect 2015 -2732 2022 -2706
rect 1960 -2736 2022 -2732
rect 1922 -2740 2022 -2736
rect 76 -2751 113 -2750
rect 74 -2759 114 -2751
rect 74 -2777 85 -2759
rect 103 -2777 114 -2759
rect 1398 -2761 1429 -2740
rect 1819 -2761 1855 -2740
rect 1241 -2762 1278 -2761
rect 74 -2825 114 -2777
rect 1240 -2771 1278 -2762
rect 1240 -2791 1249 -2771
rect 1269 -2791 1278 -2771
rect 1240 -2799 1278 -2791
rect 1344 -2767 1429 -2761
rect 1454 -2762 1491 -2761
rect 1344 -2787 1352 -2767
rect 1372 -2787 1429 -2767
rect 1344 -2795 1429 -2787
rect 1453 -2771 1491 -2762
rect 1453 -2791 1462 -2771
rect 1482 -2791 1491 -2771
rect 1344 -2796 1380 -2795
rect 1453 -2799 1491 -2791
rect 1557 -2767 1642 -2761
rect 1662 -2762 1699 -2761
rect 1557 -2787 1565 -2767
rect 1585 -2768 1642 -2767
rect 1585 -2787 1614 -2768
rect 1557 -2788 1614 -2787
rect 1635 -2788 1642 -2768
rect 1557 -2795 1642 -2788
rect 1661 -2771 1699 -2762
rect 1661 -2791 1670 -2771
rect 1690 -2791 1699 -2771
rect 1557 -2796 1593 -2795
rect 1661 -2799 1699 -2791
rect 1765 -2767 1909 -2761
rect 1765 -2787 1773 -2767
rect 1793 -2784 1829 -2767
rect 1849 -2784 1881 -2767
rect 1793 -2787 1881 -2784
rect 1901 -2787 1909 -2767
rect 1765 -2795 1909 -2787
rect 1765 -2796 1801 -2795
rect 1873 -2796 1909 -2795
rect 1975 -2762 2012 -2761
rect 1975 -2763 2013 -2762
rect 1975 -2771 2039 -2763
rect 1975 -2791 1984 -2771
rect 2004 -2785 2039 -2771
rect 2059 -2785 2062 -2765
rect 2004 -2790 2062 -2785
rect 2004 -2791 2039 -2790
rect 385 -2821 495 -2807
rect 385 -2824 428 -2821
rect 74 -2832 199 -2825
rect 385 -2829 389 -2824
rect 74 -2851 166 -2832
rect 191 -2851 199 -2832
rect 74 -2861 199 -2851
rect 307 -2851 389 -2829
rect 418 -2851 428 -2824
rect 456 -2848 463 -2821
rect 492 -2829 495 -2821
rect 1241 -2828 1278 -2799
rect 492 -2848 557 -2829
rect 1242 -2830 1278 -2828
rect 1454 -2830 1491 -2799
rect 1662 -2826 1699 -2799
rect 1975 -2803 2039 -2791
rect 456 -2851 557 -2848
rect 307 -2853 557 -2851
rect 74 -2881 114 -2861
rect 73 -2890 114 -2881
rect 73 -2908 83 -2890
rect 101 -2908 114 -2890
rect 73 -2917 114 -2908
rect 73 -2918 110 -2917
rect 307 -2932 344 -2853
rect 385 -2866 495 -2853
rect 459 -2922 490 -2921
rect 307 -2952 316 -2932
rect 336 -2952 344 -2932
rect 307 -2962 344 -2952
rect 403 -2932 490 -2922
rect 403 -2952 412 -2932
rect 432 -2952 490 -2932
rect 403 -2961 490 -2952
rect 403 -2962 440 -2961
rect 76 -2984 113 -2980
rect 73 -2989 113 -2984
rect 73 -3007 85 -2989
rect 103 -3007 113 -2989
rect 73 -3187 113 -3007
rect 459 -3014 490 -2961
rect 520 -2932 557 -2853
rect 728 -2856 1121 -2836
rect 1141 -2856 1144 -2836
rect 1242 -2852 1491 -2830
rect 1660 -2831 1701 -2826
rect 2079 -2829 2106 -2651
rect 1938 -2831 2106 -2829
rect 1660 -2837 2106 -2831
rect 728 -2861 1144 -2856
rect 1323 -2858 1434 -2852
rect 728 -2862 1069 -2861
rect 672 -2922 703 -2921
rect 520 -2952 529 -2932
rect 549 -2952 557 -2932
rect 520 -2962 557 -2952
rect 616 -2929 703 -2922
rect 616 -2932 677 -2929
rect 616 -2952 625 -2932
rect 645 -2949 677 -2932
rect 698 -2949 703 -2929
rect 645 -2952 703 -2949
rect 616 -2959 703 -2952
rect 728 -2932 765 -2862
rect 1031 -2863 1068 -2862
rect 1323 -2866 1364 -2858
rect 1323 -2886 1331 -2866
rect 1350 -2886 1364 -2866
rect 1323 -2888 1364 -2886
rect 1392 -2866 1434 -2858
rect 1392 -2886 1408 -2866
rect 1427 -2886 1434 -2866
rect 1660 -2859 1666 -2837
rect 1692 -2857 2106 -2837
rect 1692 -2859 1701 -2857
rect 1938 -2858 2106 -2857
rect 1660 -2868 1701 -2859
rect 1392 -2888 1434 -2886
rect 1323 -2903 1434 -2888
rect 880 -2922 916 -2921
rect 728 -2952 737 -2932
rect 757 -2952 765 -2932
rect 616 -2961 672 -2959
rect 616 -2962 653 -2961
rect 728 -2962 765 -2952
rect 824 -2932 972 -2922
rect 1072 -2925 1168 -2923
rect 824 -2952 833 -2932
rect 853 -2952 943 -2932
rect 963 -2952 972 -2932
rect 824 -2961 972 -2952
rect 1030 -2932 1168 -2925
rect 1030 -2952 1039 -2932
rect 1059 -2952 1168 -2932
rect 1030 -2961 1168 -2952
rect 824 -2962 861 -2961
rect 880 -3013 916 -2961
rect 935 -2962 972 -2961
rect 1031 -2962 1068 -2961
rect 351 -3015 392 -3014
rect 243 -3022 392 -3015
rect 243 -3042 361 -3022
rect 381 -3042 392 -3022
rect 243 -3050 392 -3042
rect 459 -3018 818 -3014
rect 459 -3023 781 -3018
rect 459 -3047 572 -3023
rect 596 -3042 781 -3023
rect 805 -3042 818 -3018
rect 596 -3047 818 -3042
rect 459 -3050 818 -3047
rect 880 -3050 915 -3013
rect 983 -3016 1083 -3013
rect 983 -3020 1050 -3016
rect 983 -3046 995 -3020
rect 1021 -3042 1050 -3020
rect 1076 -3042 1083 -3016
rect 1021 -3046 1083 -3042
rect 983 -3050 1083 -3046
rect 459 -3071 490 -3050
rect 880 -3071 916 -3050
rect 302 -3072 339 -3071
rect 301 -3081 339 -3072
rect 301 -3101 310 -3081
rect 330 -3101 339 -3081
rect 301 -3109 339 -3101
rect 405 -3077 490 -3071
rect 515 -3072 552 -3071
rect 405 -3097 413 -3077
rect 433 -3097 490 -3077
rect 405 -3105 490 -3097
rect 514 -3081 552 -3072
rect 514 -3101 523 -3081
rect 543 -3101 552 -3081
rect 405 -3106 441 -3105
rect 514 -3109 552 -3101
rect 618 -3077 703 -3071
rect 723 -3072 760 -3071
rect 618 -3097 626 -3077
rect 646 -3078 703 -3077
rect 646 -3097 675 -3078
rect 618 -3098 675 -3097
rect 696 -3098 703 -3078
rect 618 -3105 703 -3098
rect 722 -3081 760 -3072
rect 722 -3101 731 -3081
rect 751 -3101 760 -3081
rect 618 -3106 654 -3105
rect 722 -3109 760 -3101
rect 826 -3077 970 -3071
rect 826 -3097 834 -3077
rect 854 -3080 942 -3077
rect 854 -3097 885 -3080
rect 826 -3100 885 -3097
rect 908 -3097 942 -3080
rect 962 -3097 970 -3077
rect 908 -3100 970 -3097
rect 826 -3105 970 -3100
rect 826 -3106 862 -3105
rect 934 -3106 970 -3105
rect 1036 -3072 1073 -3071
rect 1036 -3073 1074 -3072
rect 1036 -3081 1100 -3073
rect 1036 -3101 1045 -3081
rect 1065 -3095 1100 -3081
rect 1120 -3095 1123 -3075
rect 1065 -3100 1123 -3095
rect 1065 -3101 1100 -3100
rect 302 -3138 339 -3109
rect 303 -3140 339 -3138
rect 515 -3140 552 -3109
rect 303 -3162 552 -3140
rect 723 -3141 760 -3109
rect 1036 -3113 1100 -3101
rect 1140 -3139 1167 -2961
rect 1465 -3103 1575 -3089
rect 1465 -3106 1508 -3103
rect 1465 -3111 1469 -3106
rect 999 -3141 1167 -3139
rect 723 -3144 1167 -3141
rect 384 -3168 495 -3162
rect 384 -3176 425 -3168
rect 73 -3231 112 -3187
rect 384 -3196 392 -3176
rect 411 -3196 425 -3176
rect 384 -3198 425 -3196
rect 453 -3176 495 -3168
rect 453 -3196 469 -3176
rect 488 -3196 495 -3176
rect 453 -3198 495 -3196
rect 384 -3213 495 -3198
rect 721 -3167 1167 -3144
rect 73 -3255 113 -3231
rect 413 -3255 460 -3253
rect 721 -3255 759 -3167
rect 999 -3168 1167 -3167
rect 1387 -3133 1469 -3111
rect 1498 -3133 1508 -3106
rect 1536 -3130 1543 -3103
rect 1572 -3111 1575 -3103
rect 1572 -3130 1637 -3111
rect 1536 -3133 1637 -3130
rect 1387 -3135 1637 -3133
rect 1387 -3214 1424 -3135
rect 1465 -3148 1575 -3135
rect 1539 -3204 1570 -3203
rect 1387 -3234 1396 -3214
rect 1416 -3234 1424 -3214
rect 1387 -3244 1424 -3234
rect 1483 -3214 1570 -3204
rect 1483 -3234 1492 -3214
rect 1512 -3234 1570 -3214
rect 1483 -3243 1570 -3234
rect 1483 -3244 1520 -3243
rect 73 -3288 759 -3255
rect 73 -3345 112 -3288
rect 721 -3290 759 -3288
rect 1539 -3296 1570 -3243
rect 1600 -3214 1637 -3135
rect 1808 -3122 2201 -3118
rect 1808 -3139 1827 -3122
rect 1847 -3138 2201 -3122
rect 2221 -3138 2224 -3118
rect 1847 -3139 2224 -3138
rect 1808 -3143 2224 -3139
rect 1808 -3144 2149 -3143
rect 1752 -3204 1783 -3203
rect 1600 -3234 1609 -3214
rect 1629 -3234 1637 -3214
rect 1600 -3244 1637 -3234
rect 1696 -3211 1783 -3204
rect 1696 -3214 1757 -3211
rect 1696 -3234 1705 -3214
rect 1725 -3231 1757 -3214
rect 1778 -3231 1783 -3211
rect 1725 -3234 1783 -3231
rect 1696 -3241 1783 -3234
rect 1808 -3214 1845 -3144
rect 2111 -3145 2148 -3144
rect 1960 -3204 1996 -3203
rect 1808 -3234 1817 -3214
rect 1837 -3234 1845 -3214
rect 1696 -3243 1752 -3241
rect 1696 -3244 1733 -3243
rect 1808 -3244 1845 -3234
rect 1904 -3214 2052 -3204
rect 2220 -3205 2249 -3204
rect 2152 -3207 2249 -3205
rect 1904 -3234 1913 -3214
rect 1933 -3218 2023 -3214
rect 1933 -3234 1966 -3218
rect 1904 -3243 1966 -3234
rect 1904 -3244 1941 -3243
rect 1960 -3256 1966 -3243
rect 1989 -3234 2023 -3218
rect 2043 -3234 2052 -3214
rect 1989 -3243 2052 -3234
rect 2110 -3214 2249 -3207
rect 2110 -3234 2119 -3214
rect 2139 -3234 2249 -3214
rect 2110 -3243 2249 -3234
rect 1989 -3256 1996 -3243
rect 2015 -3244 2052 -3243
rect 2111 -3244 2148 -3243
rect 1960 -3295 1996 -3256
rect 1431 -3297 1472 -3296
rect 1323 -3304 1472 -3297
rect 1323 -3324 1441 -3304
rect 1461 -3324 1472 -3304
rect 1323 -3332 1472 -3324
rect 1539 -3300 1898 -3296
rect 1539 -3305 1861 -3300
rect 1539 -3329 1652 -3305
rect 1676 -3324 1861 -3305
rect 1885 -3324 1898 -3300
rect 1676 -3329 1898 -3324
rect 1539 -3332 1898 -3329
rect 1960 -3332 1995 -3295
rect 2063 -3298 2163 -3295
rect 2063 -3302 2130 -3298
rect 2063 -3328 2075 -3302
rect 2101 -3324 2130 -3302
rect 2156 -3324 2163 -3298
rect 2101 -3328 2163 -3324
rect 2063 -3332 2163 -3328
rect 73 -3347 121 -3345
rect 73 -3365 84 -3347
rect 102 -3365 121 -3347
rect 1539 -3353 1570 -3332
rect 1960 -3353 1996 -3332
rect 1382 -3354 1419 -3353
rect 73 -3374 121 -3365
rect 74 -3375 121 -3374
rect 387 -3370 497 -3356
rect 387 -3373 430 -3370
rect 387 -3378 391 -3373
rect 309 -3400 391 -3378
rect 420 -3400 430 -3373
rect 458 -3397 465 -3370
rect 494 -3378 497 -3370
rect 1381 -3363 1419 -3354
rect 494 -3397 559 -3378
rect 1381 -3383 1390 -3363
rect 1410 -3383 1419 -3363
rect 458 -3400 559 -3397
rect 309 -3402 559 -3400
rect 77 -3438 114 -3437
rect 73 -3441 114 -3438
rect 73 -3446 115 -3441
rect 73 -3464 86 -3446
rect 104 -3464 115 -3446
rect 73 -3478 115 -3464
rect 153 -3478 200 -3474
rect 73 -3484 200 -3478
rect 73 -3513 161 -3484
rect 190 -3513 200 -3484
rect 309 -3481 346 -3402
rect 387 -3415 497 -3402
rect 461 -3471 492 -3470
rect 309 -3501 318 -3481
rect 338 -3501 346 -3481
rect 309 -3511 346 -3501
rect 405 -3481 492 -3471
rect 405 -3501 414 -3481
rect 434 -3501 492 -3481
rect 405 -3510 492 -3501
rect 405 -3511 442 -3510
rect 73 -3517 200 -3513
rect 73 -3534 112 -3517
rect 153 -3518 200 -3517
rect 73 -3552 84 -3534
rect 102 -3552 112 -3534
rect 73 -3561 112 -3552
rect 74 -3562 111 -3561
rect 461 -3563 492 -3510
rect 522 -3481 559 -3402
rect 730 -3405 1123 -3385
rect 1143 -3405 1146 -3385
rect 1381 -3391 1419 -3383
rect 1485 -3359 1570 -3353
rect 1595 -3354 1632 -3353
rect 1485 -3379 1493 -3359
rect 1513 -3379 1570 -3359
rect 1485 -3387 1570 -3379
rect 1594 -3363 1632 -3354
rect 1594 -3383 1603 -3363
rect 1623 -3383 1632 -3363
rect 1485 -3388 1521 -3387
rect 1594 -3391 1632 -3383
rect 1698 -3359 1783 -3353
rect 1803 -3354 1840 -3353
rect 1698 -3379 1706 -3359
rect 1726 -3360 1783 -3359
rect 1726 -3379 1755 -3360
rect 1698 -3380 1755 -3379
rect 1776 -3380 1783 -3360
rect 1698 -3387 1783 -3380
rect 1802 -3363 1840 -3354
rect 1802 -3383 1811 -3363
rect 1831 -3383 1840 -3363
rect 1698 -3388 1734 -3387
rect 1802 -3391 1840 -3383
rect 1906 -3359 2050 -3353
rect 1906 -3379 1914 -3359
rect 1934 -3379 2022 -3359
rect 2042 -3379 2050 -3359
rect 1906 -3387 2050 -3379
rect 1906 -3388 1942 -3387
rect 2014 -3388 2050 -3387
rect 2116 -3354 2153 -3353
rect 2116 -3355 2154 -3354
rect 2116 -3363 2180 -3355
rect 2116 -3383 2125 -3363
rect 2145 -3377 2180 -3363
rect 2200 -3377 2203 -3357
rect 2145 -3382 2203 -3377
rect 2145 -3383 2180 -3382
rect 730 -3410 1146 -3405
rect 730 -3411 1071 -3410
rect 674 -3471 705 -3470
rect 522 -3501 531 -3481
rect 551 -3501 559 -3481
rect 522 -3511 559 -3501
rect 618 -3478 705 -3471
rect 618 -3481 679 -3478
rect 618 -3501 627 -3481
rect 647 -3498 679 -3481
rect 700 -3498 705 -3478
rect 647 -3501 705 -3498
rect 618 -3508 705 -3501
rect 730 -3481 767 -3411
rect 1033 -3412 1070 -3411
rect 1382 -3420 1419 -3391
rect 1383 -3422 1419 -3420
rect 1595 -3422 1632 -3391
rect 1383 -3444 1632 -3422
rect 1803 -3423 1840 -3391
rect 2116 -3395 2180 -3383
rect 2220 -3421 2249 -3243
rect 2079 -3423 2249 -3421
rect 1800 -3430 2249 -3423
rect 1464 -3450 1575 -3444
rect 1464 -3458 1505 -3450
rect 882 -3471 918 -3470
rect 730 -3501 739 -3481
rect 759 -3501 767 -3481
rect 618 -3510 674 -3508
rect 618 -3511 655 -3510
rect 730 -3511 767 -3501
rect 826 -3481 974 -3471
rect 1074 -3474 1170 -3472
rect 826 -3501 835 -3481
rect 855 -3501 945 -3481
rect 965 -3501 974 -3481
rect 826 -3510 974 -3501
rect 1032 -3481 1170 -3474
rect 1032 -3501 1041 -3481
rect 1061 -3501 1170 -3481
rect 1464 -3478 1472 -3458
rect 1491 -3478 1505 -3458
rect 1464 -3480 1505 -3478
rect 1533 -3458 1575 -3450
rect 1533 -3478 1549 -3458
rect 1568 -3478 1575 -3458
rect 1800 -3457 1825 -3430
rect 1856 -3449 2249 -3430
rect 1856 -3457 1905 -3449
rect 2079 -3450 2249 -3449
rect 1800 -3459 1905 -3457
rect 1533 -3480 1575 -3478
rect 1464 -3495 1575 -3480
rect 1032 -3510 1170 -3501
rect 826 -3511 863 -3510
rect 882 -3562 918 -3510
rect 937 -3511 974 -3510
rect 1033 -3511 1070 -3510
rect 353 -3564 394 -3563
rect 245 -3571 394 -3564
rect 245 -3591 363 -3571
rect 383 -3591 394 -3571
rect 245 -3599 394 -3591
rect 461 -3567 820 -3563
rect 461 -3572 783 -3567
rect 461 -3596 574 -3572
rect 598 -3591 783 -3572
rect 807 -3591 820 -3567
rect 598 -3596 820 -3591
rect 461 -3599 820 -3596
rect 882 -3599 917 -3562
rect 985 -3565 1085 -3562
rect 985 -3569 1052 -3565
rect 985 -3595 997 -3569
rect 1023 -3591 1052 -3569
rect 1078 -3591 1085 -3565
rect 1023 -3595 1085 -3591
rect 985 -3599 1085 -3595
rect 461 -3620 492 -3599
rect 882 -3620 918 -3599
rect 304 -3621 341 -3620
rect 78 -3624 112 -3623
rect 77 -3633 114 -3624
rect 77 -3651 86 -3633
rect 104 -3651 114 -3633
rect 77 -3661 114 -3651
rect 303 -3630 341 -3621
rect 303 -3650 312 -3630
rect 332 -3650 341 -3630
rect 303 -3658 341 -3650
rect 407 -3626 492 -3620
rect 517 -3621 554 -3620
rect 407 -3646 415 -3626
rect 435 -3646 492 -3626
rect 407 -3654 492 -3646
rect 516 -3630 554 -3621
rect 516 -3650 525 -3630
rect 545 -3650 554 -3630
rect 407 -3655 443 -3654
rect 516 -3658 554 -3650
rect 620 -3626 705 -3620
rect 725 -3621 762 -3620
rect 620 -3646 628 -3626
rect 648 -3627 705 -3626
rect 648 -3646 677 -3627
rect 620 -3647 677 -3646
rect 698 -3647 705 -3627
rect 620 -3654 705 -3647
rect 724 -3630 762 -3621
rect 724 -3650 733 -3630
rect 753 -3650 762 -3630
rect 620 -3655 656 -3654
rect 724 -3658 762 -3650
rect 828 -3626 972 -3620
rect 828 -3646 836 -3626
rect 856 -3627 944 -3626
rect 856 -3646 887 -3627
rect 828 -3647 887 -3646
rect 912 -3646 944 -3627
rect 964 -3646 972 -3626
rect 912 -3647 972 -3646
rect 828 -3654 972 -3647
rect 828 -3655 864 -3654
rect 936 -3655 972 -3654
rect 1038 -3621 1075 -3620
rect 1038 -3622 1076 -3621
rect 1038 -3630 1102 -3622
rect 1038 -3650 1047 -3630
rect 1067 -3644 1102 -3630
rect 1122 -3644 1125 -3624
rect 1067 -3649 1125 -3644
rect 1067 -3650 1102 -3649
rect 78 -3689 112 -3661
rect 304 -3687 341 -3658
rect 305 -3689 341 -3687
rect 517 -3689 554 -3658
rect 78 -3690 250 -3689
rect 78 -3722 264 -3690
rect 305 -3711 554 -3689
rect 725 -3690 762 -3658
rect 1038 -3662 1102 -3650
rect 1142 -3688 1169 -3510
rect 1325 -3614 1435 -3600
rect 1325 -3617 1368 -3614
rect 1325 -3622 1329 -3617
rect 1001 -3690 1169 -3688
rect 725 -3696 1169 -3690
rect 78 -3754 112 -3722
rect 74 -3763 112 -3754
rect 74 -3781 84 -3763
rect 102 -3781 112 -3763
rect 74 -3787 112 -3781
rect 230 -3785 264 -3722
rect 386 -3717 497 -3711
rect 386 -3725 427 -3717
rect 386 -3745 394 -3725
rect 413 -3745 427 -3725
rect 386 -3747 427 -3745
rect 455 -3725 497 -3717
rect 455 -3745 471 -3725
rect 490 -3745 497 -3725
rect 455 -3747 497 -3745
rect 386 -3762 497 -3747
rect 724 -3716 1169 -3696
rect 724 -3785 762 -3716
rect 1001 -3717 1169 -3716
rect 1247 -3644 1329 -3622
rect 1358 -3644 1368 -3617
rect 1396 -3641 1403 -3614
rect 1432 -3622 1435 -3614
rect 1432 -3641 1497 -3622
rect 1396 -3644 1497 -3641
rect 1247 -3646 1497 -3644
rect 1247 -3725 1284 -3646
rect 1325 -3659 1435 -3646
rect 1399 -3715 1430 -3714
rect 1247 -3745 1256 -3725
rect 1276 -3745 1284 -3725
rect 1247 -3755 1284 -3745
rect 1343 -3725 1430 -3715
rect 1343 -3745 1352 -3725
rect 1372 -3745 1430 -3725
rect 1343 -3754 1430 -3745
rect 1343 -3755 1380 -3754
rect 74 -3791 111 -3787
rect 230 -3796 762 -3785
rect 229 -3812 762 -3796
rect 1399 -3807 1430 -3754
rect 1460 -3725 1497 -3646
rect 1668 -3636 2061 -3629
rect 1668 -3653 1676 -3636
rect 1708 -3649 2061 -3636
rect 2081 -3649 2084 -3629
rect 1708 -3653 2084 -3649
rect 1668 -3654 2084 -3653
rect 1668 -3655 2009 -3654
rect 1612 -3715 1643 -3714
rect 1460 -3745 1469 -3725
rect 1489 -3745 1497 -3725
rect 1460 -3755 1497 -3745
rect 1556 -3722 1643 -3715
rect 1556 -3725 1617 -3722
rect 1556 -3745 1565 -3725
rect 1585 -3742 1617 -3725
rect 1638 -3742 1643 -3722
rect 1585 -3745 1643 -3742
rect 1556 -3752 1643 -3745
rect 1668 -3725 1705 -3655
rect 1971 -3656 2008 -3655
rect 1820 -3715 1856 -3714
rect 1668 -3745 1677 -3725
rect 1697 -3745 1705 -3725
rect 1556 -3754 1612 -3752
rect 1556 -3755 1593 -3754
rect 1668 -3755 1705 -3745
rect 1764 -3725 1912 -3715
rect 2012 -3718 2108 -3716
rect 1764 -3745 1773 -3725
rect 1793 -3730 1883 -3725
rect 1793 -3745 1828 -3730
rect 1764 -3754 1828 -3745
rect 1764 -3755 1801 -3754
rect 1820 -3771 1828 -3754
rect 1849 -3745 1883 -3730
rect 1903 -3745 1912 -3725
rect 1849 -3754 1912 -3745
rect 1970 -3725 2108 -3718
rect 1970 -3745 1979 -3725
rect 1999 -3745 2108 -3725
rect 1970 -3754 2108 -3745
rect 1849 -3771 1856 -3754
rect 1875 -3755 1912 -3754
rect 1971 -3755 2008 -3754
rect 1820 -3806 1856 -3771
rect 1291 -3808 1332 -3807
rect 229 -3813 743 -3812
rect 1183 -3815 1332 -3808
rect 1183 -3835 1301 -3815
rect 1321 -3835 1332 -3815
rect 1183 -3843 1332 -3835
rect 1399 -3811 1758 -3807
rect 1399 -3816 1721 -3811
rect 1399 -3840 1512 -3816
rect 1536 -3835 1721 -3816
rect 1745 -3835 1758 -3811
rect 1536 -3840 1758 -3835
rect 1399 -3843 1758 -3840
rect 1820 -3843 1855 -3806
rect 1923 -3809 2023 -3806
rect 1923 -3813 1990 -3809
rect 1923 -3839 1935 -3813
rect 1961 -3835 1990 -3813
rect 2016 -3835 2023 -3809
rect 1961 -3839 2023 -3835
rect 1923 -3843 2023 -3839
rect 77 -3854 114 -3853
rect 75 -3862 115 -3854
rect 75 -3880 86 -3862
rect 104 -3880 115 -3862
rect 1399 -3864 1430 -3843
rect 1820 -3864 1856 -3843
rect 1242 -3865 1279 -3864
rect 75 -3928 115 -3880
rect 1241 -3874 1279 -3865
rect 1241 -3894 1250 -3874
rect 1270 -3894 1279 -3874
rect 1241 -3902 1279 -3894
rect 1345 -3870 1430 -3864
rect 1455 -3865 1492 -3864
rect 1345 -3890 1353 -3870
rect 1373 -3890 1430 -3870
rect 1345 -3898 1430 -3890
rect 1454 -3874 1492 -3865
rect 1454 -3894 1463 -3874
rect 1483 -3894 1492 -3874
rect 1345 -3899 1381 -3898
rect 1454 -3902 1492 -3894
rect 1558 -3870 1643 -3864
rect 1663 -3865 1700 -3864
rect 1558 -3890 1566 -3870
rect 1586 -3871 1643 -3870
rect 1586 -3890 1615 -3871
rect 1558 -3891 1615 -3890
rect 1636 -3891 1643 -3871
rect 1558 -3898 1643 -3891
rect 1662 -3874 1700 -3865
rect 1662 -3894 1671 -3874
rect 1691 -3894 1700 -3874
rect 1558 -3899 1594 -3898
rect 1662 -3902 1700 -3894
rect 1766 -3870 1910 -3864
rect 1766 -3890 1774 -3870
rect 1794 -3890 1882 -3870
rect 1902 -3890 1910 -3870
rect 1766 -3898 1910 -3890
rect 1766 -3899 1802 -3898
rect 1874 -3899 1910 -3898
rect 1976 -3865 2013 -3864
rect 1976 -3866 2014 -3865
rect 1976 -3874 2040 -3866
rect 1976 -3894 1985 -3874
rect 2005 -3888 2040 -3874
rect 2060 -3888 2063 -3868
rect 2005 -3893 2063 -3888
rect 2005 -3894 2040 -3893
rect 386 -3924 496 -3910
rect 386 -3927 429 -3924
rect 75 -3935 200 -3928
rect 386 -3932 390 -3927
rect 75 -3954 167 -3935
rect 192 -3954 200 -3935
rect 75 -3964 200 -3954
rect 308 -3954 390 -3932
rect 419 -3954 429 -3927
rect 457 -3951 464 -3924
rect 493 -3932 496 -3924
rect 1242 -3931 1279 -3902
rect 493 -3951 558 -3932
rect 1243 -3933 1279 -3931
rect 1455 -3933 1492 -3902
rect 1663 -3929 1700 -3902
rect 1976 -3906 2040 -3894
rect 457 -3954 558 -3951
rect 308 -3956 558 -3954
rect 75 -3984 115 -3964
rect 74 -3993 115 -3984
rect 74 -4011 84 -3993
rect 102 -4011 115 -3993
rect 74 -4020 115 -4011
rect 74 -4021 111 -4020
rect 308 -4035 345 -3956
rect 386 -3969 496 -3956
rect 460 -4025 491 -4024
rect 308 -4055 317 -4035
rect 337 -4055 345 -4035
rect 308 -4065 345 -4055
rect 404 -4035 491 -4025
rect 404 -4055 413 -4035
rect 433 -4055 491 -4035
rect 404 -4064 491 -4055
rect 404 -4065 441 -4064
rect 77 -4087 114 -4083
rect 74 -4092 114 -4087
rect 74 -4110 86 -4092
rect 104 -4110 114 -4092
rect 74 -4290 114 -4110
rect 460 -4117 491 -4064
rect 521 -4035 558 -3956
rect 729 -3959 1122 -3939
rect 1142 -3959 1145 -3939
rect 1243 -3955 1492 -3933
rect 1661 -3934 1702 -3929
rect 2080 -3932 2107 -3754
rect 1939 -3934 2107 -3932
rect 1661 -3940 2107 -3934
rect 729 -3964 1145 -3959
rect 1324 -3961 1435 -3955
rect 729 -3965 1070 -3964
rect 673 -4025 704 -4024
rect 521 -4055 530 -4035
rect 550 -4055 558 -4035
rect 521 -4065 558 -4055
rect 617 -4032 704 -4025
rect 617 -4035 678 -4032
rect 617 -4055 626 -4035
rect 646 -4052 678 -4035
rect 699 -4052 704 -4032
rect 646 -4055 704 -4052
rect 617 -4062 704 -4055
rect 729 -4035 766 -3965
rect 1032 -3966 1069 -3965
rect 1324 -3969 1365 -3961
rect 1324 -3989 1332 -3969
rect 1351 -3989 1365 -3969
rect 1324 -3991 1365 -3989
rect 1393 -3969 1435 -3961
rect 1393 -3989 1409 -3969
rect 1428 -3989 1435 -3969
rect 1661 -3962 1667 -3940
rect 1693 -3960 2107 -3940
rect 1693 -3962 1702 -3960
rect 1939 -3961 2107 -3960
rect 1661 -3971 1702 -3962
rect 1393 -3991 1435 -3989
rect 1324 -4006 1435 -3991
rect 881 -4025 917 -4024
rect 729 -4055 738 -4035
rect 758 -4055 766 -4035
rect 617 -4064 673 -4062
rect 617 -4065 654 -4064
rect 729 -4065 766 -4055
rect 825 -4035 973 -4025
rect 1073 -4028 1169 -4026
rect 825 -4055 834 -4035
rect 854 -4055 944 -4035
rect 964 -4055 973 -4035
rect 825 -4064 973 -4055
rect 1031 -4035 1169 -4028
rect 1031 -4055 1040 -4035
rect 1060 -4055 1169 -4035
rect 1031 -4064 1169 -4055
rect 825 -4065 862 -4064
rect 881 -4116 917 -4064
rect 936 -4065 973 -4064
rect 1032 -4065 1069 -4064
rect 352 -4118 393 -4117
rect 244 -4125 393 -4118
rect 244 -4145 362 -4125
rect 382 -4145 393 -4125
rect 244 -4153 393 -4145
rect 460 -4121 819 -4117
rect 460 -4126 782 -4121
rect 460 -4150 573 -4126
rect 597 -4145 782 -4126
rect 806 -4145 819 -4121
rect 597 -4150 819 -4145
rect 460 -4153 819 -4150
rect 881 -4153 916 -4116
rect 984 -4119 1084 -4116
rect 984 -4123 1051 -4119
rect 984 -4149 996 -4123
rect 1022 -4145 1051 -4123
rect 1077 -4145 1084 -4119
rect 1022 -4149 1084 -4145
rect 984 -4153 1084 -4149
rect 460 -4174 491 -4153
rect 881 -4174 917 -4153
rect 303 -4175 340 -4174
rect 302 -4184 340 -4175
rect 302 -4204 311 -4184
rect 331 -4204 340 -4184
rect 302 -4212 340 -4204
rect 406 -4180 491 -4174
rect 516 -4175 553 -4174
rect 406 -4200 414 -4180
rect 434 -4200 491 -4180
rect 406 -4208 491 -4200
rect 515 -4184 553 -4175
rect 515 -4204 524 -4184
rect 544 -4204 553 -4184
rect 406 -4209 442 -4208
rect 515 -4212 553 -4204
rect 619 -4180 704 -4174
rect 724 -4175 761 -4174
rect 619 -4200 627 -4180
rect 647 -4181 704 -4180
rect 647 -4200 676 -4181
rect 619 -4201 676 -4200
rect 697 -4201 704 -4181
rect 619 -4208 704 -4201
rect 723 -4184 761 -4175
rect 723 -4204 732 -4184
rect 752 -4204 761 -4184
rect 619 -4209 655 -4208
rect 723 -4212 761 -4204
rect 827 -4180 971 -4174
rect 827 -4200 835 -4180
rect 855 -4183 943 -4180
rect 855 -4200 886 -4183
rect 827 -4203 886 -4200
rect 909 -4200 943 -4183
rect 963 -4200 971 -4180
rect 909 -4203 971 -4200
rect 827 -4208 971 -4203
rect 827 -4209 863 -4208
rect 935 -4209 971 -4208
rect 1037 -4175 1074 -4174
rect 1037 -4176 1075 -4175
rect 1037 -4184 1101 -4176
rect 1037 -4204 1046 -4184
rect 1066 -4198 1101 -4184
rect 1121 -4198 1124 -4178
rect 1066 -4203 1124 -4198
rect 1066 -4204 1101 -4203
rect 303 -4241 340 -4212
rect 304 -4243 340 -4241
rect 516 -4243 553 -4212
rect 304 -4265 553 -4243
rect 724 -4244 761 -4212
rect 1037 -4216 1101 -4204
rect 1141 -4242 1168 -4064
rect 1000 -4244 1168 -4242
rect 724 -4247 1168 -4244
rect 385 -4271 496 -4265
rect 385 -4279 426 -4271
rect 74 -4334 113 -4290
rect 385 -4299 393 -4279
rect 412 -4299 426 -4279
rect 385 -4301 426 -4299
rect 454 -4279 496 -4271
rect 454 -4299 470 -4279
rect 489 -4299 496 -4279
rect 454 -4300 496 -4299
rect 722 -4270 1168 -4247
rect 454 -4301 497 -4300
rect 74 -4358 114 -4334
rect 385 -4340 497 -4301
rect 414 -4358 461 -4340
rect 722 -4358 760 -4270
rect 1000 -4271 1168 -4270
rect 74 -4391 760 -4358
rect 722 -4393 760 -4391
<< viali >>
rect 387 4321 416 4348
rect 461 4324 490 4351
rect 157 4208 186 4237
rect 1119 4316 1139 4336
rect 675 4223 696 4243
rect 1048 4130 1074 4156
rect 673 4074 694 4094
rect 883 4074 908 4094
rect 1098 4077 1118 4097
rect 390 3976 409 3996
rect 467 3976 486 3996
rect 1325 4077 1354 4104
rect 1399 4080 1428 4107
rect 2057 4072 2077 4092
rect 1613 3979 1634 3999
rect 1986 3886 2012 3912
rect 1611 3830 1632 3850
rect 1826 3834 1846 3851
rect 2036 3833 2056 3853
rect 163 3767 188 3786
rect 386 3767 415 3794
rect 460 3770 489 3797
rect 1118 3762 1138 3782
rect 674 3669 695 3689
rect 1328 3732 1347 3752
rect 1405 3732 1424 3752
rect 1663 3759 1689 3781
rect 1047 3576 1073 3602
rect 672 3520 693 3540
rect 882 3518 905 3538
rect 1097 3523 1117 3543
rect 389 3422 408 3442
rect 466 3422 485 3442
rect 1466 3485 1495 3512
rect 1540 3488 1569 3515
rect 1824 3479 1844 3496
rect 2198 3480 2218 3500
rect 1754 3387 1775 3407
rect 2127 3294 2153 3320
rect 388 3218 417 3245
rect 462 3221 491 3248
rect 158 3105 187 3134
rect 1120 3213 1140 3233
rect 1752 3238 1773 3258
rect 1960 3236 1987 3257
rect 2177 3241 2197 3261
rect 676 3120 697 3140
rect 1469 3140 1488 3160
rect 1546 3140 1565 3160
rect 1822 3161 1853 3188
rect 1049 3027 1075 3053
rect 674 2971 695 2991
rect 884 2971 909 2991
rect 1099 2974 1119 2994
rect 391 2873 410 2893
rect 468 2873 487 2893
rect 1326 2974 1355 3001
rect 1400 2977 1429 3004
rect 1673 2965 1705 2982
rect 2058 2969 2078 2989
rect 1614 2876 1635 2896
rect 1825 2847 1846 2888
rect 1987 2783 2013 2809
rect 1612 2727 1633 2747
rect 2037 2730 2057 2750
rect 164 2664 189 2683
rect 387 2664 416 2691
rect 461 2667 490 2694
rect 1119 2659 1139 2679
rect 675 2566 696 2586
rect 1329 2629 1348 2649
rect 1406 2629 1425 2649
rect 1664 2656 1690 2678
rect 1048 2473 1074 2499
rect 673 2417 694 2437
rect 883 2415 906 2435
rect 1098 2420 1118 2440
rect 390 2319 409 2339
rect 467 2319 486 2339
rect 1436 2395 1465 2422
rect 1510 2398 1539 2425
rect 2168 2390 2188 2410
rect 1724 2297 1745 2317
rect 2097 2204 2123 2230
rect 388 2115 417 2142
rect 462 2118 491 2145
rect 1722 2148 1743 2168
rect 1930 2148 1959 2167
rect 2147 2151 2167 2171
rect 158 2002 187 2031
rect 1120 2110 1140 2130
rect 676 2017 697 2037
rect 1439 2050 1458 2070
rect 1516 2050 1535 2070
rect 1049 1924 1075 1950
rect 674 1868 695 1888
rect 884 1868 909 1888
rect 1099 1871 1119 1891
rect 2140 1929 2188 1958
rect 391 1770 410 1790
rect 468 1770 487 1790
rect 1326 1871 1355 1898
rect 1400 1874 1429 1901
rect 2058 1866 2078 1886
rect 1614 1773 1635 1793
rect 1987 1680 2013 1706
rect 1612 1624 1633 1644
rect 1827 1628 1847 1645
rect 2037 1627 2057 1647
rect 164 1561 189 1580
rect 387 1561 416 1588
rect 461 1564 490 1591
rect 1119 1556 1139 1576
rect 675 1463 696 1483
rect 1329 1526 1348 1546
rect 1406 1526 1425 1546
rect 1664 1553 1690 1575
rect 1048 1370 1074 1396
rect 673 1314 694 1334
rect 883 1312 906 1332
rect 1098 1317 1118 1337
rect 390 1216 409 1236
rect 467 1216 486 1236
rect 1467 1279 1496 1306
rect 1541 1282 1570 1309
rect 1825 1273 1845 1290
rect 2199 1274 2219 1294
rect 1755 1181 1776 1201
rect 1964 1156 1987 1194
rect 2128 1088 2154 1114
rect 389 1012 418 1039
rect 463 1015 492 1042
rect 159 899 188 928
rect 1121 1007 1141 1027
rect 1753 1032 1774 1052
rect 2178 1035 2198 1055
rect 677 914 698 934
rect 1470 934 1489 954
rect 1547 934 1566 954
rect 1823 955 1854 982
rect 1050 821 1076 847
rect 675 765 696 785
rect 885 765 910 785
rect 1100 768 1120 788
rect 392 667 411 687
rect 469 667 488 687
rect 1327 768 1356 795
rect 1401 771 1430 798
rect 1674 759 1706 776
rect 2059 763 2079 783
rect 1615 670 1636 690
rect 1826 641 1847 682
rect 1988 577 2014 603
rect 1613 521 1634 541
rect 2038 524 2058 544
rect 165 458 190 477
rect 388 458 417 485
rect 462 461 491 488
rect 1120 453 1140 473
rect 676 360 697 380
rect 1330 423 1349 443
rect 1407 423 1426 443
rect 1665 450 1691 472
rect 1049 267 1075 293
rect 674 211 695 231
rect 884 209 907 229
rect 1099 214 1119 234
rect 391 113 410 133
rect 468 113 487 133
rect 1436 195 1465 222
rect 1510 198 1539 225
rect 2168 190 2188 210
rect 1724 97 1745 117
rect 2097 4 2123 30
rect 389 -91 418 -64
rect 463 -88 492 -61
rect 1722 -52 1743 -32
rect 2147 -49 2167 -29
rect 159 -204 188 -175
rect 1121 -96 1141 -76
rect 677 -189 698 -169
rect 1439 -150 1458 -130
rect 1516 -150 1535 -130
rect 1050 -282 1076 -256
rect 675 -338 696 -318
rect 885 -338 910 -318
rect 1100 -335 1120 -315
rect 2303 -287 2330 -247
rect 392 -436 411 -416
rect 469 -436 488 -416
rect 1327 -335 1356 -308
rect 1401 -332 1430 -305
rect 2059 -340 2079 -320
rect 1615 -433 1636 -413
rect 1988 -526 2014 -500
rect 1613 -582 1634 -562
rect 1828 -578 1848 -561
rect 2038 -579 2058 -559
rect 165 -645 190 -626
rect 388 -645 417 -618
rect 462 -642 491 -615
rect 1120 -650 1140 -630
rect 676 -743 697 -723
rect 1330 -680 1349 -660
rect 1407 -680 1426 -660
rect 1665 -653 1691 -631
rect 1049 -836 1075 -810
rect 674 -892 695 -872
rect 884 -894 907 -874
rect 1099 -889 1119 -869
rect 391 -990 410 -970
rect 468 -990 487 -970
rect 1468 -927 1497 -900
rect 1542 -924 1571 -897
rect 1826 -933 1846 -916
rect 2200 -932 2220 -912
rect 1756 -1025 1777 -1005
rect 2129 -1118 2155 -1092
rect 390 -1194 419 -1167
rect 464 -1191 493 -1164
rect 160 -1307 189 -1278
rect 1122 -1199 1142 -1179
rect 1754 -1174 1775 -1154
rect 1962 -1176 1989 -1155
rect 2179 -1171 2199 -1151
rect 678 -1292 699 -1272
rect 1471 -1272 1490 -1252
rect 1548 -1272 1567 -1252
rect 1824 -1251 1855 -1224
rect 1051 -1385 1077 -1359
rect 676 -1441 697 -1421
rect 886 -1441 911 -1421
rect 1101 -1438 1121 -1418
rect 393 -1539 412 -1519
rect 470 -1539 489 -1519
rect 1328 -1438 1357 -1411
rect 1402 -1435 1431 -1408
rect 1675 -1447 1707 -1430
rect 2060 -1443 2080 -1423
rect 1616 -1536 1637 -1516
rect 1827 -1565 1848 -1524
rect 1989 -1629 2015 -1603
rect 1614 -1685 1635 -1665
rect 2039 -1682 2059 -1662
rect 166 -1748 191 -1729
rect 389 -1748 418 -1721
rect 463 -1745 492 -1718
rect 1121 -1753 1141 -1733
rect 677 -1846 698 -1826
rect 1331 -1783 1350 -1763
rect 1408 -1783 1427 -1763
rect 1666 -1756 1692 -1734
rect 1050 -1939 1076 -1913
rect 675 -1995 696 -1975
rect 885 -1997 908 -1977
rect 1100 -1992 1120 -1972
rect 392 -2093 411 -2073
rect 469 -2093 488 -2073
rect 1438 -2017 1467 -1990
rect 1512 -2014 1541 -1987
rect 1779 -2020 1800 -2000
rect 2170 -2022 2190 -2004
rect 1726 -2115 1747 -2095
rect 1933 -2139 1960 -2107
rect 2099 -2208 2125 -2182
rect 390 -2297 419 -2270
rect 464 -2294 493 -2267
rect 1724 -2264 1745 -2244
rect 2149 -2261 2169 -2241
rect 160 -2410 189 -2381
rect 1122 -2302 1142 -2282
rect 678 -2395 699 -2375
rect 1441 -2362 1460 -2342
rect 1518 -2362 1537 -2342
rect 2142 -2343 2190 -2314
rect 1051 -2488 1077 -2462
rect 676 -2544 697 -2524
rect 886 -2544 911 -2524
rect 1101 -2541 1121 -2521
rect 393 -2642 412 -2622
rect 470 -2642 489 -2622
rect 1328 -2541 1357 -2514
rect 1402 -2538 1431 -2511
rect 2060 -2546 2080 -2526
rect 1616 -2639 1637 -2619
rect 1989 -2732 2015 -2706
rect 1614 -2788 1635 -2768
rect 1829 -2784 1849 -2767
rect 2039 -2785 2059 -2765
rect 166 -2851 191 -2832
rect 389 -2851 418 -2824
rect 463 -2848 492 -2821
rect 1121 -2856 1141 -2836
rect 677 -2949 698 -2929
rect 1331 -2886 1350 -2866
rect 1408 -2886 1427 -2866
rect 1666 -2859 1692 -2837
rect 1050 -3042 1076 -3016
rect 675 -3098 696 -3078
rect 885 -3100 908 -3080
rect 1100 -3095 1120 -3075
rect 392 -3196 411 -3176
rect 469 -3196 488 -3176
rect 1469 -3133 1498 -3106
rect 1543 -3130 1572 -3103
rect 1827 -3139 1847 -3122
rect 2201 -3138 2221 -3118
rect 1757 -3231 1778 -3211
rect 1966 -3256 1989 -3218
rect 2130 -3324 2156 -3298
rect 391 -3400 420 -3373
rect 465 -3397 494 -3370
rect 161 -3513 190 -3484
rect 1123 -3405 1143 -3385
rect 1755 -3380 1776 -3360
rect 2180 -3377 2200 -3357
rect 679 -3498 700 -3478
rect 1472 -3478 1491 -3458
rect 1549 -3478 1568 -3458
rect 1825 -3457 1856 -3430
rect 1052 -3591 1078 -3565
rect 677 -3647 698 -3627
rect 887 -3647 912 -3627
rect 1102 -3644 1122 -3624
rect 394 -3745 413 -3725
rect 471 -3745 490 -3725
rect 1329 -3644 1358 -3617
rect 1403 -3641 1432 -3614
rect 1676 -3653 1708 -3636
rect 2061 -3649 2081 -3629
rect 1617 -3742 1638 -3722
rect 1828 -3771 1849 -3730
rect 1990 -3835 2016 -3809
rect 1615 -3891 1636 -3871
rect 2040 -3888 2060 -3868
rect 167 -3954 192 -3935
rect 390 -3954 419 -3927
rect 464 -3951 493 -3924
rect 1122 -3959 1142 -3939
rect 678 -4052 699 -4032
rect 1332 -3989 1351 -3969
rect 1409 -3989 1428 -3969
rect 1667 -3962 1693 -3940
rect 1051 -4145 1077 -4119
rect 676 -4201 697 -4181
rect 886 -4203 909 -4183
rect 1101 -4198 1121 -4178
rect 393 -4299 412 -4279
rect 470 -4299 489 -4279
<< metal1 >>
rect 1114 4419 1149 4421
rect 150 4416 1149 4419
rect 149 4392 1149 4416
rect 149 4237 197 4392
rect 383 4351 493 4365
rect 383 4348 461 4351
rect 383 4321 387 4348
rect 416 4324 461 4348
rect 490 4324 493 4351
rect 1114 4341 1149 4392
rect 416 4321 493 4324
rect 383 4306 493 4321
rect 1112 4336 1149 4341
rect 1112 4316 1119 4336
rect 1139 4316 1149 4336
rect 1112 4309 1149 4316
rect 1112 4308 1147 4309
rect 149 4208 157 4237
rect 186 4208 197 4237
rect 149 4203 197 4208
rect 668 4243 700 4250
rect 668 4223 675 4243
rect 696 4223 700 4243
rect 668 4158 700 4223
rect 1038 4158 1078 4159
rect 668 4156 1080 4158
rect 668 4130 1048 4156
rect 1074 4130 1080 4156
rect 668 4122 1080 4130
rect 668 4094 700 4122
rect 1113 4102 1147 4308
rect 2051 4175 2085 4176
rect 1182 4140 2086 4175
rect 668 4074 673 4094
rect 694 4074 700 4094
rect 668 4067 700 4074
rect 875 4094 914 4100
rect 875 4074 883 4094
rect 908 4074 914 4094
rect 875 4067 914 4074
rect 1091 4097 1147 4102
rect 1091 4077 1098 4097
rect 1118 4077 1147 4097
rect 1091 4070 1147 4077
rect 1091 4069 1126 4070
rect 883 4021 914 4067
rect 382 3996 493 4018
rect 382 3976 390 3996
rect 409 3976 467 3996
rect 486 3976 493 3996
rect 882 4004 914 4021
rect 1183 4004 1220 4140
rect 1321 4107 1431 4121
rect 1321 4104 1399 4107
rect 1321 4077 1325 4104
rect 1354 4080 1399 4104
rect 1428 4080 1431 4107
rect 2051 4097 2085 4140
rect 1354 4077 1431 4080
rect 1321 4062 1431 4077
rect 2050 4092 2085 4097
rect 2050 4072 2057 4092
rect 2077 4072 2085 4092
rect 2050 4064 2085 4072
rect 882 3991 1220 4004
rect 382 3959 493 3976
rect 883 3972 1220 3991
rect 1162 3971 1220 3972
rect 1606 3999 1638 4006
rect 1606 3979 1613 3999
rect 1634 3979 1638 3999
rect 1606 3914 1638 3979
rect 1976 3914 2016 3915
rect 1606 3912 2018 3914
rect 1606 3886 1986 3912
rect 2012 3886 2018 3912
rect 1606 3878 2018 3886
rect 152 3839 1148 3865
rect 1606 3850 1638 3878
rect 154 3786 196 3839
rect 154 3767 163 3786
rect 188 3767 196 3786
rect 154 3757 196 3767
rect 382 3797 492 3811
rect 382 3794 460 3797
rect 382 3767 386 3794
rect 415 3770 460 3794
rect 489 3770 492 3797
rect 1112 3787 1146 3839
rect 1606 3830 1611 3850
rect 1632 3830 1638 3850
rect 1606 3823 1638 3830
rect 1816 3851 1854 3861
rect 2051 3858 2085 4064
rect 1816 3834 1826 3851
rect 1846 3834 1854 3851
rect 1657 3791 1698 3792
rect 415 3767 492 3770
rect 382 3752 492 3767
rect 1111 3782 1146 3787
rect 1111 3762 1118 3782
rect 1138 3762 1146 3782
rect 1656 3781 1698 3791
rect 1111 3754 1146 3762
rect 667 3689 699 3696
rect 667 3669 674 3689
rect 695 3669 699 3689
rect 667 3604 699 3669
rect 1037 3604 1077 3605
rect 667 3602 1079 3604
rect 667 3576 1047 3602
rect 1073 3576 1079 3602
rect 667 3568 1079 3576
rect 667 3540 699 3568
rect 1112 3548 1146 3754
rect 1320 3752 1431 3774
rect 1320 3732 1328 3752
rect 1347 3732 1405 3752
rect 1424 3732 1431 3752
rect 1320 3715 1431 3732
rect 1656 3759 1663 3781
rect 1689 3759 1698 3781
rect 1656 3750 1698 3759
rect 873 3545 916 3547
rect 667 3520 672 3540
rect 693 3520 699 3540
rect 667 3513 699 3520
rect 872 3538 916 3545
rect 872 3518 882 3538
rect 905 3518 916 3538
rect 872 3514 916 3518
rect 1090 3543 1146 3548
rect 1090 3523 1097 3543
rect 1117 3523 1146 3543
rect 1090 3516 1146 3523
rect 1202 3684 1235 3685
rect 1656 3684 1693 3750
rect 1202 3655 1693 3684
rect 1090 3515 1125 3516
rect 381 3442 492 3464
rect 381 3422 389 3442
rect 408 3422 466 3442
rect 485 3422 492 3442
rect 381 3405 492 3422
rect 872 3433 914 3514
rect 1202 3435 1235 3655
rect 1656 3653 1693 3655
rect 1462 3515 1572 3529
rect 1462 3512 1540 3515
rect 1462 3485 1466 3512
rect 1495 3488 1540 3512
rect 1569 3488 1572 3515
rect 1495 3485 1572 3488
rect 1462 3470 1572 3485
rect 1816 3496 1854 3834
rect 2029 3853 2085 3858
rect 2029 3833 2036 3853
rect 2056 3833 2085 3853
rect 2029 3826 2085 3833
rect 2029 3825 2064 3826
rect 2194 3505 2226 3506
rect 1816 3479 1824 3496
rect 1844 3479 1854 3496
rect 1816 3473 1854 3479
rect 2191 3500 2226 3505
rect 2191 3480 2198 3500
rect 2218 3480 2226 3500
rect 2191 3472 2226 3480
rect 1174 3433 1235 3435
rect 872 3404 1235 3433
rect 1747 3407 1779 3414
rect 872 3402 1174 3404
rect 1747 3387 1754 3407
rect 1775 3387 1779 3407
rect 1747 3322 1779 3387
rect 2117 3322 2157 3323
rect 1747 3320 2159 3322
rect 1115 3316 1150 3318
rect 151 3313 1150 3316
rect 150 3289 1150 3313
rect 150 3134 198 3289
rect 384 3248 494 3262
rect 384 3245 462 3248
rect 384 3218 388 3245
rect 417 3221 462 3245
rect 491 3221 494 3248
rect 1115 3238 1150 3289
rect 417 3218 494 3221
rect 384 3203 494 3218
rect 1113 3233 1150 3238
rect 1113 3213 1120 3233
rect 1140 3213 1150 3233
rect 1747 3294 2127 3320
rect 2153 3294 2159 3320
rect 1747 3286 2159 3294
rect 1747 3258 1779 3286
rect 1747 3238 1752 3258
rect 1773 3238 1779 3258
rect 1747 3231 1779 3238
rect 1953 3257 1995 3268
rect 2192 3266 2226 3472
rect 1953 3236 1960 3257
rect 1987 3236 1995 3257
rect 1113 3206 1150 3213
rect 1113 3205 1148 3206
rect 150 3105 158 3134
rect 187 3105 198 3134
rect 150 3100 198 3105
rect 669 3140 701 3147
rect 669 3120 676 3140
rect 697 3120 701 3140
rect 669 3055 701 3120
rect 1039 3055 1079 3056
rect 669 3053 1081 3055
rect 669 3027 1049 3053
rect 1075 3027 1081 3053
rect 669 3019 1081 3027
rect 669 2991 701 3019
rect 1114 2999 1148 3205
rect 1818 3188 1857 3195
rect 1461 3160 1572 3182
rect 1461 3140 1469 3160
rect 1488 3140 1546 3160
rect 1565 3140 1572 3160
rect 1461 3123 1572 3140
rect 1818 3161 1822 3188
rect 1853 3161 1857 3188
rect 1665 3072 1718 3076
rect 1183 3037 1718 3072
rect 669 2971 674 2991
rect 695 2971 701 2991
rect 669 2964 701 2971
rect 876 2991 915 2997
rect 876 2971 884 2991
rect 909 2971 915 2991
rect 876 2964 915 2971
rect 1092 2994 1148 2999
rect 1092 2974 1099 2994
rect 1119 2974 1148 2994
rect 1092 2967 1148 2974
rect 1092 2966 1127 2967
rect 884 2918 915 2964
rect 383 2893 494 2915
rect 383 2873 391 2893
rect 410 2873 468 2893
rect 487 2873 494 2893
rect 883 2901 915 2918
rect 1184 2901 1221 3037
rect 1322 3004 1432 3018
rect 1322 3001 1400 3004
rect 1322 2974 1326 3001
rect 1355 2977 1400 3001
rect 1429 2977 1432 3004
rect 1355 2974 1432 2977
rect 1322 2959 1432 2974
rect 1664 2990 1718 3037
rect 1664 2982 1717 2990
rect 1664 2965 1673 2982
rect 1705 2965 1717 2982
rect 1664 2962 1717 2965
rect 883 2888 1221 2901
rect 383 2856 494 2873
rect 884 2869 1221 2888
rect 1163 2868 1221 2869
rect 1607 2896 1639 2903
rect 1607 2876 1614 2896
rect 1635 2876 1639 2896
rect 1607 2811 1639 2876
rect 1818 2888 1857 3161
rect 1953 3065 1995 3236
rect 2170 3261 2226 3266
rect 2170 3241 2177 3261
rect 2197 3241 2226 3261
rect 2170 3234 2226 3241
rect 2170 3233 2205 3234
rect 1953 3031 2197 3065
rect 2160 3023 2197 3031
rect 2053 2990 2087 3001
rect 2051 2989 2087 2990
rect 2051 2969 2058 2989
rect 2078 2969 2087 2989
rect 2051 2961 2087 2969
rect 1818 2847 1825 2888
rect 1846 2847 1857 2888
rect 1818 2832 1857 2847
rect 1977 2811 2017 2812
rect 1607 2809 2019 2811
rect 1607 2783 1987 2809
rect 2013 2783 2019 2809
rect 1607 2775 2019 2783
rect 153 2736 1149 2762
rect 1607 2747 1639 2775
rect 2052 2755 2086 2961
rect 155 2683 197 2736
rect 155 2664 164 2683
rect 189 2664 197 2683
rect 155 2654 197 2664
rect 383 2694 493 2708
rect 383 2691 461 2694
rect 383 2664 387 2691
rect 416 2667 461 2691
rect 490 2667 493 2694
rect 1113 2684 1147 2736
rect 1607 2727 1612 2747
rect 1633 2727 1639 2747
rect 1607 2720 1639 2727
rect 2030 2750 2086 2755
rect 2030 2730 2037 2750
rect 2057 2730 2086 2750
rect 2030 2723 2086 2730
rect 2030 2722 2065 2723
rect 1658 2688 1699 2689
rect 416 2664 493 2667
rect 383 2649 493 2664
rect 1112 2679 1147 2684
rect 1112 2659 1119 2679
rect 1139 2659 1147 2679
rect 1657 2678 1699 2688
rect 1112 2651 1147 2659
rect 668 2586 700 2593
rect 668 2566 675 2586
rect 696 2566 700 2586
rect 668 2501 700 2566
rect 1038 2501 1078 2502
rect 668 2499 1080 2501
rect 668 2473 1048 2499
rect 1074 2473 1080 2499
rect 668 2465 1080 2473
rect 668 2437 700 2465
rect 1113 2445 1147 2651
rect 1321 2649 1432 2671
rect 1321 2629 1329 2649
rect 1348 2629 1406 2649
rect 1425 2629 1432 2649
rect 1321 2612 1432 2629
rect 1657 2656 1664 2678
rect 1690 2656 1699 2678
rect 1657 2647 1699 2656
rect 874 2442 917 2444
rect 668 2417 673 2437
rect 694 2417 700 2437
rect 668 2410 700 2417
rect 873 2435 917 2442
rect 873 2415 883 2435
rect 906 2415 917 2435
rect 873 2411 917 2415
rect 1091 2440 1147 2445
rect 1091 2420 1098 2440
rect 1118 2420 1147 2440
rect 1091 2413 1147 2420
rect 1203 2581 1236 2582
rect 1657 2581 1694 2647
rect 1203 2552 1694 2581
rect 1091 2412 1126 2413
rect 382 2339 493 2361
rect 382 2319 390 2339
rect 409 2319 467 2339
rect 486 2319 493 2339
rect 382 2303 493 2319
rect 873 2330 915 2411
rect 1203 2332 1236 2552
rect 1657 2550 1694 2552
rect 1432 2425 1542 2439
rect 1432 2422 1510 2425
rect 1432 2395 1436 2422
rect 1465 2398 1510 2422
rect 1539 2398 1542 2425
rect 1465 2395 1542 2398
rect 1432 2380 1542 2395
rect 2160 2410 2198 3023
rect 2160 2390 2168 2410
rect 2188 2390 2198 2410
rect 2160 2383 2198 2390
rect 2161 2382 2196 2383
rect 1175 2330 1236 2332
rect 873 2301 1236 2330
rect 1717 2317 1749 2324
rect 873 2299 1175 2301
rect 1717 2297 1724 2317
rect 1745 2297 1749 2317
rect 1717 2232 1749 2297
rect 2087 2232 2127 2233
rect 1717 2230 2129 2232
rect 1115 2213 1150 2215
rect 151 2210 1150 2213
rect 150 2186 1150 2210
rect 150 2031 198 2186
rect 384 2145 494 2159
rect 384 2142 462 2145
rect 384 2115 388 2142
rect 417 2118 462 2142
rect 491 2118 494 2145
rect 1115 2135 1150 2186
rect 1717 2204 2097 2230
rect 2123 2204 2129 2230
rect 1717 2196 2129 2204
rect 1717 2168 1749 2196
rect 1717 2148 1722 2168
rect 1743 2148 1749 2168
rect 1717 2141 1749 2148
rect 1923 2167 1968 2179
rect 2162 2176 2196 2382
rect 1923 2148 1930 2167
rect 1959 2148 1968 2167
rect 417 2115 494 2118
rect 384 2100 494 2115
rect 1113 2130 1150 2135
rect 1113 2110 1120 2130
rect 1140 2110 1150 2130
rect 1113 2103 1150 2110
rect 1113 2102 1148 2103
rect 150 2002 158 2031
rect 187 2002 198 2031
rect 150 1997 198 2002
rect 669 2037 701 2044
rect 669 2017 676 2037
rect 697 2017 701 2037
rect 669 1952 701 2017
rect 1039 1952 1079 1953
rect 669 1950 1081 1952
rect 669 1924 1049 1950
rect 1075 1924 1081 1950
rect 669 1916 1081 1924
rect 669 1888 701 1916
rect 1114 1896 1148 2102
rect 1431 2070 1542 2092
rect 1431 2050 1439 2070
rect 1458 2050 1516 2070
rect 1535 2050 1542 2070
rect 1431 2033 1542 2050
rect 1923 2065 1968 2148
rect 2140 2171 2196 2176
rect 2140 2151 2147 2171
rect 2167 2151 2196 2171
rect 2140 2144 2196 2151
rect 2140 2143 2175 2144
rect 2288 2065 2338 2067
rect 1923 2031 2338 2065
rect 2052 1969 2086 1970
rect 1183 1934 2087 1969
rect 2135 1958 2203 1969
rect 2135 1937 2140 1958
rect 669 1868 674 1888
rect 695 1868 701 1888
rect 669 1861 701 1868
rect 876 1888 915 1894
rect 876 1868 884 1888
rect 909 1868 915 1888
rect 876 1861 915 1868
rect 1092 1891 1148 1896
rect 1092 1871 1099 1891
rect 1119 1871 1148 1891
rect 1092 1864 1148 1871
rect 1092 1863 1127 1864
rect 884 1815 915 1861
rect 383 1790 494 1812
rect 383 1770 391 1790
rect 410 1770 468 1790
rect 487 1770 494 1790
rect 883 1798 915 1815
rect 1184 1798 1221 1934
rect 1322 1901 1432 1915
rect 1322 1898 1400 1901
rect 1322 1871 1326 1898
rect 1355 1874 1400 1898
rect 1429 1874 1432 1901
rect 2052 1891 2086 1934
rect 1355 1871 1432 1874
rect 1322 1856 1432 1871
rect 2051 1886 2086 1891
rect 2051 1866 2058 1886
rect 2078 1866 2086 1886
rect 2051 1858 2086 1866
rect 883 1785 1221 1798
rect 383 1753 494 1770
rect 884 1766 1221 1785
rect 1163 1765 1221 1766
rect 1607 1793 1639 1800
rect 1607 1773 1614 1793
rect 1635 1773 1639 1793
rect 1607 1708 1639 1773
rect 1977 1708 2017 1709
rect 1607 1706 2019 1708
rect 1607 1680 1987 1706
rect 2013 1680 2019 1706
rect 1607 1672 2019 1680
rect 153 1633 1149 1659
rect 1607 1644 1639 1672
rect 155 1580 197 1633
rect 155 1561 164 1580
rect 189 1561 197 1580
rect 155 1551 197 1561
rect 383 1591 493 1605
rect 383 1588 461 1591
rect 383 1561 387 1588
rect 416 1564 461 1588
rect 490 1564 493 1591
rect 1113 1581 1147 1633
rect 1607 1624 1612 1644
rect 1633 1624 1639 1644
rect 1607 1617 1639 1624
rect 1817 1645 1855 1655
rect 2052 1652 2086 1858
rect 1817 1628 1827 1645
rect 1847 1628 1855 1645
rect 1658 1585 1699 1586
rect 416 1561 493 1564
rect 383 1546 493 1561
rect 1112 1576 1147 1581
rect 1112 1556 1119 1576
rect 1139 1556 1147 1576
rect 1657 1575 1699 1585
rect 1112 1548 1147 1556
rect 668 1483 700 1490
rect 668 1463 675 1483
rect 696 1463 700 1483
rect 668 1398 700 1463
rect 1038 1398 1078 1399
rect 668 1396 1080 1398
rect 668 1370 1048 1396
rect 1074 1370 1080 1396
rect 668 1362 1080 1370
rect 668 1334 700 1362
rect 1113 1342 1147 1548
rect 1321 1546 1432 1568
rect 1321 1526 1329 1546
rect 1348 1526 1406 1546
rect 1425 1526 1432 1546
rect 1321 1509 1432 1526
rect 1657 1553 1664 1575
rect 1690 1553 1699 1575
rect 1657 1544 1699 1553
rect 874 1339 917 1341
rect 668 1314 673 1334
rect 694 1314 700 1334
rect 668 1307 700 1314
rect 873 1332 917 1339
rect 873 1312 883 1332
rect 906 1312 917 1332
rect 873 1308 917 1312
rect 1091 1337 1147 1342
rect 1091 1317 1098 1337
rect 1118 1317 1147 1337
rect 1091 1310 1147 1317
rect 1203 1478 1236 1479
rect 1657 1478 1694 1544
rect 1203 1449 1694 1478
rect 1091 1309 1126 1310
rect 382 1236 493 1258
rect 382 1216 390 1236
rect 409 1216 467 1236
rect 486 1216 493 1236
rect 382 1199 493 1216
rect 873 1227 915 1308
rect 1203 1229 1236 1449
rect 1657 1447 1694 1449
rect 1463 1309 1573 1323
rect 1463 1306 1541 1309
rect 1463 1279 1467 1306
rect 1496 1282 1541 1306
rect 1570 1282 1573 1309
rect 1496 1279 1573 1282
rect 1463 1264 1573 1279
rect 1817 1290 1855 1628
rect 2030 1647 2086 1652
rect 2030 1627 2037 1647
rect 2057 1627 2086 1647
rect 2030 1620 2086 1627
rect 2133 1929 2140 1937
rect 2188 1929 2203 1958
rect 2133 1920 2203 1929
rect 2030 1619 2065 1620
rect 1952 1519 1996 1523
rect 2133 1519 2183 1920
rect 2288 1903 2338 2031
rect 1952 1486 2183 1519
rect 1952 1484 2159 1486
rect 1952 1330 1996 1484
rect 1817 1273 1825 1290
rect 1845 1273 1855 1290
rect 1817 1267 1855 1273
rect 1175 1227 1236 1229
rect 873 1198 1236 1227
rect 1748 1201 1780 1208
rect 873 1196 1175 1198
rect 1748 1181 1755 1201
rect 1776 1181 1780 1201
rect 1748 1116 1780 1181
rect 1958 1194 1996 1330
rect 2195 1299 2226 1300
rect 2192 1294 2226 1299
rect 2192 1274 2199 1294
rect 2219 1274 2226 1294
rect 2192 1266 2226 1274
rect 1958 1156 1964 1194
rect 1987 1156 1996 1194
rect 1958 1146 1996 1156
rect 2193 1208 2226 1266
rect 2118 1116 2158 1117
rect 1748 1114 2160 1116
rect 1116 1110 1151 1112
rect 152 1107 1151 1110
rect 151 1083 1151 1107
rect 151 928 199 1083
rect 385 1042 495 1056
rect 385 1039 463 1042
rect 385 1012 389 1039
rect 418 1015 463 1039
rect 492 1015 495 1042
rect 1116 1032 1151 1083
rect 418 1012 495 1015
rect 385 997 495 1012
rect 1114 1027 1151 1032
rect 1114 1007 1121 1027
rect 1141 1007 1151 1027
rect 1748 1088 2128 1114
rect 2154 1088 2160 1114
rect 1748 1080 2160 1088
rect 1748 1052 1780 1080
rect 2193 1060 2229 1208
rect 1748 1032 1753 1052
rect 1774 1032 1780 1052
rect 1748 1025 1780 1032
rect 2171 1055 2229 1060
rect 2171 1035 2178 1055
rect 2198 1035 2229 1055
rect 2171 1028 2229 1035
rect 2171 1027 2206 1028
rect 1114 1000 1151 1007
rect 1114 999 1149 1000
rect 151 899 159 928
rect 188 899 199 928
rect 151 894 199 899
rect 670 934 702 941
rect 670 914 677 934
rect 698 914 702 934
rect 670 849 702 914
rect 1040 849 1080 850
rect 670 847 1082 849
rect 670 821 1050 847
rect 1076 821 1082 847
rect 670 813 1082 821
rect 670 785 702 813
rect 1115 793 1149 999
rect 1819 982 1858 989
rect 1462 954 1573 976
rect 1462 934 1470 954
rect 1489 934 1547 954
rect 1566 934 1573 954
rect 1462 917 1573 934
rect 1819 955 1823 982
rect 1854 955 1858 982
rect 1666 866 1719 870
rect 1184 831 1719 866
rect 670 765 675 785
rect 696 765 702 785
rect 670 758 702 765
rect 877 785 916 791
rect 877 765 885 785
rect 910 765 916 785
rect 877 758 916 765
rect 1093 788 1149 793
rect 1093 768 1100 788
rect 1120 768 1149 788
rect 1093 761 1149 768
rect 1093 760 1128 761
rect 885 712 916 758
rect 384 687 495 709
rect 384 667 392 687
rect 411 667 469 687
rect 488 667 495 687
rect 884 695 916 712
rect 1185 695 1222 831
rect 1323 798 1433 812
rect 1323 795 1401 798
rect 1323 768 1327 795
rect 1356 771 1401 795
rect 1430 771 1433 798
rect 1356 768 1433 771
rect 1323 753 1433 768
rect 1665 784 1719 831
rect 1665 776 1718 784
rect 1665 759 1674 776
rect 1706 759 1718 776
rect 1665 756 1718 759
rect 884 682 1222 695
rect 384 650 495 667
rect 885 663 1222 682
rect 1164 662 1222 663
rect 1608 690 1640 697
rect 1608 670 1615 690
rect 1636 670 1640 690
rect 1608 605 1640 670
rect 1819 682 1858 955
rect 2054 784 2088 795
rect 2052 783 2088 784
rect 2052 763 2059 783
rect 2079 763 2088 783
rect 2052 755 2088 763
rect 1819 641 1826 682
rect 1847 641 1858 682
rect 1819 626 1858 641
rect 1978 605 2018 606
rect 1608 603 2020 605
rect 1608 577 1988 603
rect 2014 577 2020 603
rect 1608 569 2020 577
rect 154 530 1150 556
rect 1608 541 1640 569
rect 2053 549 2087 755
rect 156 477 198 530
rect 156 458 165 477
rect 190 458 198 477
rect 156 448 198 458
rect 384 488 494 502
rect 384 485 462 488
rect 384 458 388 485
rect 417 461 462 485
rect 491 461 494 488
rect 1114 478 1148 530
rect 1608 521 1613 541
rect 1634 521 1640 541
rect 1608 514 1640 521
rect 2031 544 2087 549
rect 2031 524 2038 544
rect 2058 524 2087 544
rect 2031 517 2087 524
rect 2031 516 2066 517
rect 1659 482 1700 483
rect 417 458 494 461
rect 384 443 494 458
rect 1113 473 1148 478
rect 1113 453 1120 473
rect 1140 453 1148 473
rect 1658 472 1700 482
rect 1113 445 1148 453
rect 669 380 701 387
rect 669 360 676 380
rect 697 360 701 380
rect 669 295 701 360
rect 1039 295 1079 296
rect 669 293 1081 295
rect 669 267 1049 293
rect 1075 267 1081 293
rect 669 259 1081 267
rect 669 231 701 259
rect 1114 239 1148 445
rect 1322 443 1433 465
rect 1322 423 1330 443
rect 1349 423 1407 443
rect 1426 423 1433 443
rect 1322 406 1433 423
rect 1658 450 1665 472
rect 1691 450 1700 472
rect 1658 441 1700 450
rect 875 236 918 238
rect 669 211 674 231
rect 695 211 701 231
rect 669 204 701 211
rect 874 229 918 236
rect 874 209 884 229
rect 907 209 918 229
rect 874 205 918 209
rect 1092 234 1148 239
rect 1092 214 1099 234
rect 1119 214 1148 234
rect 1092 207 1148 214
rect 1204 375 1237 376
rect 1658 375 1695 441
rect 2290 418 2336 1903
rect 1204 346 1695 375
rect 1092 206 1127 207
rect 383 133 494 155
rect 383 113 391 133
rect 410 113 468 133
rect 487 113 494 133
rect 383 96 494 113
rect 874 124 916 205
rect 1204 126 1237 346
rect 1658 344 1695 346
rect 2288 394 2336 418
rect 1432 225 1542 239
rect 1432 222 1510 225
rect 1432 195 1436 222
rect 1465 198 1510 222
rect 1539 198 1542 225
rect 2288 216 2335 394
rect 1465 195 1542 198
rect 1432 180 1542 195
rect 2157 210 2338 216
rect 2157 190 2168 210
rect 2188 190 2338 210
rect 2157 184 2338 190
rect 2161 182 2196 184
rect 1176 124 1237 126
rect 874 95 1237 124
rect 1717 117 1749 124
rect 1717 97 1724 117
rect 1745 97 1749 117
rect 874 93 1176 95
rect 1717 32 1749 97
rect 2087 32 2127 33
rect 1717 30 2129 32
rect 1116 7 1151 9
rect 152 4 1151 7
rect 151 -20 1151 4
rect 151 -175 199 -20
rect 385 -61 495 -47
rect 385 -64 463 -61
rect 385 -91 389 -64
rect 418 -88 463 -64
rect 492 -88 495 -61
rect 1116 -71 1151 -20
rect 1717 4 2097 30
rect 2123 4 2129 30
rect 1717 -4 2129 4
rect 1717 -32 1749 -4
rect 2162 -24 2196 182
rect 1717 -52 1722 -32
rect 1743 -52 1749 -32
rect 1717 -59 1749 -52
rect 2140 -29 2196 -24
rect 2140 -49 2147 -29
rect 2167 -49 2196 -29
rect 2140 -56 2196 -49
rect 2140 -57 2175 -56
rect 418 -91 495 -88
rect 385 -106 495 -91
rect 1114 -76 1151 -71
rect 1114 -96 1121 -76
rect 1141 -96 1151 -76
rect 1114 -103 1151 -96
rect 1114 -104 1149 -103
rect 151 -204 159 -175
rect 188 -204 199 -175
rect 151 -209 199 -204
rect 670 -169 702 -162
rect 670 -189 677 -169
rect 698 -189 702 -169
rect 670 -254 702 -189
rect 1040 -254 1080 -253
rect 670 -256 1082 -254
rect 670 -282 1050 -256
rect 1076 -282 1082 -256
rect 670 -290 1082 -282
rect 670 -318 702 -290
rect 1115 -310 1149 -104
rect 1431 -130 1542 -108
rect 1431 -150 1439 -130
rect 1458 -150 1516 -130
rect 1535 -150 1542 -130
rect 1431 -167 1542 -150
rect 2053 -237 2087 -236
rect 1184 -272 2088 -237
rect 2296 -247 2343 -229
rect 670 -338 675 -318
rect 696 -338 702 -318
rect 670 -345 702 -338
rect 877 -318 916 -312
rect 877 -338 885 -318
rect 910 -338 916 -318
rect 877 -345 916 -338
rect 1093 -315 1149 -310
rect 1093 -335 1100 -315
rect 1120 -335 1149 -315
rect 1093 -342 1149 -335
rect 1093 -343 1128 -342
rect 885 -391 916 -345
rect 384 -416 495 -394
rect 384 -436 392 -416
rect 411 -436 469 -416
rect 488 -436 495 -416
rect 884 -408 916 -391
rect 1185 -408 1222 -272
rect 1323 -305 1433 -291
rect 1323 -308 1401 -305
rect 1323 -335 1327 -308
rect 1356 -332 1401 -308
rect 1430 -332 1433 -305
rect 2053 -315 2087 -272
rect 1356 -335 1433 -332
rect 1323 -350 1433 -335
rect 2052 -320 2087 -315
rect 2052 -340 2059 -320
rect 2079 -340 2087 -320
rect 2052 -348 2087 -340
rect 884 -421 1222 -408
rect 384 -453 495 -436
rect 885 -440 1222 -421
rect 1164 -441 1222 -440
rect 1608 -413 1640 -406
rect 1608 -433 1615 -413
rect 1636 -433 1640 -413
rect 1608 -498 1640 -433
rect 1978 -498 2018 -497
rect 1608 -500 2020 -498
rect 1608 -526 1988 -500
rect 2014 -526 2020 -500
rect 1608 -534 2020 -526
rect 154 -573 1150 -547
rect 1608 -562 1640 -534
rect 156 -626 198 -573
rect 156 -645 165 -626
rect 190 -645 198 -626
rect 156 -655 198 -645
rect 384 -615 494 -601
rect 384 -618 462 -615
rect 384 -645 388 -618
rect 417 -642 462 -618
rect 491 -642 494 -615
rect 1114 -625 1148 -573
rect 1608 -582 1613 -562
rect 1634 -582 1640 -562
rect 1608 -589 1640 -582
rect 1818 -561 1856 -551
rect 2053 -554 2087 -348
rect 1818 -578 1828 -561
rect 1848 -578 1856 -561
rect 1659 -621 1700 -620
rect 417 -645 494 -642
rect 384 -660 494 -645
rect 1113 -630 1148 -625
rect 1113 -650 1120 -630
rect 1140 -650 1148 -630
rect 1658 -631 1700 -621
rect 1113 -658 1148 -650
rect 669 -723 701 -716
rect 669 -743 676 -723
rect 697 -743 701 -723
rect 669 -808 701 -743
rect 1039 -808 1079 -807
rect 669 -810 1081 -808
rect 669 -836 1049 -810
rect 1075 -836 1081 -810
rect 669 -844 1081 -836
rect 669 -872 701 -844
rect 1114 -864 1148 -658
rect 1322 -660 1433 -638
rect 1322 -680 1330 -660
rect 1349 -680 1407 -660
rect 1426 -680 1433 -660
rect 1322 -697 1433 -680
rect 1658 -653 1665 -631
rect 1691 -653 1700 -631
rect 1658 -662 1700 -653
rect 875 -867 918 -865
rect 669 -892 674 -872
rect 695 -892 701 -872
rect 669 -899 701 -892
rect 874 -874 918 -867
rect 874 -894 884 -874
rect 907 -894 918 -874
rect 874 -898 918 -894
rect 1092 -869 1148 -864
rect 1092 -889 1099 -869
rect 1119 -889 1148 -869
rect 1092 -896 1148 -889
rect 1204 -728 1237 -727
rect 1658 -728 1695 -662
rect 1204 -757 1695 -728
rect 1092 -897 1127 -896
rect 383 -970 494 -948
rect 383 -990 391 -970
rect 410 -990 468 -970
rect 487 -990 494 -970
rect 383 -1007 494 -990
rect 874 -979 916 -898
rect 1204 -977 1237 -757
rect 1658 -759 1695 -757
rect 1464 -897 1574 -883
rect 1464 -900 1542 -897
rect 1464 -927 1468 -900
rect 1497 -924 1542 -900
rect 1571 -924 1574 -897
rect 1497 -927 1574 -924
rect 1464 -942 1574 -927
rect 1818 -916 1856 -578
rect 2031 -559 2087 -554
rect 2031 -579 2038 -559
rect 2058 -579 2087 -559
rect 2031 -586 2087 -579
rect 2296 -287 2303 -247
rect 2330 -287 2343 -247
rect 2031 -587 2066 -586
rect 2196 -907 2228 -906
rect 1818 -933 1826 -916
rect 1846 -933 1856 -916
rect 1818 -939 1856 -933
rect 2193 -912 2228 -907
rect 2193 -932 2200 -912
rect 2220 -932 2228 -912
rect 2193 -940 2228 -932
rect 1176 -979 1237 -977
rect 874 -1008 1237 -979
rect 1749 -1005 1781 -998
rect 874 -1010 1176 -1008
rect 1749 -1025 1756 -1005
rect 1777 -1025 1781 -1005
rect 1749 -1090 1781 -1025
rect 2119 -1090 2159 -1089
rect 1749 -1092 2161 -1090
rect 1117 -1096 1152 -1094
rect 153 -1099 1152 -1096
rect 152 -1123 1152 -1099
rect 152 -1278 200 -1123
rect 386 -1164 496 -1150
rect 386 -1167 464 -1164
rect 386 -1194 390 -1167
rect 419 -1191 464 -1167
rect 493 -1191 496 -1164
rect 1117 -1174 1152 -1123
rect 419 -1194 496 -1191
rect 386 -1209 496 -1194
rect 1115 -1179 1152 -1174
rect 1115 -1199 1122 -1179
rect 1142 -1199 1152 -1179
rect 1749 -1118 2129 -1092
rect 2155 -1118 2161 -1092
rect 1749 -1126 2161 -1118
rect 1749 -1154 1781 -1126
rect 1749 -1174 1754 -1154
rect 1775 -1174 1781 -1154
rect 1749 -1181 1781 -1174
rect 1955 -1155 1997 -1144
rect 2194 -1146 2228 -940
rect 1955 -1176 1962 -1155
rect 1989 -1176 1997 -1155
rect 1115 -1206 1152 -1199
rect 1115 -1207 1150 -1206
rect 152 -1307 160 -1278
rect 189 -1307 200 -1278
rect 152 -1312 200 -1307
rect 671 -1272 703 -1265
rect 671 -1292 678 -1272
rect 699 -1292 703 -1272
rect 671 -1357 703 -1292
rect 1041 -1357 1081 -1356
rect 671 -1359 1083 -1357
rect 671 -1385 1051 -1359
rect 1077 -1385 1083 -1359
rect 671 -1393 1083 -1385
rect 671 -1421 703 -1393
rect 1116 -1413 1150 -1207
rect 1820 -1224 1859 -1217
rect 1463 -1252 1574 -1230
rect 1463 -1272 1471 -1252
rect 1490 -1272 1548 -1252
rect 1567 -1272 1574 -1252
rect 1463 -1289 1574 -1272
rect 1820 -1251 1824 -1224
rect 1855 -1251 1859 -1224
rect 1667 -1340 1720 -1336
rect 1185 -1375 1720 -1340
rect 671 -1441 676 -1421
rect 697 -1441 703 -1421
rect 671 -1448 703 -1441
rect 878 -1421 917 -1415
rect 878 -1441 886 -1421
rect 911 -1441 917 -1421
rect 878 -1448 917 -1441
rect 1094 -1418 1150 -1413
rect 1094 -1438 1101 -1418
rect 1121 -1438 1150 -1418
rect 1094 -1445 1150 -1438
rect 1094 -1446 1129 -1445
rect 886 -1494 917 -1448
rect 385 -1519 496 -1497
rect 385 -1539 393 -1519
rect 412 -1539 470 -1519
rect 489 -1539 496 -1519
rect 885 -1511 917 -1494
rect 1186 -1511 1223 -1375
rect 1324 -1408 1434 -1394
rect 1324 -1411 1402 -1408
rect 1324 -1438 1328 -1411
rect 1357 -1435 1402 -1411
rect 1431 -1435 1434 -1408
rect 1357 -1438 1434 -1435
rect 1324 -1453 1434 -1438
rect 1666 -1422 1720 -1375
rect 1666 -1430 1719 -1422
rect 1666 -1447 1675 -1430
rect 1707 -1447 1719 -1430
rect 1666 -1450 1719 -1447
rect 885 -1524 1223 -1511
rect 385 -1556 496 -1539
rect 886 -1543 1223 -1524
rect 1165 -1544 1223 -1543
rect 1609 -1516 1641 -1509
rect 1609 -1536 1616 -1516
rect 1637 -1536 1641 -1516
rect 1609 -1601 1641 -1536
rect 1820 -1524 1859 -1251
rect 1955 -1347 1997 -1176
rect 2172 -1151 2228 -1146
rect 2172 -1171 2179 -1151
rect 2199 -1171 2228 -1151
rect 2172 -1178 2228 -1171
rect 2172 -1179 2207 -1178
rect 1955 -1381 2199 -1347
rect 2162 -1389 2199 -1381
rect 2055 -1422 2089 -1411
rect 2053 -1423 2089 -1422
rect 2053 -1443 2060 -1423
rect 2080 -1443 2089 -1423
rect 2053 -1451 2089 -1443
rect 1820 -1565 1827 -1524
rect 1848 -1565 1859 -1524
rect 1820 -1580 1859 -1565
rect 1979 -1601 2019 -1600
rect 1609 -1603 2021 -1601
rect 1609 -1629 1989 -1603
rect 2015 -1629 2021 -1603
rect 1609 -1637 2021 -1629
rect 155 -1676 1151 -1650
rect 1609 -1665 1641 -1637
rect 2054 -1657 2088 -1451
rect 157 -1729 199 -1676
rect 157 -1748 166 -1729
rect 191 -1748 199 -1729
rect 157 -1758 199 -1748
rect 385 -1718 495 -1704
rect 385 -1721 463 -1718
rect 385 -1748 389 -1721
rect 418 -1745 463 -1721
rect 492 -1745 495 -1718
rect 1115 -1728 1149 -1676
rect 1609 -1685 1614 -1665
rect 1635 -1685 1641 -1665
rect 1609 -1692 1641 -1685
rect 2032 -1662 2088 -1657
rect 2032 -1682 2039 -1662
rect 2059 -1682 2088 -1662
rect 2032 -1689 2088 -1682
rect 2032 -1690 2067 -1689
rect 1660 -1724 1701 -1723
rect 418 -1748 495 -1745
rect 385 -1763 495 -1748
rect 1114 -1733 1149 -1728
rect 1114 -1753 1121 -1733
rect 1141 -1753 1149 -1733
rect 1659 -1734 1701 -1724
rect 1114 -1761 1149 -1753
rect 670 -1826 702 -1819
rect 670 -1846 677 -1826
rect 698 -1846 702 -1826
rect 670 -1911 702 -1846
rect 1040 -1911 1080 -1910
rect 670 -1913 1082 -1911
rect 670 -1939 1050 -1913
rect 1076 -1939 1082 -1913
rect 670 -1947 1082 -1939
rect 670 -1975 702 -1947
rect 1115 -1967 1149 -1761
rect 1323 -1763 1434 -1741
rect 1323 -1783 1331 -1763
rect 1350 -1783 1408 -1763
rect 1427 -1783 1434 -1763
rect 1323 -1800 1434 -1783
rect 1659 -1756 1666 -1734
rect 1692 -1756 1701 -1734
rect 1659 -1765 1701 -1756
rect 876 -1970 919 -1968
rect 670 -1995 675 -1975
rect 696 -1995 702 -1975
rect 670 -2002 702 -1995
rect 875 -1977 919 -1970
rect 875 -1997 885 -1977
rect 908 -1997 919 -1977
rect 875 -2001 919 -1997
rect 1093 -1972 1149 -1967
rect 1093 -1992 1100 -1972
rect 1120 -1992 1149 -1972
rect 1093 -1999 1149 -1992
rect 1205 -1831 1238 -1830
rect 1659 -1831 1696 -1765
rect 2162 -1780 2200 -1389
rect 1776 -1796 2200 -1780
rect 1205 -1860 1696 -1831
rect 1093 -2000 1128 -1999
rect 384 -2073 495 -2051
rect 384 -2093 392 -2073
rect 411 -2093 469 -2073
rect 488 -2093 495 -2073
rect 384 -2109 495 -2093
rect 875 -2082 917 -2001
rect 1205 -2080 1238 -1860
rect 1659 -1862 1696 -1860
rect 1775 -1821 2200 -1796
rect 1434 -1987 1544 -1973
rect 1434 -1990 1512 -1987
rect 1434 -2017 1438 -1990
rect 1467 -2014 1512 -1990
rect 1541 -2014 1544 -1987
rect 1467 -2017 1544 -2014
rect 1434 -2032 1544 -2017
rect 1775 -2000 1809 -1821
rect 2296 -1864 2343 -287
rect 1775 -2020 1779 -2000
rect 1800 -2020 1809 -2000
rect 1775 -2026 1809 -2020
rect 1928 -1889 2257 -1886
rect 2296 -1889 2340 -1864
rect 1928 -1919 2340 -1889
rect 1177 -2082 1238 -2080
rect 875 -2111 1238 -2082
rect 1719 -2095 1751 -2088
rect 875 -2113 1177 -2111
rect 1719 -2115 1726 -2095
rect 1747 -2115 1751 -2095
rect 1719 -2180 1751 -2115
rect 1928 -2107 1963 -1919
rect 2230 -1921 2340 -1919
rect 2156 -2004 2206 -1997
rect 2156 -2018 2170 -2004
rect 2162 -2022 2170 -2018
rect 2190 -2018 2206 -2004
rect 2190 -2022 2200 -2018
rect 2162 -2029 2200 -2022
rect 2163 -2030 2198 -2029
rect 1928 -2139 1933 -2107
rect 1960 -2139 1963 -2107
rect 1928 -2157 1963 -2139
rect 2089 -2180 2129 -2179
rect 1719 -2182 2131 -2180
rect 1117 -2199 1152 -2197
rect 153 -2202 1152 -2199
rect 152 -2226 1152 -2202
rect 152 -2381 200 -2226
rect 386 -2267 496 -2253
rect 386 -2270 464 -2267
rect 386 -2297 390 -2270
rect 419 -2294 464 -2270
rect 493 -2294 496 -2267
rect 1117 -2277 1152 -2226
rect 1719 -2208 2099 -2182
rect 2125 -2208 2131 -2182
rect 1719 -2216 2131 -2208
rect 1719 -2244 1751 -2216
rect 2164 -2236 2198 -2030
rect 1719 -2264 1724 -2244
rect 1745 -2264 1751 -2244
rect 1719 -2271 1751 -2264
rect 2142 -2241 2198 -2236
rect 2142 -2261 2149 -2241
rect 2169 -2261 2198 -2241
rect 2142 -2268 2198 -2261
rect 2142 -2269 2177 -2268
rect 419 -2297 496 -2294
rect 386 -2312 496 -2297
rect 1115 -2282 1152 -2277
rect 1115 -2302 1122 -2282
rect 1142 -2302 1152 -2282
rect 1115 -2309 1152 -2302
rect 2137 -2307 2207 -2297
rect 1115 -2310 1150 -2309
rect 152 -2410 160 -2381
rect 189 -2410 200 -2381
rect 152 -2415 200 -2410
rect 671 -2375 703 -2368
rect 671 -2395 678 -2375
rect 699 -2395 703 -2375
rect 671 -2460 703 -2395
rect 1041 -2460 1081 -2459
rect 671 -2462 1083 -2460
rect 671 -2488 1051 -2462
rect 1077 -2488 1083 -2462
rect 671 -2496 1083 -2488
rect 671 -2524 703 -2496
rect 1116 -2516 1150 -2310
rect 2135 -2314 2207 -2307
rect 1433 -2342 1544 -2320
rect 1433 -2362 1441 -2342
rect 1460 -2362 1518 -2342
rect 1537 -2362 1544 -2342
rect 1433 -2379 1544 -2362
rect 2135 -2343 2142 -2314
rect 2190 -2343 2207 -2314
rect 2135 -2352 2207 -2343
rect 2054 -2443 2088 -2442
rect 1185 -2478 2089 -2443
rect 671 -2544 676 -2524
rect 697 -2544 703 -2524
rect 671 -2551 703 -2544
rect 878 -2524 917 -2518
rect 878 -2544 886 -2524
rect 911 -2544 917 -2524
rect 878 -2551 917 -2544
rect 1094 -2521 1150 -2516
rect 1094 -2541 1101 -2521
rect 1121 -2541 1150 -2521
rect 1094 -2548 1150 -2541
rect 1094 -2549 1129 -2548
rect 886 -2597 917 -2551
rect 385 -2622 496 -2600
rect 385 -2642 393 -2622
rect 412 -2642 470 -2622
rect 489 -2642 496 -2622
rect 885 -2614 917 -2597
rect 1186 -2614 1223 -2478
rect 1324 -2511 1434 -2497
rect 1324 -2514 1402 -2511
rect 1324 -2541 1328 -2514
rect 1357 -2538 1402 -2514
rect 1431 -2538 1434 -2511
rect 2054 -2521 2088 -2478
rect 1357 -2541 1434 -2538
rect 1324 -2556 1434 -2541
rect 2053 -2526 2088 -2521
rect 2053 -2546 2060 -2526
rect 2080 -2546 2088 -2526
rect 2053 -2554 2088 -2546
rect 885 -2627 1223 -2614
rect 385 -2659 496 -2642
rect 886 -2646 1223 -2627
rect 1165 -2647 1223 -2646
rect 1609 -2619 1641 -2612
rect 1609 -2639 1616 -2619
rect 1637 -2639 1641 -2619
rect 1609 -2704 1641 -2639
rect 1979 -2704 2019 -2703
rect 1609 -2706 2021 -2704
rect 1609 -2732 1989 -2706
rect 2015 -2732 2021 -2706
rect 1609 -2740 2021 -2732
rect 155 -2779 1151 -2753
rect 1609 -2768 1641 -2740
rect 157 -2832 199 -2779
rect 157 -2851 166 -2832
rect 191 -2851 199 -2832
rect 157 -2861 199 -2851
rect 385 -2821 495 -2807
rect 385 -2824 463 -2821
rect 385 -2851 389 -2824
rect 418 -2848 463 -2824
rect 492 -2848 495 -2821
rect 1115 -2831 1149 -2779
rect 1609 -2788 1614 -2768
rect 1635 -2788 1641 -2768
rect 1609 -2795 1641 -2788
rect 1819 -2767 1857 -2757
rect 2054 -2760 2088 -2554
rect 1819 -2784 1829 -2767
rect 1849 -2784 1857 -2767
rect 1660 -2827 1701 -2826
rect 418 -2851 495 -2848
rect 385 -2866 495 -2851
rect 1114 -2836 1149 -2831
rect 1114 -2856 1121 -2836
rect 1141 -2856 1149 -2836
rect 1659 -2837 1701 -2827
rect 1114 -2864 1149 -2856
rect 670 -2929 702 -2922
rect 670 -2949 677 -2929
rect 698 -2949 702 -2929
rect 670 -3014 702 -2949
rect 1040 -3014 1080 -3013
rect 670 -3016 1082 -3014
rect 670 -3042 1050 -3016
rect 1076 -3042 1082 -3016
rect 670 -3050 1082 -3042
rect 670 -3078 702 -3050
rect 1115 -3070 1149 -2864
rect 1323 -2866 1434 -2844
rect 1323 -2886 1331 -2866
rect 1350 -2886 1408 -2866
rect 1427 -2886 1434 -2866
rect 1323 -2903 1434 -2886
rect 1659 -2859 1666 -2837
rect 1692 -2859 1701 -2837
rect 1659 -2868 1701 -2859
rect 876 -3073 919 -3071
rect 670 -3098 675 -3078
rect 696 -3098 702 -3078
rect 670 -3105 702 -3098
rect 875 -3080 919 -3073
rect 875 -3100 885 -3080
rect 908 -3100 919 -3080
rect 875 -3104 919 -3100
rect 1093 -3075 1149 -3070
rect 1093 -3095 1100 -3075
rect 1120 -3095 1149 -3075
rect 1093 -3102 1149 -3095
rect 1205 -2934 1238 -2933
rect 1659 -2934 1696 -2868
rect 1205 -2963 1696 -2934
rect 1093 -3103 1128 -3102
rect 384 -3176 495 -3154
rect 384 -3196 392 -3176
rect 411 -3196 469 -3176
rect 488 -3196 495 -3176
rect 384 -3213 495 -3196
rect 875 -3185 917 -3104
rect 1205 -3183 1238 -2963
rect 1659 -2965 1696 -2963
rect 1465 -3103 1575 -3089
rect 1465 -3106 1543 -3103
rect 1465 -3133 1469 -3106
rect 1498 -3130 1543 -3106
rect 1572 -3130 1575 -3103
rect 1498 -3133 1575 -3130
rect 1465 -3148 1575 -3133
rect 1819 -3122 1857 -2784
rect 2032 -2765 2088 -2760
rect 2032 -2785 2039 -2765
rect 2059 -2785 2088 -2765
rect 2032 -2792 2088 -2785
rect 2032 -2793 2067 -2792
rect 1954 -2893 1998 -2889
rect 2135 -2893 2185 -2352
rect 1954 -2926 2185 -2893
rect 1954 -2928 2161 -2926
rect 1954 -3082 1998 -2928
rect 1819 -3139 1827 -3122
rect 1847 -3139 1857 -3122
rect 1819 -3145 1857 -3139
rect 1177 -3185 1238 -3183
rect 875 -3214 1238 -3185
rect 1750 -3211 1782 -3204
rect 875 -3216 1177 -3214
rect 1750 -3231 1757 -3211
rect 1778 -3231 1782 -3211
rect 1750 -3296 1782 -3231
rect 1960 -3218 1998 -3082
rect 2197 -3113 2228 -3112
rect 2194 -3118 2228 -3113
rect 2194 -3138 2201 -3118
rect 2221 -3138 2228 -3118
rect 2194 -3146 2228 -3138
rect 1960 -3256 1966 -3218
rect 1989 -3256 1998 -3218
rect 1960 -3266 1998 -3256
rect 2195 -3204 2228 -3146
rect 2120 -3296 2160 -3295
rect 1750 -3298 2162 -3296
rect 1118 -3302 1153 -3300
rect 154 -3305 1153 -3302
rect 153 -3329 1153 -3305
rect 153 -3484 201 -3329
rect 387 -3370 497 -3356
rect 387 -3373 465 -3370
rect 387 -3400 391 -3373
rect 420 -3397 465 -3373
rect 494 -3397 497 -3370
rect 1118 -3380 1153 -3329
rect 420 -3400 497 -3397
rect 387 -3415 497 -3400
rect 1116 -3385 1153 -3380
rect 1116 -3405 1123 -3385
rect 1143 -3405 1153 -3385
rect 1750 -3324 2130 -3298
rect 2156 -3324 2162 -3298
rect 1750 -3332 2162 -3324
rect 1750 -3360 1782 -3332
rect 2195 -3352 2231 -3204
rect 1750 -3380 1755 -3360
rect 1776 -3380 1782 -3360
rect 1750 -3387 1782 -3380
rect 2173 -3357 2231 -3352
rect 2173 -3377 2180 -3357
rect 2200 -3377 2231 -3357
rect 2173 -3384 2231 -3377
rect 2173 -3385 2208 -3384
rect 1116 -3412 1153 -3405
rect 1116 -3413 1151 -3412
rect 153 -3513 161 -3484
rect 190 -3513 201 -3484
rect 153 -3518 201 -3513
rect 672 -3478 704 -3471
rect 672 -3498 679 -3478
rect 700 -3498 704 -3478
rect 672 -3563 704 -3498
rect 1042 -3563 1082 -3562
rect 672 -3565 1084 -3563
rect 672 -3591 1052 -3565
rect 1078 -3591 1084 -3565
rect 672 -3599 1084 -3591
rect 672 -3627 704 -3599
rect 1117 -3619 1151 -3413
rect 1821 -3430 1860 -3423
rect 1464 -3458 1575 -3436
rect 1464 -3478 1472 -3458
rect 1491 -3478 1549 -3458
rect 1568 -3478 1575 -3458
rect 1464 -3495 1575 -3478
rect 1821 -3457 1825 -3430
rect 1856 -3457 1860 -3430
rect 1668 -3546 1721 -3542
rect 1186 -3581 1721 -3546
rect 672 -3647 677 -3627
rect 698 -3647 704 -3627
rect 672 -3654 704 -3647
rect 879 -3627 918 -3621
rect 879 -3647 887 -3627
rect 912 -3647 918 -3627
rect 879 -3654 918 -3647
rect 1095 -3624 1151 -3619
rect 1095 -3644 1102 -3624
rect 1122 -3644 1151 -3624
rect 1095 -3651 1151 -3644
rect 1095 -3652 1130 -3651
rect 887 -3700 918 -3654
rect 386 -3725 497 -3703
rect 386 -3745 394 -3725
rect 413 -3745 471 -3725
rect 490 -3745 497 -3725
rect 886 -3717 918 -3700
rect 1187 -3717 1224 -3581
rect 1325 -3614 1435 -3600
rect 1325 -3617 1403 -3614
rect 1325 -3644 1329 -3617
rect 1358 -3641 1403 -3617
rect 1432 -3641 1435 -3614
rect 1358 -3644 1435 -3641
rect 1325 -3659 1435 -3644
rect 1667 -3628 1721 -3581
rect 1667 -3636 1720 -3628
rect 1667 -3653 1676 -3636
rect 1708 -3653 1720 -3636
rect 1667 -3656 1720 -3653
rect 886 -3730 1224 -3717
rect 386 -3762 497 -3745
rect 887 -3749 1224 -3730
rect 1166 -3750 1224 -3749
rect 1610 -3722 1642 -3715
rect 1610 -3742 1617 -3722
rect 1638 -3742 1642 -3722
rect 1610 -3807 1642 -3742
rect 1821 -3730 1860 -3457
rect 2056 -3628 2090 -3617
rect 2054 -3629 2090 -3628
rect 2054 -3649 2061 -3629
rect 2081 -3649 2090 -3629
rect 2054 -3657 2090 -3649
rect 1821 -3771 1828 -3730
rect 1849 -3771 1860 -3730
rect 1821 -3786 1860 -3771
rect 1980 -3807 2020 -3806
rect 1610 -3809 2022 -3807
rect 1610 -3835 1990 -3809
rect 2016 -3835 2022 -3809
rect 1610 -3843 2022 -3835
rect 156 -3882 1152 -3856
rect 1610 -3871 1642 -3843
rect 2055 -3863 2089 -3657
rect 158 -3935 200 -3882
rect 158 -3954 167 -3935
rect 192 -3954 200 -3935
rect 158 -3964 200 -3954
rect 386 -3924 496 -3910
rect 386 -3927 464 -3924
rect 386 -3954 390 -3927
rect 419 -3951 464 -3927
rect 493 -3951 496 -3924
rect 1116 -3934 1150 -3882
rect 1610 -3891 1615 -3871
rect 1636 -3891 1642 -3871
rect 1610 -3898 1642 -3891
rect 2033 -3868 2089 -3863
rect 2033 -3888 2040 -3868
rect 2060 -3888 2089 -3868
rect 2033 -3895 2089 -3888
rect 2033 -3896 2068 -3895
rect 1661 -3930 1702 -3929
rect 419 -3954 496 -3951
rect 386 -3969 496 -3954
rect 1115 -3939 1150 -3934
rect 1115 -3959 1122 -3939
rect 1142 -3959 1150 -3939
rect 1660 -3940 1702 -3930
rect 1115 -3967 1150 -3959
rect 671 -4032 703 -4025
rect 671 -4052 678 -4032
rect 699 -4052 703 -4032
rect 671 -4117 703 -4052
rect 1041 -4117 1081 -4116
rect 671 -4119 1083 -4117
rect 671 -4145 1051 -4119
rect 1077 -4145 1083 -4119
rect 671 -4153 1083 -4145
rect 671 -4181 703 -4153
rect 1116 -4173 1150 -3967
rect 1324 -3969 1435 -3947
rect 1324 -3989 1332 -3969
rect 1351 -3989 1409 -3969
rect 1428 -3989 1435 -3969
rect 1324 -4006 1435 -3989
rect 1660 -3962 1667 -3940
rect 1693 -3962 1702 -3940
rect 1660 -3971 1702 -3962
rect 877 -4176 920 -4174
rect 671 -4201 676 -4181
rect 697 -4201 703 -4181
rect 671 -4208 703 -4201
rect 876 -4183 920 -4176
rect 876 -4203 886 -4183
rect 909 -4203 920 -4183
rect 876 -4207 920 -4203
rect 1094 -4178 1150 -4173
rect 1094 -4198 1101 -4178
rect 1121 -4198 1150 -4178
rect 1094 -4205 1150 -4198
rect 1206 -4037 1239 -4036
rect 1660 -4037 1697 -3971
rect 1206 -4066 1697 -4037
rect 1094 -4206 1129 -4205
rect 385 -4279 496 -4257
rect 385 -4299 393 -4279
rect 412 -4299 470 -4279
rect 489 -4299 496 -4279
rect 385 -4316 496 -4299
rect 876 -4288 918 -4207
rect 1206 -4286 1239 -4066
rect 1660 -4068 1697 -4066
rect 1178 -4288 1239 -4286
rect 876 -4317 1239 -4288
rect 876 -4319 1178 -4317
<< labels >>
rlabel locali 254 4132 276 4147 1 d0
rlabel metal1 423 4355 451 4360 1 vdd
rlabel metal1 420 3962 454 3968 1 gnd
rlabel locali 1191 3884 1219 3905 1 d1
rlabel metal1 1358 3718 1392 3724 1 gnd
rlabel metal1 1361 4111 1389 4116 1 vdd
rlabel locali 253 3578 275 3593 1 d0
rlabel metal1 422 3801 450 3806 1 vdd
rlabel metal1 419 3408 453 3414 1 gnd
rlabel locali 74 4417 102 4425 1 vref
rlabel locali 255 3029 277 3044 1 d0
rlabel metal1 424 3252 452 3257 1 vdd
rlabel metal1 421 2859 455 2865 1 gnd
rlabel locali 1192 2781 1220 2802 1 d1
rlabel metal1 1359 2615 1393 2621 1 gnd
rlabel metal1 1362 3008 1390 3013 1 vdd
rlabel locali 254 2475 276 2490 1 d0
rlabel metal1 423 2698 451 2703 1 vdd
rlabel metal1 420 2305 454 2311 1 gnd
rlabel metal1 1502 3519 1530 3524 1 vdd
rlabel metal1 1499 3126 1533 3132 1 gnd
rlabel locali 1330 3291 1351 3310 1 d2
rlabel locali 255 1926 277 1941 1 d0
rlabel metal1 424 2149 452 2154 1 vdd
rlabel metal1 421 1756 455 1762 1 gnd
rlabel locali 1192 1678 1220 1699 1 d1
rlabel metal1 1359 1512 1393 1518 1 gnd
rlabel metal1 1362 1905 1390 1910 1 vdd
rlabel locali 254 1372 276 1387 1 d0
rlabel metal1 423 1595 451 1600 1 vdd
rlabel metal1 420 1202 454 1208 1 gnd
rlabel locali 256 823 278 838 1 d0
rlabel metal1 425 1046 453 1051 1 vdd
rlabel metal1 422 653 456 659 1 gnd
rlabel locali 1193 575 1221 596 1 d1
rlabel metal1 1360 409 1394 415 1 gnd
rlabel metal1 1363 802 1391 807 1 vdd
rlabel locali 255 269 277 284 1 d0
rlabel metal1 424 492 452 497 1 vdd
rlabel metal1 421 99 455 105 1 gnd
rlabel metal1 1503 1313 1531 1318 1 vdd
rlabel metal1 1500 920 1534 926 1 gnd
rlabel locali 1331 1085 1352 1104 1 d2
rlabel metal1 1472 2429 1500 2434 1 vdd
rlabel metal1 1469 2036 1503 2042 1 gnd
rlabel locali 1302 2205 1328 2222 1 d3
rlabel locali 1304 -2207 1330 -2190 1 d3
rlabel metal1 1471 -2376 1505 -2370 1 gnd
rlabel metal1 1474 -1983 1502 -1978 1 vdd
rlabel locali 1333 -3327 1354 -3308 1 d2
rlabel metal1 1502 -3492 1536 -3486 1 gnd
rlabel metal1 1505 -3099 1533 -3094 1 vdd
rlabel metal1 423 -4313 457 -4307 1 gnd
rlabel metal1 426 -3920 454 -3915 1 vdd
rlabel locali 257 -4143 279 -4128 1 d0
rlabel metal1 1365 -3610 1393 -3605 1 vdd
rlabel metal1 1362 -4003 1396 -3997 1 gnd
rlabel locali 1195 -3837 1223 -3816 1 d1
rlabel metal1 424 -3759 458 -3753 1 gnd
rlabel metal1 427 -3366 455 -3361 1 vdd
rlabel locali 258 -3589 280 -3574 1 d0
rlabel metal1 422 -3210 456 -3204 1 gnd
rlabel metal1 425 -2817 453 -2812 1 vdd
rlabel locali 256 -3040 278 -3025 1 d0
rlabel metal1 1364 -2507 1392 -2502 1 vdd
rlabel metal1 1361 -2900 1395 -2894 1 gnd
rlabel locali 1194 -2734 1222 -2713 1 d1
rlabel metal1 423 -2656 457 -2650 1 gnd
rlabel metal1 426 -2263 454 -2258 1 vdd
rlabel locali 257 -2486 279 -2471 1 d0
rlabel locali 1332 -1121 1353 -1102 1 d2
rlabel metal1 1501 -1286 1535 -1280 1 gnd
rlabel metal1 1504 -893 1532 -888 1 vdd
rlabel metal1 422 -2107 456 -2101 1 gnd
rlabel metal1 425 -1714 453 -1709 1 vdd
rlabel locali 256 -1937 278 -1922 1 d0
rlabel metal1 1364 -1404 1392 -1399 1 vdd
rlabel metal1 1361 -1797 1395 -1791 1 gnd
rlabel locali 1194 -1631 1222 -1610 1 d1
rlabel metal1 423 -1553 457 -1547 1 gnd
rlabel metal1 426 -1160 454 -1155 1 vdd
rlabel locali 257 -1383 279 -1368 1 d0
rlabel metal1 421 -1004 455 -998 1 gnd
rlabel metal1 424 -611 452 -606 1 vdd
rlabel locali 255 -834 277 -819 1 d0
rlabel metal1 1363 -301 1391 -296 1 vdd
rlabel metal1 1360 -694 1394 -688 1 gnd
rlabel locali 1193 -528 1221 -507 1 d1
rlabel metal1 422 -450 456 -444 1 gnd
rlabel metal1 425 -57 453 -52 1 vdd
rlabel locali 256 -280 278 -265 1 d0
rlabel locali 1933 41 1955 56 1 vout
rlabel metal1 1472 229 1500 234 1 vdd
rlabel metal1 1469 -164 1503 -158 1 gnd
rlabel locali 1296 -2 1331 24 1 d4
<< end >>
