* SPICE3 file created from 6bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_404_5408# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X1 a_1932_3702# a_1719_3702# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X2 a_130_5209# a_135_4823# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3 vref a_116_7550# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4 vdd a_4395_4156# a_4187_4156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X5 vdd a_4390_5137# a_4182_5137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X6 a_838_2470# a_417_2470# a_141_2370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X7 a_3126_4527# a_4187_4156# a_4138_4346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X8 a_4130_6129# a_4126_6306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9 a_408_4012# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X10 a_3118_6310# a_3371_6297# a_3059_7048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X11 gnd a_3383_4337# a_3175_4337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X12 vdd d0 a_4399_3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X13 a_3126_4527# a_4187_4156# a_4142_4169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X14 a_4153_1410# a_4163_667# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X15 a_133_4327# a_622_4427# a_830_4427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X16 gnd a_4410_1220# a_4202_1220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X17 a_155_311# a_641_95# a_849_95# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X18 a_1441_329# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X19 a_2153_n386# a_2880_3905# a_2835_3918# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X20 a_1818_868# a_1436_1310# a_844_1076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X21 a_2930_1926# a_3183_1913# a_2831_4095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X22 a_3095_994# a_3190_1401# a_3141_1591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X23 vdd d0 a_4403_2199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X24 a_629_2055# a_416_2055# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X25 a_1429_2289# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X26 vdd a_4410_1220# a_4202_1220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X27 gnd a_3403_420# a_3195_420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X28 a_1654_329# a_1441_329# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X29 vdd a_3348_981# a_3140_981# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X30 a_3079_3131# a_3336_2941# a_2930_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X31 a_4131_6544# a_4384_6531# a_3118_6310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X32 a_2906_6020# a_3120_4898# a_3075_4911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X33 a_3133_3374# a_3386_3361# a_3083_2954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X34 vdd a_3403_420# a_3195_420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X35 a_143_2271# a_629_2055# a_837_2055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X36 a_1409_6206# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X37 a_4146_3608# a_4142_3785# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X38 a_2041_3702# a_1932_3702# a_2140_3702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X39 a_4127_6721# a_4384_6531# a_3118_6310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X40 vout a_1831_n386# a_2140_3702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X41 vdd a_4403_2199# a_4195_2199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X42 a_416_2055# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X43 a_141_2370# a_143_2271# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X44 a_3129_3551# a_3386_3361# a_3083_2954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X45 a_4125_7110# a_4378_7097# a_3109_7468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X46 a_4142_3785# a_4145_3193# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X47 a_3133_3374# a_4191_3595# a_4146_3608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X48 a_3075_4911# a_3170_5318# a_3125_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X49 a_143_2271# a_150_1887# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X50 a_4126_6306# a_4138_5565# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X51 gnd a_4390_5137# a_4182_5137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X52 a_1617_7187# a_1404_7187# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X53 a_1692_2709# a_1479_2709# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X54 a_1798_4785# a_1416_5227# a_824_4993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X55 a_2831_4095# a_2975_1913# a_2926_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X56 a_3134_2570# a_4195_2199# a_4150_2212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X57 a_4151_2627# a_4404_2614# a_3138_2393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X58 a_844_1076# a_423_1076# a_150_1292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X59 gnd d2 a_3316_6858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X60 a_622_4427# a_409_4427# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X61 a_2906_6020# a_3163_5830# a_2835_3918# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X62 a_2930_1926# a_3128_2941# a_3079_3131# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X63 gnd a_4383_6116# a_4175_6116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X64 a_4147_2804# a_4404_2614# a_3138_2393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X65 a_1404_7187# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X66 a_604_6953# a_391_6953# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X67 vdd a_3088_3905# a_2880_3905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X68 a_4122_7702# a_4125_7110# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X69 a_123_6188# a_609_5972# a_817_5972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X70 gnd d0 a_4416_654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X71 a_1781_6626# a_1409_6206# a_817_5972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X72 a_4163_667# a_4416_654# a_3150_433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X73 a_824_4993# a_403_4993# a_130_5209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X74 vdd a_4383_6116# a_4175_6116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X75 gnd d0 a_4411_1635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X76 a_1837_5694# a_1624_5694# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X77 a_429_510# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X78 vdd d0 a_4416_654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X79 a_3129_3551# a_4190_3180# a_4141_3370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X80 a_4159_844# a_4416_654# a_3150_433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X81 a_1644_1777# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X82 gnd a_3316_6858# a_3108_6858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X83 a_428_95# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X84 vdd d0 a_4411_1635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X85 a_829_4012# a_1634_4246# a_1793_4666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X86 a_4121_7287# a_4131_6544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X87 a_155_906# a_636_1076# a_844_1076# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X88 a_153_692# a_153_410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X89 gnd a_3371_6297# a_3163_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X90 a_4154_1825# a_4157_1233# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X91 a_391_6953# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X92 a_3129_3551# a_4190_3180# a_4145_3193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X93 a_136_3351# a_625_3451# a_833_3451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X94 a_1806_2828# a_1424_3270# a_833_3451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X95 a_3075_4911# a_3170_5318# a_3121_5508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X96 a_1624_5694# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X97 a_617_5408# a_404_5408# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X98 a_849_95# a_428_95# a_162_110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X99 a_2835_3918# a_2955_5830# a_2910_5843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X100 a_850_510# a_429_510# a_153_692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X101 a_1801_2709# a_1692_2709# a_1900_2709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X102 a_3109_7468# a_4170_7097# a_4125_7110# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X103 a_630_2470# a_417_2470# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X104 a_813_7368# a_392_7368# a_116_7268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X105 a_4143_4584# a_4396_4571# a_3130_4350# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X106 a_1786_6745# a_1404_7187# a_813_7368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X107 a_3145_1414# a_3398_1401# a_3095_994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X108 a_2910_5843# a_3108_6858# a_3063_6871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X109 a_641_95# a_428_95# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X110 a_128_5590# a_617_5408# a_825_5408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X111 a_1459_6626# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X112 a_1491_749# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X113 a_1912_749# a_1491_749# a_1813_749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X114 a_4139_4761# a_4396_4571# a_3130_4350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X115 a_3071_5088# a_3328_4898# a_2906_6020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X116 a_610_6387# a_397_6387# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X117 a_4134_5742# a_4137_5150# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X118 a_404_5408# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X119 a_143_2866# a_141_2652# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X120 a_624_3036# a_411_3036# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X121 a_3063_6871# a_3158_7278# a_3113_7291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X122 a_135_4228# a_621_4012# a_829_4012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X123 a_3138_2393# a_3391_2380# a_3079_3131# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X124 a_133_4609# a_133_4327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X125 a_4142_3785# a_4399_3595# a_3133_3374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X126 a_3121_5508# a_3378_5318# a_3075_4911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X127 a_408_4012# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X128 a_642_510# a_429_510# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X129 a_3134_2570# a_3391_2380# a_3079_3131# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X130 a_4138_4346# a_4146_3608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X131 gnd d2 a_3328_4898# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X132 a_411_3036# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X133 gnd d4 a_3088_3905# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X134 vdd d0 a_4390_5137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X135 a_3114_6487# a_3371_6297# a_3059_7048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X136 a_1441_329# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X137 a_1793_4666# a_1421_4246# a_829_4012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X138 a_1880_6626# a_1459_6626# a_1781_6626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X139 a_1900_2709# a_1857_1777# a_2041_3702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X140 a_1654_329# a_1441_329# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X141 a_136_3351# a_138_3252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X142 a_4158_429# a_162_110# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X143 a_818_6387# a_1622_6206# a_1781_6626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X144 a_604_6953# a_391_6953# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X145 gnd a_3328_4898# a_3120_4898# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X146 a_2045_5694# a_1624_5694# a_1892_4666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X147 a_397_6387# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X148 a_4150_2212# a_4403_2199# a_3134_2570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X149 a_1409_6206# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X150 a_150_1887# a_629_2055# a_837_2055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X151 a_4145_3193# a_4398_3180# a_3129_3551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X152 a_121_6569# a_121_6287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X153 a_136_3633# a_136_3351# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X154 a_123_6188# a_130_5804# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X155 a_1637_3270# a_1424_3270# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X156 a_844_1076# a_1649_1310# a_1818_868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X157 a_3063_6871# a_3158_7278# a_3109_7468# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X158 a_4141_3370# a_4398_3180# a_3129_3551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X159 gnd a_4399_3595# a_4191_3595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X160 a_391_6953# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X161 a_3121_5508# a_4182_5137# a_4137_5150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X162 a_3125_5331# a_3378_5318# a_3075_4911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X163 a_1798_4785# a_1416_5227# a_825_5408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X164 vout a_1831_n386# a_2153_n386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X165 a_838_2470# a_417_2470# a_141_2652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X166 gnd d2 a_3336_2941# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X167 a_4121_7287# a_4378_7097# a_3109_7468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X168 a_1798_4785# a_1684_4666# a_1892_4666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X169 a_813_7368# a_1617_7187# a_1786_6745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X170 a_1424_3270# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X171 a_622_4427# a_409_4427# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X172 gnd d0 a_4390_5137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X173 a_3141_1591# a_4202_1220# a_4153_1410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X174 a_636_1076# a_423_1076# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X175 a_818_6387# a_397_6387# a_121_6569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X176 a_1781_6626# a_1409_6206# a_818_6387# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X177 a_3141_1591# a_4202_1220# a_4157_1233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X178 a_4142_4169# a_4138_4346# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X179 gnd a_3336_2941# a_3128_2941# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X180 a_1818_868# a_1436_1310# a_845_1491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X181 a_123_6783# a_604_6953# a_812_6953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X182 gnd a_3391_2380# a_3183_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X183 a_423_1076# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X184 a_838_2470# a_1642_2289# a_1801_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X185 vdd a_3391_2380# a_3183_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X186 a_637_1491# a_424_1491# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X187 a_3126_4527# a_3383_4337# a_3071_5088# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X188 a_1892_4666# a_1471_4666# a_1793_4666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X189 gnd d3 a_3163_5830# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X190 a_4125_7110# a_4121_7287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X191 a_428_95# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X192 a_849_95# a_428_95# a_155_311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X193 a_3095_994# a_3190_1401# a_3145_1414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X194 a_1801_2709# a_1429_2289# a_838_2470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X195 a_3121_5508# a_4182_5137# a_4133_5327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X196 a_833_3451# a_412_3451# a_136_3351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X197 a_153_692# a_642_510# a_850_510# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X198 a_4158_429# a_4415_239# a_3146_610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X199 vdd d0 a_4415_239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X200 a_1719_3702# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X201 vdd d2 a_3316_6858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X202 a_2044_n386# a_1831_n386# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X203 a_138_3847# a_136_3633# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X204 vdd a_3371_6297# a_3163_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X205 a_616_4993# a_403_4993# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X206 a_813_7368# a_392_7368# a_116_7550# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X207 a_1459_6626# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X208 a_128_5308# a_617_5408# a_825_5408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X209 a_1912_749# a_1491_749# a_1818_868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X210 a_424_1491# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X211 a_1491_749# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X212 a_153_410# a_155_311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X213 gnd a_3163_5830# a_2955_5830# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X214 vdd d1 a_3366_7278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X215 a_817_5972# a_396_5972# a_123_6188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X216 a_2926_2103# a_3183_1913# a_2831_4095# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X217 a_1831_n386# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X218 a_624_3036# a_411_3036# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X219 vdd a_3316_6858# a_3108_6858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X220 gnd d3 a_3183_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X221 a_138_3847# a_621_4012# a_829_4012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X222 a_403_4993# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X223 gnd d0 a_4384_6531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X224 gnd d2 a_3348_981# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X225 a_138_3252# a_624_3036# a_832_3036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X226 gnd d1 a_3386_3361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X227 vdd a_3366_7278# a_3158_7278# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X228 a_3059_7048# a_3163_6297# a_3114_6487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X229 a_2153_n386# a_2880_3905# a_2831_4095# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X230 a_411_3036# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X231 a_138_3252# a_143_2866# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X232 vdd d0 a_4384_6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X233 a_1818_868# a_1704_749# a_1912_749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X234 vdd d1 a_3386_3361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X235 a_3130_4350# a_3383_4337# a_3071_5088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X236 a_1793_4666# a_1421_4246# a_830_4427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X237 a_1880_6626# a_1459_6626# a_1786_6745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X238 a_1912_749# a_1857_1777# a_2041_3702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X239 a_116_7550# a_116_7268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X240 gnd d0 a_4415_239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X241 a_4162_252# a_4415_239# a_3146_610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X242 gnd a_3348_981# a_3140_981# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X243 a_4162_252# a_4158_429# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X244 a_641_95# a_428_95# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X245 a_2831_4095# a_2975_1913# a_2930_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X246 a_121_6569# a_610_6387# a_818_6387# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X247 a_817_5972# a_1622_6206# a_1781_6626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X248 a_417_2470# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X249 a_1892_4666# a_1837_5694# a_2045_5694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X250 a_2930_1926# a_3128_2941# a_3083_2954# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X251 a_4159_844# a_4162_252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X252 a_1479_2709# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X253 gnd d1 a_3366_7278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X254 a_3118_6310# a_4176_6531# a_4127_6721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X255 a_3083_2954# a_3178_3361# a_3129_3551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X256 a_118_7169# a_604_6953# a_812_6953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X257 a_837_2055# a_416_2055# a_150_1887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X258 a_845_1491# a_424_1491# a_148_1391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X259 a_621_4012# a_408_4012# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X260 a_3118_6310# a_4176_6531# a_4131_6544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X261 a_4146_2389# a_4403_2199# a_3134_2570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X262 a_3083_2954# a_3178_3361# a_3133_3374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X263 a_3141_1591# a_3398_1401# a_3095_994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X264 gnd a_3366_7278# a_3158_7278# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X265 gnd d0 a_4410_1220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X266 a_1793_4666# a_1684_4666# a_1892_4666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X267 gnd a_3088_3905# a_2880_3905# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X268 a_1629_5227# a_1416_5227# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X269 a_4138_5565# a_4134_5742# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X270 a_636_1076# a_423_1076# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X271 a_4150_2212# a_4146_2389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X272 a_1642_2289# a_1429_2289# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X273 vdd d0 a_4410_1220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X274 a_148_1673# a_637_1491# a_845_1491# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X275 a_1900_2709# a_1479_2709# a_1801_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X276 a_4130_6129# a_4383_6116# a_3114_6487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X277 a_4138_5565# a_4391_5552# a_3125_5331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X278 a_2831_4095# a_3088_3905# a_2153_n386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X279 a_817_5972# a_396_5972# a_130_5804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X280 gnd d0 a_4396_4571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X281 a_1622_6206# a_1409_6206# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X282 gnd d1 a_3398_1401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X283 a_1416_5227# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X284 a_2906_6020# a_3120_4898# a_3071_5088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X285 a_616_4993# a_403_4993# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X286 a_4126_6306# a_4383_6116# a_3114_6487# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X287 a_1813_749# a_1441_329# a_849_95# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X288 a_4134_5742# a_4391_5552# a_3125_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X289 gnd a_4379_7512# a_4171_7512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X290 a_423_1076# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X291 a_1429_2289# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X292 vdd d0 a_4396_4571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X293 a_3063_6871# a_3316_6858# a_2910_5843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X294 a_1892_4666# a_1471_4666# a_1798_4785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X295 vdd a_4379_7512# a_4171_7512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X296 a_4145_3193# a_4141_3370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X297 a_148_1391# a_150_1292# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X298 gnd d1 a_3391_2380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X299 a_833_3451# a_412_3451# a_136_3633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X300 gnd a_4396_4571# a_4188_4571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X301 gnd a_3398_1401# a_3190_1401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X302 a_4131_6544# a_4127_6721# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X303 a_1637_3270# a_1424_3270# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X304 a_1719_3702# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X305 a_403_4993# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X306 a_4158_1648# a_4411_1635# a_3145_1414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X307 a_4133_5327# a_4143_4584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X308 a_4127_6721# a_4130_6129# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X309 vdd d1 a_3391_2380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X310 vdd a_4396_4571# a_4188_4571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X311 a_148_1673# a_148_1391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X312 a_4154_1825# a_4411_1635# a_3145_1414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X313 a_605_7368# a_392_7368# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X314 a_3130_4350# a_4188_4571# a_4139_4761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X315 a_1617_7187# a_1404_7187# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X316 a_2044_n386# a_1831_n386# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X317 a_130_5209# a_616_4993# a_824_4993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X318 a_825_5408# a_404_5408# a_128_5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X319 a_155_906# a_153_692# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X320 a_1424_3270# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X321 vdd a_4399_3595# a_4191_3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X322 gnd d1 a_3403_420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X323 a_3130_4350# a_4188_4571# a_4143_4584# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X324 a_3091_1171# a_3348_981# a_2926_2103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X325 vdd d2 a_3348_981# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X326 a_3150_433# a_3403_420# a_3091_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X327 a_833_3451# a_1637_3270# a_1806_2828# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X328 gnd a_4122_7702# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X329 gnd a_4416_654# a_4208_654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X330 gnd d1 a_3371_6297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X331 vdd d1 a_3403_420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X332 a_829_4012# a_408_4012# a_138_3847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X333 a_392_7368# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X334 a_3146_610# a_3403_420# a_3091_1171# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X335 a_3079_3131# a_3183_2380# a_3134_2570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X336 a_1404_7187# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X337 a_143_2866# a_624_3036# a_832_3036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X338 a_128_5590# a_128_5308# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X339 a_1831_n386# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X340 gnd d0 a_4398_3180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X341 vdd a_4416_654# a_4208_654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X342 a_4157_1233# a_4153_1410# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X343 a_1813_749# a_1704_749# a_1912_749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X344 a_3079_3131# a_3183_2380# a_3138_2393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X345 a_141_2652# a_141_2370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X346 vdd d0 a_4398_3180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X347 a_141_2652# a_630_2470# a_838_2470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X348 a_4142_4169# a_4395_4156# a_3126_4527# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X349 a_1634_4246# a_1421_4246# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X350 a_1672_6626# a_1459_6626# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X351 a_3059_7048# a_3163_6297# a_3118_6310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X352 vdd d2 a_3336_2941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X353 a_3091_1171# a_3195_420# a_3146_610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X354 a_2041_3702# a_1644_1777# a_1912_749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X355 gnd a_4398_3180# a_4190_3180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X356 a_4138_4346# a_4395_4156# a_3126_4527# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X357 a_153_410# a_642_510# a_850_510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X358 gnd a_4391_5552# a_4183_5552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X359 a_1479_2709# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X360 a_3075_4911# a_3328_4898# a_2906_6020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X361 a_1837_5694# a_1624_5694# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X362 a_3091_1171# a_3195_420# a_3150_433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X363 vdd a_4398_3180# a_4190_3180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X364 gnd a_3183_1913# a_2975_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X365 a_4137_5150# a_4133_5327# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X366 vdd a_4391_5552# a_4183_5552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X367 a_3150_433# a_4208_654# a_4159_844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X368 a_837_2055# a_416_2055# a_143_2271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X369 gnd d0 a_4378_7097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X370 a_150_1887# a_148_1673# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X371 a_621_4012# a_408_4012# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X372 a_1421_4246# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X373 a_409_4427# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X374 vdd a_3336_2941# a_3128_2941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X375 a_133_4327# a_135_4228# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X376 gnd a_4384_6531# a_4176_6531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X377 a_2926_2103# a_3140_981# a_3095_994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X378 a_3150_433# a_4208_654# a_4163_667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X379 gnd a_3386_3361# a_3178_3361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X380 a_1649_1310# a_1436_1310# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X381 a_135_4228# a_138_3847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X382 gnd d0 a_4404_2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X383 a_1624_5694# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X384 gnd a_4411_1635# a_4203_1635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X385 vdd a_4384_6531# a_4176_6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X386 a_2153_n386# a_2044_n386# vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X387 vdd a_3386_3361# a_3178_3361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X388 a_1629_5227# a_1416_5227# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X389 gnd a_4378_7097# a_4170_7097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X390 a_1857_1777# a_1644_1777# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X391 vdd d3 a_3163_5830# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X392 vdd d0 a_4404_2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X393 vdd a_4411_1635# a_4203_1635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X394 vdd d1 a_3383_4337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X395 a_1786_6745# a_1404_7187# a_812_6953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X396 a_1900_2709# a_1479_2709# a_1806_2828# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X397 a_2926_2103# a_3140_981# a_3091_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X398 a_1436_1310# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X399 a_825_5408# a_1629_5227# a_1798_4785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X400 gnd a_4404_2614# a_4196_2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X401 a_1786_6745# a_1672_6626# a_1880_6626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X402 a_610_6387# a_397_6387# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X403 a_1622_6206# a_1409_6206# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X404 a_1416_5227# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X405 a_1704_749# a_1491_749# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X406 a_1813_749# a_1441_329# a_850_510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X407 a_830_4427# a_409_4427# a_133_4327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X408 vdd a_3163_5830# a_2955_5830# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X409 a_150_1292# a_155_906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X410 vdd a_4404_2614# a_4196_2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X411 a_417_2470# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X412 a_3083_2954# a_3336_2941# a_2930_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X413 a_118_7169# a_123_6783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X414 a_812_6953# a_391_6953# a_118_7169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X415 a_121_6287# a_123_6188# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X416 gnd d0 a_4399_3595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X417 vdd d3 a_3183_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X418 a_3138_2393# a_4196_2614# a_4147_2804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X419 a_135_4823# a_616_4993# a_824_4993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X420 a_2045_5694# a_1624_5694# a_1880_6626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X421 a_397_6387# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X422 a_4151_2627# a_4147_2804# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X423 a_3138_2393# a_4196_2614# a_4151_2627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X424 a_3071_5088# a_3175_4337# a_3130_4350# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X425 a_1684_4666# a_1471_4666# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X426 gnd d0 a_4379_7512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X427 a_4147_2804# a_4150_2212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X428 a_625_3451# a_412_3451# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X429 a_2140_3702# a_1719_3702# a_2041_3702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X430 a_605_7368# a_392_7368# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X431 vdd d0 a_4379_7512# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X432 a_850_510# a_1654_329# a_1813_749# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X433 vdd d2 a_3328_4898# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X434 a_825_5408# a_404_5408# a_128_5590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X435 gnd d1 a_3383_4337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X436 a_1471_4666# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X437 a_2910_5843# a_3163_5830# a_2835_3918# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X438 a_3133_3374# a_4191_3595# a_4142_3785# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X439 a_116_7550# a_605_7368# a_813_7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X440 a_609_5972# a_396_5972# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X441 a_412_3451# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X442 a_812_6953# a_1617_7187# a_1786_6745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X443 a_135_4823# a_133_4609# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X444 a_3059_7048# a_3316_6858# a_2910_5843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X445 vdd d1 a_3378_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X446 a_829_4012# a_408_4012# a_135_4228# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X447 a_392_7368# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X448 vdd a_3328_4898# a_3120_4898# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X449 a_3113_7291# a_4171_7512# a_4122_7702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X450 a_4146_2389# a_4158_1648# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X451 a_832_3036# a_411_3036# a_143_2866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X452 a_3109_7468# a_3366_7278# a_3063_6871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X453 a_396_5972# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X454 a_3113_7291# a_4171_7512# gnd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X455 a_1932_3702# a_1719_3702# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X456 vdd d1 a_3371_6297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X457 vdd a_3378_5318# a_3170_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X458 a_3071_5088# a_3175_4337# a_3126_4527# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X459 a_837_2055# a_1642_2289# a_1801_2709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X460 a_1634_4246# a_1421_4246# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X461 a_1672_6626# a_1459_6626# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X462 vdd d1 a_3398_1401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X463 a_2041_3702# a_1644_1777# a_1900_2709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X464 a_2835_3918# a_2955_5830# a_2906_6020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X465 vdd a_4415_239# a_4207_239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X466 a_3095_994# a_3348_981# a_2926_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X467 a_818_6387# a_397_6387# a_121_6287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X468 a_128_5308# a_130_5209# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X469 gnd d0 a_4403_2199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X470 a_123_6783# a_121_6569# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X471 a_133_4609# a_622_4427# a_830_4427# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X472 a_4143_4584# a_4139_4761# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X473 a_1421_4246# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X474 a_409_4427# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X475 gnd d0 a_4383_6116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X476 a_429_510# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X477 vdd a_3398_1401# a_3190_1401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X478 a_812_6953# a_391_6953# a_123_6783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X479 gnd d0 a_4391_5552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X480 a_162_110# a_641_95# a_849_95# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X481 vdd d4 a_3088_3905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X482 a_4139_4761# a_4142_4169# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X483 gnd d1 a_3378_5318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X484 a_629_2055# a_416_2055# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X485 a_637_1491# a_424_1491# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X486 gnd a_4403_2199# a_4195_2199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X487 vdd d0 a_4383_6116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X488 vdd d0 a_4391_5552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X489 a_155_311# a_162_110# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X490 a_1801_2709# a_1429_2289# a_837_2055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X491 a_832_3036# a_1637_3270# a_1806_2828# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X492 vdd d0 a_4378_7097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X493 a_1857_1777# a_1644_1777# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X494 a_1806_2828# a_1424_3270# a_832_3036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X495 a_3113_7291# a_3366_7278# a_3063_6871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X496 a_3134_2570# a_4195_2199# a_4146_2389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X497 a_2045_5694# a_1932_3702# a_2140_3702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X498 a_2835_3918# a_3088_3905# a_2153_n386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X499 a_850_510# a_429_510# a_153_410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X500 a_4133_5327# a_4390_5137# a_3121_5508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X501 gnd a_3378_5318# a_3170_5318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X502 a_3146_610# a_4207_239# a_4162_252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X503 a_416_2055# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X504 a_630_2470# a_417_2470# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X505 a_824_4993# a_1629_5227# a_1798_4785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X506 a_424_1491# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X507 a_116_7268# a_118_7169# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X508 a_2140_3702# a_2044_n386# vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X509 a_1781_6626# a_1672_6626# a_1880_6626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X510 a_141_2370# a_630_2470# a_838_2470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X511 vdd a_4378_7097# a_4170_7097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X512 gnd a_4415_239# a_4207_239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X513 a_1692_2709# a_1479_2709# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X514 a_4146_3608# a_4399_3595# a_3133_3374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X515 a_3114_6487# a_4175_6116# a_4126_6306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X516 a_1704_749# a_1491_749# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X517 a_830_4427# a_409_4427# a_133_4609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X518 a_3125_5331# a_4183_5552# a_4134_5742# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X519 a_609_5972# a_396_5972# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X520 a_4157_1233# a_4410_1220# a_3141_1591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X521 a_844_1076# a_423_1076# a_155_906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X522 a_3114_6487# a_4175_6116# a_4130_6129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X523 a_121_6287# a_610_6387# a_818_6387# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X524 a_3125_5331# a_4183_5552# a_4138_5565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X525 gnd a_4379_7512# a_3113_7291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X526 a_4153_1410# a_4410_1220# a_3141_1591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X527 a_2910_5843# a_3108_6858# a_3059_7048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X528 a_1684_4666# a_1471_4666# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X529 a_4122_7702# a_4379_7512# a_3113_7291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X530 a_642_510# a_429_510# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X531 a_396_5972# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X532 a_625_3451# a_412_3451# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X533 a_1644_1777# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X534 a_3145_1414# a_4203_1635# a_4154_1825# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X535 a_130_5804# a_128_5590# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X536 a_845_1491# a_424_1491# a_148_1673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X537 a_2140_3702# a_1719_3702# a_2045_5694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X538 a_849_95# a_1654_329# a_1813_749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X539 a_830_4427# a_1634_4246# a_1793_4666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X540 a_3109_7468# a_4170_7097# a_4121_7287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X541 a_150_1292# a_636_1076# a_844_1076# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X542 a_1649_1310# a_1436_1310# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X543 vdd a_3383_4337# a_3175_4337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X544 a_4163_667# a_4159_844# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X545 a_4137_5150# a_4390_5137# a_3121_5508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X546 a_3145_1414# a_4203_1635# a_4158_1648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X547 a_136_3633# a_625_3451# a_833_3451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X548 a_3146_610# a_4207_239# a_4158_429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X549 gnd d0 a_4395_4156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X550 a_1471_4666# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X551 a_4141_3370# a_4151_2627# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X552 a_1880_6626# a_1837_5694# a_2045_5694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X553 a_824_4993# a_403_4993# a_135_4823# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X554 a_116_7268# a_605_7368# a_813_7368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X555 a_617_5408# a_404_5408# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X556 a_412_3451# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X557 a_4158_1648# a_4154_1825# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X558 a_1806_2828# a_1692_2709# a_1900_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X559 vdd d0 a_4395_4156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X560 a_1642_2289# a_1429_2289# vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X561 a_1436_1310# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X562 a_148_1391# a_637_1491# a_845_1491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X563 a_130_5804# a_609_5972# a_817_5972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X564 vdd a_3183_1913# a_2975_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X565 a_845_1491# a_1649_1310# a_1818_868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
X566 a_832_3036# a_411_3036# a_138_3252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X567 gnd a_4395_4156# a_4187_4156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.50
C0 gnd d0 2.57fF
C1 vdd gnd 3.37fF
C2 a_2140_3702# a_2153_n386# 3.90fF
C3 gnd SUB 22.11fF
C4 vdd SUB 85.51fF
C5 a_162_110# SUB 6.03fF
C6 d0 SUB 8.45fF
C7 a_849_95# SUB 2.20fF
C8 d1 SUB 5.40fF
C9 a_3146_610# SUB 2.33fF
C10 a_3150_433# SUB 2.20fF
C11 a_1813_749# SUB 2.04fF
C12 d2 SUB 2.56fF
C13 a_844_1076# SUB 2.20fF
C14 a_3095_994# SUB 2.04fF
C15 a_3141_1591# SUB 2.33fF
C16 a_3145_1414# SUB 2.20fF
C17 a_1912_749# SUB 2.78fF
C18 a_2926_2103# SUB 2.02fF
C19 a_3134_2570# SUB 2.33fF
C20 a_3138_2393# SUB 2.20fF
C21 a_1801_2709# SUB 2.04fF
C22 a_1900_2709# SUB 2.02fF
C23 a_2930_1926# SUB 2.78fF
C24 a_832_3036# SUB 2.20fF
C25 a_3083_2954# SUB 2.04fF
C26 a_3129_3551# SUB 2.33fF
C27 a_3133_3374# SUB 2.20fF
C28 a_2041_3702# SUB 3.86fF
C29 a_2140_3702# SUB 4.80fF
C30 a_2153_n386# SUB 5.58fF
C31 a_2831_4095# SUB 2.93fF
C32 a_829_4012# SUB 2.20fF
C33 a_3126_4527# SUB 2.33fF
C34 a_830_4427# SUB 2.33fF
C35 a_3130_4350# SUB 2.20fF
C36 a_1793_4666# SUB 2.04fF
C37 a_824_4993# SUB 2.20fF
C38 a_3075_4911# SUB 2.04fF
C39 a_3121_5508# SUB 2.33fF
C40 a_3125_5331# SUB 2.20fF
C41 a_1892_4666# SUB 2.78fF
C42 a_2045_5694# SUB 2.93fF
C43 a_2835_3918# SUB 3.86fF
C44 a_2906_6020# SUB 2.02fF
C45 a_817_5972# SUB 2.20fF
C46 a_3114_6487# SUB 2.33fF
C47 a_818_6387# SUB 2.33fF
C48 a_3118_6310# SUB 2.20fF
C49 a_1781_6626# SUB 2.04fF
C50 a_1880_6626# SUB 2.02fF
C51 a_2910_5843# SUB 2.78fF
C52 a_812_6953# SUB 2.20fF
C53 a_3063_6871# SUB 2.04fF
C54 a_3109_7468# SUB 2.33fF
C55 a_813_7368# SUB 2.33fF
C56 a_3113_7291# SUB 2.20fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0 0.1ps 0.1ps 5us 10us)
Vd1 d1 0 pulse(0 1.8 0 0.1ps 0.1ps 10us 20us)
Vd2 d2 0 pulse(0 1.8 0 0.1ps 0.1ps 20us 40us)
Vd3 d3 0 pulse(0 1.8 0 0.1ps 0.1ps 40us 80us)
Vd4 d4 0 pulse(0 1.8 0 0.1ps 0.1ps 80us 160us)
Vd5 d5 0 pulse(0 1.8 0 0.1ps 0.1ps 160us 320us)


.tran 1us 320us
.control
run
plot V(vout)
.endc
.end
