magic
tech sky130A
timestamp 1633153601
<< nwell >>
rect 752 11541 1563 11765
rect 1800 11537 2611 11761
rect 752 10862 1563 11086
rect 3247 10857 4058 11081
rect 752 10094 1563 10318
rect 1800 10090 2611 10314
rect 752 9415 1563 9639
rect 3290 9412 4101 9636
rect 753 8574 1564 8798
rect 1801 8570 2612 8794
rect 753 7895 1564 8119
rect 3248 7890 4059 8114
rect 753 7127 1564 7351
rect 1801 7123 2612 7347
rect 753 6448 1564 6672
rect 4356 6439 5167 6663
rect 750 5533 1561 5757
rect 1798 5529 2609 5753
rect 750 4854 1561 5078
rect 3245 4849 4056 5073
rect 750 4086 1561 4310
rect 1798 4082 2609 4306
rect 750 3407 1561 3631
rect 3288 3404 4099 3628
rect 751 2566 1562 2790
rect 1799 2562 2610 2786
rect 751 1887 1562 2111
rect 3246 1882 4057 2106
rect 751 1119 1562 1343
rect 1799 1115 2610 1339
rect 751 440 1562 664
<< nmos >>
rect 816 11440 866 11482
rect 1029 11440 1079 11482
rect 1237 11440 1287 11482
rect 1445 11440 1495 11482
rect 1864 11436 1914 11478
rect 2077 11436 2127 11478
rect 2285 11436 2335 11478
rect 2493 11436 2543 11478
rect 816 10761 866 10803
rect 1029 10761 1079 10803
rect 1237 10761 1287 10803
rect 1445 10761 1495 10803
rect 3311 10756 3361 10798
rect 3524 10756 3574 10798
rect 3732 10756 3782 10798
rect 3940 10756 3990 10798
rect 816 9993 866 10035
rect 1029 9993 1079 10035
rect 1237 9993 1287 10035
rect 1445 9993 1495 10035
rect 1864 9989 1914 10031
rect 2077 9989 2127 10031
rect 2285 9989 2335 10031
rect 2493 9989 2543 10031
rect 816 9314 866 9356
rect 1029 9314 1079 9356
rect 1237 9314 1287 9356
rect 1445 9314 1495 9356
rect 3354 9311 3404 9353
rect 3567 9311 3617 9353
rect 3775 9311 3825 9353
rect 3983 9311 4033 9353
rect 817 8473 867 8515
rect 1030 8473 1080 8515
rect 1238 8473 1288 8515
rect 1446 8473 1496 8515
rect 1865 8469 1915 8511
rect 2078 8469 2128 8511
rect 2286 8469 2336 8511
rect 2494 8469 2544 8511
rect 817 7794 867 7836
rect 1030 7794 1080 7836
rect 1238 7794 1288 7836
rect 1446 7794 1496 7836
rect 3312 7789 3362 7831
rect 3525 7789 3575 7831
rect 3733 7789 3783 7831
rect 3941 7789 3991 7831
rect 817 7026 867 7068
rect 1030 7026 1080 7068
rect 1238 7026 1288 7068
rect 1446 7026 1496 7068
rect 1865 7022 1915 7064
rect 2078 7022 2128 7064
rect 2286 7022 2336 7064
rect 2494 7022 2544 7064
rect 817 6347 867 6389
rect 1030 6347 1080 6389
rect 1238 6347 1288 6389
rect 1446 6347 1496 6389
rect 4420 6338 4470 6380
rect 4633 6338 4683 6380
rect 4841 6338 4891 6380
rect 5049 6338 5099 6380
rect 814 5432 864 5474
rect 1027 5432 1077 5474
rect 1235 5432 1285 5474
rect 1443 5432 1493 5474
rect 1862 5428 1912 5470
rect 2075 5428 2125 5470
rect 2283 5428 2333 5470
rect 2491 5428 2541 5470
rect 814 4753 864 4795
rect 1027 4753 1077 4795
rect 1235 4753 1285 4795
rect 1443 4753 1493 4795
rect 3309 4748 3359 4790
rect 3522 4748 3572 4790
rect 3730 4748 3780 4790
rect 3938 4748 3988 4790
rect 814 3985 864 4027
rect 1027 3985 1077 4027
rect 1235 3985 1285 4027
rect 1443 3985 1493 4027
rect 1862 3981 1912 4023
rect 2075 3981 2125 4023
rect 2283 3981 2333 4023
rect 2491 3981 2541 4023
rect 814 3306 864 3348
rect 1027 3306 1077 3348
rect 1235 3306 1285 3348
rect 1443 3306 1493 3348
rect 3352 3303 3402 3345
rect 3565 3303 3615 3345
rect 3773 3303 3823 3345
rect 3981 3303 4031 3345
rect 815 2465 865 2507
rect 1028 2465 1078 2507
rect 1236 2465 1286 2507
rect 1444 2465 1494 2507
rect 1863 2461 1913 2503
rect 2076 2461 2126 2503
rect 2284 2461 2334 2503
rect 2492 2461 2542 2503
rect 815 1786 865 1828
rect 1028 1786 1078 1828
rect 1236 1786 1286 1828
rect 1444 1786 1494 1828
rect 3310 1781 3360 1823
rect 3523 1781 3573 1823
rect 3731 1781 3781 1823
rect 3939 1781 3989 1823
rect 815 1018 865 1060
rect 1028 1018 1078 1060
rect 1236 1018 1286 1060
rect 1444 1018 1494 1060
rect 1863 1014 1913 1056
rect 2076 1014 2126 1056
rect 2284 1014 2334 1056
rect 2492 1014 2542 1056
rect 815 339 865 381
rect 1028 339 1078 381
rect 1236 339 1286 381
rect 1444 339 1494 381
<< pmos >>
rect 816 11559 866 11659
rect 1029 11559 1079 11659
rect 1237 11559 1287 11659
rect 1445 11559 1495 11659
rect 1864 11555 1914 11655
rect 2077 11555 2127 11655
rect 2285 11555 2335 11655
rect 2493 11555 2543 11655
rect 816 10880 866 10980
rect 1029 10880 1079 10980
rect 1237 10880 1287 10980
rect 1445 10880 1495 10980
rect 3311 10875 3361 10975
rect 3524 10875 3574 10975
rect 3732 10875 3782 10975
rect 3940 10875 3990 10975
rect 816 10112 866 10212
rect 1029 10112 1079 10212
rect 1237 10112 1287 10212
rect 1445 10112 1495 10212
rect 1864 10108 1914 10208
rect 2077 10108 2127 10208
rect 2285 10108 2335 10208
rect 2493 10108 2543 10208
rect 816 9433 866 9533
rect 1029 9433 1079 9533
rect 1237 9433 1287 9533
rect 1445 9433 1495 9533
rect 3354 9430 3404 9530
rect 3567 9430 3617 9530
rect 3775 9430 3825 9530
rect 3983 9430 4033 9530
rect 817 8592 867 8692
rect 1030 8592 1080 8692
rect 1238 8592 1288 8692
rect 1446 8592 1496 8692
rect 1865 8588 1915 8688
rect 2078 8588 2128 8688
rect 2286 8588 2336 8688
rect 2494 8588 2544 8688
rect 817 7913 867 8013
rect 1030 7913 1080 8013
rect 1238 7913 1288 8013
rect 1446 7913 1496 8013
rect 3312 7908 3362 8008
rect 3525 7908 3575 8008
rect 3733 7908 3783 8008
rect 3941 7908 3991 8008
rect 817 7145 867 7245
rect 1030 7145 1080 7245
rect 1238 7145 1288 7245
rect 1446 7145 1496 7245
rect 1865 7141 1915 7241
rect 2078 7141 2128 7241
rect 2286 7141 2336 7241
rect 2494 7141 2544 7241
rect 817 6466 867 6566
rect 1030 6466 1080 6566
rect 1238 6466 1288 6566
rect 1446 6466 1496 6566
rect 4420 6457 4470 6557
rect 4633 6457 4683 6557
rect 4841 6457 4891 6557
rect 5049 6457 5099 6557
rect 814 5551 864 5651
rect 1027 5551 1077 5651
rect 1235 5551 1285 5651
rect 1443 5551 1493 5651
rect 1862 5547 1912 5647
rect 2075 5547 2125 5647
rect 2283 5547 2333 5647
rect 2491 5547 2541 5647
rect 814 4872 864 4972
rect 1027 4872 1077 4972
rect 1235 4872 1285 4972
rect 1443 4872 1493 4972
rect 3309 4867 3359 4967
rect 3522 4867 3572 4967
rect 3730 4867 3780 4967
rect 3938 4867 3988 4967
rect 814 4104 864 4204
rect 1027 4104 1077 4204
rect 1235 4104 1285 4204
rect 1443 4104 1493 4204
rect 1862 4100 1912 4200
rect 2075 4100 2125 4200
rect 2283 4100 2333 4200
rect 2491 4100 2541 4200
rect 814 3425 864 3525
rect 1027 3425 1077 3525
rect 1235 3425 1285 3525
rect 1443 3425 1493 3525
rect 3352 3422 3402 3522
rect 3565 3422 3615 3522
rect 3773 3422 3823 3522
rect 3981 3422 4031 3522
rect 815 2584 865 2684
rect 1028 2584 1078 2684
rect 1236 2584 1286 2684
rect 1444 2584 1494 2684
rect 1863 2580 1913 2680
rect 2076 2580 2126 2680
rect 2284 2580 2334 2680
rect 2492 2580 2542 2680
rect 815 1905 865 2005
rect 1028 1905 1078 2005
rect 1236 1905 1286 2005
rect 1444 1905 1494 2005
rect 3310 1900 3360 2000
rect 3523 1900 3573 2000
rect 3731 1900 3781 2000
rect 3939 1900 3989 2000
rect 815 1137 865 1237
rect 1028 1137 1078 1237
rect 1236 1137 1286 1237
rect 1444 1137 1494 1237
rect 1863 1133 1913 1233
rect 2076 1133 2126 1233
rect 2284 1133 2334 1233
rect 2492 1133 2542 1233
rect 815 458 865 558
rect 1028 458 1078 558
rect 1236 458 1286 558
rect 1444 458 1494 558
<< ndiff >>
rect 767 11472 816 11482
rect 767 11452 778 11472
rect 798 11452 816 11472
rect 767 11440 816 11452
rect 866 11476 910 11482
rect 866 11456 881 11476
rect 901 11456 910 11476
rect 866 11440 910 11456
rect 980 11472 1029 11482
rect 980 11452 991 11472
rect 1011 11452 1029 11472
rect 980 11440 1029 11452
rect 1079 11476 1123 11482
rect 1079 11456 1094 11476
rect 1114 11456 1123 11476
rect 1079 11440 1123 11456
rect 1188 11472 1237 11482
rect 1188 11452 1199 11472
rect 1219 11452 1237 11472
rect 1188 11440 1237 11452
rect 1287 11476 1331 11482
rect 1287 11456 1302 11476
rect 1322 11456 1331 11476
rect 1287 11440 1331 11456
rect 1401 11476 1445 11482
rect 1401 11456 1410 11476
rect 1430 11456 1445 11476
rect 1401 11440 1445 11456
rect 1495 11472 1544 11482
rect 1495 11452 1513 11472
rect 1533 11452 1544 11472
rect 1495 11440 1544 11452
rect 1815 11468 1864 11478
rect 1815 11448 1826 11468
rect 1846 11448 1864 11468
rect 1815 11436 1864 11448
rect 1914 11472 1958 11478
rect 1914 11452 1929 11472
rect 1949 11452 1958 11472
rect 1914 11436 1958 11452
rect 2028 11468 2077 11478
rect 2028 11448 2039 11468
rect 2059 11448 2077 11468
rect 2028 11436 2077 11448
rect 2127 11472 2171 11478
rect 2127 11452 2142 11472
rect 2162 11452 2171 11472
rect 2127 11436 2171 11452
rect 2236 11468 2285 11478
rect 2236 11448 2247 11468
rect 2267 11448 2285 11468
rect 2236 11436 2285 11448
rect 2335 11472 2379 11478
rect 2335 11452 2350 11472
rect 2370 11452 2379 11472
rect 2335 11436 2379 11452
rect 2449 11472 2493 11478
rect 2449 11452 2458 11472
rect 2478 11452 2493 11472
rect 2449 11436 2493 11452
rect 2543 11468 2592 11478
rect 2543 11448 2561 11468
rect 2581 11448 2592 11468
rect 2543 11436 2592 11448
rect 767 10793 816 10803
rect 767 10773 778 10793
rect 798 10773 816 10793
rect 767 10761 816 10773
rect 866 10797 910 10803
rect 866 10777 881 10797
rect 901 10777 910 10797
rect 866 10761 910 10777
rect 980 10793 1029 10803
rect 980 10773 991 10793
rect 1011 10773 1029 10793
rect 980 10761 1029 10773
rect 1079 10797 1123 10803
rect 1079 10777 1094 10797
rect 1114 10777 1123 10797
rect 1079 10761 1123 10777
rect 1188 10793 1237 10803
rect 1188 10773 1199 10793
rect 1219 10773 1237 10793
rect 1188 10761 1237 10773
rect 1287 10797 1331 10803
rect 1287 10777 1302 10797
rect 1322 10777 1331 10797
rect 1287 10761 1331 10777
rect 1401 10797 1445 10803
rect 1401 10777 1410 10797
rect 1430 10777 1445 10797
rect 1401 10761 1445 10777
rect 1495 10793 1544 10803
rect 1495 10773 1513 10793
rect 1533 10773 1544 10793
rect 1495 10761 1544 10773
rect 3262 10788 3311 10798
rect 3262 10768 3273 10788
rect 3293 10768 3311 10788
rect 3262 10756 3311 10768
rect 3361 10792 3405 10798
rect 3361 10772 3376 10792
rect 3396 10772 3405 10792
rect 3361 10756 3405 10772
rect 3475 10788 3524 10798
rect 3475 10768 3486 10788
rect 3506 10768 3524 10788
rect 3475 10756 3524 10768
rect 3574 10792 3618 10798
rect 3574 10772 3589 10792
rect 3609 10772 3618 10792
rect 3574 10756 3618 10772
rect 3683 10788 3732 10798
rect 3683 10768 3694 10788
rect 3714 10768 3732 10788
rect 3683 10756 3732 10768
rect 3782 10792 3826 10798
rect 3782 10772 3797 10792
rect 3817 10772 3826 10792
rect 3782 10756 3826 10772
rect 3896 10792 3940 10798
rect 3896 10772 3905 10792
rect 3925 10772 3940 10792
rect 3896 10756 3940 10772
rect 3990 10788 4039 10798
rect 3990 10768 4008 10788
rect 4028 10768 4039 10788
rect 3990 10756 4039 10768
rect 767 10025 816 10035
rect 767 10005 778 10025
rect 798 10005 816 10025
rect 767 9993 816 10005
rect 866 10029 910 10035
rect 866 10009 881 10029
rect 901 10009 910 10029
rect 866 9993 910 10009
rect 980 10025 1029 10035
rect 980 10005 991 10025
rect 1011 10005 1029 10025
rect 980 9993 1029 10005
rect 1079 10029 1123 10035
rect 1079 10009 1094 10029
rect 1114 10009 1123 10029
rect 1079 9993 1123 10009
rect 1188 10025 1237 10035
rect 1188 10005 1199 10025
rect 1219 10005 1237 10025
rect 1188 9993 1237 10005
rect 1287 10029 1331 10035
rect 1287 10009 1302 10029
rect 1322 10009 1331 10029
rect 1287 9993 1331 10009
rect 1401 10029 1445 10035
rect 1401 10009 1410 10029
rect 1430 10009 1445 10029
rect 1401 9993 1445 10009
rect 1495 10025 1544 10035
rect 1495 10005 1513 10025
rect 1533 10005 1544 10025
rect 1495 9993 1544 10005
rect 1815 10021 1864 10031
rect 1815 10001 1826 10021
rect 1846 10001 1864 10021
rect 1815 9989 1864 10001
rect 1914 10025 1958 10031
rect 1914 10005 1929 10025
rect 1949 10005 1958 10025
rect 1914 9989 1958 10005
rect 2028 10021 2077 10031
rect 2028 10001 2039 10021
rect 2059 10001 2077 10021
rect 2028 9989 2077 10001
rect 2127 10025 2171 10031
rect 2127 10005 2142 10025
rect 2162 10005 2171 10025
rect 2127 9989 2171 10005
rect 2236 10021 2285 10031
rect 2236 10001 2247 10021
rect 2267 10001 2285 10021
rect 2236 9989 2285 10001
rect 2335 10025 2379 10031
rect 2335 10005 2350 10025
rect 2370 10005 2379 10025
rect 2335 9989 2379 10005
rect 2449 10025 2493 10031
rect 2449 10005 2458 10025
rect 2478 10005 2493 10025
rect 2449 9989 2493 10005
rect 2543 10021 2592 10031
rect 2543 10001 2561 10021
rect 2581 10001 2592 10021
rect 2543 9989 2592 10001
rect 767 9346 816 9356
rect 767 9326 778 9346
rect 798 9326 816 9346
rect 767 9314 816 9326
rect 866 9350 910 9356
rect 866 9330 881 9350
rect 901 9330 910 9350
rect 866 9314 910 9330
rect 980 9346 1029 9356
rect 980 9326 991 9346
rect 1011 9326 1029 9346
rect 980 9314 1029 9326
rect 1079 9350 1123 9356
rect 1079 9330 1094 9350
rect 1114 9330 1123 9350
rect 1079 9314 1123 9330
rect 1188 9346 1237 9356
rect 1188 9326 1199 9346
rect 1219 9326 1237 9346
rect 1188 9314 1237 9326
rect 1287 9350 1331 9356
rect 1287 9330 1302 9350
rect 1322 9330 1331 9350
rect 1287 9314 1331 9330
rect 1401 9350 1445 9356
rect 1401 9330 1410 9350
rect 1430 9330 1445 9350
rect 1401 9314 1445 9330
rect 1495 9346 1544 9356
rect 1495 9326 1513 9346
rect 1533 9326 1544 9346
rect 1495 9314 1544 9326
rect 3305 9343 3354 9353
rect 3305 9323 3316 9343
rect 3336 9323 3354 9343
rect 3305 9311 3354 9323
rect 3404 9347 3448 9353
rect 3404 9327 3419 9347
rect 3439 9327 3448 9347
rect 3404 9311 3448 9327
rect 3518 9343 3567 9353
rect 3518 9323 3529 9343
rect 3549 9323 3567 9343
rect 3518 9311 3567 9323
rect 3617 9347 3661 9353
rect 3617 9327 3632 9347
rect 3652 9327 3661 9347
rect 3617 9311 3661 9327
rect 3726 9343 3775 9353
rect 3726 9323 3737 9343
rect 3757 9323 3775 9343
rect 3726 9311 3775 9323
rect 3825 9347 3869 9353
rect 3825 9327 3840 9347
rect 3860 9327 3869 9347
rect 3825 9311 3869 9327
rect 3939 9347 3983 9353
rect 3939 9327 3948 9347
rect 3968 9327 3983 9347
rect 3939 9311 3983 9327
rect 4033 9343 4082 9353
rect 4033 9323 4051 9343
rect 4071 9323 4082 9343
rect 4033 9311 4082 9323
rect 768 8505 817 8515
rect 768 8485 779 8505
rect 799 8485 817 8505
rect 768 8473 817 8485
rect 867 8509 911 8515
rect 867 8489 882 8509
rect 902 8489 911 8509
rect 867 8473 911 8489
rect 981 8505 1030 8515
rect 981 8485 992 8505
rect 1012 8485 1030 8505
rect 981 8473 1030 8485
rect 1080 8509 1124 8515
rect 1080 8489 1095 8509
rect 1115 8489 1124 8509
rect 1080 8473 1124 8489
rect 1189 8505 1238 8515
rect 1189 8485 1200 8505
rect 1220 8485 1238 8505
rect 1189 8473 1238 8485
rect 1288 8509 1332 8515
rect 1288 8489 1303 8509
rect 1323 8489 1332 8509
rect 1288 8473 1332 8489
rect 1402 8509 1446 8515
rect 1402 8489 1411 8509
rect 1431 8489 1446 8509
rect 1402 8473 1446 8489
rect 1496 8505 1545 8515
rect 1496 8485 1514 8505
rect 1534 8485 1545 8505
rect 1496 8473 1545 8485
rect 1816 8501 1865 8511
rect 1816 8481 1827 8501
rect 1847 8481 1865 8501
rect 1816 8469 1865 8481
rect 1915 8505 1959 8511
rect 1915 8485 1930 8505
rect 1950 8485 1959 8505
rect 1915 8469 1959 8485
rect 2029 8501 2078 8511
rect 2029 8481 2040 8501
rect 2060 8481 2078 8501
rect 2029 8469 2078 8481
rect 2128 8505 2172 8511
rect 2128 8485 2143 8505
rect 2163 8485 2172 8505
rect 2128 8469 2172 8485
rect 2237 8501 2286 8511
rect 2237 8481 2248 8501
rect 2268 8481 2286 8501
rect 2237 8469 2286 8481
rect 2336 8505 2380 8511
rect 2336 8485 2351 8505
rect 2371 8485 2380 8505
rect 2336 8469 2380 8485
rect 2450 8505 2494 8511
rect 2450 8485 2459 8505
rect 2479 8485 2494 8505
rect 2450 8469 2494 8485
rect 2544 8501 2593 8511
rect 2544 8481 2562 8501
rect 2582 8481 2593 8501
rect 2544 8469 2593 8481
rect 768 7826 817 7836
rect 768 7806 779 7826
rect 799 7806 817 7826
rect 768 7794 817 7806
rect 867 7830 911 7836
rect 867 7810 882 7830
rect 902 7810 911 7830
rect 867 7794 911 7810
rect 981 7826 1030 7836
rect 981 7806 992 7826
rect 1012 7806 1030 7826
rect 981 7794 1030 7806
rect 1080 7830 1124 7836
rect 1080 7810 1095 7830
rect 1115 7810 1124 7830
rect 1080 7794 1124 7810
rect 1189 7826 1238 7836
rect 1189 7806 1200 7826
rect 1220 7806 1238 7826
rect 1189 7794 1238 7806
rect 1288 7830 1332 7836
rect 1288 7810 1303 7830
rect 1323 7810 1332 7830
rect 1288 7794 1332 7810
rect 1402 7830 1446 7836
rect 1402 7810 1411 7830
rect 1431 7810 1446 7830
rect 1402 7794 1446 7810
rect 1496 7826 1545 7836
rect 1496 7806 1514 7826
rect 1534 7806 1545 7826
rect 1496 7794 1545 7806
rect 3263 7821 3312 7831
rect 3263 7801 3274 7821
rect 3294 7801 3312 7821
rect 3263 7789 3312 7801
rect 3362 7825 3406 7831
rect 3362 7805 3377 7825
rect 3397 7805 3406 7825
rect 3362 7789 3406 7805
rect 3476 7821 3525 7831
rect 3476 7801 3487 7821
rect 3507 7801 3525 7821
rect 3476 7789 3525 7801
rect 3575 7825 3619 7831
rect 3575 7805 3590 7825
rect 3610 7805 3619 7825
rect 3575 7789 3619 7805
rect 3684 7821 3733 7831
rect 3684 7801 3695 7821
rect 3715 7801 3733 7821
rect 3684 7789 3733 7801
rect 3783 7825 3827 7831
rect 3783 7805 3798 7825
rect 3818 7805 3827 7825
rect 3783 7789 3827 7805
rect 3897 7825 3941 7831
rect 3897 7805 3906 7825
rect 3926 7805 3941 7825
rect 3897 7789 3941 7805
rect 3991 7821 4040 7831
rect 3991 7801 4009 7821
rect 4029 7801 4040 7821
rect 3991 7789 4040 7801
rect 768 7058 817 7068
rect 768 7038 779 7058
rect 799 7038 817 7058
rect 768 7026 817 7038
rect 867 7062 911 7068
rect 867 7042 882 7062
rect 902 7042 911 7062
rect 867 7026 911 7042
rect 981 7058 1030 7068
rect 981 7038 992 7058
rect 1012 7038 1030 7058
rect 981 7026 1030 7038
rect 1080 7062 1124 7068
rect 1080 7042 1095 7062
rect 1115 7042 1124 7062
rect 1080 7026 1124 7042
rect 1189 7058 1238 7068
rect 1189 7038 1200 7058
rect 1220 7038 1238 7058
rect 1189 7026 1238 7038
rect 1288 7062 1332 7068
rect 1288 7042 1303 7062
rect 1323 7042 1332 7062
rect 1288 7026 1332 7042
rect 1402 7062 1446 7068
rect 1402 7042 1411 7062
rect 1431 7042 1446 7062
rect 1402 7026 1446 7042
rect 1496 7058 1545 7068
rect 1496 7038 1514 7058
rect 1534 7038 1545 7058
rect 1496 7026 1545 7038
rect 1816 7054 1865 7064
rect 1816 7034 1827 7054
rect 1847 7034 1865 7054
rect 1816 7022 1865 7034
rect 1915 7058 1959 7064
rect 1915 7038 1930 7058
rect 1950 7038 1959 7058
rect 1915 7022 1959 7038
rect 2029 7054 2078 7064
rect 2029 7034 2040 7054
rect 2060 7034 2078 7054
rect 2029 7022 2078 7034
rect 2128 7058 2172 7064
rect 2128 7038 2143 7058
rect 2163 7038 2172 7058
rect 2128 7022 2172 7038
rect 2237 7054 2286 7064
rect 2237 7034 2248 7054
rect 2268 7034 2286 7054
rect 2237 7022 2286 7034
rect 2336 7058 2380 7064
rect 2336 7038 2351 7058
rect 2371 7038 2380 7058
rect 2336 7022 2380 7038
rect 2450 7058 2494 7064
rect 2450 7038 2459 7058
rect 2479 7038 2494 7058
rect 2450 7022 2494 7038
rect 2544 7054 2593 7064
rect 2544 7034 2562 7054
rect 2582 7034 2593 7054
rect 2544 7022 2593 7034
rect 768 6379 817 6389
rect 768 6359 779 6379
rect 799 6359 817 6379
rect 768 6347 817 6359
rect 867 6383 911 6389
rect 867 6363 882 6383
rect 902 6363 911 6383
rect 867 6347 911 6363
rect 981 6379 1030 6389
rect 981 6359 992 6379
rect 1012 6359 1030 6379
rect 981 6347 1030 6359
rect 1080 6383 1124 6389
rect 1080 6363 1095 6383
rect 1115 6363 1124 6383
rect 1080 6347 1124 6363
rect 1189 6379 1238 6389
rect 1189 6359 1200 6379
rect 1220 6359 1238 6379
rect 1189 6347 1238 6359
rect 1288 6383 1332 6389
rect 1288 6363 1303 6383
rect 1323 6363 1332 6383
rect 1288 6347 1332 6363
rect 1402 6383 1446 6389
rect 1402 6363 1411 6383
rect 1431 6363 1446 6383
rect 1402 6347 1446 6363
rect 1496 6379 1545 6389
rect 1496 6359 1514 6379
rect 1534 6359 1545 6379
rect 1496 6347 1545 6359
rect 4371 6370 4420 6380
rect 4371 6350 4382 6370
rect 4402 6350 4420 6370
rect 4371 6338 4420 6350
rect 4470 6374 4514 6380
rect 4470 6354 4485 6374
rect 4505 6354 4514 6374
rect 4470 6338 4514 6354
rect 4584 6370 4633 6380
rect 4584 6350 4595 6370
rect 4615 6350 4633 6370
rect 4584 6338 4633 6350
rect 4683 6374 4727 6380
rect 4683 6354 4698 6374
rect 4718 6354 4727 6374
rect 4683 6338 4727 6354
rect 4792 6370 4841 6380
rect 4792 6350 4803 6370
rect 4823 6350 4841 6370
rect 4792 6338 4841 6350
rect 4891 6374 4935 6380
rect 4891 6354 4906 6374
rect 4926 6354 4935 6374
rect 4891 6338 4935 6354
rect 5005 6374 5049 6380
rect 5005 6354 5014 6374
rect 5034 6354 5049 6374
rect 5005 6338 5049 6354
rect 5099 6370 5148 6380
rect 5099 6350 5117 6370
rect 5137 6350 5148 6370
rect 5099 6338 5148 6350
rect 765 5464 814 5474
rect 765 5444 776 5464
rect 796 5444 814 5464
rect 765 5432 814 5444
rect 864 5468 908 5474
rect 864 5448 879 5468
rect 899 5448 908 5468
rect 864 5432 908 5448
rect 978 5464 1027 5474
rect 978 5444 989 5464
rect 1009 5444 1027 5464
rect 978 5432 1027 5444
rect 1077 5468 1121 5474
rect 1077 5448 1092 5468
rect 1112 5448 1121 5468
rect 1077 5432 1121 5448
rect 1186 5464 1235 5474
rect 1186 5444 1197 5464
rect 1217 5444 1235 5464
rect 1186 5432 1235 5444
rect 1285 5468 1329 5474
rect 1285 5448 1300 5468
rect 1320 5448 1329 5468
rect 1285 5432 1329 5448
rect 1399 5468 1443 5474
rect 1399 5448 1408 5468
rect 1428 5448 1443 5468
rect 1399 5432 1443 5448
rect 1493 5464 1542 5474
rect 1493 5444 1511 5464
rect 1531 5444 1542 5464
rect 1493 5432 1542 5444
rect 1813 5460 1862 5470
rect 1813 5440 1824 5460
rect 1844 5440 1862 5460
rect 1813 5428 1862 5440
rect 1912 5464 1956 5470
rect 1912 5444 1927 5464
rect 1947 5444 1956 5464
rect 1912 5428 1956 5444
rect 2026 5460 2075 5470
rect 2026 5440 2037 5460
rect 2057 5440 2075 5460
rect 2026 5428 2075 5440
rect 2125 5464 2169 5470
rect 2125 5444 2140 5464
rect 2160 5444 2169 5464
rect 2125 5428 2169 5444
rect 2234 5460 2283 5470
rect 2234 5440 2245 5460
rect 2265 5440 2283 5460
rect 2234 5428 2283 5440
rect 2333 5464 2377 5470
rect 2333 5444 2348 5464
rect 2368 5444 2377 5464
rect 2333 5428 2377 5444
rect 2447 5464 2491 5470
rect 2447 5444 2456 5464
rect 2476 5444 2491 5464
rect 2447 5428 2491 5444
rect 2541 5460 2590 5470
rect 2541 5440 2559 5460
rect 2579 5440 2590 5460
rect 2541 5428 2590 5440
rect 765 4785 814 4795
rect 765 4765 776 4785
rect 796 4765 814 4785
rect 765 4753 814 4765
rect 864 4789 908 4795
rect 864 4769 879 4789
rect 899 4769 908 4789
rect 864 4753 908 4769
rect 978 4785 1027 4795
rect 978 4765 989 4785
rect 1009 4765 1027 4785
rect 978 4753 1027 4765
rect 1077 4789 1121 4795
rect 1077 4769 1092 4789
rect 1112 4769 1121 4789
rect 1077 4753 1121 4769
rect 1186 4785 1235 4795
rect 1186 4765 1197 4785
rect 1217 4765 1235 4785
rect 1186 4753 1235 4765
rect 1285 4789 1329 4795
rect 1285 4769 1300 4789
rect 1320 4769 1329 4789
rect 1285 4753 1329 4769
rect 1399 4789 1443 4795
rect 1399 4769 1408 4789
rect 1428 4769 1443 4789
rect 1399 4753 1443 4769
rect 1493 4785 1542 4795
rect 1493 4765 1511 4785
rect 1531 4765 1542 4785
rect 1493 4753 1542 4765
rect 3260 4780 3309 4790
rect 3260 4760 3271 4780
rect 3291 4760 3309 4780
rect 3260 4748 3309 4760
rect 3359 4784 3403 4790
rect 3359 4764 3374 4784
rect 3394 4764 3403 4784
rect 3359 4748 3403 4764
rect 3473 4780 3522 4790
rect 3473 4760 3484 4780
rect 3504 4760 3522 4780
rect 3473 4748 3522 4760
rect 3572 4784 3616 4790
rect 3572 4764 3587 4784
rect 3607 4764 3616 4784
rect 3572 4748 3616 4764
rect 3681 4780 3730 4790
rect 3681 4760 3692 4780
rect 3712 4760 3730 4780
rect 3681 4748 3730 4760
rect 3780 4784 3824 4790
rect 3780 4764 3795 4784
rect 3815 4764 3824 4784
rect 3780 4748 3824 4764
rect 3894 4784 3938 4790
rect 3894 4764 3903 4784
rect 3923 4764 3938 4784
rect 3894 4748 3938 4764
rect 3988 4780 4037 4790
rect 3988 4760 4006 4780
rect 4026 4760 4037 4780
rect 3988 4748 4037 4760
rect 765 4017 814 4027
rect 765 3997 776 4017
rect 796 3997 814 4017
rect 765 3985 814 3997
rect 864 4021 908 4027
rect 864 4001 879 4021
rect 899 4001 908 4021
rect 864 3985 908 4001
rect 978 4017 1027 4027
rect 978 3997 989 4017
rect 1009 3997 1027 4017
rect 978 3985 1027 3997
rect 1077 4021 1121 4027
rect 1077 4001 1092 4021
rect 1112 4001 1121 4021
rect 1077 3985 1121 4001
rect 1186 4017 1235 4027
rect 1186 3997 1197 4017
rect 1217 3997 1235 4017
rect 1186 3985 1235 3997
rect 1285 4021 1329 4027
rect 1285 4001 1300 4021
rect 1320 4001 1329 4021
rect 1285 3985 1329 4001
rect 1399 4021 1443 4027
rect 1399 4001 1408 4021
rect 1428 4001 1443 4021
rect 1399 3985 1443 4001
rect 1493 4017 1542 4027
rect 1493 3997 1511 4017
rect 1531 3997 1542 4017
rect 1493 3985 1542 3997
rect 1813 4013 1862 4023
rect 1813 3993 1824 4013
rect 1844 3993 1862 4013
rect 1813 3981 1862 3993
rect 1912 4017 1956 4023
rect 1912 3997 1927 4017
rect 1947 3997 1956 4017
rect 1912 3981 1956 3997
rect 2026 4013 2075 4023
rect 2026 3993 2037 4013
rect 2057 3993 2075 4013
rect 2026 3981 2075 3993
rect 2125 4017 2169 4023
rect 2125 3997 2140 4017
rect 2160 3997 2169 4017
rect 2125 3981 2169 3997
rect 2234 4013 2283 4023
rect 2234 3993 2245 4013
rect 2265 3993 2283 4013
rect 2234 3981 2283 3993
rect 2333 4017 2377 4023
rect 2333 3997 2348 4017
rect 2368 3997 2377 4017
rect 2333 3981 2377 3997
rect 2447 4017 2491 4023
rect 2447 3997 2456 4017
rect 2476 3997 2491 4017
rect 2447 3981 2491 3997
rect 2541 4013 2590 4023
rect 2541 3993 2559 4013
rect 2579 3993 2590 4013
rect 2541 3981 2590 3993
rect 765 3338 814 3348
rect 765 3318 776 3338
rect 796 3318 814 3338
rect 765 3306 814 3318
rect 864 3342 908 3348
rect 864 3322 879 3342
rect 899 3322 908 3342
rect 864 3306 908 3322
rect 978 3338 1027 3348
rect 978 3318 989 3338
rect 1009 3318 1027 3338
rect 978 3306 1027 3318
rect 1077 3342 1121 3348
rect 1077 3322 1092 3342
rect 1112 3322 1121 3342
rect 1077 3306 1121 3322
rect 1186 3338 1235 3348
rect 1186 3318 1197 3338
rect 1217 3318 1235 3338
rect 1186 3306 1235 3318
rect 1285 3342 1329 3348
rect 1285 3322 1300 3342
rect 1320 3322 1329 3342
rect 1285 3306 1329 3322
rect 1399 3342 1443 3348
rect 1399 3322 1408 3342
rect 1428 3322 1443 3342
rect 1399 3306 1443 3322
rect 1493 3338 1542 3348
rect 1493 3318 1511 3338
rect 1531 3318 1542 3338
rect 1493 3306 1542 3318
rect 3303 3335 3352 3345
rect 3303 3315 3314 3335
rect 3334 3315 3352 3335
rect 3303 3303 3352 3315
rect 3402 3339 3446 3345
rect 3402 3319 3417 3339
rect 3437 3319 3446 3339
rect 3402 3303 3446 3319
rect 3516 3335 3565 3345
rect 3516 3315 3527 3335
rect 3547 3315 3565 3335
rect 3516 3303 3565 3315
rect 3615 3339 3659 3345
rect 3615 3319 3630 3339
rect 3650 3319 3659 3339
rect 3615 3303 3659 3319
rect 3724 3335 3773 3345
rect 3724 3315 3735 3335
rect 3755 3315 3773 3335
rect 3724 3303 3773 3315
rect 3823 3339 3867 3345
rect 3823 3319 3838 3339
rect 3858 3319 3867 3339
rect 3823 3303 3867 3319
rect 3937 3339 3981 3345
rect 3937 3319 3946 3339
rect 3966 3319 3981 3339
rect 3937 3303 3981 3319
rect 4031 3335 4080 3345
rect 4031 3315 4049 3335
rect 4069 3315 4080 3335
rect 4031 3303 4080 3315
rect 766 2497 815 2507
rect 766 2477 777 2497
rect 797 2477 815 2497
rect 766 2465 815 2477
rect 865 2501 909 2507
rect 865 2481 880 2501
rect 900 2481 909 2501
rect 865 2465 909 2481
rect 979 2497 1028 2507
rect 979 2477 990 2497
rect 1010 2477 1028 2497
rect 979 2465 1028 2477
rect 1078 2501 1122 2507
rect 1078 2481 1093 2501
rect 1113 2481 1122 2501
rect 1078 2465 1122 2481
rect 1187 2497 1236 2507
rect 1187 2477 1198 2497
rect 1218 2477 1236 2497
rect 1187 2465 1236 2477
rect 1286 2501 1330 2507
rect 1286 2481 1301 2501
rect 1321 2481 1330 2501
rect 1286 2465 1330 2481
rect 1400 2501 1444 2507
rect 1400 2481 1409 2501
rect 1429 2481 1444 2501
rect 1400 2465 1444 2481
rect 1494 2497 1543 2507
rect 1494 2477 1512 2497
rect 1532 2477 1543 2497
rect 1494 2465 1543 2477
rect 1814 2493 1863 2503
rect 1814 2473 1825 2493
rect 1845 2473 1863 2493
rect 1814 2461 1863 2473
rect 1913 2497 1957 2503
rect 1913 2477 1928 2497
rect 1948 2477 1957 2497
rect 1913 2461 1957 2477
rect 2027 2493 2076 2503
rect 2027 2473 2038 2493
rect 2058 2473 2076 2493
rect 2027 2461 2076 2473
rect 2126 2497 2170 2503
rect 2126 2477 2141 2497
rect 2161 2477 2170 2497
rect 2126 2461 2170 2477
rect 2235 2493 2284 2503
rect 2235 2473 2246 2493
rect 2266 2473 2284 2493
rect 2235 2461 2284 2473
rect 2334 2497 2378 2503
rect 2334 2477 2349 2497
rect 2369 2477 2378 2497
rect 2334 2461 2378 2477
rect 2448 2497 2492 2503
rect 2448 2477 2457 2497
rect 2477 2477 2492 2497
rect 2448 2461 2492 2477
rect 2542 2493 2591 2503
rect 2542 2473 2560 2493
rect 2580 2473 2591 2493
rect 2542 2461 2591 2473
rect 766 1818 815 1828
rect 766 1798 777 1818
rect 797 1798 815 1818
rect 766 1786 815 1798
rect 865 1822 909 1828
rect 865 1802 880 1822
rect 900 1802 909 1822
rect 865 1786 909 1802
rect 979 1818 1028 1828
rect 979 1798 990 1818
rect 1010 1798 1028 1818
rect 979 1786 1028 1798
rect 1078 1822 1122 1828
rect 1078 1802 1093 1822
rect 1113 1802 1122 1822
rect 1078 1786 1122 1802
rect 1187 1818 1236 1828
rect 1187 1798 1198 1818
rect 1218 1798 1236 1818
rect 1187 1786 1236 1798
rect 1286 1822 1330 1828
rect 1286 1802 1301 1822
rect 1321 1802 1330 1822
rect 1286 1786 1330 1802
rect 1400 1822 1444 1828
rect 1400 1802 1409 1822
rect 1429 1802 1444 1822
rect 1400 1786 1444 1802
rect 1494 1818 1543 1828
rect 1494 1798 1512 1818
rect 1532 1798 1543 1818
rect 1494 1786 1543 1798
rect 3261 1813 3310 1823
rect 3261 1793 3272 1813
rect 3292 1793 3310 1813
rect 3261 1781 3310 1793
rect 3360 1817 3404 1823
rect 3360 1797 3375 1817
rect 3395 1797 3404 1817
rect 3360 1781 3404 1797
rect 3474 1813 3523 1823
rect 3474 1793 3485 1813
rect 3505 1793 3523 1813
rect 3474 1781 3523 1793
rect 3573 1817 3617 1823
rect 3573 1797 3588 1817
rect 3608 1797 3617 1817
rect 3573 1781 3617 1797
rect 3682 1813 3731 1823
rect 3682 1793 3693 1813
rect 3713 1793 3731 1813
rect 3682 1781 3731 1793
rect 3781 1817 3825 1823
rect 3781 1797 3796 1817
rect 3816 1797 3825 1817
rect 3781 1781 3825 1797
rect 3895 1817 3939 1823
rect 3895 1797 3904 1817
rect 3924 1797 3939 1817
rect 3895 1781 3939 1797
rect 3989 1813 4038 1823
rect 3989 1793 4007 1813
rect 4027 1793 4038 1813
rect 3989 1781 4038 1793
rect 766 1050 815 1060
rect 766 1030 777 1050
rect 797 1030 815 1050
rect 766 1018 815 1030
rect 865 1054 909 1060
rect 865 1034 880 1054
rect 900 1034 909 1054
rect 865 1018 909 1034
rect 979 1050 1028 1060
rect 979 1030 990 1050
rect 1010 1030 1028 1050
rect 979 1018 1028 1030
rect 1078 1054 1122 1060
rect 1078 1034 1093 1054
rect 1113 1034 1122 1054
rect 1078 1018 1122 1034
rect 1187 1050 1236 1060
rect 1187 1030 1198 1050
rect 1218 1030 1236 1050
rect 1187 1018 1236 1030
rect 1286 1054 1330 1060
rect 1286 1034 1301 1054
rect 1321 1034 1330 1054
rect 1286 1018 1330 1034
rect 1400 1054 1444 1060
rect 1400 1034 1409 1054
rect 1429 1034 1444 1054
rect 1400 1018 1444 1034
rect 1494 1050 1543 1060
rect 1494 1030 1512 1050
rect 1532 1030 1543 1050
rect 1494 1018 1543 1030
rect 1814 1046 1863 1056
rect 1814 1026 1825 1046
rect 1845 1026 1863 1046
rect 1814 1014 1863 1026
rect 1913 1050 1957 1056
rect 1913 1030 1928 1050
rect 1948 1030 1957 1050
rect 1913 1014 1957 1030
rect 2027 1046 2076 1056
rect 2027 1026 2038 1046
rect 2058 1026 2076 1046
rect 2027 1014 2076 1026
rect 2126 1050 2170 1056
rect 2126 1030 2141 1050
rect 2161 1030 2170 1050
rect 2126 1014 2170 1030
rect 2235 1046 2284 1056
rect 2235 1026 2246 1046
rect 2266 1026 2284 1046
rect 2235 1014 2284 1026
rect 2334 1050 2378 1056
rect 2334 1030 2349 1050
rect 2369 1030 2378 1050
rect 2334 1014 2378 1030
rect 2448 1050 2492 1056
rect 2448 1030 2457 1050
rect 2477 1030 2492 1050
rect 2448 1014 2492 1030
rect 2542 1046 2591 1056
rect 2542 1026 2560 1046
rect 2580 1026 2591 1046
rect 2542 1014 2591 1026
rect 766 371 815 381
rect 766 351 777 371
rect 797 351 815 371
rect 766 339 815 351
rect 865 375 909 381
rect 865 355 880 375
rect 900 355 909 375
rect 865 339 909 355
rect 979 371 1028 381
rect 979 351 990 371
rect 1010 351 1028 371
rect 979 339 1028 351
rect 1078 375 1122 381
rect 1078 355 1093 375
rect 1113 355 1122 375
rect 1078 339 1122 355
rect 1187 371 1236 381
rect 1187 351 1198 371
rect 1218 351 1236 371
rect 1187 339 1236 351
rect 1286 375 1330 381
rect 1286 355 1301 375
rect 1321 355 1330 375
rect 1286 339 1330 355
rect 1400 375 1444 381
rect 1400 355 1409 375
rect 1429 355 1444 375
rect 1400 339 1444 355
rect 1494 371 1543 381
rect 1494 351 1512 371
rect 1532 351 1543 371
rect 1494 339 1543 351
<< pdiff >>
rect 772 11621 816 11659
rect 772 11601 784 11621
rect 804 11601 816 11621
rect 772 11559 816 11601
rect 866 11621 908 11659
rect 866 11601 880 11621
rect 900 11601 908 11621
rect 866 11559 908 11601
rect 985 11621 1029 11659
rect 985 11601 997 11621
rect 1017 11601 1029 11621
rect 985 11559 1029 11601
rect 1079 11621 1121 11659
rect 1079 11601 1093 11621
rect 1113 11601 1121 11621
rect 1079 11559 1121 11601
rect 1193 11621 1237 11659
rect 1193 11601 1205 11621
rect 1225 11601 1237 11621
rect 1193 11559 1237 11601
rect 1287 11621 1329 11659
rect 1287 11601 1301 11621
rect 1321 11601 1329 11621
rect 1287 11559 1329 11601
rect 1403 11621 1445 11659
rect 1403 11601 1411 11621
rect 1431 11601 1445 11621
rect 1403 11559 1445 11601
rect 1495 11628 1540 11659
rect 1495 11621 1539 11628
rect 1495 11601 1507 11621
rect 1527 11601 1539 11621
rect 1495 11559 1539 11601
rect 1820 11617 1864 11655
rect 1820 11597 1832 11617
rect 1852 11597 1864 11617
rect 1820 11555 1864 11597
rect 1914 11617 1956 11655
rect 1914 11597 1928 11617
rect 1948 11597 1956 11617
rect 1914 11555 1956 11597
rect 2033 11617 2077 11655
rect 2033 11597 2045 11617
rect 2065 11597 2077 11617
rect 2033 11555 2077 11597
rect 2127 11617 2169 11655
rect 2127 11597 2141 11617
rect 2161 11597 2169 11617
rect 2127 11555 2169 11597
rect 2241 11617 2285 11655
rect 2241 11597 2253 11617
rect 2273 11597 2285 11617
rect 2241 11555 2285 11597
rect 2335 11617 2377 11655
rect 2335 11597 2349 11617
rect 2369 11597 2377 11617
rect 2335 11555 2377 11597
rect 2451 11617 2493 11655
rect 2451 11597 2459 11617
rect 2479 11597 2493 11617
rect 2451 11555 2493 11597
rect 2543 11624 2588 11655
rect 2543 11617 2587 11624
rect 2543 11597 2555 11617
rect 2575 11597 2587 11617
rect 2543 11555 2587 11597
rect 772 10942 816 10980
rect 772 10922 784 10942
rect 804 10922 816 10942
rect 772 10880 816 10922
rect 866 10942 908 10980
rect 866 10922 880 10942
rect 900 10922 908 10942
rect 866 10880 908 10922
rect 985 10942 1029 10980
rect 985 10922 997 10942
rect 1017 10922 1029 10942
rect 985 10880 1029 10922
rect 1079 10942 1121 10980
rect 1079 10922 1093 10942
rect 1113 10922 1121 10942
rect 1079 10880 1121 10922
rect 1193 10942 1237 10980
rect 1193 10922 1205 10942
rect 1225 10922 1237 10942
rect 1193 10880 1237 10922
rect 1287 10942 1329 10980
rect 1287 10922 1301 10942
rect 1321 10922 1329 10942
rect 1287 10880 1329 10922
rect 1403 10942 1445 10980
rect 1403 10922 1411 10942
rect 1431 10922 1445 10942
rect 1403 10880 1445 10922
rect 1495 10949 1540 10980
rect 1495 10942 1539 10949
rect 1495 10922 1507 10942
rect 1527 10922 1539 10942
rect 1495 10880 1539 10922
rect 3267 10937 3311 10975
rect 3267 10917 3279 10937
rect 3299 10917 3311 10937
rect 3267 10875 3311 10917
rect 3361 10937 3403 10975
rect 3361 10917 3375 10937
rect 3395 10917 3403 10937
rect 3361 10875 3403 10917
rect 3480 10937 3524 10975
rect 3480 10917 3492 10937
rect 3512 10917 3524 10937
rect 3480 10875 3524 10917
rect 3574 10937 3616 10975
rect 3574 10917 3588 10937
rect 3608 10917 3616 10937
rect 3574 10875 3616 10917
rect 3688 10937 3732 10975
rect 3688 10917 3700 10937
rect 3720 10917 3732 10937
rect 3688 10875 3732 10917
rect 3782 10937 3824 10975
rect 3782 10917 3796 10937
rect 3816 10917 3824 10937
rect 3782 10875 3824 10917
rect 3898 10937 3940 10975
rect 3898 10917 3906 10937
rect 3926 10917 3940 10937
rect 3898 10875 3940 10917
rect 3990 10944 4035 10975
rect 3990 10937 4034 10944
rect 3990 10917 4002 10937
rect 4022 10917 4034 10937
rect 3990 10875 4034 10917
rect 772 10174 816 10212
rect 772 10154 784 10174
rect 804 10154 816 10174
rect 772 10112 816 10154
rect 866 10174 908 10212
rect 866 10154 880 10174
rect 900 10154 908 10174
rect 866 10112 908 10154
rect 985 10174 1029 10212
rect 985 10154 997 10174
rect 1017 10154 1029 10174
rect 985 10112 1029 10154
rect 1079 10174 1121 10212
rect 1079 10154 1093 10174
rect 1113 10154 1121 10174
rect 1079 10112 1121 10154
rect 1193 10174 1237 10212
rect 1193 10154 1205 10174
rect 1225 10154 1237 10174
rect 1193 10112 1237 10154
rect 1287 10174 1329 10212
rect 1287 10154 1301 10174
rect 1321 10154 1329 10174
rect 1287 10112 1329 10154
rect 1403 10174 1445 10212
rect 1403 10154 1411 10174
rect 1431 10154 1445 10174
rect 1403 10112 1445 10154
rect 1495 10181 1540 10212
rect 1495 10174 1539 10181
rect 1495 10154 1507 10174
rect 1527 10154 1539 10174
rect 1495 10112 1539 10154
rect 1820 10170 1864 10208
rect 1820 10150 1832 10170
rect 1852 10150 1864 10170
rect 1820 10108 1864 10150
rect 1914 10170 1956 10208
rect 1914 10150 1928 10170
rect 1948 10150 1956 10170
rect 1914 10108 1956 10150
rect 2033 10170 2077 10208
rect 2033 10150 2045 10170
rect 2065 10150 2077 10170
rect 2033 10108 2077 10150
rect 2127 10170 2169 10208
rect 2127 10150 2141 10170
rect 2161 10150 2169 10170
rect 2127 10108 2169 10150
rect 2241 10170 2285 10208
rect 2241 10150 2253 10170
rect 2273 10150 2285 10170
rect 2241 10108 2285 10150
rect 2335 10170 2377 10208
rect 2335 10150 2349 10170
rect 2369 10150 2377 10170
rect 2335 10108 2377 10150
rect 2451 10170 2493 10208
rect 2451 10150 2459 10170
rect 2479 10150 2493 10170
rect 2451 10108 2493 10150
rect 2543 10177 2588 10208
rect 2543 10170 2587 10177
rect 2543 10150 2555 10170
rect 2575 10150 2587 10170
rect 2543 10108 2587 10150
rect 772 9495 816 9533
rect 772 9475 784 9495
rect 804 9475 816 9495
rect 772 9433 816 9475
rect 866 9495 908 9533
rect 866 9475 880 9495
rect 900 9475 908 9495
rect 866 9433 908 9475
rect 985 9495 1029 9533
rect 985 9475 997 9495
rect 1017 9475 1029 9495
rect 985 9433 1029 9475
rect 1079 9495 1121 9533
rect 1079 9475 1093 9495
rect 1113 9475 1121 9495
rect 1079 9433 1121 9475
rect 1193 9495 1237 9533
rect 1193 9475 1205 9495
rect 1225 9475 1237 9495
rect 1193 9433 1237 9475
rect 1287 9495 1329 9533
rect 1287 9475 1301 9495
rect 1321 9475 1329 9495
rect 1287 9433 1329 9475
rect 1403 9495 1445 9533
rect 1403 9475 1411 9495
rect 1431 9475 1445 9495
rect 1403 9433 1445 9475
rect 1495 9502 1540 9533
rect 1495 9495 1539 9502
rect 1495 9475 1507 9495
rect 1527 9475 1539 9495
rect 1495 9433 1539 9475
rect 3310 9492 3354 9530
rect 3310 9472 3322 9492
rect 3342 9472 3354 9492
rect 3310 9430 3354 9472
rect 3404 9492 3446 9530
rect 3404 9472 3418 9492
rect 3438 9472 3446 9492
rect 3404 9430 3446 9472
rect 3523 9492 3567 9530
rect 3523 9472 3535 9492
rect 3555 9472 3567 9492
rect 3523 9430 3567 9472
rect 3617 9492 3659 9530
rect 3617 9472 3631 9492
rect 3651 9472 3659 9492
rect 3617 9430 3659 9472
rect 3731 9492 3775 9530
rect 3731 9472 3743 9492
rect 3763 9472 3775 9492
rect 3731 9430 3775 9472
rect 3825 9492 3867 9530
rect 3825 9472 3839 9492
rect 3859 9472 3867 9492
rect 3825 9430 3867 9472
rect 3941 9492 3983 9530
rect 3941 9472 3949 9492
rect 3969 9472 3983 9492
rect 3941 9430 3983 9472
rect 4033 9499 4078 9530
rect 4033 9492 4077 9499
rect 4033 9472 4045 9492
rect 4065 9472 4077 9492
rect 4033 9430 4077 9472
rect 773 8654 817 8692
rect 773 8634 785 8654
rect 805 8634 817 8654
rect 773 8592 817 8634
rect 867 8654 909 8692
rect 867 8634 881 8654
rect 901 8634 909 8654
rect 867 8592 909 8634
rect 986 8654 1030 8692
rect 986 8634 998 8654
rect 1018 8634 1030 8654
rect 986 8592 1030 8634
rect 1080 8654 1122 8692
rect 1080 8634 1094 8654
rect 1114 8634 1122 8654
rect 1080 8592 1122 8634
rect 1194 8654 1238 8692
rect 1194 8634 1206 8654
rect 1226 8634 1238 8654
rect 1194 8592 1238 8634
rect 1288 8654 1330 8692
rect 1288 8634 1302 8654
rect 1322 8634 1330 8654
rect 1288 8592 1330 8634
rect 1404 8654 1446 8692
rect 1404 8634 1412 8654
rect 1432 8634 1446 8654
rect 1404 8592 1446 8634
rect 1496 8661 1541 8692
rect 1496 8654 1540 8661
rect 1496 8634 1508 8654
rect 1528 8634 1540 8654
rect 1496 8592 1540 8634
rect 1821 8650 1865 8688
rect 1821 8630 1833 8650
rect 1853 8630 1865 8650
rect 1821 8588 1865 8630
rect 1915 8650 1957 8688
rect 1915 8630 1929 8650
rect 1949 8630 1957 8650
rect 1915 8588 1957 8630
rect 2034 8650 2078 8688
rect 2034 8630 2046 8650
rect 2066 8630 2078 8650
rect 2034 8588 2078 8630
rect 2128 8650 2170 8688
rect 2128 8630 2142 8650
rect 2162 8630 2170 8650
rect 2128 8588 2170 8630
rect 2242 8650 2286 8688
rect 2242 8630 2254 8650
rect 2274 8630 2286 8650
rect 2242 8588 2286 8630
rect 2336 8650 2378 8688
rect 2336 8630 2350 8650
rect 2370 8630 2378 8650
rect 2336 8588 2378 8630
rect 2452 8650 2494 8688
rect 2452 8630 2460 8650
rect 2480 8630 2494 8650
rect 2452 8588 2494 8630
rect 2544 8657 2589 8688
rect 2544 8650 2588 8657
rect 2544 8630 2556 8650
rect 2576 8630 2588 8650
rect 2544 8588 2588 8630
rect 773 7975 817 8013
rect 773 7955 785 7975
rect 805 7955 817 7975
rect 773 7913 817 7955
rect 867 7975 909 8013
rect 867 7955 881 7975
rect 901 7955 909 7975
rect 867 7913 909 7955
rect 986 7975 1030 8013
rect 986 7955 998 7975
rect 1018 7955 1030 7975
rect 986 7913 1030 7955
rect 1080 7975 1122 8013
rect 1080 7955 1094 7975
rect 1114 7955 1122 7975
rect 1080 7913 1122 7955
rect 1194 7975 1238 8013
rect 1194 7955 1206 7975
rect 1226 7955 1238 7975
rect 1194 7913 1238 7955
rect 1288 7975 1330 8013
rect 1288 7955 1302 7975
rect 1322 7955 1330 7975
rect 1288 7913 1330 7955
rect 1404 7975 1446 8013
rect 1404 7955 1412 7975
rect 1432 7955 1446 7975
rect 1404 7913 1446 7955
rect 1496 7982 1541 8013
rect 1496 7975 1540 7982
rect 1496 7955 1508 7975
rect 1528 7955 1540 7975
rect 1496 7913 1540 7955
rect 3268 7970 3312 8008
rect 3268 7950 3280 7970
rect 3300 7950 3312 7970
rect 3268 7908 3312 7950
rect 3362 7970 3404 8008
rect 3362 7950 3376 7970
rect 3396 7950 3404 7970
rect 3362 7908 3404 7950
rect 3481 7970 3525 8008
rect 3481 7950 3493 7970
rect 3513 7950 3525 7970
rect 3481 7908 3525 7950
rect 3575 7970 3617 8008
rect 3575 7950 3589 7970
rect 3609 7950 3617 7970
rect 3575 7908 3617 7950
rect 3689 7970 3733 8008
rect 3689 7950 3701 7970
rect 3721 7950 3733 7970
rect 3689 7908 3733 7950
rect 3783 7970 3825 8008
rect 3783 7950 3797 7970
rect 3817 7950 3825 7970
rect 3783 7908 3825 7950
rect 3899 7970 3941 8008
rect 3899 7950 3907 7970
rect 3927 7950 3941 7970
rect 3899 7908 3941 7950
rect 3991 7977 4036 8008
rect 3991 7970 4035 7977
rect 3991 7950 4003 7970
rect 4023 7950 4035 7970
rect 3991 7908 4035 7950
rect 773 7207 817 7245
rect 773 7187 785 7207
rect 805 7187 817 7207
rect 773 7145 817 7187
rect 867 7207 909 7245
rect 867 7187 881 7207
rect 901 7187 909 7207
rect 867 7145 909 7187
rect 986 7207 1030 7245
rect 986 7187 998 7207
rect 1018 7187 1030 7207
rect 986 7145 1030 7187
rect 1080 7207 1122 7245
rect 1080 7187 1094 7207
rect 1114 7187 1122 7207
rect 1080 7145 1122 7187
rect 1194 7207 1238 7245
rect 1194 7187 1206 7207
rect 1226 7187 1238 7207
rect 1194 7145 1238 7187
rect 1288 7207 1330 7245
rect 1288 7187 1302 7207
rect 1322 7187 1330 7207
rect 1288 7145 1330 7187
rect 1404 7207 1446 7245
rect 1404 7187 1412 7207
rect 1432 7187 1446 7207
rect 1404 7145 1446 7187
rect 1496 7214 1541 7245
rect 1496 7207 1540 7214
rect 1496 7187 1508 7207
rect 1528 7187 1540 7207
rect 1496 7145 1540 7187
rect 1821 7203 1865 7241
rect 1821 7183 1833 7203
rect 1853 7183 1865 7203
rect 1821 7141 1865 7183
rect 1915 7203 1957 7241
rect 1915 7183 1929 7203
rect 1949 7183 1957 7203
rect 1915 7141 1957 7183
rect 2034 7203 2078 7241
rect 2034 7183 2046 7203
rect 2066 7183 2078 7203
rect 2034 7141 2078 7183
rect 2128 7203 2170 7241
rect 2128 7183 2142 7203
rect 2162 7183 2170 7203
rect 2128 7141 2170 7183
rect 2242 7203 2286 7241
rect 2242 7183 2254 7203
rect 2274 7183 2286 7203
rect 2242 7141 2286 7183
rect 2336 7203 2378 7241
rect 2336 7183 2350 7203
rect 2370 7183 2378 7203
rect 2336 7141 2378 7183
rect 2452 7203 2494 7241
rect 2452 7183 2460 7203
rect 2480 7183 2494 7203
rect 2452 7141 2494 7183
rect 2544 7210 2589 7241
rect 2544 7203 2588 7210
rect 2544 7183 2556 7203
rect 2576 7183 2588 7203
rect 2544 7141 2588 7183
rect 773 6528 817 6566
rect 773 6508 785 6528
rect 805 6508 817 6528
rect 773 6466 817 6508
rect 867 6528 909 6566
rect 867 6508 881 6528
rect 901 6508 909 6528
rect 867 6466 909 6508
rect 986 6528 1030 6566
rect 986 6508 998 6528
rect 1018 6508 1030 6528
rect 986 6466 1030 6508
rect 1080 6528 1122 6566
rect 1080 6508 1094 6528
rect 1114 6508 1122 6528
rect 1080 6466 1122 6508
rect 1194 6528 1238 6566
rect 1194 6508 1206 6528
rect 1226 6508 1238 6528
rect 1194 6466 1238 6508
rect 1288 6528 1330 6566
rect 1288 6508 1302 6528
rect 1322 6508 1330 6528
rect 1288 6466 1330 6508
rect 1404 6528 1446 6566
rect 1404 6508 1412 6528
rect 1432 6508 1446 6528
rect 1404 6466 1446 6508
rect 1496 6535 1541 6566
rect 1496 6528 1540 6535
rect 1496 6508 1508 6528
rect 1528 6508 1540 6528
rect 1496 6466 1540 6508
rect 4376 6519 4420 6557
rect 4376 6499 4388 6519
rect 4408 6499 4420 6519
rect 4376 6457 4420 6499
rect 4470 6519 4512 6557
rect 4470 6499 4484 6519
rect 4504 6499 4512 6519
rect 4470 6457 4512 6499
rect 4589 6519 4633 6557
rect 4589 6499 4601 6519
rect 4621 6499 4633 6519
rect 4589 6457 4633 6499
rect 4683 6519 4725 6557
rect 4683 6499 4697 6519
rect 4717 6499 4725 6519
rect 4683 6457 4725 6499
rect 4797 6519 4841 6557
rect 4797 6499 4809 6519
rect 4829 6499 4841 6519
rect 4797 6457 4841 6499
rect 4891 6519 4933 6557
rect 4891 6499 4905 6519
rect 4925 6499 4933 6519
rect 4891 6457 4933 6499
rect 5007 6519 5049 6557
rect 5007 6499 5015 6519
rect 5035 6499 5049 6519
rect 5007 6457 5049 6499
rect 5099 6526 5144 6557
rect 5099 6519 5143 6526
rect 5099 6499 5111 6519
rect 5131 6499 5143 6519
rect 5099 6457 5143 6499
rect 770 5613 814 5651
rect 770 5593 782 5613
rect 802 5593 814 5613
rect 770 5551 814 5593
rect 864 5613 906 5651
rect 864 5593 878 5613
rect 898 5593 906 5613
rect 864 5551 906 5593
rect 983 5613 1027 5651
rect 983 5593 995 5613
rect 1015 5593 1027 5613
rect 983 5551 1027 5593
rect 1077 5613 1119 5651
rect 1077 5593 1091 5613
rect 1111 5593 1119 5613
rect 1077 5551 1119 5593
rect 1191 5613 1235 5651
rect 1191 5593 1203 5613
rect 1223 5593 1235 5613
rect 1191 5551 1235 5593
rect 1285 5613 1327 5651
rect 1285 5593 1299 5613
rect 1319 5593 1327 5613
rect 1285 5551 1327 5593
rect 1401 5613 1443 5651
rect 1401 5593 1409 5613
rect 1429 5593 1443 5613
rect 1401 5551 1443 5593
rect 1493 5620 1538 5651
rect 1493 5613 1537 5620
rect 1493 5593 1505 5613
rect 1525 5593 1537 5613
rect 1493 5551 1537 5593
rect 1818 5609 1862 5647
rect 1818 5589 1830 5609
rect 1850 5589 1862 5609
rect 1818 5547 1862 5589
rect 1912 5609 1954 5647
rect 1912 5589 1926 5609
rect 1946 5589 1954 5609
rect 1912 5547 1954 5589
rect 2031 5609 2075 5647
rect 2031 5589 2043 5609
rect 2063 5589 2075 5609
rect 2031 5547 2075 5589
rect 2125 5609 2167 5647
rect 2125 5589 2139 5609
rect 2159 5589 2167 5609
rect 2125 5547 2167 5589
rect 2239 5609 2283 5647
rect 2239 5589 2251 5609
rect 2271 5589 2283 5609
rect 2239 5547 2283 5589
rect 2333 5609 2375 5647
rect 2333 5589 2347 5609
rect 2367 5589 2375 5609
rect 2333 5547 2375 5589
rect 2449 5609 2491 5647
rect 2449 5589 2457 5609
rect 2477 5589 2491 5609
rect 2449 5547 2491 5589
rect 2541 5616 2586 5647
rect 2541 5609 2585 5616
rect 2541 5589 2553 5609
rect 2573 5589 2585 5609
rect 2541 5547 2585 5589
rect 770 4934 814 4972
rect 770 4914 782 4934
rect 802 4914 814 4934
rect 770 4872 814 4914
rect 864 4934 906 4972
rect 864 4914 878 4934
rect 898 4914 906 4934
rect 864 4872 906 4914
rect 983 4934 1027 4972
rect 983 4914 995 4934
rect 1015 4914 1027 4934
rect 983 4872 1027 4914
rect 1077 4934 1119 4972
rect 1077 4914 1091 4934
rect 1111 4914 1119 4934
rect 1077 4872 1119 4914
rect 1191 4934 1235 4972
rect 1191 4914 1203 4934
rect 1223 4914 1235 4934
rect 1191 4872 1235 4914
rect 1285 4934 1327 4972
rect 1285 4914 1299 4934
rect 1319 4914 1327 4934
rect 1285 4872 1327 4914
rect 1401 4934 1443 4972
rect 1401 4914 1409 4934
rect 1429 4914 1443 4934
rect 1401 4872 1443 4914
rect 1493 4941 1538 4972
rect 1493 4934 1537 4941
rect 1493 4914 1505 4934
rect 1525 4914 1537 4934
rect 1493 4872 1537 4914
rect 3265 4929 3309 4967
rect 3265 4909 3277 4929
rect 3297 4909 3309 4929
rect 3265 4867 3309 4909
rect 3359 4929 3401 4967
rect 3359 4909 3373 4929
rect 3393 4909 3401 4929
rect 3359 4867 3401 4909
rect 3478 4929 3522 4967
rect 3478 4909 3490 4929
rect 3510 4909 3522 4929
rect 3478 4867 3522 4909
rect 3572 4929 3614 4967
rect 3572 4909 3586 4929
rect 3606 4909 3614 4929
rect 3572 4867 3614 4909
rect 3686 4929 3730 4967
rect 3686 4909 3698 4929
rect 3718 4909 3730 4929
rect 3686 4867 3730 4909
rect 3780 4929 3822 4967
rect 3780 4909 3794 4929
rect 3814 4909 3822 4929
rect 3780 4867 3822 4909
rect 3896 4929 3938 4967
rect 3896 4909 3904 4929
rect 3924 4909 3938 4929
rect 3896 4867 3938 4909
rect 3988 4936 4033 4967
rect 3988 4929 4032 4936
rect 3988 4909 4000 4929
rect 4020 4909 4032 4929
rect 3988 4867 4032 4909
rect 770 4166 814 4204
rect 770 4146 782 4166
rect 802 4146 814 4166
rect 770 4104 814 4146
rect 864 4166 906 4204
rect 864 4146 878 4166
rect 898 4146 906 4166
rect 864 4104 906 4146
rect 983 4166 1027 4204
rect 983 4146 995 4166
rect 1015 4146 1027 4166
rect 983 4104 1027 4146
rect 1077 4166 1119 4204
rect 1077 4146 1091 4166
rect 1111 4146 1119 4166
rect 1077 4104 1119 4146
rect 1191 4166 1235 4204
rect 1191 4146 1203 4166
rect 1223 4146 1235 4166
rect 1191 4104 1235 4146
rect 1285 4166 1327 4204
rect 1285 4146 1299 4166
rect 1319 4146 1327 4166
rect 1285 4104 1327 4146
rect 1401 4166 1443 4204
rect 1401 4146 1409 4166
rect 1429 4146 1443 4166
rect 1401 4104 1443 4146
rect 1493 4173 1538 4204
rect 1493 4166 1537 4173
rect 1493 4146 1505 4166
rect 1525 4146 1537 4166
rect 1493 4104 1537 4146
rect 1818 4162 1862 4200
rect 1818 4142 1830 4162
rect 1850 4142 1862 4162
rect 1818 4100 1862 4142
rect 1912 4162 1954 4200
rect 1912 4142 1926 4162
rect 1946 4142 1954 4162
rect 1912 4100 1954 4142
rect 2031 4162 2075 4200
rect 2031 4142 2043 4162
rect 2063 4142 2075 4162
rect 2031 4100 2075 4142
rect 2125 4162 2167 4200
rect 2125 4142 2139 4162
rect 2159 4142 2167 4162
rect 2125 4100 2167 4142
rect 2239 4162 2283 4200
rect 2239 4142 2251 4162
rect 2271 4142 2283 4162
rect 2239 4100 2283 4142
rect 2333 4162 2375 4200
rect 2333 4142 2347 4162
rect 2367 4142 2375 4162
rect 2333 4100 2375 4142
rect 2449 4162 2491 4200
rect 2449 4142 2457 4162
rect 2477 4142 2491 4162
rect 2449 4100 2491 4142
rect 2541 4169 2586 4200
rect 2541 4162 2585 4169
rect 2541 4142 2553 4162
rect 2573 4142 2585 4162
rect 2541 4100 2585 4142
rect 770 3487 814 3525
rect 770 3467 782 3487
rect 802 3467 814 3487
rect 770 3425 814 3467
rect 864 3487 906 3525
rect 864 3467 878 3487
rect 898 3467 906 3487
rect 864 3425 906 3467
rect 983 3487 1027 3525
rect 983 3467 995 3487
rect 1015 3467 1027 3487
rect 983 3425 1027 3467
rect 1077 3487 1119 3525
rect 1077 3467 1091 3487
rect 1111 3467 1119 3487
rect 1077 3425 1119 3467
rect 1191 3487 1235 3525
rect 1191 3467 1203 3487
rect 1223 3467 1235 3487
rect 1191 3425 1235 3467
rect 1285 3487 1327 3525
rect 1285 3467 1299 3487
rect 1319 3467 1327 3487
rect 1285 3425 1327 3467
rect 1401 3487 1443 3525
rect 1401 3467 1409 3487
rect 1429 3467 1443 3487
rect 1401 3425 1443 3467
rect 1493 3494 1538 3525
rect 1493 3487 1537 3494
rect 1493 3467 1505 3487
rect 1525 3467 1537 3487
rect 1493 3425 1537 3467
rect 3308 3484 3352 3522
rect 3308 3464 3320 3484
rect 3340 3464 3352 3484
rect 3308 3422 3352 3464
rect 3402 3484 3444 3522
rect 3402 3464 3416 3484
rect 3436 3464 3444 3484
rect 3402 3422 3444 3464
rect 3521 3484 3565 3522
rect 3521 3464 3533 3484
rect 3553 3464 3565 3484
rect 3521 3422 3565 3464
rect 3615 3484 3657 3522
rect 3615 3464 3629 3484
rect 3649 3464 3657 3484
rect 3615 3422 3657 3464
rect 3729 3484 3773 3522
rect 3729 3464 3741 3484
rect 3761 3464 3773 3484
rect 3729 3422 3773 3464
rect 3823 3484 3865 3522
rect 3823 3464 3837 3484
rect 3857 3464 3865 3484
rect 3823 3422 3865 3464
rect 3939 3484 3981 3522
rect 3939 3464 3947 3484
rect 3967 3464 3981 3484
rect 3939 3422 3981 3464
rect 4031 3491 4076 3522
rect 4031 3484 4075 3491
rect 4031 3464 4043 3484
rect 4063 3464 4075 3484
rect 4031 3422 4075 3464
rect 771 2646 815 2684
rect 771 2626 783 2646
rect 803 2626 815 2646
rect 771 2584 815 2626
rect 865 2646 907 2684
rect 865 2626 879 2646
rect 899 2626 907 2646
rect 865 2584 907 2626
rect 984 2646 1028 2684
rect 984 2626 996 2646
rect 1016 2626 1028 2646
rect 984 2584 1028 2626
rect 1078 2646 1120 2684
rect 1078 2626 1092 2646
rect 1112 2626 1120 2646
rect 1078 2584 1120 2626
rect 1192 2646 1236 2684
rect 1192 2626 1204 2646
rect 1224 2626 1236 2646
rect 1192 2584 1236 2626
rect 1286 2646 1328 2684
rect 1286 2626 1300 2646
rect 1320 2626 1328 2646
rect 1286 2584 1328 2626
rect 1402 2646 1444 2684
rect 1402 2626 1410 2646
rect 1430 2626 1444 2646
rect 1402 2584 1444 2626
rect 1494 2653 1539 2684
rect 1494 2646 1538 2653
rect 1494 2626 1506 2646
rect 1526 2626 1538 2646
rect 1494 2584 1538 2626
rect 1819 2642 1863 2680
rect 1819 2622 1831 2642
rect 1851 2622 1863 2642
rect 1819 2580 1863 2622
rect 1913 2642 1955 2680
rect 1913 2622 1927 2642
rect 1947 2622 1955 2642
rect 1913 2580 1955 2622
rect 2032 2642 2076 2680
rect 2032 2622 2044 2642
rect 2064 2622 2076 2642
rect 2032 2580 2076 2622
rect 2126 2642 2168 2680
rect 2126 2622 2140 2642
rect 2160 2622 2168 2642
rect 2126 2580 2168 2622
rect 2240 2642 2284 2680
rect 2240 2622 2252 2642
rect 2272 2622 2284 2642
rect 2240 2580 2284 2622
rect 2334 2642 2376 2680
rect 2334 2622 2348 2642
rect 2368 2622 2376 2642
rect 2334 2580 2376 2622
rect 2450 2642 2492 2680
rect 2450 2622 2458 2642
rect 2478 2622 2492 2642
rect 2450 2580 2492 2622
rect 2542 2649 2587 2680
rect 2542 2642 2586 2649
rect 2542 2622 2554 2642
rect 2574 2622 2586 2642
rect 2542 2580 2586 2622
rect 771 1967 815 2005
rect 771 1947 783 1967
rect 803 1947 815 1967
rect 771 1905 815 1947
rect 865 1967 907 2005
rect 865 1947 879 1967
rect 899 1947 907 1967
rect 865 1905 907 1947
rect 984 1967 1028 2005
rect 984 1947 996 1967
rect 1016 1947 1028 1967
rect 984 1905 1028 1947
rect 1078 1967 1120 2005
rect 1078 1947 1092 1967
rect 1112 1947 1120 1967
rect 1078 1905 1120 1947
rect 1192 1967 1236 2005
rect 1192 1947 1204 1967
rect 1224 1947 1236 1967
rect 1192 1905 1236 1947
rect 1286 1967 1328 2005
rect 1286 1947 1300 1967
rect 1320 1947 1328 1967
rect 1286 1905 1328 1947
rect 1402 1967 1444 2005
rect 1402 1947 1410 1967
rect 1430 1947 1444 1967
rect 1402 1905 1444 1947
rect 1494 1974 1539 2005
rect 1494 1967 1538 1974
rect 1494 1947 1506 1967
rect 1526 1947 1538 1967
rect 1494 1905 1538 1947
rect 3266 1962 3310 2000
rect 3266 1942 3278 1962
rect 3298 1942 3310 1962
rect 3266 1900 3310 1942
rect 3360 1962 3402 2000
rect 3360 1942 3374 1962
rect 3394 1942 3402 1962
rect 3360 1900 3402 1942
rect 3479 1962 3523 2000
rect 3479 1942 3491 1962
rect 3511 1942 3523 1962
rect 3479 1900 3523 1942
rect 3573 1962 3615 2000
rect 3573 1942 3587 1962
rect 3607 1942 3615 1962
rect 3573 1900 3615 1942
rect 3687 1962 3731 2000
rect 3687 1942 3699 1962
rect 3719 1942 3731 1962
rect 3687 1900 3731 1942
rect 3781 1962 3823 2000
rect 3781 1942 3795 1962
rect 3815 1942 3823 1962
rect 3781 1900 3823 1942
rect 3897 1962 3939 2000
rect 3897 1942 3905 1962
rect 3925 1942 3939 1962
rect 3897 1900 3939 1942
rect 3989 1969 4034 2000
rect 3989 1962 4033 1969
rect 3989 1942 4001 1962
rect 4021 1942 4033 1962
rect 3989 1900 4033 1942
rect 771 1199 815 1237
rect 771 1179 783 1199
rect 803 1179 815 1199
rect 771 1137 815 1179
rect 865 1199 907 1237
rect 865 1179 879 1199
rect 899 1179 907 1199
rect 865 1137 907 1179
rect 984 1199 1028 1237
rect 984 1179 996 1199
rect 1016 1179 1028 1199
rect 984 1137 1028 1179
rect 1078 1199 1120 1237
rect 1078 1179 1092 1199
rect 1112 1179 1120 1199
rect 1078 1137 1120 1179
rect 1192 1199 1236 1237
rect 1192 1179 1204 1199
rect 1224 1179 1236 1199
rect 1192 1137 1236 1179
rect 1286 1199 1328 1237
rect 1286 1179 1300 1199
rect 1320 1179 1328 1199
rect 1286 1137 1328 1179
rect 1402 1199 1444 1237
rect 1402 1179 1410 1199
rect 1430 1179 1444 1199
rect 1402 1137 1444 1179
rect 1494 1206 1539 1237
rect 1494 1199 1538 1206
rect 1494 1179 1506 1199
rect 1526 1179 1538 1199
rect 1494 1137 1538 1179
rect 1819 1195 1863 1233
rect 1819 1175 1831 1195
rect 1851 1175 1863 1195
rect 1819 1133 1863 1175
rect 1913 1195 1955 1233
rect 1913 1175 1927 1195
rect 1947 1175 1955 1195
rect 1913 1133 1955 1175
rect 2032 1195 2076 1233
rect 2032 1175 2044 1195
rect 2064 1175 2076 1195
rect 2032 1133 2076 1175
rect 2126 1195 2168 1233
rect 2126 1175 2140 1195
rect 2160 1175 2168 1195
rect 2126 1133 2168 1175
rect 2240 1195 2284 1233
rect 2240 1175 2252 1195
rect 2272 1175 2284 1195
rect 2240 1133 2284 1175
rect 2334 1195 2376 1233
rect 2334 1175 2348 1195
rect 2368 1175 2376 1195
rect 2334 1133 2376 1175
rect 2450 1195 2492 1233
rect 2450 1175 2458 1195
rect 2478 1175 2492 1195
rect 2450 1133 2492 1175
rect 2542 1202 2587 1233
rect 2542 1195 2586 1202
rect 2542 1175 2554 1195
rect 2574 1175 2586 1195
rect 2542 1133 2586 1175
rect 771 520 815 558
rect 771 500 783 520
rect 803 500 815 520
rect 771 458 815 500
rect 865 520 907 558
rect 865 500 879 520
rect 899 500 907 520
rect 865 458 907 500
rect 984 520 1028 558
rect 984 500 996 520
rect 1016 500 1028 520
rect 984 458 1028 500
rect 1078 520 1120 558
rect 1078 500 1092 520
rect 1112 500 1120 520
rect 1078 458 1120 500
rect 1192 520 1236 558
rect 1192 500 1204 520
rect 1224 500 1236 520
rect 1192 458 1236 500
rect 1286 520 1328 558
rect 1286 500 1300 520
rect 1320 500 1328 520
rect 1286 458 1328 500
rect 1402 520 1444 558
rect 1402 500 1410 520
rect 1430 500 1444 520
rect 1402 458 1444 500
rect 1494 527 1539 558
rect 1494 520 1538 527
rect 1494 500 1506 520
rect 1526 500 1538 520
rect 1494 458 1538 500
<< ndiffc >>
rect 458 11775 476 11793
rect 460 11676 478 11694
rect 458 11519 476 11537
rect 778 11452 798 11472
rect 881 11456 901 11476
rect 991 11452 1011 11472
rect 1094 11456 1114 11476
rect 1199 11452 1219 11472
rect 1302 11456 1322 11476
rect 1410 11456 1430 11476
rect 1513 11452 1533 11472
rect 1826 11448 1846 11468
rect 460 11420 478 11438
rect 1929 11452 1949 11472
rect 2039 11448 2059 11468
rect 2142 11452 2162 11472
rect 2247 11448 2267 11468
rect 2350 11452 2370 11472
rect 2458 11452 2478 11472
rect 2561 11448 2581 11468
rect 458 11124 476 11142
rect 460 11025 478 11043
rect 458 10869 476 10887
rect 460 10770 478 10788
rect 778 10773 798 10793
rect 881 10777 901 10797
rect 991 10773 1011 10793
rect 1094 10777 1114 10797
rect 1199 10773 1219 10793
rect 1302 10777 1322 10797
rect 1410 10777 1430 10797
rect 1513 10773 1533 10793
rect 3273 10768 3293 10788
rect 3376 10772 3396 10792
rect 3486 10768 3506 10788
rect 3589 10772 3609 10792
rect 3694 10768 3714 10788
rect 3797 10772 3817 10792
rect 3905 10772 3925 10792
rect 4008 10768 4028 10788
rect 458 10328 476 10346
rect 460 10229 478 10247
rect 458 10072 476 10090
rect 778 10005 798 10025
rect 881 10009 901 10029
rect 991 10005 1011 10025
rect 1094 10009 1114 10029
rect 1199 10005 1219 10025
rect 1302 10009 1322 10029
rect 1410 10009 1430 10029
rect 1513 10005 1533 10025
rect 1826 10001 1846 10021
rect 460 9973 478 9991
rect 1929 10005 1949 10025
rect 2039 10001 2059 10021
rect 2142 10005 2162 10025
rect 2247 10001 2267 10021
rect 2350 10005 2370 10025
rect 2458 10005 2478 10025
rect 2561 10001 2581 10021
rect 458 9677 476 9695
rect 460 9578 478 9596
rect 458 9422 476 9440
rect 460 9323 478 9341
rect 778 9326 798 9346
rect 881 9330 901 9350
rect 991 9326 1011 9346
rect 1094 9330 1114 9350
rect 1199 9326 1219 9346
rect 1302 9330 1322 9350
rect 1410 9330 1430 9350
rect 1513 9326 1533 9346
rect 3316 9323 3336 9343
rect 3419 9327 3439 9347
rect 3529 9323 3549 9343
rect 3632 9327 3652 9347
rect 3737 9323 3757 9343
rect 3840 9327 3860 9347
rect 3948 9327 3968 9347
rect 4051 9323 4071 9343
rect 459 8808 477 8826
rect 461 8709 479 8727
rect 459 8552 477 8570
rect 779 8485 799 8505
rect 882 8489 902 8509
rect 992 8485 1012 8505
rect 1095 8489 1115 8509
rect 1200 8485 1220 8505
rect 1303 8489 1323 8509
rect 1411 8489 1431 8509
rect 1514 8485 1534 8505
rect 1827 8481 1847 8501
rect 461 8453 479 8471
rect 1930 8485 1950 8505
rect 2040 8481 2060 8501
rect 2143 8485 2163 8505
rect 2248 8481 2268 8501
rect 2351 8485 2371 8505
rect 2459 8485 2479 8505
rect 2562 8481 2582 8501
rect 459 8157 477 8175
rect 461 8058 479 8076
rect 459 7902 477 7920
rect 461 7803 479 7821
rect 779 7806 799 7826
rect 882 7810 902 7830
rect 992 7806 1012 7826
rect 1095 7810 1115 7830
rect 1200 7806 1220 7826
rect 1303 7810 1323 7830
rect 1411 7810 1431 7830
rect 1514 7806 1534 7826
rect 3274 7801 3294 7821
rect 3377 7805 3397 7825
rect 3487 7801 3507 7821
rect 3590 7805 3610 7825
rect 3695 7801 3715 7821
rect 3798 7805 3818 7825
rect 3906 7805 3926 7825
rect 4009 7801 4029 7821
rect 459 7361 477 7379
rect 461 7262 479 7280
rect 459 7105 477 7123
rect 779 7038 799 7058
rect 882 7042 902 7062
rect 992 7038 1012 7058
rect 1095 7042 1115 7062
rect 1200 7038 1220 7058
rect 1303 7042 1323 7062
rect 1411 7042 1431 7062
rect 1514 7038 1534 7058
rect 1827 7034 1847 7054
rect 461 7006 479 7024
rect 1930 7038 1950 7058
rect 2040 7034 2060 7054
rect 2143 7038 2163 7058
rect 2248 7034 2268 7054
rect 2351 7038 2371 7058
rect 2459 7038 2479 7058
rect 2562 7034 2582 7054
rect 459 6710 477 6728
rect 461 6611 479 6629
rect 459 6455 477 6473
rect 461 6356 479 6374
rect 779 6359 799 6379
rect 882 6363 902 6383
rect 992 6359 1012 6379
rect 1095 6363 1115 6383
rect 1200 6359 1220 6379
rect 1303 6363 1323 6383
rect 1411 6363 1431 6383
rect 1514 6359 1534 6379
rect 4382 6350 4402 6370
rect 4485 6354 4505 6374
rect 4595 6350 4615 6370
rect 4698 6354 4718 6374
rect 4803 6350 4823 6370
rect 4906 6354 4926 6374
rect 5014 6354 5034 6374
rect 5117 6350 5137 6370
rect 456 5767 474 5785
rect 458 5668 476 5686
rect 456 5511 474 5529
rect 776 5444 796 5464
rect 879 5448 899 5468
rect 989 5444 1009 5464
rect 1092 5448 1112 5468
rect 1197 5444 1217 5464
rect 1300 5448 1320 5468
rect 1408 5448 1428 5468
rect 1511 5444 1531 5464
rect 1824 5440 1844 5460
rect 458 5412 476 5430
rect 1927 5444 1947 5464
rect 2037 5440 2057 5460
rect 2140 5444 2160 5464
rect 2245 5440 2265 5460
rect 2348 5444 2368 5464
rect 2456 5444 2476 5464
rect 2559 5440 2579 5460
rect 456 5116 474 5134
rect 458 5017 476 5035
rect 456 4861 474 4879
rect 458 4762 476 4780
rect 776 4765 796 4785
rect 879 4769 899 4789
rect 989 4765 1009 4785
rect 1092 4769 1112 4789
rect 1197 4765 1217 4785
rect 1300 4769 1320 4789
rect 1408 4769 1428 4789
rect 1511 4765 1531 4785
rect 3271 4760 3291 4780
rect 3374 4764 3394 4784
rect 3484 4760 3504 4780
rect 3587 4764 3607 4784
rect 3692 4760 3712 4780
rect 3795 4764 3815 4784
rect 3903 4764 3923 4784
rect 4006 4760 4026 4780
rect 456 4320 474 4338
rect 458 4221 476 4239
rect 456 4064 474 4082
rect 776 3997 796 4017
rect 879 4001 899 4021
rect 989 3997 1009 4017
rect 1092 4001 1112 4021
rect 1197 3997 1217 4017
rect 1300 4001 1320 4021
rect 1408 4001 1428 4021
rect 1511 3997 1531 4017
rect 1824 3993 1844 4013
rect 458 3965 476 3983
rect 1927 3997 1947 4017
rect 2037 3993 2057 4013
rect 2140 3997 2160 4017
rect 2245 3993 2265 4013
rect 2348 3997 2368 4017
rect 2456 3997 2476 4017
rect 2559 3993 2579 4013
rect 456 3669 474 3687
rect 458 3570 476 3588
rect 456 3414 474 3432
rect 458 3315 476 3333
rect 776 3318 796 3338
rect 879 3322 899 3342
rect 989 3318 1009 3338
rect 1092 3322 1112 3342
rect 1197 3318 1217 3338
rect 1300 3322 1320 3342
rect 1408 3322 1428 3342
rect 1511 3318 1531 3338
rect 3314 3315 3334 3335
rect 3417 3319 3437 3339
rect 3527 3315 3547 3335
rect 3630 3319 3650 3339
rect 3735 3315 3755 3335
rect 3838 3319 3858 3339
rect 3946 3319 3966 3339
rect 4049 3315 4069 3335
rect 457 2800 475 2818
rect 459 2701 477 2719
rect 457 2544 475 2562
rect 777 2477 797 2497
rect 880 2481 900 2501
rect 990 2477 1010 2497
rect 1093 2481 1113 2501
rect 1198 2477 1218 2497
rect 1301 2481 1321 2501
rect 1409 2481 1429 2501
rect 1512 2477 1532 2497
rect 1825 2473 1845 2493
rect 459 2445 477 2463
rect 1928 2477 1948 2497
rect 2038 2473 2058 2493
rect 2141 2477 2161 2497
rect 2246 2473 2266 2493
rect 2349 2477 2369 2497
rect 2457 2477 2477 2497
rect 2560 2473 2580 2493
rect 457 2149 475 2167
rect 459 2050 477 2068
rect 457 1894 475 1912
rect 459 1795 477 1813
rect 777 1798 797 1818
rect 880 1802 900 1822
rect 990 1798 1010 1818
rect 1093 1802 1113 1822
rect 1198 1798 1218 1818
rect 1301 1802 1321 1822
rect 1409 1802 1429 1822
rect 1512 1798 1532 1818
rect 3272 1793 3292 1813
rect 3375 1797 3395 1817
rect 3485 1793 3505 1813
rect 3588 1797 3608 1817
rect 3693 1793 3713 1813
rect 3796 1797 3816 1817
rect 3904 1797 3924 1817
rect 4007 1793 4027 1813
rect 457 1353 475 1371
rect 459 1254 477 1272
rect 457 1097 475 1115
rect 777 1030 797 1050
rect 880 1034 900 1054
rect 990 1030 1010 1050
rect 1093 1034 1113 1054
rect 1198 1030 1218 1050
rect 1301 1034 1321 1054
rect 1409 1034 1429 1054
rect 1512 1030 1532 1050
rect 1825 1026 1845 1046
rect 459 998 477 1016
rect 1928 1030 1948 1050
rect 2038 1026 2058 1046
rect 2141 1030 2161 1050
rect 2246 1026 2266 1046
rect 2349 1030 2369 1050
rect 2457 1030 2477 1050
rect 2560 1026 2580 1046
rect 457 702 475 720
rect 459 603 477 621
rect 457 447 475 465
rect 459 348 477 366
rect 777 351 797 371
rect 880 355 900 375
rect 990 351 1010 371
rect 1093 355 1113 375
rect 1198 351 1218 371
rect 1301 355 1321 375
rect 1409 355 1429 375
rect 1512 351 1532 371
<< pdiffc >>
rect 784 11601 804 11621
rect 880 11601 900 11621
rect 997 11601 1017 11621
rect 1093 11601 1113 11621
rect 1205 11601 1225 11621
rect 1301 11601 1321 11621
rect 1411 11601 1431 11621
rect 1507 11601 1527 11621
rect 1832 11597 1852 11617
rect 1928 11597 1948 11617
rect 2045 11597 2065 11617
rect 2141 11597 2161 11617
rect 2253 11597 2273 11617
rect 2349 11597 2369 11617
rect 2459 11597 2479 11617
rect 2555 11597 2575 11617
rect 784 10922 804 10942
rect 880 10922 900 10942
rect 997 10922 1017 10942
rect 1093 10922 1113 10942
rect 1205 10922 1225 10942
rect 1301 10922 1321 10942
rect 1411 10922 1431 10942
rect 1507 10922 1527 10942
rect 3279 10917 3299 10937
rect 3375 10917 3395 10937
rect 3492 10917 3512 10937
rect 3588 10917 3608 10937
rect 3700 10917 3720 10937
rect 3796 10917 3816 10937
rect 3906 10917 3926 10937
rect 4002 10917 4022 10937
rect 784 10154 804 10174
rect 880 10154 900 10174
rect 997 10154 1017 10174
rect 1093 10154 1113 10174
rect 1205 10154 1225 10174
rect 1301 10154 1321 10174
rect 1411 10154 1431 10174
rect 1507 10154 1527 10174
rect 1832 10150 1852 10170
rect 1928 10150 1948 10170
rect 2045 10150 2065 10170
rect 2141 10150 2161 10170
rect 2253 10150 2273 10170
rect 2349 10150 2369 10170
rect 2459 10150 2479 10170
rect 2555 10150 2575 10170
rect 784 9475 804 9495
rect 880 9475 900 9495
rect 997 9475 1017 9495
rect 1093 9475 1113 9495
rect 1205 9475 1225 9495
rect 1301 9475 1321 9495
rect 1411 9475 1431 9495
rect 1507 9475 1527 9495
rect 3322 9472 3342 9492
rect 3418 9472 3438 9492
rect 3535 9472 3555 9492
rect 3631 9472 3651 9492
rect 3743 9472 3763 9492
rect 3839 9472 3859 9492
rect 3949 9472 3969 9492
rect 4045 9472 4065 9492
rect 785 8634 805 8654
rect 881 8634 901 8654
rect 998 8634 1018 8654
rect 1094 8634 1114 8654
rect 1206 8634 1226 8654
rect 1302 8634 1322 8654
rect 1412 8634 1432 8654
rect 1508 8634 1528 8654
rect 1833 8630 1853 8650
rect 1929 8630 1949 8650
rect 2046 8630 2066 8650
rect 2142 8630 2162 8650
rect 2254 8630 2274 8650
rect 2350 8630 2370 8650
rect 2460 8630 2480 8650
rect 2556 8630 2576 8650
rect 785 7955 805 7975
rect 881 7955 901 7975
rect 998 7955 1018 7975
rect 1094 7955 1114 7975
rect 1206 7955 1226 7975
rect 1302 7955 1322 7975
rect 1412 7955 1432 7975
rect 1508 7955 1528 7975
rect 3280 7950 3300 7970
rect 3376 7950 3396 7970
rect 3493 7950 3513 7970
rect 3589 7950 3609 7970
rect 3701 7950 3721 7970
rect 3797 7950 3817 7970
rect 3907 7950 3927 7970
rect 4003 7950 4023 7970
rect 785 7187 805 7207
rect 881 7187 901 7207
rect 998 7187 1018 7207
rect 1094 7187 1114 7207
rect 1206 7187 1226 7207
rect 1302 7187 1322 7207
rect 1412 7187 1432 7207
rect 1508 7187 1528 7207
rect 1833 7183 1853 7203
rect 1929 7183 1949 7203
rect 2046 7183 2066 7203
rect 2142 7183 2162 7203
rect 2254 7183 2274 7203
rect 2350 7183 2370 7203
rect 2460 7183 2480 7203
rect 2556 7183 2576 7203
rect 785 6508 805 6528
rect 881 6508 901 6528
rect 998 6508 1018 6528
rect 1094 6508 1114 6528
rect 1206 6508 1226 6528
rect 1302 6508 1322 6528
rect 1412 6508 1432 6528
rect 1508 6508 1528 6528
rect 4388 6499 4408 6519
rect 4484 6499 4504 6519
rect 4601 6499 4621 6519
rect 4697 6499 4717 6519
rect 4809 6499 4829 6519
rect 4905 6499 4925 6519
rect 5015 6499 5035 6519
rect 5111 6499 5131 6519
rect 782 5593 802 5613
rect 878 5593 898 5613
rect 995 5593 1015 5613
rect 1091 5593 1111 5613
rect 1203 5593 1223 5613
rect 1299 5593 1319 5613
rect 1409 5593 1429 5613
rect 1505 5593 1525 5613
rect 1830 5589 1850 5609
rect 1926 5589 1946 5609
rect 2043 5589 2063 5609
rect 2139 5589 2159 5609
rect 2251 5589 2271 5609
rect 2347 5589 2367 5609
rect 2457 5589 2477 5609
rect 2553 5589 2573 5609
rect 782 4914 802 4934
rect 878 4914 898 4934
rect 995 4914 1015 4934
rect 1091 4914 1111 4934
rect 1203 4914 1223 4934
rect 1299 4914 1319 4934
rect 1409 4914 1429 4934
rect 1505 4914 1525 4934
rect 3277 4909 3297 4929
rect 3373 4909 3393 4929
rect 3490 4909 3510 4929
rect 3586 4909 3606 4929
rect 3698 4909 3718 4929
rect 3794 4909 3814 4929
rect 3904 4909 3924 4929
rect 4000 4909 4020 4929
rect 782 4146 802 4166
rect 878 4146 898 4166
rect 995 4146 1015 4166
rect 1091 4146 1111 4166
rect 1203 4146 1223 4166
rect 1299 4146 1319 4166
rect 1409 4146 1429 4166
rect 1505 4146 1525 4166
rect 1830 4142 1850 4162
rect 1926 4142 1946 4162
rect 2043 4142 2063 4162
rect 2139 4142 2159 4162
rect 2251 4142 2271 4162
rect 2347 4142 2367 4162
rect 2457 4142 2477 4162
rect 2553 4142 2573 4162
rect 782 3467 802 3487
rect 878 3467 898 3487
rect 995 3467 1015 3487
rect 1091 3467 1111 3487
rect 1203 3467 1223 3487
rect 1299 3467 1319 3487
rect 1409 3467 1429 3487
rect 1505 3467 1525 3487
rect 3320 3464 3340 3484
rect 3416 3464 3436 3484
rect 3533 3464 3553 3484
rect 3629 3464 3649 3484
rect 3741 3464 3761 3484
rect 3837 3464 3857 3484
rect 3947 3464 3967 3484
rect 4043 3464 4063 3484
rect 783 2626 803 2646
rect 879 2626 899 2646
rect 996 2626 1016 2646
rect 1092 2626 1112 2646
rect 1204 2626 1224 2646
rect 1300 2626 1320 2646
rect 1410 2626 1430 2646
rect 1506 2626 1526 2646
rect 1831 2622 1851 2642
rect 1927 2622 1947 2642
rect 2044 2622 2064 2642
rect 2140 2622 2160 2642
rect 2252 2622 2272 2642
rect 2348 2622 2368 2642
rect 2458 2622 2478 2642
rect 2554 2622 2574 2642
rect 783 1947 803 1967
rect 879 1947 899 1967
rect 996 1947 1016 1967
rect 1092 1947 1112 1967
rect 1204 1947 1224 1967
rect 1300 1947 1320 1967
rect 1410 1947 1430 1967
rect 1506 1947 1526 1967
rect 3278 1942 3298 1962
rect 3374 1942 3394 1962
rect 3491 1942 3511 1962
rect 3587 1942 3607 1962
rect 3699 1942 3719 1962
rect 3795 1942 3815 1962
rect 3905 1942 3925 1962
rect 4001 1942 4021 1962
rect 783 1179 803 1199
rect 879 1179 899 1199
rect 996 1179 1016 1199
rect 1092 1179 1112 1199
rect 1204 1179 1224 1199
rect 1300 1179 1320 1199
rect 1410 1179 1430 1199
rect 1506 1179 1526 1199
rect 1831 1175 1851 1195
rect 1927 1175 1947 1195
rect 2044 1175 2064 1195
rect 2140 1175 2160 1195
rect 2252 1175 2272 1195
rect 2348 1175 2368 1195
rect 2458 1175 2478 1195
rect 2554 1175 2574 1195
rect 783 500 803 520
rect 879 500 899 520
rect 996 500 1016 520
rect 1092 500 1112 520
rect 1204 500 1224 520
rect 1300 500 1320 520
rect 1410 500 1430 520
rect 1506 500 1526 520
<< psubdiff >>
rect 852 11385 963 11399
rect 852 11355 893 11385
rect 921 11355 963 11385
rect 852 11340 963 11355
rect 1900 11381 2011 11395
rect 1900 11351 1941 11381
rect 1969 11351 2011 11381
rect 1900 11336 2011 11351
rect 852 10706 963 10720
rect 852 10676 893 10706
rect 921 10676 963 10706
rect 852 10663 963 10676
rect 3347 10701 3458 10715
rect 3347 10671 3388 10701
rect 3416 10671 3458 10701
rect 3347 10656 3458 10671
rect 852 9938 963 9952
rect 852 9908 893 9938
rect 921 9908 963 9938
rect 852 9893 963 9908
rect 1900 9934 2011 9948
rect 1900 9904 1941 9934
rect 1969 9904 2011 9934
rect 1900 9889 2011 9904
rect 852 9259 963 9273
rect 852 9229 893 9259
rect 921 9229 963 9259
rect 852 9214 963 9229
rect 3390 9256 3501 9270
rect 3390 9226 3431 9256
rect 3459 9226 3501 9256
rect 3390 9211 3501 9226
rect 853 8418 964 8432
rect 853 8388 894 8418
rect 922 8388 964 8418
rect 853 8373 964 8388
rect 1901 8414 2012 8428
rect 1901 8384 1942 8414
rect 1970 8384 2012 8414
rect 1901 8369 2012 8384
rect 853 7739 964 7753
rect 853 7709 894 7739
rect 922 7709 964 7739
rect 853 7696 964 7709
rect 3348 7734 3459 7748
rect 3348 7704 3389 7734
rect 3417 7704 3459 7734
rect 3348 7689 3459 7704
rect 853 6971 964 6985
rect 853 6941 894 6971
rect 922 6941 964 6971
rect 853 6926 964 6941
rect 1901 6967 2012 6981
rect 1901 6937 1942 6967
rect 1970 6937 2012 6967
rect 1901 6922 2012 6937
rect 853 6292 964 6306
rect 853 6262 894 6292
rect 922 6262 964 6292
rect 853 6247 964 6262
rect 4456 6283 4567 6297
rect 4456 6253 4497 6283
rect 4525 6253 4567 6283
rect 4456 6238 4567 6253
rect 850 5377 961 5391
rect 850 5347 891 5377
rect 919 5347 961 5377
rect 850 5332 961 5347
rect 1898 5373 2009 5387
rect 1898 5343 1939 5373
rect 1967 5343 2009 5373
rect 1898 5328 2009 5343
rect 850 4698 961 4712
rect 850 4668 891 4698
rect 919 4668 961 4698
rect 850 4655 961 4668
rect 3345 4693 3456 4707
rect 3345 4663 3386 4693
rect 3414 4663 3456 4693
rect 3345 4648 3456 4663
rect 850 3930 961 3944
rect 850 3900 891 3930
rect 919 3900 961 3930
rect 850 3885 961 3900
rect 1898 3926 2009 3940
rect 1898 3896 1939 3926
rect 1967 3896 2009 3926
rect 1898 3881 2009 3896
rect 850 3251 961 3265
rect 850 3221 891 3251
rect 919 3221 961 3251
rect 850 3206 961 3221
rect 3388 3248 3499 3262
rect 3388 3218 3429 3248
rect 3457 3218 3499 3248
rect 3388 3203 3499 3218
rect 851 2410 962 2424
rect 851 2380 892 2410
rect 920 2380 962 2410
rect 851 2365 962 2380
rect 1899 2406 2010 2420
rect 1899 2376 1940 2406
rect 1968 2376 2010 2406
rect 1899 2361 2010 2376
rect 851 1731 962 1745
rect 851 1701 892 1731
rect 920 1701 962 1731
rect 851 1688 962 1701
rect 3346 1726 3457 1740
rect 3346 1696 3387 1726
rect 3415 1696 3457 1726
rect 3346 1681 3457 1696
rect 851 963 962 977
rect 851 933 892 963
rect 920 933 962 963
rect 851 918 962 933
rect 1899 959 2010 973
rect 1899 929 1940 959
rect 1968 929 2010 959
rect 1899 914 2010 929
rect 851 284 962 298
rect 851 254 892 284
rect 920 254 962 284
rect 851 239 962 254
<< nsubdiff >>
rect 853 11732 963 11746
rect 853 11702 896 11732
rect 924 11702 963 11732
rect 853 11687 963 11702
rect 1901 11728 2011 11742
rect 1901 11698 1944 11728
rect 1972 11698 2011 11728
rect 1901 11683 2011 11698
rect 853 11053 963 11067
rect 853 11023 896 11053
rect 924 11023 963 11053
rect 853 11008 963 11023
rect 3348 11048 3458 11062
rect 3348 11018 3391 11048
rect 3419 11018 3458 11048
rect 3348 11003 3458 11018
rect 853 10285 963 10299
rect 853 10255 896 10285
rect 924 10255 963 10285
rect 853 10240 963 10255
rect 1901 10281 2011 10295
rect 1901 10251 1944 10281
rect 1972 10251 2011 10281
rect 1901 10236 2011 10251
rect 853 9606 963 9620
rect 853 9576 896 9606
rect 924 9576 963 9606
rect 853 9561 963 9576
rect 3391 9603 3501 9617
rect 3391 9573 3434 9603
rect 3462 9573 3501 9603
rect 3391 9558 3501 9573
rect 854 8765 964 8779
rect 854 8735 897 8765
rect 925 8735 964 8765
rect 854 8720 964 8735
rect 1902 8761 2012 8775
rect 1902 8731 1945 8761
rect 1973 8731 2012 8761
rect 1902 8716 2012 8731
rect 854 8086 964 8100
rect 854 8056 897 8086
rect 925 8056 964 8086
rect 854 8041 964 8056
rect 3349 8081 3459 8095
rect 3349 8051 3392 8081
rect 3420 8051 3459 8081
rect 3349 8036 3459 8051
rect 854 7318 964 7332
rect 854 7288 897 7318
rect 925 7288 964 7318
rect 854 7273 964 7288
rect 1902 7314 2012 7328
rect 1902 7284 1945 7314
rect 1973 7284 2012 7314
rect 1902 7269 2012 7284
rect 854 6639 964 6653
rect 854 6609 897 6639
rect 925 6609 964 6639
rect 854 6594 964 6609
rect 4457 6630 4567 6644
rect 4457 6600 4500 6630
rect 4528 6600 4567 6630
rect 4457 6585 4567 6600
rect 851 5724 961 5738
rect 851 5694 894 5724
rect 922 5694 961 5724
rect 851 5679 961 5694
rect 1899 5720 2009 5734
rect 1899 5690 1942 5720
rect 1970 5690 2009 5720
rect 1899 5675 2009 5690
rect 851 5045 961 5059
rect 851 5015 894 5045
rect 922 5015 961 5045
rect 851 5000 961 5015
rect 3346 5040 3456 5054
rect 3346 5010 3389 5040
rect 3417 5010 3456 5040
rect 3346 4995 3456 5010
rect 851 4277 961 4291
rect 851 4247 894 4277
rect 922 4247 961 4277
rect 851 4232 961 4247
rect 1899 4273 2009 4287
rect 1899 4243 1942 4273
rect 1970 4243 2009 4273
rect 1899 4228 2009 4243
rect 851 3598 961 3612
rect 851 3568 894 3598
rect 922 3568 961 3598
rect 851 3553 961 3568
rect 3389 3595 3499 3609
rect 3389 3565 3432 3595
rect 3460 3565 3499 3595
rect 3389 3550 3499 3565
rect 852 2757 962 2771
rect 852 2727 895 2757
rect 923 2727 962 2757
rect 852 2712 962 2727
rect 1900 2753 2010 2767
rect 1900 2723 1943 2753
rect 1971 2723 2010 2753
rect 1900 2708 2010 2723
rect 852 2078 962 2092
rect 852 2048 895 2078
rect 923 2048 962 2078
rect 852 2033 962 2048
rect 3347 2073 3457 2087
rect 3347 2043 3390 2073
rect 3418 2043 3457 2073
rect 3347 2028 3457 2043
rect 852 1310 962 1324
rect 852 1280 895 1310
rect 923 1280 962 1310
rect 852 1265 962 1280
rect 1900 1306 2010 1320
rect 1900 1276 1943 1306
rect 1971 1276 2010 1306
rect 1900 1261 2010 1276
rect 852 631 962 645
rect 852 601 895 631
rect 923 601 962 631
rect 852 586 962 601
<< psubdiffcont >>
rect 893 11355 921 11385
rect 1941 11351 1969 11381
rect 893 10676 921 10706
rect 3388 10671 3416 10701
rect 893 9908 921 9938
rect 1941 9904 1969 9934
rect 893 9229 921 9259
rect 3431 9226 3459 9256
rect 894 8388 922 8418
rect 1942 8384 1970 8414
rect 894 7709 922 7739
rect 3389 7704 3417 7734
rect 894 6941 922 6971
rect 1942 6937 1970 6967
rect 894 6262 922 6292
rect 4497 6253 4525 6283
rect 891 5347 919 5377
rect 1939 5343 1967 5373
rect 891 4668 919 4698
rect 3386 4663 3414 4693
rect 891 3900 919 3930
rect 1939 3896 1967 3926
rect 891 3221 919 3251
rect 3429 3218 3457 3248
rect 892 2380 920 2410
rect 1940 2376 1968 2406
rect 892 1701 920 1731
rect 3387 1696 3415 1726
rect 892 933 920 963
rect 1940 929 1968 959
rect 892 254 920 284
<< nsubdiffcont >>
rect 896 11702 924 11732
rect 1944 11698 1972 11728
rect 896 11023 924 11053
rect 3391 11018 3419 11048
rect 896 10255 924 10285
rect 1944 10251 1972 10281
rect 896 9576 924 9606
rect 3434 9573 3462 9603
rect 897 8735 925 8765
rect 1945 8731 1973 8761
rect 897 8056 925 8086
rect 3392 8051 3420 8081
rect 897 7288 925 7318
rect 1945 7284 1973 7314
rect 897 6609 925 6639
rect 4500 6600 4528 6630
rect 894 5694 922 5724
rect 1942 5690 1970 5720
rect 894 5015 922 5045
rect 3389 5010 3417 5040
rect 894 4247 922 4277
rect 1942 4243 1970 4273
rect 894 3568 922 3598
rect 3432 3565 3460 3595
rect 895 2727 923 2757
rect 1943 2723 1971 2753
rect 895 2048 923 2078
rect 3390 2043 3418 2073
rect 895 1280 923 1310
rect 1943 1276 1971 1306
rect 895 601 923 631
<< poly >>
rect 816 11659 866 11672
rect 1029 11659 1079 11672
rect 1237 11659 1287 11672
rect 1445 11659 1495 11672
rect 1864 11655 1914 11668
rect 2077 11655 2127 11668
rect 2285 11655 2335 11668
rect 2493 11655 2543 11668
rect 816 11531 866 11559
rect 816 11511 829 11531
rect 849 11511 866 11531
rect 816 11482 866 11511
rect 1029 11530 1079 11559
rect 1029 11506 1040 11530
rect 1064 11506 1079 11530
rect 1029 11482 1079 11506
rect 1237 11535 1287 11559
rect 1237 11511 1249 11535
rect 1273 11511 1287 11535
rect 1237 11482 1287 11511
rect 1445 11533 1495 11559
rect 1445 11507 1463 11533
rect 1489 11507 1495 11533
rect 1445 11482 1495 11507
rect 1864 11527 1914 11555
rect 1864 11507 1877 11527
rect 1897 11507 1914 11527
rect 1864 11478 1914 11507
rect 2077 11526 2127 11555
rect 2077 11502 2088 11526
rect 2112 11502 2127 11526
rect 2077 11478 2127 11502
rect 2285 11531 2335 11555
rect 2285 11507 2297 11531
rect 2321 11507 2335 11531
rect 2285 11478 2335 11507
rect 2493 11529 2543 11555
rect 2493 11503 2511 11529
rect 2537 11503 2543 11529
rect 2493 11478 2543 11503
rect 816 11424 866 11440
rect 1029 11424 1079 11440
rect 1237 11424 1287 11440
rect 1445 11424 1495 11440
rect 1864 11420 1914 11436
rect 2077 11420 2127 11436
rect 2285 11420 2335 11436
rect 2493 11420 2543 11436
rect 816 10980 866 10993
rect 1029 10980 1079 10993
rect 1237 10980 1287 10993
rect 1445 10980 1495 10993
rect 3311 10975 3361 10988
rect 3524 10975 3574 10988
rect 3732 10975 3782 10988
rect 3940 10975 3990 10988
rect 816 10852 866 10880
rect 816 10832 829 10852
rect 849 10832 866 10852
rect 816 10803 866 10832
rect 1029 10851 1079 10880
rect 1029 10827 1040 10851
rect 1064 10827 1079 10851
rect 1029 10803 1079 10827
rect 1237 10856 1287 10880
rect 1237 10832 1249 10856
rect 1273 10832 1287 10856
rect 1237 10803 1287 10832
rect 1445 10854 1495 10880
rect 1445 10828 1463 10854
rect 1489 10828 1495 10854
rect 1445 10803 1495 10828
rect 3311 10847 3361 10875
rect 3311 10827 3324 10847
rect 3344 10827 3361 10847
rect 3311 10798 3361 10827
rect 3524 10846 3574 10875
rect 3524 10822 3535 10846
rect 3559 10822 3574 10846
rect 3524 10798 3574 10822
rect 3732 10851 3782 10875
rect 3732 10827 3744 10851
rect 3768 10827 3782 10851
rect 3732 10798 3782 10827
rect 3940 10849 3990 10875
rect 3940 10823 3958 10849
rect 3984 10823 3990 10849
rect 3940 10798 3990 10823
rect 816 10745 866 10761
rect 1029 10745 1079 10761
rect 1237 10745 1287 10761
rect 1445 10745 1495 10761
rect 3311 10740 3361 10756
rect 3524 10740 3574 10756
rect 3732 10740 3782 10756
rect 3940 10740 3990 10756
rect 816 10212 866 10225
rect 1029 10212 1079 10225
rect 1237 10212 1287 10225
rect 1445 10212 1495 10225
rect 1864 10208 1914 10221
rect 2077 10208 2127 10221
rect 2285 10208 2335 10221
rect 2493 10208 2543 10221
rect 816 10084 866 10112
rect 816 10064 829 10084
rect 849 10064 866 10084
rect 816 10035 866 10064
rect 1029 10083 1079 10112
rect 1029 10059 1040 10083
rect 1064 10059 1079 10083
rect 1029 10035 1079 10059
rect 1237 10088 1287 10112
rect 1237 10064 1249 10088
rect 1273 10064 1287 10088
rect 1237 10035 1287 10064
rect 1445 10086 1495 10112
rect 1445 10060 1463 10086
rect 1489 10060 1495 10086
rect 1445 10035 1495 10060
rect 1864 10080 1914 10108
rect 1864 10060 1877 10080
rect 1897 10060 1914 10080
rect 1864 10031 1914 10060
rect 2077 10079 2127 10108
rect 2077 10055 2088 10079
rect 2112 10055 2127 10079
rect 2077 10031 2127 10055
rect 2285 10084 2335 10108
rect 2285 10060 2297 10084
rect 2321 10060 2335 10084
rect 2285 10031 2335 10060
rect 2493 10082 2543 10108
rect 2493 10056 2511 10082
rect 2537 10056 2543 10082
rect 2493 10031 2543 10056
rect 816 9977 866 9993
rect 1029 9977 1079 9993
rect 1237 9977 1287 9993
rect 1445 9977 1495 9993
rect 1864 9973 1914 9989
rect 2077 9973 2127 9989
rect 2285 9973 2335 9989
rect 2493 9973 2543 9989
rect 816 9533 866 9546
rect 1029 9533 1079 9546
rect 1237 9533 1287 9546
rect 1445 9533 1495 9546
rect 3354 9530 3404 9543
rect 3567 9530 3617 9543
rect 3775 9530 3825 9543
rect 3983 9530 4033 9543
rect 816 9405 866 9433
rect 816 9385 829 9405
rect 849 9385 866 9405
rect 816 9356 866 9385
rect 1029 9404 1079 9433
rect 1029 9380 1040 9404
rect 1064 9380 1079 9404
rect 1029 9356 1079 9380
rect 1237 9409 1287 9433
rect 1237 9385 1249 9409
rect 1273 9385 1287 9409
rect 1237 9356 1287 9385
rect 1445 9407 1495 9433
rect 1445 9381 1463 9407
rect 1489 9381 1495 9407
rect 1445 9356 1495 9381
rect 3354 9402 3404 9430
rect 3354 9382 3367 9402
rect 3387 9382 3404 9402
rect 3354 9353 3404 9382
rect 3567 9401 3617 9430
rect 3567 9377 3578 9401
rect 3602 9377 3617 9401
rect 3567 9353 3617 9377
rect 3775 9406 3825 9430
rect 3775 9382 3787 9406
rect 3811 9382 3825 9406
rect 3775 9353 3825 9382
rect 3983 9404 4033 9430
rect 3983 9378 4001 9404
rect 4027 9378 4033 9404
rect 3983 9353 4033 9378
rect 816 9298 866 9314
rect 1029 9298 1079 9314
rect 1237 9298 1287 9314
rect 1445 9298 1495 9314
rect 3354 9295 3404 9311
rect 3567 9295 3617 9311
rect 3775 9295 3825 9311
rect 3983 9295 4033 9311
rect 817 8692 867 8705
rect 1030 8692 1080 8705
rect 1238 8692 1288 8705
rect 1446 8692 1496 8705
rect 1865 8688 1915 8701
rect 2078 8688 2128 8701
rect 2286 8688 2336 8701
rect 2494 8688 2544 8701
rect 817 8564 867 8592
rect 817 8544 830 8564
rect 850 8544 867 8564
rect 817 8515 867 8544
rect 1030 8563 1080 8592
rect 1030 8539 1041 8563
rect 1065 8539 1080 8563
rect 1030 8515 1080 8539
rect 1238 8568 1288 8592
rect 1238 8544 1250 8568
rect 1274 8544 1288 8568
rect 1238 8515 1288 8544
rect 1446 8566 1496 8592
rect 1446 8540 1464 8566
rect 1490 8540 1496 8566
rect 1446 8515 1496 8540
rect 1865 8560 1915 8588
rect 1865 8540 1878 8560
rect 1898 8540 1915 8560
rect 1865 8511 1915 8540
rect 2078 8559 2128 8588
rect 2078 8535 2089 8559
rect 2113 8535 2128 8559
rect 2078 8511 2128 8535
rect 2286 8564 2336 8588
rect 2286 8540 2298 8564
rect 2322 8540 2336 8564
rect 2286 8511 2336 8540
rect 2494 8562 2544 8588
rect 2494 8536 2512 8562
rect 2538 8536 2544 8562
rect 2494 8511 2544 8536
rect 817 8457 867 8473
rect 1030 8457 1080 8473
rect 1238 8457 1288 8473
rect 1446 8457 1496 8473
rect 1865 8453 1915 8469
rect 2078 8453 2128 8469
rect 2286 8453 2336 8469
rect 2494 8453 2544 8469
rect 817 8013 867 8026
rect 1030 8013 1080 8026
rect 1238 8013 1288 8026
rect 1446 8013 1496 8026
rect 3312 8008 3362 8021
rect 3525 8008 3575 8021
rect 3733 8008 3783 8021
rect 3941 8008 3991 8021
rect 817 7885 867 7913
rect 817 7865 830 7885
rect 850 7865 867 7885
rect 817 7836 867 7865
rect 1030 7884 1080 7913
rect 1030 7860 1041 7884
rect 1065 7860 1080 7884
rect 1030 7836 1080 7860
rect 1238 7889 1288 7913
rect 1238 7865 1250 7889
rect 1274 7865 1288 7889
rect 1238 7836 1288 7865
rect 1446 7887 1496 7913
rect 1446 7861 1464 7887
rect 1490 7861 1496 7887
rect 1446 7836 1496 7861
rect 3312 7880 3362 7908
rect 3312 7860 3325 7880
rect 3345 7860 3362 7880
rect 3312 7831 3362 7860
rect 3525 7879 3575 7908
rect 3525 7855 3536 7879
rect 3560 7855 3575 7879
rect 3525 7831 3575 7855
rect 3733 7884 3783 7908
rect 3733 7860 3745 7884
rect 3769 7860 3783 7884
rect 3733 7831 3783 7860
rect 3941 7882 3991 7908
rect 3941 7856 3959 7882
rect 3985 7856 3991 7882
rect 3941 7831 3991 7856
rect 817 7778 867 7794
rect 1030 7778 1080 7794
rect 1238 7778 1288 7794
rect 1446 7778 1496 7794
rect 3312 7773 3362 7789
rect 3525 7773 3575 7789
rect 3733 7773 3783 7789
rect 3941 7773 3991 7789
rect 817 7245 867 7258
rect 1030 7245 1080 7258
rect 1238 7245 1288 7258
rect 1446 7245 1496 7258
rect 1865 7241 1915 7254
rect 2078 7241 2128 7254
rect 2286 7241 2336 7254
rect 2494 7241 2544 7254
rect 817 7117 867 7145
rect 817 7097 830 7117
rect 850 7097 867 7117
rect 817 7068 867 7097
rect 1030 7116 1080 7145
rect 1030 7092 1041 7116
rect 1065 7092 1080 7116
rect 1030 7068 1080 7092
rect 1238 7121 1288 7145
rect 1238 7097 1250 7121
rect 1274 7097 1288 7121
rect 1238 7068 1288 7097
rect 1446 7119 1496 7145
rect 1446 7093 1464 7119
rect 1490 7093 1496 7119
rect 1446 7068 1496 7093
rect 1865 7113 1915 7141
rect 1865 7093 1878 7113
rect 1898 7093 1915 7113
rect 1865 7064 1915 7093
rect 2078 7112 2128 7141
rect 2078 7088 2089 7112
rect 2113 7088 2128 7112
rect 2078 7064 2128 7088
rect 2286 7117 2336 7141
rect 2286 7093 2298 7117
rect 2322 7093 2336 7117
rect 2286 7064 2336 7093
rect 2494 7115 2544 7141
rect 2494 7089 2512 7115
rect 2538 7089 2544 7115
rect 2494 7064 2544 7089
rect 817 7010 867 7026
rect 1030 7010 1080 7026
rect 1238 7010 1288 7026
rect 1446 7010 1496 7026
rect 1865 7006 1915 7022
rect 2078 7006 2128 7022
rect 2286 7006 2336 7022
rect 2494 7006 2544 7022
rect 817 6566 867 6579
rect 1030 6566 1080 6579
rect 1238 6566 1288 6579
rect 1446 6566 1496 6579
rect 4420 6557 4470 6570
rect 4633 6557 4683 6570
rect 4841 6557 4891 6570
rect 5049 6557 5099 6570
rect 817 6438 867 6466
rect 817 6418 830 6438
rect 850 6418 867 6438
rect 817 6389 867 6418
rect 1030 6437 1080 6466
rect 1030 6413 1041 6437
rect 1065 6413 1080 6437
rect 1030 6389 1080 6413
rect 1238 6442 1288 6466
rect 1238 6418 1250 6442
rect 1274 6418 1288 6442
rect 1238 6389 1288 6418
rect 1446 6440 1496 6466
rect 1446 6414 1464 6440
rect 1490 6414 1496 6440
rect 1446 6389 1496 6414
rect 4420 6429 4470 6457
rect 4420 6409 4433 6429
rect 4453 6409 4470 6429
rect 4420 6380 4470 6409
rect 4633 6428 4683 6457
rect 4633 6404 4644 6428
rect 4668 6404 4683 6428
rect 4633 6380 4683 6404
rect 4841 6433 4891 6457
rect 4841 6409 4853 6433
rect 4877 6409 4891 6433
rect 4841 6380 4891 6409
rect 5049 6431 5099 6457
rect 5049 6405 5067 6431
rect 5093 6405 5099 6431
rect 5049 6380 5099 6405
rect 817 6331 867 6347
rect 1030 6331 1080 6347
rect 1238 6331 1288 6347
rect 1446 6331 1496 6347
rect 4420 6322 4470 6338
rect 4633 6322 4683 6338
rect 4841 6322 4891 6338
rect 5049 6322 5099 6338
rect 814 5651 864 5664
rect 1027 5651 1077 5664
rect 1235 5651 1285 5664
rect 1443 5651 1493 5664
rect 1862 5647 1912 5660
rect 2075 5647 2125 5660
rect 2283 5647 2333 5660
rect 2491 5647 2541 5660
rect 814 5523 864 5551
rect 814 5503 827 5523
rect 847 5503 864 5523
rect 814 5474 864 5503
rect 1027 5522 1077 5551
rect 1027 5498 1038 5522
rect 1062 5498 1077 5522
rect 1027 5474 1077 5498
rect 1235 5527 1285 5551
rect 1235 5503 1247 5527
rect 1271 5503 1285 5527
rect 1235 5474 1285 5503
rect 1443 5525 1493 5551
rect 1443 5499 1461 5525
rect 1487 5499 1493 5525
rect 1443 5474 1493 5499
rect 1862 5519 1912 5547
rect 1862 5499 1875 5519
rect 1895 5499 1912 5519
rect 1862 5470 1912 5499
rect 2075 5518 2125 5547
rect 2075 5494 2086 5518
rect 2110 5494 2125 5518
rect 2075 5470 2125 5494
rect 2283 5523 2333 5547
rect 2283 5499 2295 5523
rect 2319 5499 2333 5523
rect 2283 5470 2333 5499
rect 2491 5521 2541 5547
rect 2491 5495 2509 5521
rect 2535 5495 2541 5521
rect 2491 5470 2541 5495
rect 814 5416 864 5432
rect 1027 5416 1077 5432
rect 1235 5416 1285 5432
rect 1443 5416 1493 5432
rect 1862 5412 1912 5428
rect 2075 5412 2125 5428
rect 2283 5412 2333 5428
rect 2491 5412 2541 5428
rect 814 4972 864 4985
rect 1027 4972 1077 4985
rect 1235 4972 1285 4985
rect 1443 4972 1493 4985
rect 3309 4967 3359 4980
rect 3522 4967 3572 4980
rect 3730 4967 3780 4980
rect 3938 4967 3988 4980
rect 814 4844 864 4872
rect 814 4824 827 4844
rect 847 4824 864 4844
rect 814 4795 864 4824
rect 1027 4843 1077 4872
rect 1027 4819 1038 4843
rect 1062 4819 1077 4843
rect 1027 4795 1077 4819
rect 1235 4848 1285 4872
rect 1235 4824 1247 4848
rect 1271 4824 1285 4848
rect 1235 4795 1285 4824
rect 1443 4846 1493 4872
rect 1443 4820 1461 4846
rect 1487 4820 1493 4846
rect 1443 4795 1493 4820
rect 3309 4839 3359 4867
rect 3309 4819 3322 4839
rect 3342 4819 3359 4839
rect 3309 4790 3359 4819
rect 3522 4838 3572 4867
rect 3522 4814 3533 4838
rect 3557 4814 3572 4838
rect 3522 4790 3572 4814
rect 3730 4843 3780 4867
rect 3730 4819 3742 4843
rect 3766 4819 3780 4843
rect 3730 4790 3780 4819
rect 3938 4841 3988 4867
rect 3938 4815 3956 4841
rect 3982 4815 3988 4841
rect 3938 4790 3988 4815
rect 814 4737 864 4753
rect 1027 4737 1077 4753
rect 1235 4737 1285 4753
rect 1443 4737 1493 4753
rect 3309 4732 3359 4748
rect 3522 4732 3572 4748
rect 3730 4732 3780 4748
rect 3938 4732 3988 4748
rect 814 4204 864 4217
rect 1027 4204 1077 4217
rect 1235 4204 1285 4217
rect 1443 4204 1493 4217
rect 1862 4200 1912 4213
rect 2075 4200 2125 4213
rect 2283 4200 2333 4213
rect 2491 4200 2541 4213
rect 814 4076 864 4104
rect 814 4056 827 4076
rect 847 4056 864 4076
rect 814 4027 864 4056
rect 1027 4075 1077 4104
rect 1027 4051 1038 4075
rect 1062 4051 1077 4075
rect 1027 4027 1077 4051
rect 1235 4080 1285 4104
rect 1235 4056 1247 4080
rect 1271 4056 1285 4080
rect 1235 4027 1285 4056
rect 1443 4078 1493 4104
rect 1443 4052 1461 4078
rect 1487 4052 1493 4078
rect 1443 4027 1493 4052
rect 1862 4072 1912 4100
rect 1862 4052 1875 4072
rect 1895 4052 1912 4072
rect 1862 4023 1912 4052
rect 2075 4071 2125 4100
rect 2075 4047 2086 4071
rect 2110 4047 2125 4071
rect 2075 4023 2125 4047
rect 2283 4076 2333 4100
rect 2283 4052 2295 4076
rect 2319 4052 2333 4076
rect 2283 4023 2333 4052
rect 2491 4074 2541 4100
rect 2491 4048 2509 4074
rect 2535 4048 2541 4074
rect 2491 4023 2541 4048
rect 814 3969 864 3985
rect 1027 3969 1077 3985
rect 1235 3969 1285 3985
rect 1443 3969 1493 3985
rect 1862 3965 1912 3981
rect 2075 3965 2125 3981
rect 2283 3965 2333 3981
rect 2491 3965 2541 3981
rect 814 3525 864 3538
rect 1027 3525 1077 3538
rect 1235 3525 1285 3538
rect 1443 3525 1493 3538
rect 3352 3522 3402 3535
rect 3565 3522 3615 3535
rect 3773 3522 3823 3535
rect 3981 3522 4031 3535
rect 814 3397 864 3425
rect 814 3377 827 3397
rect 847 3377 864 3397
rect 814 3348 864 3377
rect 1027 3396 1077 3425
rect 1027 3372 1038 3396
rect 1062 3372 1077 3396
rect 1027 3348 1077 3372
rect 1235 3401 1285 3425
rect 1235 3377 1247 3401
rect 1271 3377 1285 3401
rect 1235 3348 1285 3377
rect 1443 3399 1493 3425
rect 1443 3373 1461 3399
rect 1487 3373 1493 3399
rect 1443 3348 1493 3373
rect 3352 3394 3402 3422
rect 3352 3374 3365 3394
rect 3385 3374 3402 3394
rect 3352 3345 3402 3374
rect 3565 3393 3615 3422
rect 3565 3369 3576 3393
rect 3600 3369 3615 3393
rect 3565 3345 3615 3369
rect 3773 3398 3823 3422
rect 3773 3374 3785 3398
rect 3809 3374 3823 3398
rect 3773 3345 3823 3374
rect 3981 3396 4031 3422
rect 3981 3370 3999 3396
rect 4025 3370 4031 3396
rect 3981 3345 4031 3370
rect 814 3290 864 3306
rect 1027 3290 1077 3306
rect 1235 3290 1285 3306
rect 1443 3290 1493 3306
rect 3352 3287 3402 3303
rect 3565 3287 3615 3303
rect 3773 3287 3823 3303
rect 3981 3287 4031 3303
rect 815 2684 865 2697
rect 1028 2684 1078 2697
rect 1236 2684 1286 2697
rect 1444 2684 1494 2697
rect 1863 2680 1913 2693
rect 2076 2680 2126 2693
rect 2284 2680 2334 2693
rect 2492 2680 2542 2693
rect 815 2556 865 2584
rect 815 2536 828 2556
rect 848 2536 865 2556
rect 815 2507 865 2536
rect 1028 2555 1078 2584
rect 1028 2531 1039 2555
rect 1063 2531 1078 2555
rect 1028 2507 1078 2531
rect 1236 2560 1286 2584
rect 1236 2536 1248 2560
rect 1272 2536 1286 2560
rect 1236 2507 1286 2536
rect 1444 2558 1494 2584
rect 1444 2532 1462 2558
rect 1488 2532 1494 2558
rect 1444 2507 1494 2532
rect 1863 2552 1913 2580
rect 1863 2532 1876 2552
rect 1896 2532 1913 2552
rect 1863 2503 1913 2532
rect 2076 2551 2126 2580
rect 2076 2527 2087 2551
rect 2111 2527 2126 2551
rect 2076 2503 2126 2527
rect 2284 2556 2334 2580
rect 2284 2532 2296 2556
rect 2320 2532 2334 2556
rect 2284 2503 2334 2532
rect 2492 2554 2542 2580
rect 2492 2528 2510 2554
rect 2536 2528 2542 2554
rect 2492 2503 2542 2528
rect 815 2449 865 2465
rect 1028 2449 1078 2465
rect 1236 2449 1286 2465
rect 1444 2449 1494 2465
rect 1863 2445 1913 2461
rect 2076 2445 2126 2461
rect 2284 2445 2334 2461
rect 2492 2445 2542 2461
rect 815 2005 865 2018
rect 1028 2005 1078 2018
rect 1236 2005 1286 2018
rect 1444 2005 1494 2018
rect 3310 2000 3360 2013
rect 3523 2000 3573 2013
rect 3731 2000 3781 2013
rect 3939 2000 3989 2013
rect 815 1877 865 1905
rect 815 1857 828 1877
rect 848 1857 865 1877
rect 815 1828 865 1857
rect 1028 1876 1078 1905
rect 1028 1852 1039 1876
rect 1063 1852 1078 1876
rect 1028 1828 1078 1852
rect 1236 1881 1286 1905
rect 1236 1857 1248 1881
rect 1272 1857 1286 1881
rect 1236 1828 1286 1857
rect 1444 1879 1494 1905
rect 1444 1853 1462 1879
rect 1488 1853 1494 1879
rect 1444 1828 1494 1853
rect 3310 1872 3360 1900
rect 3310 1852 3323 1872
rect 3343 1852 3360 1872
rect 3310 1823 3360 1852
rect 3523 1871 3573 1900
rect 3523 1847 3534 1871
rect 3558 1847 3573 1871
rect 3523 1823 3573 1847
rect 3731 1876 3781 1900
rect 3731 1852 3743 1876
rect 3767 1852 3781 1876
rect 3731 1823 3781 1852
rect 3939 1874 3989 1900
rect 3939 1848 3957 1874
rect 3983 1848 3989 1874
rect 3939 1823 3989 1848
rect 815 1770 865 1786
rect 1028 1770 1078 1786
rect 1236 1770 1286 1786
rect 1444 1770 1494 1786
rect 3310 1765 3360 1781
rect 3523 1765 3573 1781
rect 3731 1765 3781 1781
rect 3939 1765 3989 1781
rect 815 1237 865 1250
rect 1028 1237 1078 1250
rect 1236 1237 1286 1250
rect 1444 1237 1494 1250
rect 1863 1233 1913 1246
rect 2076 1233 2126 1246
rect 2284 1233 2334 1246
rect 2492 1233 2542 1246
rect 815 1109 865 1137
rect 815 1089 828 1109
rect 848 1089 865 1109
rect 815 1060 865 1089
rect 1028 1108 1078 1137
rect 1028 1084 1039 1108
rect 1063 1084 1078 1108
rect 1028 1060 1078 1084
rect 1236 1113 1286 1137
rect 1236 1089 1248 1113
rect 1272 1089 1286 1113
rect 1236 1060 1286 1089
rect 1444 1111 1494 1137
rect 1444 1085 1462 1111
rect 1488 1085 1494 1111
rect 1444 1060 1494 1085
rect 1863 1105 1913 1133
rect 1863 1085 1876 1105
rect 1896 1085 1913 1105
rect 1863 1056 1913 1085
rect 2076 1104 2126 1133
rect 2076 1080 2087 1104
rect 2111 1080 2126 1104
rect 2076 1056 2126 1080
rect 2284 1109 2334 1133
rect 2284 1085 2296 1109
rect 2320 1085 2334 1109
rect 2284 1056 2334 1085
rect 2492 1107 2542 1133
rect 2492 1081 2510 1107
rect 2536 1081 2542 1107
rect 2492 1056 2542 1081
rect 815 1002 865 1018
rect 1028 1002 1078 1018
rect 1236 1002 1286 1018
rect 1444 1002 1494 1018
rect 1863 998 1913 1014
rect 2076 998 2126 1014
rect 2284 998 2334 1014
rect 2492 998 2542 1014
rect 815 558 865 571
rect 1028 558 1078 571
rect 1236 558 1286 571
rect 1444 558 1494 571
rect 815 430 865 458
rect 815 410 828 430
rect 848 410 865 430
rect 815 381 865 410
rect 1028 429 1078 458
rect 1028 405 1039 429
rect 1063 405 1078 429
rect 1028 381 1078 405
rect 1236 434 1286 458
rect 1236 410 1248 434
rect 1272 410 1286 434
rect 1236 381 1286 410
rect 1444 432 1494 458
rect 1444 406 1462 432
rect 1488 406 1494 432
rect 1444 381 1494 406
rect 815 323 865 339
rect 1028 323 1078 339
rect 1236 323 1286 339
rect 1444 323 1494 339
<< polycont >>
rect 829 11511 849 11531
rect 1040 11506 1064 11530
rect 1249 11511 1273 11535
rect 1463 11507 1489 11533
rect 1877 11507 1897 11527
rect 2088 11502 2112 11526
rect 2297 11507 2321 11531
rect 2511 11503 2537 11529
rect 829 10832 849 10852
rect 1040 10827 1064 10851
rect 1249 10832 1273 10856
rect 1463 10828 1489 10854
rect 3324 10827 3344 10847
rect 3535 10822 3559 10846
rect 3744 10827 3768 10851
rect 3958 10823 3984 10849
rect 829 10064 849 10084
rect 1040 10059 1064 10083
rect 1249 10064 1273 10088
rect 1463 10060 1489 10086
rect 1877 10060 1897 10080
rect 2088 10055 2112 10079
rect 2297 10060 2321 10084
rect 2511 10056 2537 10082
rect 829 9385 849 9405
rect 1040 9380 1064 9404
rect 1249 9385 1273 9409
rect 1463 9381 1489 9407
rect 3367 9382 3387 9402
rect 3578 9377 3602 9401
rect 3787 9382 3811 9406
rect 4001 9378 4027 9404
rect 830 8544 850 8564
rect 1041 8539 1065 8563
rect 1250 8544 1274 8568
rect 1464 8540 1490 8566
rect 1878 8540 1898 8560
rect 2089 8535 2113 8559
rect 2298 8540 2322 8564
rect 2512 8536 2538 8562
rect 830 7865 850 7885
rect 1041 7860 1065 7884
rect 1250 7865 1274 7889
rect 1464 7861 1490 7887
rect 3325 7860 3345 7880
rect 3536 7855 3560 7879
rect 3745 7860 3769 7884
rect 3959 7856 3985 7882
rect 830 7097 850 7117
rect 1041 7092 1065 7116
rect 1250 7097 1274 7121
rect 1464 7093 1490 7119
rect 1878 7093 1898 7113
rect 2089 7088 2113 7112
rect 2298 7093 2322 7117
rect 2512 7089 2538 7115
rect 830 6418 850 6438
rect 1041 6413 1065 6437
rect 1250 6418 1274 6442
rect 1464 6414 1490 6440
rect 4433 6409 4453 6429
rect 4644 6404 4668 6428
rect 4853 6409 4877 6433
rect 5067 6405 5093 6431
rect 827 5503 847 5523
rect 1038 5498 1062 5522
rect 1247 5503 1271 5527
rect 1461 5499 1487 5525
rect 1875 5499 1895 5519
rect 2086 5494 2110 5518
rect 2295 5499 2319 5523
rect 2509 5495 2535 5521
rect 827 4824 847 4844
rect 1038 4819 1062 4843
rect 1247 4824 1271 4848
rect 1461 4820 1487 4846
rect 3322 4819 3342 4839
rect 3533 4814 3557 4838
rect 3742 4819 3766 4843
rect 3956 4815 3982 4841
rect 827 4056 847 4076
rect 1038 4051 1062 4075
rect 1247 4056 1271 4080
rect 1461 4052 1487 4078
rect 1875 4052 1895 4072
rect 2086 4047 2110 4071
rect 2295 4052 2319 4076
rect 2509 4048 2535 4074
rect 827 3377 847 3397
rect 1038 3372 1062 3396
rect 1247 3377 1271 3401
rect 1461 3373 1487 3399
rect 3365 3374 3385 3394
rect 3576 3369 3600 3393
rect 3785 3374 3809 3398
rect 3999 3370 4025 3396
rect 828 2536 848 2556
rect 1039 2531 1063 2555
rect 1248 2536 1272 2560
rect 1462 2532 1488 2558
rect 1876 2532 1896 2552
rect 2087 2527 2111 2551
rect 2296 2532 2320 2556
rect 2510 2528 2536 2554
rect 828 1857 848 1877
rect 1039 1852 1063 1876
rect 1248 1857 1272 1881
rect 1462 1853 1488 1879
rect 3323 1852 3343 1872
rect 3534 1847 3558 1871
rect 3743 1852 3767 1876
rect 3957 1848 3983 1874
rect 828 1089 848 1109
rect 1039 1084 1063 1108
rect 1248 1089 1272 1113
rect 1462 1085 1488 1111
rect 1876 1085 1896 1105
rect 2087 1080 2111 1104
rect 2296 1085 2320 1109
rect 2510 1081 2536 1107
rect 828 410 848 430
rect 1039 405 1063 429
rect 1248 410 1272 434
rect 1462 406 1488 432
<< ndiffres >>
rect 437 11793 494 11812
rect 437 11790 458 11793
rect 343 11775 458 11790
rect 476 11775 494 11793
rect 343 11752 494 11775
rect 343 11716 385 11752
rect 342 11715 442 11716
rect 342 11694 498 11715
rect 342 11676 460 11694
rect 478 11676 498 11694
rect 342 11672 498 11676
rect 437 11656 498 11672
rect 437 11537 494 11556
rect 437 11534 458 11537
rect 343 11519 458 11534
rect 476 11519 494 11537
rect 343 11496 494 11519
rect 343 11460 385 11496
rect 342 11459 442 11460
rect 342 11438 498 11459
rect 342 11420 460 11438
rect 478 11420 498 11438
rect 342 11416 498 11420
rect 437 11400 498 11416
rect 437 11142 494 11161
rect 437 11139 458 11142
rect 343 11124 458 11139
rect 476 11124 494 11142
rect 343 11101 494 11124
rect 343 11065 385 11101
rect 342 11064 442 11065
rect 342 11043 498 11064
rect 342 11025 460 11043
rect 478 11025 498 11043
rect 342 11021 498 11025
rect 437 11005 498 11021
rect 437 10887 494 10906
rect 437 10884 458 10887
rect 343 10869 458 10884
rect 476 10869 494 10887
rect 343 10846 494 10869
rect 343 10810 385 10846
rect 342 10809 442 10810
rect 342 10788 498 10809
rect 342 10770 460 10788
rect 478 10770 498 10788
rect 342 10766 498 10770
rect 437 10750 498 10766
rect 437 10346 494 10365
rect 437 10343 458 10346
rect 343 10328 458 10343
rect 476 10328 494 10346
rect 343 10305 494 10328
rect 343 10269 385 10305
rect 342 10268 442 10269
rect 342 10247 498 10268
rect 342 10229 460 10247
rect 478 10229 498 10247
rect 342 10225 498 10229
rect 437 10209 498 10225
rect 437 10090 494 10109
rect 437 10087 458 10090
rect 343 10072 458 10087
rect 476 10072 494 10090
rect 343 10049 494 10072
rect 343 10013 385 10049
rect 342 10012 442 10013
rect 342 9991 498 10012
rect 342 9973 460 9991
rect 478 9973 498 9991
rect 342 9969 498 9973
rect 437 9953 498 9969
rect 437 9695 494 9714
rect 437 9692 458 9695
rect 343 9677 458 9692
rect 476 9677 494 9695
rect 343 9654 494 9677
rect 343 9618 385 9654
rect 342 9617 442 9618
rect 342 9596 498 9617
rect 342 9578 460 9596
rect 478 9578 498 9596
rect 342 9574 498 9578
rect 437 9558 498 9574
rect 437 9440 494 9459
rect 437 9437 458 9440
rect 343 9422 458 9437
rect 476 9422 494 9440
rect 343 9399 494 9422
rect 343 9363 385 9399
rect 342 9362 442 9363
rect 342 9341 498 9362
rect 342 9323 460 9341
rect 478 9323 498 9341
rect 342 9319 498 9323
rect 437 9303 498 9319
rect 438 8826 495 8845
rect 438 8823 459 8826
rect 344 8808 459 8823
rect 477 8808 495 8826
rect 344 8785 495 8808
rect 344 8749 386 8785
rect 343 8748 443 8749
rect 343 8727 499 8748
rect 343 8709 461 8727
rect 479 8709 499 8727
rect 343 8705 499 8709
rect 438 8689 499 8705
rect 438 8570 495 8589
rect 438 8567 459 8570
rect 344 8552 459 8567
rect 477 8552 495 8570
rect 344 8529 495 8552
rect 344 8493 386 8529
rect 343 8492 443 8493
rect 343 8471 499 8492
rect 343 8453 461 8471
rect 479 8453 499 8471
rect 343 8449 499 8453
rect 438 8433 499 8449
rect 438 8175 495 8194
rect 438 8172 459 8175
rect 344 8157 459 8172
rect 477 8157 495 8175
rect 344 8134 495 8157
rect 344 8098 386 8134
rect 343 8097 443 8098
rect 343 8076 499 8097
rect 343 8058 461 8076
rect 479 8058 499 8076
rect 343 8054 499 8058
rect 438 8038 499 8054
rect 438 7920 495 7939
rect 438 7917 459 7920
rect 344 7902 459 7917
rect 477 7902 495 7920
rect 344 7879 495 7902
rect 344 7843 386 7879
rect 343 7842 443 7843
rect 343 7821 499 7842
rect 343 7803 461 7821
rect 479 7803 499 7821
rect 343 7799 499 7803
rect 438 7783 499 7799
rect 438 7379 495 7398
rect 438 7376 459 7379
rect 344 7361 459 7376
rect 477 7361 495 7379
rect 344 7338 495 7361
rect 344 7302 386 7338
rect 343 7301 443 7302
rect 343 7280 499 7301
rect 343 7262 461 7280
rect 479 7262 499 7280
rect 343 7258 499 7262
rect 438 7242 499 7258
rect 438 7123 495 7142
rect 438 7120 459 7123
rect 344 7105 459 7120
rect 477 7105 495 7123
rect 344 7082 495 7105
rect 344 7046 386 7082
rect 343 7045 443 7046
rect 343 7024 499 7045
rect 343 7006 461 7024
rect 479 7006 499 7024
rect 343 7002 499 7006
rect 438 6986 499 7002
rect 438 6728 495 6747
rect 438 6725 459 6728
rect 344 6710 459 6725
rect 477 6710 495 6728
rect 344 6687 495 6710
rect 344 6651 386 6687
rect 343 6650 443 6651
rect 343 6629 499 6650
rect 343 6611 461 6629
rect 479 6611 499 6629
rect 343 6607 499 6611
rect 438 6591 499 6607
rect 438 6473 495 6492
rect 438 6470 459 6473
rect 344 6455 459 6470
rect 477 6455 495 6473
rect 344 6432 495 6455
rect 344 6396 386 6432
rect 343 6395 443 6396
rect 343 6374 499 6395
rect 343 6356 461 6374
rect 479 6356 499 6374
rect 343 6352 499 6356
rect 438 6336 499 6352
rect 435 5785 492 5804
rect 435 5782 456 5785
rect 341 5767 456 5782
rect 474 5767 492 5785
rect 341 5744 492 5767
rect 341 5708 383 5744
rect 340 5707 440 5708
rect 340 5686 496 5707
rect 340 5668 458 5686
rect 476 5668 496 5686
rect 340 5664 496 5668
rect 435 5648 496 5664
rect 435 5529 492 5548
rect 435 5526 456 5529
rect 341 5511 456 5526
rect 474 5511 492 5529
rect 341 5488 492 5511
rect 341 5452 383 5488
rect 340 5451 440 5452
rect 340 5430 496 5451
rect 340 5412 458 5430
rect 476 5412 496 5430
rect 340 5408 496 5412
rect 435 5392 496 5408
rect 435 5134 492 5153
rect 435 5131 456 5134
rect 341 5116 456 5131
rect 474 5116 492 5134
rect 341 5093 492 5116
rect 341 5057 383 5093
rect 340 5056 440 5057
rect 340 5035 496 5056
rect 340 5017 458 5035
rect 476 5017 496 5035
rect 340 5013 496 5017
rect 435 4997 496 5013
rect 435 4879 492 4898
rect 435 4876 456 4879
rect 341 4861 456 4876
rect 474 4861 492 4879
rect 341 4838 492 4861
rect 341 4802 383 4838
rect 340 4801 440 4802
rect 340 4780 496 4801
rect 340 4762 458 4780
rect 476 4762 496 4780
rect 340 4758 496 4762
rect 435 4742 496 4758
rect 435 4338 492 4357
rect 435 4335 456 4338
rect 341 4320 456 4335
rect 474 4320 492 4338
rect 341 4297 492 4320
rect 341 4261 383 4297
rect 340 4260 440 4261
rect 340 4239 496 4260
rect 340 4221 458 4239
rect 476 4221 496 4239
rect 340 4217 496 4221
rect 435 4201 496 4217
rect 435 4082 492 4101
rect 435 4079 456 4082
rect 341 4064 456 4079
rect 474 4064 492 4082
rect 341 4041 492 4064
rect 341 4005 383 4041
rect 340 4004 440 4005
rect 340 3983 496 4004
rect 340 3965 458 3983
rect 476 3965 496 3983
rect 340 3961 496 3965
rect 435 3945 496 3961
rect 435 3687 492 3706
rect 435 3684 456 3687
rect 341 3669 456 3684
rect 474 3669 492 3687
rect 341 3646 492 3669
rect 341 3610 383 3646
rect 340 3609 440 3610
rect 340 3588 496 3609
rect 340 3570 458 3588
rect 476 3570 496 3588
rect 340 3566 496 3570
rect 435 3550 496 3566
rect 435 3432 492 3451
rect 435 3429 456 3432
rect 341 3414 456 3429
rect 474 3414 492 3432
rect 341 3391 492 3414
rect 341 3355 383 3391
rect 340 3354 440 3355
rect 340 3333 496 3354
rect 340 3315 458 3333
rect 476 3315 496 3333
rect 340 3311 496 3315
rect 435 3295 496 3311
rect 436 2818 493 2837
rect 436 2815 457 2818
rect 342 2800 457 2815
rect 475 2800 493 2818
rect 342 2777 493 2800
rect 342 2741 384 2777
rect 341 2740 441 2741
rect 341 2719 497 2740
rect 341 2701 459 2719
rect 477 2701 497 2719
rect 341 2697 497 2701
rect 436 2681 497 2697
rect 436 2562 493 2581
rect 436 2559 457 2562
rect 342 2544 457 2559
rect 475 2544 493 2562
rect 342 2521 493 2544
rect 342 2485 384 2521
rect 341 2484 441 2485
rect 341 2463 497 2484
rect 341 2445 459 2463
rect 477 2445 497 2463
rect 341 2441 497 2445
rect 436 2425 497 2441
rect 436 2167 493 2186
rect 436 2164 457 2167
rect 342 2149 457 2164
rect 475 2149 493 2167
rect 342 2126 493 2149
rect 342 2090 384 2126
rect 341 2089 441 2090
rect 341 2068 497 2089
rect 341 2050 459 2068
rect 477 2050 497 2068
rect 341 2046 497 2050
rect 436 2030 497 2046
rect 436 1912 493 1931
rect 436 1909 457 1912
rect 342 1894 457 1909
rect 475 1894 493 1912
rect 342 1871 493 1894
rect 342 1835 384 1871
rect 341 1834 441 1835
rect 341 1813 497 1834
rect 341 1795 459 1813
rect 477 1795 497 1813
rect 341 1791 497 1795
rect 436 1775 497 1791
rect 436 1371 493 1390
rect 436 1368 457 1371
rect 342 1353 457 1368
rect 475 1353 493 1371
rect 342 1330 493 1353
rect 342 1294 384 1330
rect 341 1293 441 1294
rect 341 1272 497 1293
rect 341 1254 459 1272
rect 477 1254 497 1272
rect 341 1250 497 1254
rect 436 1234 497 1250
rect 436 1115 493 1134
rect 436 1112 457 1115
rect 342 1097 457 1112
rect 475 1097 493 1115
rect 342 1074 493 1097
rect 342 1038 384 1074
rect 341 1037 441 1038
rect 341 1016 497 1037
rect 341 998 459 1016
rect 477 998 497 1016
rect 341 994 497 998
rect 436 978 497 994
rect 436 720 493 739
rect 436 717 457 720
rect 342 702 457 717
rect 475 702 493 720
rect 342 679 493 702
rect 342 643 384 679
rect 341 642 441 643
rect 341 621 497 642
rect 341 603 459 621
rect 477 603 497 621
rect 341 599 497 603
rect 436 583 497 599
rect 436 465 493 484
rect 436 462 457 465
rect 342 447 457 462
rect 475 447 493 465
rect 342 424 493 447
rect 342 388 384 424
rect 341 387 441 388
rect 341 366 497 387
rect 341 348 459 366
rect 477 348 497 366
rect 341 344 497 348
rect 436 328 497 344
<< locali >>
rect 436 11793 495 11983
rect 2813 11974 2878 11985
rect 2813 11926 2826 11974
rect 2863 11926 2878 11974
rect 2813 11913 2878 11926
rect 3026 11876 3737 11878
rect 2399 11875 3737 11876
rect 1349 11874 1421 11875
rect 1348 11866 1447 11874
rect 1348 11863 1400 11866
rect 1348 11828 1356 11863
rect 1381 11828 1400 11863
rect 1425 11855 1447 11866
rect 2398 11867 3737 11875
rect 2398 11864 2450 11867
rect 1425 11854 2292 11855
rect 1425 11828 2293 11854
rect 1348 11818 2293 11828
rect 1348 11816 1447 11818
rect 436 11775 458 11793
rect 476 11775 495 11793
rect 436 11753 495 11775
rect 703 11789 1235 11794
rect 703 11769 1589 11789
rect 1609 11769 1612 11789
rect 2248 11785 2293 11818
rect 2398 11829 2406 11864
rect 2431 11829 2450 11864
rect 2475 11829 3737 11867
rect 2398 11820 3737 11829
rect 2398 11817 2487 11820
rect 3026 11818 3737 11820
rect 703 11765 1612 11769
rect 703 11718 746 11765
rect 1196 11764 1612 11765
rect 2244 11765 2637 11785
rect 2657 11765 2660 11785
rect 1196 11763 1537 11764
rect 853 11732 963 11746
rect 853 11729 896 11732
rect 853 11724 857 11729
rect 691 11717 746 11718
rect 435 11694 746 11717
rect 435 11676 460 11694
rect 478 11682 746 11694
rect 775 11702 857 11724
rect 886 11702 896 11729
rect 924 11705 931 11732
rect 960 11724 963 11732
rect 960 11705 1025 11724
rect 924 11702 1025 11705
rect 775 11700 1025 11702
rect 478 11676 500 11682
rect 435 11537 500 11676
rect 775 11621 812 11700
rect 853 11687 963 11700
rect 927 11631 958 11632
rect 775 11601 784 11621
rect 804 11601 812 11621
rect 435 11519 458 11537
rect 476 11519 500 11537
rect 435 11502 500 11519
rect 655 11583 723 11596
rect 775 11591 812 11601
rect 871 11621 958 11631
rect 871 11601 880 11621
rect 900 11601 958 11621
rect 871 11592 958 11601
rect 871 11591 908 11592
rect 655 11541 662 11583
rect 711 11541 723 11583
rect 655 11538 723 11541
rect 927 11539 958 11592
rect 988 11621 1025 11700
rect 1140 11631 1171 11632
rect 988 11601 997 11621
rect 1017 11601 1025 11621
rect 988 11591 1025 11601
rect 1084 11624 1171 11631
rect 1084 11621 1145 11624
rect 1084 11601 1093 11621
rect 1113 11604 1145 11621
rect 1166 11604 1171 11624
rect 1113 11601 1171 11604
rect 1084 11594 1171 11601
rect 1196 11621 1233 11763
rect 1499 11762 1536 11763
rect 2244 11760 2660 11765
rect 2244 11759 2585 11760
rect 1901 11728 2011 11742
rect 1901 11725 1944 11728
rect 1901 11720 1905 11725
rect 1823 11698 1905 11720
rect 1934 11698 1944 11725
rect 1972 11701 1979 11728
rect 2008 11720 2011 11728
rect 2008 11701 2073 11720
rect 1972 11698 2073 11701
rect 1823 11696 2073 11698
rect 1348 11631 1384 11632
rect 1196 11601 1205 11621
rect 1225 11601 1233 11621
rect 1084 11592 1140 11594
rect 1084 11591 1121 11592
rect 1196 11591 1233 11601
rect 1292 11621 1440 11631
rect 1540 11628 1636 11630
rect 1292 11601 1301 11621
rect 1321 11601 1411 11621
rect 1431 11601 1440 11621
rect 1292 11595 1440 11601
rect 1292 11592 1356 11595
rect 1292 11591 1329 11592
rect 1348 11565 1356 11592
rect 1377 11592 1440 11595
rect 1498 11621 1636 11628
rect 1498 11601 1507 11621
rect 1527 11601 1636 11621
rect 1498 11592 1636 11601
rect 1823 11617 1860 11696
rect 1901 11683 2011 11696
rect 1975 11627 2006 11628
rect 1823 11597 1832 11617
rect 1852 11597 1860 11617
rect 1377 11565 1384 11592
rect 1403 11591 1440 11592
rect 1499 11591 1536 11592
rect 1348 11540 1384 11565
rect 819 11538 860 11539
rect 655 11531 860 11538
rect 655 11520 829 11531
rect 655 11487 663 11520
rect 656 11478 663 11487
rect 712 11511 829 11520
rect 849 11511 860 11531
rect 712 11503 860 11511
rect 927 11535 1286 11539
rect 927 11530 1249 11535
rect 927 11506 1040 11530
rect 1064 11511 1249 11530
rect 1273 11511 1286 11535
rect 1064 11506 1286 11511
rect 927 11503 1286 11506
rect 1348 11503 1383 11540
rect 1451 11537 1551 11540
rect 1451 11533 1518 11537
rect 1451 11507 1463 11533
rect 1489 11511 1518 11533
rect 1544 11511 1551 11537
rect 1489 11507 1551 11511
rect 1451 11503 1551 11507
rect 712 11487 723 11503
rect 712 11478 720 11487
rect 927 11482 958 11503
rect 1348 11482 1384 11503
rect 770 11481 807 11482
rect 435 11438 500 11457
rect 435 11420 460 11438
rect 478 11420 500 11438
rect 435 11219 500 11420
rect 656 11294 720 11478
rect 769 11472 807 11481
rect 769 11452 778 11472
rect 798 11452 807 11472
rect 769 11444 807 11452
rect 873 11476 958 11482
rect 983 11481 1020 11482
rect 873 11456 881 11476
rect 901 11456 958 11476
rect 873 11448 958 11456
rect 982 11472 1020 11481
rect 982 11452 991 11472
rect 1011 11452 1020 11472
rect 873 11447 909 11448
rect 982 11444 1020 11452
rect 1086 11476 1171 11482
rect 1191 11481 1228 11482
rect 1086 11456 1094 11476
rect 1114 11475 1171 11476
rect 1114 11456 1143 11475
rect 1086 11455 1143 11456
rect 1164 11455 1171 11475
rect 1086 11448 1171 11455
rect 1190 11472 1228 11481
rect 1190 11452 1199 11472
rect 1219 11452 1228 11472
rect 1086 11447 1122 11448
rect 1190 11444 1228 11452
rect 1294 11476 1438 11482
rect 1294 11456 1302 11476
rect 1322 11456 1410 11476
rect 1430 11456 1438 11476
rect 1294 11448 1438 11456
rect 1294 11447 1330 11448
rect 1402 11447 1438 11448
rect 1504 11481 1541 11482
rect 1504 11480 1542 11481
rect 1504 11472 1568 11480
rect 1504 11452 1513 11472
rect 1533 11458 1568 11472
rect 1588 11458 1591 11478
rect 1533 11453 1591 11458
rect 1533 11452 1568 11453
rect 770 11415 807 11444
rect 771 11413 807 11415
rect 983 11413 1020 11444
rect 771 11391 1020 11413
rect 852 11385 963 11391
rect 852 11377 893 11385
rect 852 11357 860 11377
rect 879 11357 893 11377
rect 852 11355 893 11357
rect 921 11377 963 11385
rect 921 11357 937 11377
rect 956 11357 963 11377
rect 921 11355 963 11357
rect 852 11340 963 11355
rect 656 11284 724 11294
rect 656 11251 673 11284
rect 713 11251 724 11284
rect 656 11239 724 11251
rect 656 11237 720 11239
rect 1191 11220 1228 11444
rect 1504 11440 1568 11452
rect 1608 11222 1635 11592
rect 1823 11587 1860 11597
rect 1919 11617 2006 11627
rect 1919 11597 1928 11617
rect 1948 11597 2006 11617
rect 1919 11588 2006 11597
rect 1919 11587 1956 11588
rect 1699 11574 1769 11579
rect 1694 11568 1769 11574
rect 1694 11535 1702 11568
rect 1755 11535 1769 11568
rect 1975 11535 2006 11588
rect 2036 11617 2073 11696
rect 2188 11627 2219 11628
rect 2036 11597 2045 11617
rect 2065 11597 2073 11617
rect 2036 11587 2073 11597
rect 2132 11620 2219 11627
rect 2132 11617 2193 11620
rect 2132 11597 2141 11617
rect 2161 11600 2193 11617
rect 2214 11600 2219 11620
rect 2161 11597 2219 11600
rect 2132 11590 2219 11597
rect 2244 11617 2281 11759
rect 2547 11758 2584 11759
rect 2396 11627 2432 11628
rect 2244 11597 2253 11617
rect 2273 11597 2281 11617
rect 2132 11588 2188 11590
rect 2132 11587 2169 11588
rect 2244 11587 2281 11597
rect 2340 11617 2488 11627
rect 2588 11624 2684 11626
rect 2340 11597 2349 11617
rect 2369 11597 2459 11617
rect 2479 11597 2488 11617
rect 2340 11591 2488 11597
rect 2340 11588 2404 11591
rect 2340 11587 2377 11588
rect 2396 11561 2404 11588
rect 2425 11588 2488 11591
rect 2546 11617 2684 11624
rect 2546 11597 2555 11617
rect 2575 11597 2684 11617
rect 2546 11588 2684 11597
rect 2425 11561 2432 11588
rect 2451 11587 2488 11588
rect 2547 11587 2584 11588
rect 2396 11536 2432 11561
rect 1694 11534 1777 11535
rect 1867 11534 1908 11535
rect 1694 11527 1908 11534
rect 1694 11510 1877 11527
rect 1694 11477 1707 11510
rect 1760 11507 1877 11510
rect 1897 11507 1908 11527
rect 1760 11499 1908 11507
rect 1975 11531 2334 11535
rect 1975 11526 2297 11531
rect 1975 11502 2088 11526
rect 2112 11507 2297 11526
rect 2321 11507 2334 11531
rect 2112 11502 2334 11507
rect 1975 11499 2334 11502
rect 2396 11499 2431 11536
rect 2499 11533 2599 11536
rect 2499 11529 2566 11533
rect 2499 11503 2511 11529
rect 2537 11507 2566 11529
rect 2592 11507 2599 11533
rect 2537 11503 2599 11507
rect 2499 11499 2599 11503
rect 1760 11477 1777 11499
rect 1975 11478 2006 11499
rect 2396 11478 2432 11499
rect 1818 11477 1855 11478
rect 1694 11463 1777 11477
rect 1467 11220 1635 11222
rect 1191 11219 1635 11220
rect 435 11189 1635 11219
rect 1705 11253 1777 11463
rect 1817 11468 1855 11477
rect 1817 11448 1826 11468
rect 1846 11448 1855 11468
rect 1817 11440 1855 11448
rect 1921 11472 2006 11478
rect 2031 11477 2068 11478
rect 1921 11452 1929 11472
rect 1949 11452 2006 11472
rect 1921 11444 2006 11452
rect 2030 11468 2068 11477
rect 2030 11448 2039 11468
rect 2059 11448 2068 11468
rect 1921 11443 1957 11444
rect 2030 11440 2068 11448
rect 2134 11472 2219 11478
rect 2239 11477 2276 11478
rect 2134 11452 2142 11472
rect 2162 11471 2219 11472
rect 2162 11452 2191 11471
rect 2134 11451 2191 11452
rect 2212 11451 2219 11471
rect 2134 11444 2219 11451
rect 2238 11468 2276 11477
rect 2238 11448 2247 11468
rect 2267 11448 2276 11468
rect 2134 11443 2170 11444
rect 2238 11440 2276 11448
rect 2342 11472 2486 11478
rect 2342 11452 2350 11472
rect 2370 11452 2458 11472
rect 2478 11452 2486 11472
rect 2342 11444 2486 11452
rect 2342 11443 2378 11444
rect 2450 11443 2486 11444
rect 2552 11477 2589 11478
rect 2552 11476 2590 11477
rect 2552 11468 2616 11476
rect 2552 11448 2561 11468
rect 2581 11454 2616 11468
rect 2636 11454 2639 11474
rect 2581 11449 2639 11454
rect 2581 11448 2616 11449
rect 1818 11411 1855 11440
rect 1819 11409 1855 11411
rect 2031 11409 2068 11440
rect 1819 11387 2068 11409
rect 1900 11381 2011 11387
rect 1900 11373 1941 11381
rect 1900 11353 1908 11373
rect 1927 11353 1941 11373
rect 1900 11351 1941 11353
rect 1969 11373 2011 11381
rect 1969 11353 1985 11373
rect 2004 11353 2011 11373
rect 1969 11351 2011 11353
rect 1900 11336 2011 11351
rect 1705 11214 1724 11253
rect 1769 11214 1777 11253
rect 1705 11197 1777 11214
rect 2239 11241 2276 11440
rect 2552 11436 2616 11448
rect 2239 11235 2280 11241
rect 2656 11237 2683 11588
rect 2978 11575 3073 11601
rect 2814 11553 2878 11572
rect 2814 11514 2827 11553
rect 2861 11514 2878 11553
rect 2814 11495 2878 11514
rect 2515 11235 2683 11237
rect 2239 11209 2683 11235
rect 435 11142 500 11189
rect 435 11124 458 11142
rect 476 11124 500 11142
rect 1348 11169 1383 11171
rect 1348 11167 1452 11169
rect 2241 11167 2280 11209
rect 2515 11208 2683 11209
rect 1348 11160 2282 11167
rect 1348 11159 1399 11160
rect 1348 11139 1351 11159
rect 1376 11140 1399 11159
rect 1431 11140 2282 11160
rect 1376 11139 2282 11140
rect 1348 11132 2282 11139
rect 1621 11131 2282 11132
rect 435 11103 500 11124
rect 712 11114 752 11117
rect 712 11110 1615 11114
rect 712 11090 1589 11110
rect 1609 11090 1615 11110
rect 712 11087 1615 11090
rect 436 11043 501 11063
rect 436 11025 460 11043
rect 478 11025 501 11043
rect 436 10998 501 11025
rect 712 10998 752 11087
rect 1196 11085 1612 11087
rect 1196 11084 1537 11085
rect 853 11053 963 11067
rect 853 11050 896 11053
rect 853 11045 857 11050
rect 435 10963 752 10998
rect 775 11023 857 11045
rect 886 11023 896 11050
rect 924 11026 931 11053
rect 960 11045 963 11053
rect 960 11026 1025 11045
rect 924 11023 1025 11026
rect 775 11021 1025 11023
rect 436 10887 501 10963
rect 775 10942 812 11021
rect 853 11008 963 11021
rect 927 10952 958 10953
rect 775 10922 784 10942
rect 804 10922 812 10942
rect 775 10912 812 10922
rect 871 10942 958 10952
rect 871 10922 880 10942
rect 900 10922 958 10942
rect 871 10913 958 10922
rect 871 10912 908 10913
rect 436 10869 458 10887
rect 476 10869 501 10887
rect 436 10848 501 10869
rect 649 10867 714 10876
rect 649 10830 659 10867
rect 699 10859 714 10867
rect 927 10860 958 10913
rect 988 10942 1025 11021
rect 1140 10952 1171 10953
rect 988 10922 997 10942
rect 1017 10922 1025 10942
rect 988 10912 1025 10922
rect 1084 10945 1171 10952
rect 1084 10942 1145 10945
rect 1084 10922 1093 10942
rect 1113 10925 1145 10942
rect 1166 10925 1171 10945
rect 1113 10922 1171 10925
rect 1084 10915 1171 10922
rect 1196 10942 1233 11084
rect 1499 11083 1536 11084
rect 2816 11024 2878 11495
rect 2978 11534 3004 11575
rect 3040 11534 3073 11575
rect 2978 11238 3073 11534
rect 2978 11194 2993 11238
rect 3053 11194 3073 11238
rect 2978 11174 3073 11194
rect 3690 11105 3733 11818
rect 3690 11085 4084 11105
rect 4104 11085 4107 11105
rect 3691 11080 4107 11085
rect 3691 11079 4032 11080
rect 3348 11048 3458 11062
rect 3348 11045 3391 11048
rect 3348 11040 3352 11045
rect 2811 10972 2886 11024
rect 3270 11018 3352 11040
rect 3381 11018 3391 11045
rect 3419 11021 3426 11048
rect 3455 11040 3458 11048
rect 3455 11021 3520 11040
rect 3419 11018 3520 11021
rect 3270 11016 3520 11018
rect 3180 10972 3226 10973
rect 1348 10952 1384 10953
rect 1196 10922 1205 10942
rect 1225 10922 1233 10942
rect 1084 10913 1140 10915
rect 1084 10912 1121 10913
rect 1196 10912 1233 10922
rect 1292 10942 1440 10952
rect 1540 10949 1636 10951
rect 1292 10922 1301 10942
rect 1321 10922 1411 10942
rect 1431 10922 1440 10942
rect 1292 10916 1440 10922
rect 1292 10913 1356 10916
rect 1292 10912 1329 10913
rect 1348 10886 1356 10913
rect 1377 10913 1440 10916
rect 1498 10942 1636 10949
rect 1498 10922 1507 10942
rect 1527 10922 1636 10942
rect 1498 10913 1636 10922
rect 2811 10937 3226 10972
rect 1377 10886 1384 10913
rect 1403 10912 1440 10913
rect 1499 10912 1536 10913
rect 1348 10861 1384 10886
rect 819 10859 860 10860
rect 699 10852 860 10859
rect 699 10832 829 10852
rect 849 10832 860 10852
rect 699 10830 860 10832
rect 649 10824 860 10830
rect 927 10856 1286 10860
rect 927 10851 1249 10856
rect 927 10827 1040 10851
rect 1064 10832 1249 10851
rect 1273 10832 1286 10856
rect 1064 10827 1286 10832
rect 927 10824 1286 10827
rect 1348 10824 1383 10861
rect 1451 10858 1551 10861
rect 1451 10854 1518 10858
rect 1451 10828 1463 10854
rect 1489 10832 1518 10854
rect 1544 10832 1551 10858
rect 1489 10828 1551 10832
rect 1451 10824 1551 10828
rect 649 10811 716 10824
rect 441 10788 497 10808
rect 441 10770 460 10788
rect 478 10770 497 10788
rect 441 10657 497 10770
rect 649 10790 663 10811
rect 699 10790 716 10811
rect 927 10803 958 10824
rect 1348 10803 1384 10824
rect 770 10802 807 10803
rect 649 10783 716 10790
rect 769 10793 807 10802
rect 441 10519 496 10657
rect 649 10631 714 10783
rect 769 10773 778 10793
rect 798 10773 807 10793
rect 769 10765 807 10773
rect 873 10797 958 10803
rect 983 10802 1020 10803
rect 873 10777 881 10797
rect 901 10777 958 10797
rect 873 10769 958 10777
rect 982 10793 1020 10802
rect 982 10773 991 10793
rect 1011 10773 1020 10793
rect 873 10768 909 10769
rect 982 10765 1020 10773
rect 1086 10797 1171 10803
rect 1191 10802 1228 10803
rect 1086 10777 1094 10797
rect 1114 10796 1171 10797
rect 1114 10777 1143 10796
rect 1086 10776 1143 10777
rect 1164 10776 1171 10796
rect 1086 10769 1171 10776
rect 1190 10793 1228 10802
rect 1190 10773 1199 10793
rect 1219 10773 1228 10793
rect 1086 10768 1122 10769
rect 1190 10765 1228 10773
rect 1294 10797 1438 10803
rect 1294 10777 1302 10797
rect 1322 10777 1410 10797
rect 1430 10777 1438 10797
rect 1294 10769 1438 10777
rect 1294 10768 1330 10769
rect 1402 10768 1438 10769
rect 1504 10802 1541 10803
rect 1504 10801 1542 10802
rect 1504 10793 1568 10801
rect 1504 10773 1513 10793
rect 1533 10779 1568 10793
rect 1588 10779 1591 10799
rect 1533 10774 1591 10779
rect 1533 10773 1568 10774
rect 770 10736 807 10765
rect 771 10734 807 10736
rect 983 10734 1020 10765
rect 771 10712 1020 10734
rect 852 10706 963 10712
rect 852 10698 893 10706
rect 852 10678 860 10698
rect 879 10678 893 10698
rect 852 10676 893 10678
rect 921 10698 963 10706
rect 921 10678 937 10698
rect 956 10678 963 10698
rect 921 10676 963 10678
rect 852 10663 963 10676
rect 1191 10666 1228 10765
rect 1504 10761 1568 10773
rect 642 10621 763 10631
rect 642 10619 711 10621
rect 642 10578 655 10619
rect 692 10580 711 10619
rect 748 10580 763 10621
rect 692 10578 763 10580
rect 642 10560 763 10578
rect 434 10516 498 10519
rect 854 10516 958 10522
rect 1189 10516 1230 10666
rect 1608 10658 1635 10913
rect 1697 10903 1777 10914
rect 1697 10877 1714 10903
rect 1754 10877 1777 10903
rect 1697 10850 1777 10877
rect 1697 10824 1718 10850
rect 1758 10824 1777 10850
rect 1697 10805 1777 10824
rect 1697 10779 1721 10805
rect 1761 10779 1777 10805
rect 1697 10728 1777 10779
rect 434 10513 1230 10516
rect 1609 10527 1635 10658
rect 1609 10513 1637 10527
rect 434 10478 1637 10513
rect 1699 10520 1769 10728
rect 2811 10653 2886 10937
rect 3180 10854 3226 10937
rect 3270 10937 3307 11016
rect 3348 11003 3458 11016
rect 3422 10947 3453 10948
rect 3270 10917 3279 10937
rect 3299 10917 3307 10937
rect 3270 10907 3307 10917
rect 3366 10937 3453 10947
rect 3366 10917 3375 10937
rect 3395 10917 3453 10937
rect 3366 10908 3453 10917
rect 3366 10907 3403 10908
rect 3422 10855 3453 10908
rect 3483 10937 3520 11016
rect 3635 10947 3666 10948
rect 3483 10917 3492 10937
rect 3512 10917 3520 10937
rect 3483 10907 3520 10917
rect 3579 10940 3666 10947
rect 3579 10937 3640 10940
rect 3579 10917 3588 10937
rect 3608 10920 3640 10937
rect 3661 10920 3666 10940
rect 3608 10917 3666 10920
rect 3579 10910 3666 10917
rect 3691 10937 3728 11079
rect 3994 11078 4031 11079
rect 3843 10947 3879 10948
rect 3691 10917 3700 10937
rect 3720 10917 3728 10937
rect 3579 10908 3635 10910
rect 3579 10907 3616 10908
rect 3691 10907 3728 10917
rect 3787 10937 3935 10947
rect 4035 10944 4131 10946
rect 3787 10917 3796 10937
rect 3816 10917 3906 10937
rect 3926 10917 3935 10937
rect 3787 10911 3935 10917
rect 3787 10908 3851 10911
rect 3787 10907 3824 10908
rect 3843 10881 3851 10908
rect 3872 10908 3935 10911
rect 3993 10937 4131 10944
rect 3993 10917 4002 10937
rect 4022 10917 4131 10937
rect 3993 10908 4131 10917
rect 3872 10881 3879 10908
rect 3898 10907 3935 10908
rect 3994 10907 4031 10908
rect 3843 10856 3879 10881
rect 3314 10854 3355 10855
rect 3180 10847 3355 10854
rect 2978 10821 3064 10840
rect 2978 10780 2993 10821
rect 3047 10780 3064 10821
rect 3180 10827 3324 10847
rect 3344 10827 3355 10847
rect 3180 10819 3355 10827
rect 3422 10851 3781 10855
rect 3422 10846 3744 10851
rect 3422 10822 3535 10846
rect 3559 10827 3744 10846
rect 3768 10827 3781 10851
rect 3559 10822 3781 10827
rect 3422 10819 3781 10822
rect 3843 10819 3878 10856
rect 3946 10853 4046 10856
rect 3946 10849 4013 10853
rect 3946 10823 3958 10849
rect 3984 10827 4013 10849
rect 4039 10827 4046 10853
rect 3984 10823 4046 10827
rect 3946 10819 4046 10823
rect 3180 10815 3226 10819
rect 3422 10798 3453 10819
rect 3843 10798 3879 10819
rect 3265 10797 3302 10798
rect 2978 10744 3064 10780
rect 3264 10788 3302 10797
rect 3264 10768 3273 10788
rect 3293 10768 3302 10788
rect 3264 10760 3302 10768
rect 3368 10792 3453 10798
rect 3478 10797 3515 10798
rect 3368 10772 3376 10792
rect 3396 10772 3453 10792
rect 3368 10764 3453 10772
rect 3477 10788 3515 10797
rect 3477 10768 3486 10788
rect 3506 10768 3515 10788
rect 3368 10763 3404 10764
rect 3477 10760 3515 10768
rect 3581 10792 3666 10798
rect 3686 10797 3723 10798
rect 3581 10772 3589 10792
rect 3609 10791 3666 10792
rect 3609 10772 3638 10791
rect 3581 10771 3638 10772
rect 3659 10771 3666 10791
rect 3581 10764 3666 10771
rect 3685 10788 3723 10797
rect 3685 10768 3694 10788
rect 3714 10768 3723 10788
rect 3581 10763 3617 10764
rect 3685 10760 3723 10768
rect 3789 10792 3933 10798
rect 3789 10772 3797 10792
rect 3817 10772 3905 10792
rect 3925 10772 3933 10792
rect 3789 10764 3933 10772
rect 3789 10763 3825 10764
rect 434 10417 498 10478
rect 854 10476 958 10478
rect 1189 10476 1230 10478
rect 1699 10475 1720 10520
rect 1700 10454 1720 10475
rect 1750 10475 1769 10520
rect 2806 10611 2886 10653
rect 1750 10454 1767 10475
rect 1700 10435 1767 10454
rect 1349 10427 1421 10428
rect 1348 10419 1447 10427
rect 436 10346 495 10417
rect 1348 10416 1400 10419
rect 1348 10381 1356 10416
rect 1381 10381 1400 10416
rect 1425 10408 1447 10419
rect 1425 10407 2292 10408
rect 1425 10381 2293 10407
rect 1348 10371 2293 10381
rect 1348 10369 1447 10371
rect 436 10328 458 10346
rect 476 10328 495 10346
rect 436 10306 495 10328
rect 703 10342 1235 10347
rect 703 10322 1589 10342
rect 1609 10322 1612 10342
rect 2248 10338 2293 10371
rect 703 10318 1612 10322
rect 703 10271 746 10318
rect 1196 10317 1612 10318
rect 2244 10318 2637 10338
rect 2657 10318 2660 10338
rect 1196 10316 1537 10317
rect 853 10285 963 10299
rect 853 10282 896 10285
rect 853 10277 857 10282
rect 691 10270 746 10271
rect 435 10247 746 10270
rect 435 10229 460 10247
rect 478 10235 746 10247
rect 775 10255 857 10277
rect 886 10255 896 10282
rect 924 10258 931 10285
rect 960 10277 963 10285
rect 960 10258 1025 10277
rect 924 10255 1025 10258
rect 775 10253 1025 10255
rect 478 10229 500 10235
rect 435 10090 500 10229
rect 775 10174 812 10253
rect 853 10240 963 10253
rect 927 10184 958 10185
rect 775 10154 784 10174
rect 804 10154 812 10174
rect 435 10072 458 10090
rect 476 10072 500 10090
rect 435 10055 500 10072
rect 655 10136 723 10149
rect 775 10144 812 10154
rect 871 10174 958 10184
rect 871 10154 880 10174
rect 900 10154 958 10174
rect 871 10145 958 10154
rect 871 10144 908 10145
rect 655 10094 662 10136
rect 711 10094 723 10136
rect 655 10091 723 10094
rect 927 10092 958 10145
rect 988 10174 1025 10253
rect 1140 10184 1171 10185
rect 988 10154 997 10174
rect 1017 10154 1025 10174
rect 988 10144 1025 10154
rect 1084 10177 1171 10184
rect 1084 10174 1145 10177
rect 1084 10154 1093 10174
rect 1113 10157 1145 10174
rect 1166 10157 1171 10177
rect 1113 10154 1171 10157
rect 1084 10147 1171 10154
rect 1196 10174 1233 10316
rect 1499 10315 1536 10316
rect 2244 10313 2660 10318
rect 2244 10312 2585 10313
rect 1901 10281 2011 10295
rect 1901 10278 1944 10281
rect 1901 10273 1905 10278
rect 1823 10251 1905 10273
rect 1934 10251 1944 10278
rect 1972 10254 1979 10281
rect 2008 10273 2011 10281
rect 2008 10254 2073 10273
rect 1972 10251 2073 10254
rect 1823 10249 2073 10251
rect 1348 10184 1384 10185
rect 1196 10154 1205 10174
rect 1225 10154 1233 10174
rect 1084 10145 1140 10147
rect 1084 10144 1121 10145
rect 1196 10144 1233 10154
rect 1292 10174 1440 10184
rect 1540 10181 1636 10183
rect 1292 10154 1301 10174
rect 1321 10154 1411 10174
rect 1431 10154 1440 10174
rect 1292 10148 1440 10154
rect 1292 10145 1356 10148
rect 1292 10144 1329 10145
rect 1348 10118 1356 10145
rect 1377 10145 1440 10148
rect 1498 10174 1636 10181
rect 1498 10154 1507 10174
rect 1527 10154 1636 10174
rect 1498 10145 1636 10154
rect 1823 10170 1860 10249
rect 1901 10236 2011 10249
rect 1975 10180 2006 10181
rect 1823 10150 1832 10170
rect 1852 10150 1860 10170
rect 1377 10118 1384 10145
rect 1403 10144 1440 10145
rect 1499 10144 1536 10145
rect 1348 10093 1384 10118
rect 819 10091 860 10092
rect 655 10084 860 10091
rect 655 10073 829 10084
rect 655 10040 663 10073
rect 656 10031 663 10040
rect 712 10064 829 10073
rect 849 10064 860 10084
rect 712 10056 860 10064
rect 927 10088 1286 10092
rect 927 10083 1249 10088
rect 927 10059 1040 10083
rect 1064 10064 1249 10083
rect 1273 10064 1286 10088
rect 1064 10059 1286 10064
rect 927 10056 1286 10059
rect 1348 10056 1383 10093
rect 1451 10090 1551 10093
rect 1451 10086 1518 10090
rect 1451 10060 1463 10086
rect 1489 10064 1518 10086
rect 1544 10064 1551 10090
rect 1489 10060 1551 10064
rect 1451 10056 1551 10060
rect 712 10040 723 10056
rect 712 10031 720 10040
rect 927 10035 958 10056
rect 1348 10035 1384 10056
rect 770 10034 807 10035
rect 435 9991 500 10010
rect 435 9973 460 9991
rect 478 9973 500 9991
rect 435 9772 500 9973
rect 656 9847 720 10031
rect 769 10025 807 10034
rect 769 10005 778 10025
rect 798 10005 807 10025
rect 769 9997 807 10005
rect 873 10029 958 10035
rect 983 10034 1020 10035
rect 873 10009 881 10029
rect 901 10009 958 10029
rect 873 10001 958 10009
rect 982 10025 1020 10034
rect 982 10005 991 10025
rect 1011 10005 1020 10025
rect 873 10000 909 10001
rect 982 9997 1020 10005
rect 1086 10029 1171 10035
rect 1191 10034 1228 10035
rect 1086 10009 1094 10029
rect 1114 10028 1171 10029
rect 1114 10009 1143 10028
rect 1086 10008 1143 10009
rect 1164 10008 1171 10028
rect 1086 10001 1171 10008
rect 1190 10025 1228 10034
rect 1190 10005 1199 10025
rect 1219 10005 1228 10025
rect 1086 10000 1122 10001
rect 1190 9997 1228 10005
rect 1294 10029 1438 10035
rect 1294 10009 1302 10029
rect 1322 10009 1410 10029
rect 1430 10009 1438 10029
rect 1294 10001 1438 10009
rect 1294 10000 1330 10001
rect 1402 10000 1438 10001
rect 1504 10034 1541 10035
rect 1504 10033 1542 10034
rect 1504 10025 1568 10033
rect 1504 10005 1513 10025
rect 1533 10011 1568 10025
rect 1588 10011 1591 10031
rect 1533 10006 1591 10011
rect 1533 10005 1568 10006
rect 770 9968 807 9997
rect 771 9966 807 9968
rect 983 9966 1020 9997
rect 771 9944 1020 9966
rect 852 9938 963 9944
rect 852 9930 893 9938
rect 852 9910 860 9930
rect 879 9910 893 9930
rect 852 9908 893 9910
rect 921 9930 963 9938
rect 921 9910 937 9930
rect 956 9910 963 9930
rect 921 9908 963 9910
rect 852 9893 963 9908
rect 656 9837 724 9847
rect 656 9804 673 9837
rect 713 9804 724 9837
rect 656 9792 724 9804
rect 656 9790 720 9792
rect 1191 9773 1228 9997
rect 1504 9993 1568 10005
rect 1608 9775 1635 10145
rect 1823 10140 1860 10150
rect 1919 10170 2006 10180
rect 1919 10150 1928 10170
rect 1948 10150 2006 10170
rect 1919 10141 2006 10150
rect 1919 10140 1956 10141
rect 1699 10127 1769 10132
rect 1694 10121 1769 10127
rect 1694 10088 1702 10121
rect 1755 10088 1769 10121
rect 1975 10088 2006 10141
rect 2036 10170 2073 10249
rect 2188 10180 2219 10181
rect 2036 10150 2045 10170
rect 2065 10150 2073 10170
rect 2036 10140 2073 10150
rect 2132 10173 2219 10180
rect 2132 10170 2193 10173
rect 2132 10150 2141 10170
rect 2161 10153 2193 10170
rect 2214 10153 2219 10173
rect 2161 10150 2219 10153
rect 2132 10143 2219 10150
rect 2244 10170 2281 10312
rect 2547 10311 2584 10312
rect 2396 10180 2432 10181
rect 2244 10150 2253 10170
rect 2273 10150 2281 10170
rect 2132 10141 2188 10143
rect 2132 10140 2169 10141
rect 2244 10140 2281 10150
rect 2340 10170 2488 10180
rect 2588 10177 2684 10179
rect 2340 10150 2349 10170
rect 2369 10150 2459 10170
rect 2479 10150 2488 10170
rect 2340 10144 2488 10150
rect 2340 10141 2404 10144
rect 2340 10140 2377 10141
rect 2396 10114 2404 10141
rect 2425 10141 2488 10144
rect 2546 10170 2684 10177
rect 2546 10150 2555 10170
rect 2575 10150 2684 10170
rect 2546 10141 2684 10150
rect 2425 10114 2432 10141
rect 2451 10140 2488 10141
rect 2547 10140 2584 10141
rect 2396 10089 2432 10114
rect 1694 10087 1777 10088
rect 1867 10087 1908 10088
rect 1694 10080 1908 10087
rect 1694 10063 1877 10080
rect 1694 10030 1707 10063
rect 1760 10060 1877 10063
rect 1897 10060 1908 10080
rect 1760 10052 1908 10060
rect 1975 10084 2334 10088
rect 1975 10079 2297 10084
rect 1975 10055 2088 10079
rect 2112 10060 2297 10079
rect 2321 10060 2334 10084
rect 2112 10055 2334 10060
rect 1975 10052 2334 10055
rect 2396 10052 2431 10089
rect 2499 10086 2599 10089
rect 2499 10082 2566 10086
rect 2499 10056 2511 10082
rect 2537 10060 2566 10082
rect 2592 10060 2599 10086
rect 2537 10056 2599 10060
rect 2499 10052 2599 10056
rect 1760 10030 1777 10052
rect 1975 10031 2006 10052
rect 2396 10031 2432 10052
rect 1818 10030 1855 10031
rect 1694 10016 1777 10030
rect 1467 9773 1635 9775
rect 1191 9772 1635 9773
rect 435 9742 1635 9772
rect 1705 9806 1777 10016
rect 1817 10021 1855 10030
rect 1817 10001 1826 10021
rect 1846 10001 1855 10021
rect 1817 9993 1855 10001
rect 1921 10025 2006 10031
rect 2031 10030 2068 10031
rect 1921 10005 1929 10025
rect 1949 10005 2006 10025
rect 1921 9997 2006 10005
rect 2030 10021 2068 10030
rect 2030 10001 2039 10021
rect 2059 10001 2068 10021
rect 1921 9996 1957 9997
rect 2030 9993 2068 10001
rect 2134 10025 2219 10031
rect 2239 10030 2276 10031
rect 2134 10005 2142 10025
rect 2162 10024 2219 10025
rect 2162 10005 2191 10024
rect 2134 10004 2191 10005
rect 2212 10004 2219 10024
rect 2134 9997 2219 10004
rect 2238 10021 2276 10030
rect 2238 10001 2247 10021
rect 2267 10001 2276 10021
rect 2134 9996 2170 9997
rect 2238 9993 2276 10001
rect 2342 10025 2486 10031
rect 2342 10005 2350 10025
rect 2370 10005 2458 10025
rect 2478 10005 2486 10025
rect 2342 9997 2486 10005
rect 2342 9996 2378 9997
rect 2450 9996 2486 9997
rect 2552 10030 2589 10031
rect 2552 10029 2590 10030
rect 2552 10021 2616 10029
rect 2552 10001 2561 10021
rect 2581 10007 2616 10021
rect 2636 10007 2639 10027
rect 2581 10002 2639 10007
rect 2581 10001 2616 10002
rect 1818 9964 1855 9993
rect 1819 9962 1855 9964
rect 2031 9962 2068 9993
rect 1819 9940 2068 9962
rect 1900 9934 2011 9940
rect 1900 9926 1941 9934
rect 1900 9906 1908 9926
rect 1927 9906 1941 9926
rect 1900 9904 1941 9906
rect 1969 9926 2011 9934
rect 1969 9906 1985 9926
rect 2004 9906 2011 9926
rect 1969 9904 2011 9906
rect 1900 9889 2011 9904
rect 1705 9767 1724 9806
rect 1769 9767 1777 9806
rect 1705 9750 1777 9767
rect 2239 9794 2276 9993
rect 2552 9989 2616 10001
rect 2239 9788 2280 9794
rect 2656 9790 2683 10141
rect 2806 10011 2885 10611
rect 2982 10159 3061 10744
rect 3265 10731 3302 10760
rect 3266 10729 3302 10731
rect 3478 10729 3515 10760
rect 3266 10707 3515 10729
rect 3347 10701 3458 10707
rect 3347 10693 3388 10701
rect 3347 10673 3355 10693
rect 3374 10673 3388 10693
rect 3347 10671 3388 10673
rect 3416 10693 3458 10701
rect 3416 10673 3432 10693
rect 3451 10673 3458 10693
rect 3416 10671 3458 10673
rect 3347 10656 3458 10671
rect 3686 10645 3723 10760
rect 3679 10533 3726 10645
rect 3847 10605 3877 10764
rect 3897 10763 3933 10764
rect 3999 10797 4036 10798
rect 3999 10796 4037 10797
rect 3999 10788 4063 10796
rect 3999 10768 4008 10788
rect 4028 10774 4063 10788
rect 4083 10774 4086 10794
rect 4028 10769 4086 10774
rect 4028 10768 4063 10769
rect 3999 10756 4063 10768
rect 3847 10601 3933 10605
rect 3847 10583 3862 10601
rect 3914 10583 3933 10601
rect 3847 10574 3933 10583
rect 4103 10535 4130 10908
rect 3962 10533 4130 10535
rect 3679 10507 4130 10533
rect 3679 10429 3726 10507
rect 3962 10506 4130 10507
rect 3624 10428 3726 10429
rect 3623 10420 3726 10428
rect 3623 10417 3675 10420
rect 3623 10382 3631 10417
rect 3656 10382 3675 10417
rect 3700 10382 3726 10420
rect 3623 10376 3726 10382
rect 3886 10421 3922 10425
rect 3886 10398 3894 10421
rect 3918 10398 3922 10421
rect 3886 10377 3922 10398
rect 3623 10372 3722 10376
rect 3886 10354 3894 10377
rect 3918 10354 3922 10377
rect 2515 9788 2683 9790
rect 2239 9762 2683 9788
rect 435 9695 500 9742
rect 435 9677 458 9695
rect 476 9677 500 9695
rect 1348 9722 1383 9724
rect 1348 9720 1452 9722
rect 2241 9720 2280 9762
rect 2515 9761 2683 9762
rect 1348 9713 2282 9720
rect 1348 9712 1399 9713
rect 1348 9692 1351 9712
rect 1376 9693 1399 9712
rect 1431 9693 2282 9713
rect 1376 9692 2282 9693
rect 1348 9685 2282 9692
rect 1621 9684 2282 9685
rect 435 9656 500 9677
rect 712 9667 752 9670
rect 712 9663 1615 9667
rect 712 9643 1589 9663
rect 1609 9643 1615 9663
rect 712 9640 1615 9643
rect 436 9596 501 9616
rect 436 9578 460 9596
rect 478 9578 501 9596
rect 436 9551 501 9578
rect 712 9551 752 9640
rect 1196 9638 1612 9640
rect 1196 9637 1537 9638
rect 853 9606 963 9620
rect 853 9603 896 9606
rect 853 9598 857 9603
rect 435 9516 752 9551
rect 775 9576 857 9598
rect 886 9576 896 9603
rect 924 9579 931 9606
rect 960 9598 963 9606
rect 960 9579 1025 9598
rect 924 9576 1025 9579
rect 775 9574 1025 9576
rect 436 9440 501 9516
rect 775 9495 812 9574
rect 853 9561 963 9574
rect 927 9505 958 9506
rect 775 9475 784 9495
rect 804 9475 812 9495
rect 775 9465 812 9475
rect 871 9495 958 9505
rect 871 9475 880 9495
rect 900 9475 958 9495
rect 871 9466 958 9475
rect 871 9465 908 9466
rect 436 9422 458 9440
rect 476 9422 501 9440
rect 436 9401 501 9422
rect 649 9420 714 9429
rect 649 9383 659 9420
rect 699 9412 714 9420
rect 927 9413 958 9466
rect 988 9495 1025 9574
rect 1140 9505 1171 9506
rect 988 9475 997 9495
rect 1017 9475 1025 9495
rect 988 9465 1025 9475
rect 1084 9498 1171 9505
rect 1084 9495 1145 9498
rect 1084 9475 1093 9495
rect 1113 9478 1145 9495
rect 1166 9478 1171 9498
rect 1113 9475 1171 9478
rect 1084 9468 1171 9475
rect 1196 9495 1233 9637
rect 1499 9636 1536 9637
rect 1348 9505 1384 9506
rect 1196 9475 1205 9495
rect 1225 9475 1233 9495
rect 1084 9466 1140 9468
rect 1084 9465 1121 9466
rect 1196 9465 1233 9475
rect 1292 9495 1440 9505
rect 1540 9502 1636 9504
rect 1292 9475 1301 9495
rect 1321 9475 1411 9495
rect 1431 9475 1440 9495
rect 1292 9469 1440 9475
rect 1292 9466 1356 9469
rect 1292 9465 1329 9466
rect 1348 9439 1356 9466
rect 1377 9466 1440 9469
rect 1498 9495 1636 9502
rect 1498 9475 1507 9495
rect 1527 9475 1636 9495
rect 1498 9466 1636 9475
rect 1377 9439 1384 9466
rect 1403 9465 1440 9466
rect 1499 9465 1536 9466
rect 1348 9414 1384 9439
rect 819 9412 860 9413
rect 699 9405 860 9412
rect 699 9385 829 9405
rect 849 9385 860 9405
rect 699 9383 860 9385
rect 649 9377 860 9383
rect 927 9409 1286 9413
rect 927 9404 1249 9409
rect 927 9380 1040 9404
rect 1064 9385 1249 9404
rect 1273 9385 1286 9409
rect 1064 9380 1286 9385
rect 927 9377 1286 9380
rect 1348 9377 1383 9414
rect 1451 9411 1551 9414
rect 1451 9407 1518 9411
rect 1451 9381 1463 9407
rect 1489 9385 1518 9407
rect 1544 9385 1551 9411
rect 1489 9381 1551 9385
rect 1451 9377 1551 9381
rect 649 9364 716 9377
rect 441 9341 497 9361
rect 441 9323 460 9341
rect 478 9323 497 9341
rect 441 9210 497 9323
rect 649 9343 663 9364
rect 699 9343 716 9364
rect 927 9356 958 9377
rect 1348 9356 1384 9377
rect 770 9355 807 9356
rect 649 9336 716 9343
rect 769 9346 807 9355
rect 441 9081 496 9210
rect 649 9184 714 9336
rect 769 9326 778 9346
rect 798 9326 807 9346
rect 769 9318 807 9326
rect 873 9350 958 9356
rect 983 9355 1020 9356
rect 873 9330 881 9350
rect 901 9330 958 9350
rect 873 9322 958 9330
rect 982 9346 1020 9355
rect 982 9326 991 9346
rect 1011 9326 1020 9346
rect 873 9321 909 9322
rect 982 9318 1020 9326
rect 1086 9350 1171 9356
rect 1191 9355 1228 9356
rect 1086 9330 1094 9350
rect 1114 9349 1171 9350
rect 1114 9330 1143 9349
rect 1086 9329 1143 9330
rect 1164 9329 1171 9349
rect 1086 9322 1171 9329
rect 1190 9346 1228 9355
rect 1190 9326 1199 9346
rect 1219 9326 1228 9346
rect 1086 9321 1122 9322
rect 1190 9318 1228 9326
rect 1294 9350 1438 9356
rect 1294 9330 1302 9350
rect 1322 9330 1410 9350
rect 1430 9330 1438 9350
rect 1294 9322 1438 9330
rect 1294 9321 1330 9322
rect 1402 9321 1438 9322
rect 1504 9355 1541 9356
rect 1504 9354 1542 9355
rect 1504 9346 1568 9354
rect 1504 9326 1513 9346
rect 1533 9332 1568 9346
rect 1588 9332 1591 9352
rect 1533 9327 1591 9332
rect 1533 9326 1568 9327
rect 770 9289 807 9318
rect 771 9287 807 9289
rect 983 9287 1020 9318
rect 771 9265 1020 9287
rect 852 9259 963 9265
rect 852 9251 893 9259
rect 852 9231 860 9251
rect 879 9231 893 9251
rect 852 9229 893 9231
rect 921 9251 963 9259
rect 921 9231 937 9251
rect 956 9231 963 9251
rect 921 9229 963 9231
rect 852 9214 963 9229
rect 1191 9219 1228 9318
rect 1504 9314 1568 9326
rect 854 9205 958 9214
rect 642 9174 763 9184
rect 642 9172 711 9174
rect 642 9131 655 9172
rect 692 9133 711 9172
rect 748 9133 763 9174
rect 692 9131 763 9133
rect 642 9113 763 9131
rect 435 9069 496 9081
rect 1189 9069 1230 9219
rect 1608 9211 1635 9466
rect 1697 9456 1777 9467
rect 1697 9430 1714 9456
rect 1754 9430 1777 9456
rect 1697 9403 1777 9430
rect 1697 9377 1718 9403
rect 1758 9377 1777 9403
rect 1697 9358 1777 9377
rect 1697 9332 1721 9358
rect 1761 9332 1777 9358
rect 1697 9281 1777 9332
rect 435 9066 1230 9069
rect 1609 9080 1635 9211
rect 1699 9125 1769 9281
rect 1698 9109 1774 9125
rect 1609 9066 1637 9080
rect 435 9031 1637 9066
rect 1698 9072 1713 9109
rect 1757 9072 1774 9109
rect 1698 9052 1774 9072
rect 2812 9102 2882 10011
rect 2981 9446 3062 10159
rect 3886 10045 3922 10354
rect 3810 10016 3923 10045
rect 3810 9660 3841 10016
rect 3880 9761 4871 9786
rect 3880 9756 3940 9761
rect 3880 9735 3899 9756
rect 3919 9740 3940 9756
rect 3960 9740 4871 9761
rect 3919 9735 4871 9740
rect 3880 9727 4871 9735
rect 3885 9704 3991 9727
rect 3885 9701 3990 9704
rect 3734 9640 4127 9660
rect 4147 9640 4150 9660
rect 3734 9635 4150 9640
rect 3734 9634 4075 9635
rect 3391 9603 3501 9617
rect 3391 9600 3434 9603
rect 3391 9595 3395 9600
rect 3313 9573 3395 9595
rect 3424 9573 3434 9600
rect 3462 9576 3469 9603
rect 3498 9595 3501 9603
rect 3498 9576 3563 9595
rect 3462 9573 3563 9576
rect 3313 9571 3563 9573
rect 3313 9492 3350 9571
rect 3391 9558 3501 9571
rect 3465 9502 3496 9503
rect 3313 9472 3322 9492
rect 3342 9472 3350 9492
rect 3313 9462 3350 9472
rect 3409 9492 3496 9502
rect 3409 9472 3418 9492
rect 3438 9472 3496 9492
rect 3409 9463 3496 9472
rect 3409 9462 3446 9463
rect 2979 9410 3071 9446
rect 3465 9410 3496 9463
rect 3526 9492 3563 9571
rect 3678 9502 3709 9503
rect 3526 9472 3535 9492
rect 3555 9472 3563 9492
rect 3526 9462 3563 9472
rect 3622 9495 3709 9502
rect 3622 9492 3683 9495
rect 3622 9472 3631 9492
rect 3651 9475 3683 9492
rect 3704 9475 3709 9495
rect 3651 9472 3709 9475
rect 3622 9465 3709 9472
rect 3734 9492 3771 9634
rect 4037 9633 4074 9634
rect 3886 9502 3922 9503
rect 3734 9472 3743 9492
rect 3763 9472 3771 9492
rect 3622 9463 3678 9465
rect 3622 9462 3659 9463
rect 3734 9462 3771 9472
rect 3830 9492 3978 9502
rect 4078 9499 4174 9501
rect 3830 9472 3839 9492
rect 3859 9472 3949 9492
rect 3969 9472 3978 9492
rect 3830 9466 3978 9472
rect 3830 9463 3894 9466
rect 3830 9462 3867 9463
rect 3886 9436 3894 9463
rect 3915 9463 3978 9466
rect 4036 9492 4174 9499
rect 4036 9472 4045 9492
rect 4065 9472 4174 9492
rect 4036 9463 4174 9472
rect 3915 9436 3922 9463
rect 3941 9462 3978 9463
rect 4037 9462 4074 9463
rect 3886 9411 3922 9436
rect 2979 9409 3315 9410
rect 3357 9409 3398 9410
rect 2979 9402 3398 9409
rect 2979 9382 3367 9402
rect 3387 9382 3398 9402
rect 2979 9374 3398 9382
rect 3465 9406 3824 9410
rect 3465 9401 3787 9406
rect 3465 9377 3578 9401
rect 3602 9382 3787 9401
rect 3811 9382 3824 9406
rect 3602 9377 3824 9382
rect 3465 9374 3824 9377
rect 3886 9374 3921 9411
rect 3989 9408 4089 9411
rect 3989 9404 4056 9408
rect 3989 9378 4001 9404
rect 4027 9382 4056 9404
rect 4082 9382 4089 9408
rect 4027 9378 4089 9382
rect 3989 9374 4089 9378
rect 2979 9370 3315 9374
rect 2812 9052 2884 9102
rect 435 8956 496 9031
rect 854 9029 958 9031
rect 1189 9029 1230 9031
rect 1698 8986 1708 9052
rect 1762 8986 1774 9052
rect 1698 8962 1774 8986
rect 437 8826 496 8956
rect 1350 8907 1422 8908
rect 1349 8899 1448 8907
rect 1349 8896 1401 8899
rect 1349 8861 1357 8896
rect 1382 8861 1401 8896
rect 1426 8888 1448 8899
rect 1426 8887 2293 8888
rect 1426 8861 2294 8887
rect 1349 8851 2294 8861
rect 1349 8849 1448 8851
rect 437 8808 459 8826
rect 477 8808 496 8826
rect 437 8786 496 8808
rect 704 8822 1236 8827
rect 704 8802 1590 8822
rect 1610 8802 1613 8822
rect 2249 8818 2294 8851
rect 704 8798 1613 8802
rect 704 8751 747 8798
rect 1197 8797 1613 8798
rect 2245 8798 2638 8818
rect 2658 8798 2661 8818
rect 1197 8796 1538 8797
rect 854 8765 964 8779
rect 854 8762 897 8765
rect 854 8757 858 8762
rect 692 8750 747 8751
rect 436 8727 747 8750
rect 436 8709 461 8727
rect 479 8715 747 8727
rect 776 8735 858 8757
rect 887 8735 897 8762
rect 925 8738 932 8765
rect 961 8757 964 8765
rect 961 8738 1026 8757
rect 925 8735 1026 8738
rect 776 8733 1026 8735
rect 479 8709 501 8715
rect 436 8570 501 8709
rect 776 8654 813 8733
rect 854 8720 964 8733
rect 928 8664 959 8665
rect 776 8634 785 8654
rect 805 8634 813 8654
rect 436 8552 459 8570
rect 477 8552 501 8570
rect 436 8535 501 8552
rect 656 8616 724 8629
rect 776 8624 813 8634
rect 872 8654 959 8664
rect 872 8634 881 8654
rect 901 8634 959 8654
rect 872 8625 959 8634
rect 872 8624 909 8625
rect 656 8574 663 8616
rect 712 8574 724 8616
rect 656 8571 724 8574
rect 928 8572 959 8625
rect 989 8654 1026 8733
rect 1141 8664 1172 8665
rect 989 8634 998 8654
rect 1018 8634 1026 8654
rect 989 8624 1026 8634
rect 1085 8657 1172 8664
rect 1085 8654 1146 8657
rect 1085 8634 1094 8654
rect 1114 8637 1146 8654
rect 1167 8637 1172 8657
rect 1114 8634 1172 8637
rect 1085 8627 1172 8634
rect 1197 8654 1234 8796
rect 1500 8795 1537 8796
rect 2245 8793 2661 8798
rect 2245 8792 2586 8793
rect 1902 8761 2012 8775
rect 1902 8758 1945 8761
rect 1902 8753 1906 8758
rect 1824 8731 1906 8753
rect 1935 8731 1945 8758
rect 1973 8734 1980 8761
rect 2009 8753 2012 8761
rect 2009 8734 2074 8753
rect 1973 8731 2074 8734
rect 1824 8729 2074 8731
rect 1349 8664 1385 8665
rect 1197 8634 1206 8654
rect 1226 8634 1234 8654
rect 1085 8625 1141 8627
rect 1085 8624 1122 8625
rect 1197 8624 1234 8634
rect 1293 8654 1441 8664
rect 1541 8661 1637 8663
rect 1293 8634 1302 8654
rect 1322 8634 1412 8654
rect 1432 8634 1441 8654
rect 1293 8628 1441 8634
rect 1293 8625 1357 8628
rect 1293 8624 1330 8625
rect 1349 8598 1357 8625
rect 1378 8625 1441 8628
rect 1499 8654 1637 8661
rect 1499 8634 1508 8654
rect 1528 8634 1637 8654
rect 1499 8625 1637 8634
rect 1824 8650 1861 8729
rect 1902 8716 2012 8729
rect 1976 8660 2007 8661
rect 1824 8630 1833 8650
rect 1853 8630 1861 8650
rect 1378 8598 1385 8625
rect 1404 8624 1441 8625
rect 1500 8624 1537 8625
rect 1349 8573 1385 8598
rect 820 8571 861 8572
rect 656 8564 861 8571
rect 656 8553 830 8564
rect 656 8520 664 8553
rect 657 8511 664 8520
rect 713 8544 830 8553
rect 850 8544 861 8564
rect 713 8536 861 8544
rect 928 8568 1287 8572
rect 928 8563 1250 8568
rect 928 8539 1041 8563
rect 1065 8544 1250 8563
rect 1274 8544 1287 8568
rect 1065 8539 1287 8544
rect 928 8536 1287 8539
rect 1349 8536 1384 8573
rect 1452 8570 1552 8573
rect 1452 8566 1519 8570
rect 1452 8540 1464 8566
rect 1490 8544 1519 8566
rect 1545 8544 1552 8570
rect 1490 8540 1552 8544
rect 1452 8536 1552 8540
rect 713 8520 724 8536
rect 713 8511 721 8520
rect 928 8515 959 8536
rect 1349 8515 1385 8536
rect 771 8514 808 8515
rect 436 8471 501 8490
rect 436 8453 461 8471
rect 479 8453 501 8471
rect 436 8252 501 8453
rect 657 8327 721 8511
rect 770 8505 808 8514
rect 770 8485 779 8505
rect 799 8485 808 8505
rect 770 8477 808 8485
rect 874 8509 959 8515
rect 984 8514 1021 8515
rect 874 8489 882 8509
rect 902 8489 959 8509
rect 874 8481 959 8489
rect 983 8505 1021 8514
rect 983 8485 992 8505
rect 1012 8485 1021 8505
rect 874 8480 910 8481
rect 983 8477 1021 8485
rect 1087 8509 1172 8515
rect 1192 8514 1229 8515
rect 1087 8489 1095 8509
rect 1115 8508 1172 8509
rect 1115 8489 1144 8508
rect 1087 8488 1144 8489
rect 1165 8488 1172 8508
rect 1087 8481 1172 8488
rect 1191 8505 1229 8514
rect 1191 8485 1200 8505
rect 1220 8485 1229 8505
rect 1087 8480 1123 8481
rect 1191 8477 1229 8485
rect 1295 8509 1439 8515
rect 1295 8489 1303 8509
rect 1323 8489 1411 8509
rect 1431 8489 1439 8509
rect 1295 8481 1439 8489
rect 1295 8480 1331 8481
rect 1403 8480 1439 8481
rect 1505 8514 1542 8515
rect 1505 8513 1543 8514
rect 1505 8505 1569 8513
rect 1505 8485 1514 8505
rect 1534 8491 1569 8505
rect 1589 8491 1592 8511
rect 1534 8486 1592 8491
rect 1534 8485 1569 8486
rect 771 8448 808 8477
rect 772 8446 808 8448
rect 984 8446 1021 8477
rect 772 8424 1021 8446
rect 853 8418 964 8424
rect 853 8410 894 8418
rect 853 8390 861 8410
rect 880 8390 894 8410
rect 853 8388 894 8390
rect 922 8410 964 8418
rect 922 8390 938 8410
rect 957 8390 964 8410
rect 922 8388 964 8390
rect 853 8373 964 8388
rect 657 8317 725 8327
rect 657 8284 674 8317
rect 714 8284 725 8317
rect 657 8272 725 8284
rect 657 8270 721 8272
rect 1192 8253 1229 8477
rect 1505 8473 1569 8485
rect 1609 8255 1636 8625
rect 1824 8620 1861 8630
rect 1920 8650 2007 8660
rect 1920 8630 1929 8650
rect 1949 8630 2007 8650
rect 1920 8621 2007 8630
rect 1920 8620 1957 8621
rect 1700 8607 1770 8612
rect 1695 8601 1770 8607
rect 1695 8568 1703 8601
rect 1756 8568 1770 8601
rect 1976 8568 2007 8621
rect 2037 8650 2074 8729
rect 2189 8660 2220 8661
rect 2037 8630 2046 8650
rect 2066 8630 2074 8650
rect 2037 8620 2074 8630
rect 2133 8653 2220 8660
rect 2133 8650 2194 8653
rect 2133 8630 2142 8650
rect 2162 8633 2194 8650
rect 2215 8633 2220 8653
rect 2162 8630 2220 8633
rect 2133 8623 2220 8630
rect 2245 8650 2282 8792
rect 2548 8791 2585 8792
rect 2397 8660 2433 8661
rect 2245 8630 2254 8650
rect 2274 8630 2282 8650
rect 2133 8621 2189 8623
rect 2133 8620 2170 8621
rect 2245 8620 2282 8630
rect 2341 8650 2489 8660
rect 2589 8657 2685 8659
rect 2341 8630 2350 8650
rect 2370 8630 2460 8650
rect 2480 8630 2489 8650
rect 2341 8624 2489 8630
rect 2341 8621 2405 8624
rect 2341 8620 2378 8621
rect 2397 8594 2405 8621
rect 2426 8621 2489 8624
rect 2547 8650 2685 8657
rect 2547 8630 2556 8650
rect 2576 8630 2685 8650
rect 2547 8621 2685 8630
rect 2426 8594 2433 8621
rect 2452 8620 2489 8621
rect 2548 8620 2585 8621
rect 2397 8569 2433 8594
rect 1695 8567 1778 8568
rect 1868 8567 1909 8568
rect 1695 8560 1909 8567
rect 1695 8543 1878 8560
rect 1695 8510 1708 8543
rect 1761 8540 1878 8543
rect 1898 8540 1909 8560
rect 1761 8532 1909 8540
rect 1976 8564 2335 8568
rect 1976 8559 2298 8564
rect 1976 8535 2089 8559
rect 2113 8540 2298 8559
rect 2322 8540 2335 8564
rect 2113 8535 2335 8540
rect 1976 8532 2335 8535
rect 2397 8532 2432 8569
rect 2500 8566 2600 8569
rect 2500 8562 2567 8566
rect 2500 8536 2512 8562
rect 2538 8540 2567 8562
rect 2593 8540 2600 8566
rect 2538 8536 2600 8540
rect 2500 8532 2600 8536
rect 1761 8510 1778 8532
rect 1976 8511 2007 8532
rect 2397 8511 2433 8532
rect 1819 8510 1856 8511
rect 1695 8496 1778 8510
rect 1468 8253 1636 8255
rect 1192 8252 1636 8253
rect 436 8222 1636 8252
rect 1706 8286 1778 8496
rect 1818 8501 1856 8510
rect 1818 8481 1827 8501
rect 1847 8481 1856 8501
rect 1818 8473 1856 8481
rect 1922 8505 2007 8511
rect 2032 8510 2069 8511
rect 1922 8485 1930 8505
rect 1950 8485 2007 8505
rect 1922 8477 2007 8485
rect 2031 8501 2069 8510
rect 2031 8481 2040 8501
rect 2060 8481 2069 8501
rect 1922 8476 1958 8477
rect 2031 8473 2069 8481
rect 2135 8505 2220 8511
rect 2240 8510 2277 8511
rect 2135 8485 2143 8505
rect 2163 8504 2220 8505
rect 2163 8485 2192 8504
rect 2135 8484 2192 8485
rect 2213 8484 2220 8504
rect 2135 8477 2220 8484
rect 2239 8501 2277 8510
rect 2239 8481 2248 8501
rect 2268 8481 2277 8501
rect 2135 8476 2171 8477
rect 2239 8473 2277 8481
rect 2343 8505 2487 8511
rect 2343 8485 2351 8505
rect 2371 8485 2459 8505
rect 2479 8485 2487 8505
rect 2343 8477 2487 8485
rect 2343 8476 2379 8477
rect 2451 8476 2487 8477
rect 2553 8510 2590 8511
rect 2553 8509 2591 8510
rect 2553 8501 2617 8509
rect 2553 8481 2562 8501
rect 2582 8487 2617 8501
rect 2637 8487 2640 8507
rect 2582 8482 2640 8487
rect 2582 8481 2617 8482
rect 1819 8444 1856 8473
rect 1820 8442 1856 8444
rect 2032 8442 2069 8473
rect 1820 8420 2069 8442
rect 1901 8414 2012 8420
rect 1901 8406 1942 8414
rect 1901 8386 1909 8406
rect 1928 8386 1942 8406
rect 1901 8384 1942 8386
rect 1970 8406 2012 8414
rect 1970 8386 1986 8406
rect 2005 8386 2012 8406
rect 1970 8384 2012 8386
rect 1901 8369 2012 8384
rect 1706 8247 1725 8286
rect 1770 8247 1778 8286
rect 1706 8230 1778 8247
rect 2240 8274 2277 8473
rect 2553 8469 2617 8481
rect 2240 8268 2281 8274
rect 2657 8270 2684 8621
rect 2813 8573 2884 9052
rect 2813 8489 2882 8573
rect 2516 8268 2684 8270
rect 2240 8242 2684 8268
rect 436 8175 501 8222
rect 436 8157 459 8175
rect 477 8157 501 8175
rect 1349 8202 1384 8204
rect 1349 8200 1453 8202
rect 2242 8200 2281 8242
rect 2516 8241 2684 8242
rect 1349 8193 2283 8200
rect 1349 8192 1400 8193
rect 1349 8172 1352 8192
rect 1377 8173 1400 8192
rect 1432 8173 2283 8193
rect 1377 8172 2283 8173
rect 1349 8165 2283 8172
rect 1622 8164 2283 8165
rect 436 8136 501 8157
rect 713 8147 753 8150
rect 713 8143 1616 8147
rect 713 8123 1590 8143
rect 1610 8123 1616 8143
rect 713 8120 1616 8123
rect 437 8076 502 8096
rect 437 8058 461 8076
rect 479 8058 502 8076
rect 437 8031 502 8058
rect 713 8031 753 8120
rect 1197 8118 1613 8120
rect 1197 8117 1538 8118
rect 854 8086 964 8100
rect 854 8083 897 8086
rect 854 8078 858 8083
rect 436 7996 753 8031
rect 776 8056 858 8078
rect 887 8056 897 8083
rect 925 8059 932 8086
rect 961 8078 964 8086
rect 961 8059 1026 8078
rect 925 8056 1026 8059
rect 776 8054 1026 8056
rect 437 7920 502 7996
rect 776 7975 813 8054
rect 854 8041 964 8054
rect 928 7985 959 7986
rect 776 7955 785 7975
rect 805 7955 813 7975
rect 776 7945 813 7955
rect 872 7975 959 7985
rect 872 7955 881 7975
rect 901 7955 959 7975
rect 872 7946 959 7955
rect 872 7945 909 7946
rect 437 7902 459 7920
rect 477 7902 502 7920
rect 437 7881 502 7902
rect 650 7900 715 7909
rect 650 7863 660 7900
rect 700 7892 715 7900
rect 928 7893 959 7946
rect 989 7975 1026 8054
rect 1141 7985 1172 7986
rect 989 7955 998 7975
rect 1018 7955 1026 7975
rect 989 7945 1026 7955
rect 1085 7978 1172 7985
rect 1085 7975 1146 7978
rect 1085 7955 1094 7975
rect 1114 7958 1146 7975
rect 1167 7958 1172 7978
rect 1114 7955 1172 7958
rect 1085 7948 1172 7955
rect 1197 7975 1234 8117
rect 1500 8116 1537 8117
rect 1349 7985 1385 7986
rect 1197 7955 1206 7975
rect 1226 7955 1234 7975
rect 1085 7946 1141 7948
rect 1085 7945 1122 7946
rect 1197 7945 1234 7955
rect 1293 7975 1441 7985
rect 1541 7982 1637 7984
rect 1293 7955 1302 7975
rect 1322 7955 1412 7975
rect 1432 7955 1441 7975
rect 1293 7949 1441 7955
rect 1293 7946 1357 7949
rect 1293 7945 1330 7946
rect 1349 7919 1357 7946
rect 1378 7946 1441 7949
rect 1499 7975 1637 7982
rect 1499 7955 1508 7975
rect 1528 7955 1637 7975
rect 2817 7973 2879 8489
rect 1499 7946 1637 7955
rect 1378 7919 1385 7946
rect 1404 7945 1441 7946
rect 1500 7945 1537 7946
rect 1349 7894 1385 7919
rect 820 7892 861 7893
rect 700 7885 861 7892
rect 700 7865 830 7885
rect 850 7865 861 7885
rect 700 7863 861 7865
rect 650 7857 861 7863
rect 928 7889 1287 7893
rect 928 7884 1250 7889
rect 928 7860 1041 7884
rect 1065 7865 1250 7884
rect 1274 7865 1287 7889
rect 1065 7860 1287 7865
rect 928 7857 1287 7860
rect 1349 7857 1384 7894
rect 1452 7891 1552 7894
rect 1452 7887 1519 7891
rect 1452 7861 1464 7887
rect 1490 7865 1519 7887
rect 1545 7865 1552 7891
rect 1490 7861 1552 7865
rect 1452 7857 1552 7861
rect 650 7844 717 7857
rect 442 7821 498 7841
rect 442 7803 461 7821
rect 479 7803 498 7821
rect 442 7690 498 7803
rect 650 7823 664 7844
rect 700 7823 717 7844
rect 928 7836 959 7857
rect 1349 7836 1385 7857
rect 771 7835 808 7836
rect 650 7816 717 7823
rect 770 7826 808 7835
rect 442 7552 497 7690
rect 650 7664 715 7816
rect 770 7806 779 7826
rect 799 7806 808 7826
rect 770 7798 808 7806
rect 874 7830 959 7836
rect 984 7835 1021 7836
rect 874 7810 882 7830
rect 902 7810 959 7830
rect 874 7802 959 7810
rect 983 7826 1021 7835
rect 983 7806 992 7826
rect 1012 7806 1021 7826
rect 874 7801 910 7802
rect 983 7798 1021 7806
rect 1087 7830 1172 7836
rect 1192 7835 1229 7836
rect 1087 7810 1095 7830
rect 1115 7829 1172 7830
rect 1115 7810 1144 7829
rect 1087 7809 1144 7810
rect 1165 7809 1172 7829
rect 1087 7802 1172 7809
rect 1191 7826 1229 7835
rect 1191 7806 1200 7826
rect 1220 7806 1229 7826
rect 1087 7801 1123 7802
rect 1191 7798 1229 7806
rect 1295 7830 1439 7836
rect 1295 7810 1303 7830
rect 1323 7810 1411 7830
rect 1431 7810 1439 7830
rect 1295 7802 1439 7810
rect 1295 7801 1331 7802
rect 1403 7801 1439 7802
rect 1505 7835 1542 7836
rect 1505 7834 1543 7835
rect 1505 7826 1569 7834
rect 1505 7806 1514 7826
rect 1534 7812 1569 7826
rect 1589 7812 1592 7832
rect 1534 7807 1592 7812
rect 1534 7806 1569 7807
rect 771 7769 808 7798
rect 772 7767 808 7769
rect 984 7767 1021 7798
rect 772 7745 1021 7767
rect 853 7739 964 7745
rect 853 7731 894 7739
rect 853 7711 861 7731
rect 880 7711 894 7731
rect 853 7709 894 7711
rect 922 7731 964 7739
rect 922 7711 938 7731
rect 957 7711 964 7731
rect 922 7709 964 7711
rect 853 7696 964 7709
rect 1192 7699 1229 7798
rect 1505 7794 1569 7806
rect 643 7654 764 7664
rect 643 7652 712 7654
rect 643 7611 656 7652
rect 693 7613 712 7652
rect 749 7613 764 7654
rect 693 7611 764 7613
rect 643 7593 764 7611
rect 435 7549 499 7552
rect 855 7549 959 7555
rect 1190 7549 1231 7699
rect 1609 7691 1636 7946
rect 1698 7936 1778 7947
rect 1698 7910 1715 7936
rect 1755 7910 1778 7936
rect 1698 7883 1778 7910
rect 1698 7857 1719 7883
rect 1759 7857 1778 7883
rect 1698 7838 1778 7857
rect 1698 7812 1722 7838
rect 1762 7812 1778 7838
rect 1698 7761 1778 7812
rect 2801 7938 2879 7973
rect 2801 7876 2883 7938
rect 2801 7853 2829 7876
rect 2855 7853 2883 7876
rect 2801 7833 2883 7853
rect 435 7546 1231 7549
rect 1610 7560 1636 7691
rect 1610 7546 1638 7560
rect 435 7511 1638 7546
rect 1700 7553 1770 7761
rect 435 7450 499 7511
rect 855 7509 959 7511
rect 1190 7509 1231 7511
rect 1700 7508 1721 7553
rect 1701 7487 1721 7508
rect 1751 7508 1770 7553
rect 1751 7487 1768 7508
rect 1701 7468 1768 7487
rect 1350 7460 1422 7461
rect 1349 7452 1448 7460
rect 437 7379 496 7450
rect 1349 7449 1401 7452
rect 1349 7414 1357 7449
rect 1382 7414 1401 7449
rect 1426 7441 1448 7452
rect 1426 7440 2293 7441
rect 1426 7414 2294 7440
rect 1349 7404 2294 7414
rect 1349 7402 1448 7404
rect 437 7361 459 7379
rect 477 7361 496 7379
rect 437 7339 496 7361
rect 704 7375 1236 7380
rect 704 7355 1590 7375
rect 1610 7355 1613 7375
rect 2249 7371 2294 7404
rect 704 7351 1613 7355
rect 704 7304 747 7351
rect 1197 7350 1613 7351
rect 2245 7351 2638 7371
rect 2658 7351 2661 7371
rect 1197 7349 1538 7350
rect 854 7318 964 7332
rect 854 7315 897 7318
rect 854 7310 858 7315
rect 692 7303 747 7304
rect 436 7280 747 7303
rect 436 7262 461 7280
rect 479 7268 747 7280
rect 776 7288 858 7310
rect 887 7288 897 7315
rect 925 7291 932 7318
rect 961 7310 964 7318
rect 961 7291 1026 7310
rect 925 7288 1026 7291
rect 776 7286 1026 7288
rect 479 7262 501 7268
rect 436 7123 501 7262
rect 776 7207 813 7286
rect 854 7273 964 7286
rect 928 7217 959 7218
rect 776 7187 785 7207
rect 805 7187 813 7207
rect 436 7105 459 7123
rect 477 7105 501 7123
rect 436 7088 501 7105
rect 656 7169 724 7182
rect 776 7177 813 7187
rect 872 7207 959 7217
rect 872 7187 881 7207
rect 901 7187 959 7207
rect 872 7178 959 7187
rect 872 7177 909 7178
rect 656 7127 663 7169
rect 712 7127 724 7169
rect 656 7124 724 7127
rect 928 7125 959 7178
rect 989 7207 1026 7286
rect 1141 7217 1172 7218
rect 989 7187 998 7207
rect 1018 7187 1026 7207
rect 989 7177 1026 7187
rect 1085 7210 1172 7217
rect 1085 7207 1146 7210
rect 1085 7187 1094 7207
rect 1114 7190 1146 7207
rect 1167 7190 1172 7210
rect 1114 7187 1172 7190
rect 1085 7180 1172 7187
rect 1197 7207 1234 7349
rect 1500 7348 1537 7349
rect 2245 7346 2661 7351
rect 2245 7345 2586 7346
rect 1902 7314 2012 7328
rect 1902 7311 1945 7314
rect 1902 7306 1906 7311
rect 1824 7284 1906 7306
rect 1935 7284 1945 7311
rect 1973 7287 1980 7314
rect 2009 7306 2012 7314
rect 2009 7287 2074 7306
rect 1973 7284 2074 7287
rect 1824 7282 2074 7284
rect 1349 7217 1385 7218
rect 1197 7187 1206 7207
rect 1226 7187 1234 7207
rect 1085 7178 1141 7180
rect 1085 7177 1122 7178
rect 1197 7177 1234 7187
rect 1293 7207 1441 7217
rect 1541 7214 1637 7216
rect 1293 7187 1302 7207
rect 1322 7187 1412 7207
rect 1432 7187 1441 7207
rect 1293 7181 1441 7187
rect 1293 7178 1357 7181
rect 1293 7177 1330 7178
rect 1349 7151 1357 7178
rect 1378 7178 1441 7181
rect 1499 7207 1637 7214
rect 1499 7187 1508 7207
rect 1528 7187 1637 7207
rect 1499 7178 1637 7187
rect 1824 7203 1861 7282
rect 1902 7269 2012 7282
rect 1976 7213 2007 7214
rect 1824 7183 1833 7203
rect 1853 7183 1861 7203
rect 1378 7151 1385 7178
rect 1404 7177 1441 7178
rect 1500 7177 1537 7178
rect 1349 7126 1385 7151
rect 820 7124 861 7125
rect 656 7117 861 7124
rect 656 7106 830 7117
rect 656 7073 664 7106
rect 657 7064 664 7073
rect 713 7097 830 7106
rect 850 7097 861 7117
rect 713 7089 861 7097
rect 928 7121 1287 7125
rect 928 7116 1250 7121
rect 928 7092 1041 7116
rect 1065 7097 1250 7116
rect 1274 7097 1287 7121
rect 1065 7092 1287 7097
rect 928 7089 1287 7092
rect 1349 7089 1384 7126
rect 1452 7123 1552 7126
rect 1452 7119 1519 7123
rect 1452 7093 1464 7119
rect 1490 7097 1519 7119
rect 1545 7097 1552 7123
rect 1490 7093 1552 7097
rect 1452 7089 1552 7093
rect 713 7073 724 7089
rect 713 7064 721 7073
rect 928 7068 959 7089
rect 1349 7068 1385 7089
rect 771 7067 808 7068
rect 436 7024 501 7043
rect 436 7006 461 7024
rect 479 7006 501 7024
rect 436 6805 501 7006
rect 657 6880 721 7064
rect 770 7058 808 7067
rect 770 7038 779 7058
rect 799 7038 808 7058
rect 770 7030 808 7038
rect 874 7062 959 7068
rect 984 7067 1021 7068
rect 874 7042 882 7062
rect 902 7042 959 7062
rect 874 7034 959 7042
rect 983 7058 1021 7067
rect 983 7038 992 7058
rect 1012 7038 1021 7058
rect 874 7033 910 7034
rect 983 7030 1021 7038
rect 1087 7062 1172 7068
rect 1192 7067 1229 7068
rect 1087 7042 1095 7062
rect 1115 7061 1172 7062
rect 1115 7042 1144 7061
rect 1087 7041 1144 7042
rect 1165 7041 1172 7061
rect 1087 7034 1172 7041
rect 1191 7058 1229 7067
rect 1191 7038 1200 7058
rect 1220 7038 1229 7058
rect 1087 7033 1123 7034
rect 1191 7030 1229 7038
rect 1295 7062 1439 7068
rect 1295 7042 1303 7062
rect 1323 7042 1411 7062
rect 1431 7042 1439 7062
rect 1295 7034 1439 7042
rect 1295 7033 1331 7034
rect 1403 7033 1439 7034
rect 1505 7067 1542 7068
rect 1505 7066 1543 7067
rect 1505 7058 1569 7066
rect 1505 7038 1514 7058
rect 1534 7044 1569 7058
rect 1589 7044 1592 7064
rect 1534 7039 1592 7044
rect 1534 7038 1569 7039
rect 771 7001 808 7030
rect 772 6999 808 7001
rect 984 6999 1021 7030
rect 772 6977 1021 6999
rect 853 6971 964 6977
rect 853 6963 894 6971
rect 853 6943 861 6963
rect 880 6943 894 6963
rect 853 6941 894 6943
rect 922 6963 964 6971
rect 922 6943 938 6963
rect 957 6943 964 6963
rect 922 6941 964 6943
rect 853 6926 964 6941
rect 657 6870 725 6880
rect 657 6837 674 6870
rect 714 6837 725 6870
rect 657 6825 725 6837
rect 657 6823 721 6825
rect 1192 6806 1229 7030
rect 1505 7026 1569 7038
rect 1609 6808 1636 7178
rect 1824 7173 1861 7183
rect 1920 7203 2007 7213
rect 1920 7183 1929 7203
rect 1949 7183 2007 7203
rect 1920 7174 2007 7183
rect 1920 7173 1957 7174
rect 1700 7160 1770 7165
rect 1695 7154 1770 7160
rect 1695 7121 1703 7154
rect 1756 7121 1770 7154
rect 1976 7121 2007 7174
rect 2037 7203 2074 7282
rect 2189 7213 2220 7214
rect 2037 7183 2046 7203
rect 2066 7183 2074 7203
rect 2037 7173 2074 7183
rect 2133 7206 2220 7213
rect 2133 7203 2194 7206
rect 2133 7183 2142 7203
rect 2162 7186 2194 7203
rect 2215 7186 2220 7206
rect 2162 7183 2220 7186
rect 2133 7176 2220 7183
rect 2245 7203 2282 7345
rect 2548 7344 2585 7345
rect 2397 7213 2433 7214
rect 2245 7183 2254 7203
rect 2274 7183 2282 7203
rect 2133 7174 2189 7176
rect 2133 7173 2170 7174
rect 2245 7173 2282 7183
rect 2341 7203 2489 7213
rect 2589 7210 2685 7212
rect 2341 7183 2350 7203
rect 2370 7183 2460 7203
rect 2480 7183 2489 7203
rect 2341 7177 2489 7183
rect 2341 7174 2405 7177
rect 2341 7173 2378 7174
rect 2397 7147 2405 7174
rect 2426 7174 2489 7177
rect 2547 7203 2685 7210
rect 2547 7183 2556 7203
rect 2576 7183 2685 7203
rect 2547 7174 2685 7183
rect 2426 7147 2433 7174
rect 2452 7173 2489 7174
rect 2548 7173 2585 7174
rect 2397 7122 2433 7147
rect 1695 7120 1778 7121
rect 1868 7120 1909 7121
rect 1695 7113 1909 7120
rect 1695 7096 1878 7113
rect 1695 7063 1708 7096
rect 1761 7093 1878 7096
rect 1898 7093 1909 7113
rect 1761 7085 1909 7093
rect 1976 7117 2335 7121
rect 1976 7112 2298 7117
rect 1976 7088 2089 7112
rect 2113 7093 2298 7112
rect 2322 7093 2335 7117
rect 2113 7088 2335 7093
rect 1976 7085 2335 7088
rect 2397 7085 2432 7122
rect 2500 7119 2600 7122
rect 2500 7115 2567 7119
rect 2500 7089 2512 7115
rect 2538 7093 2567 7115
rect 2593 7093 2600 7119
rect 2538 7089 2600 7093
rect 2500 7085 2600 7089
rect 1761 7063 1778 7085
rect 1976 7064 2007 7085
rect 2397 7064 2433 7085
rect 1819 7063 1856 7064
rect 1695 7049 1778 7063
rect 1468 6806 1636 6808
rect 1192 6805 1636 6806
rect 436 6775 1636 6805
rect 1706 6839 1778 7049
rect 1818 7054 1856 7063
rect 1818 7034 1827 7054
rect 1847 7034 1856 7054
rect 1818 7026 1856 7034
rect 1922 7058 2007 7064
rect 2032 7063 2069 7064
rect 1922 7038 1930 7058
rect 1950 7038 2007 7058
rect 1922 7030 2007 7038
rect 2031 7054 2069 7063
rect 2031 7034 2040 7054
rect 2060 7034 2069 7054
rect 1922 7029 1958 7030
rect 2031 7026 2069 7034
rect 2135 7058 2220 7064
rect 2240 7063 2277 7064
rect 2135 7038 2143 7058
rect 2163 7057 2220 7058
rect 2163 7038 2192 7057
rect 2135 7037 2192 7038
rect 2213 7037 2220 7057
rect 2135 7030 2220 7037
rect 2239 7054 2277 7063
rect 2239 7034 2248 7054
rect 2268 7034 2277 7054
rect 2135 7029 2171 7030
rect 2239 7026 2277 7034
rect 2343 7058 2487 7064
rect 2343 7038 2351 7058
rect 2371 7038 2459 7058
rect 2479 7038 2487 7058
rect 2343 7030 2487 7038
rect 2343 7029 2379 7030
rect 2451 7029 2487 7030
rect 2553 7063 2590 7064
rect 2553 7062 2591 7063
rect 2553 7054 2617 7062
rect 2553 7034 2562 7054
rect 2582 7040 2617 7054
rect 2637 7040 2640 7060
rect 2582 7035 2640 7040
rect 2582 7034 2617 7035
rect 1819 6997 1856 7026
rect 1820 6995 1856 6997
rect 2032 6995 2069 7026
rect 1820 6973 2069 6995
rect 1901 6967 2012 6973
rect 1901 6959 1942 6967
rect 1901 6939 1909 6959
rect 1928 6939 1942 6959
rect 1901 6937 1942 6939
rect 1970 6959 2012 6967
rect 1970 6939 1986 6959
rect 2005 6939 2012 6959
rect 1970 6937 2012 6939
rect 1901 6922 2012 6937
rect 1706 6800 1725 6839
rect 1770 6800 1778 6839
rect 1706 6783 1778 6800
rect 2240 6827 2277 7026
rect 2553 7022 2617 7034
rect 2240 6821 2281 6827
rect 2657 6823 2684 7174
rect 2516 6821 2684 6823
rect 2240 6795 2684 6821
rect 436 6728 501 6775
rect 436 6710 459 6728
rect 477 6710 501 6728
rect 1349 6755 1384 6757
rect 1349 6753 1453 6755
rect 2242 6753 2281 6795
rect 2516 6794 2684 6795
rect 1349 6746 2283 6753
rect 1349 6745 1400 6746
rect 1349 6725 1352 6745
rect 1377 6726 1400 6745
rect 1432 6726 2283 6746
rect 1377 6725 2283 6726
rect 1349 6718 2283 6725
rect 1622 6717 2283 6718
rect 436 6689 501 6710
rect 713 6700 753 6703
rect 713 6696 1616 6700
rect 713 6676 1590 6696
rect 1610 6676 1616 6696
rect 713 6673 1616 6676
rect 437 6629 502 6649
rect 437 6611 461 6629
rect 479 6611 502 6629
rect 437 6584 502 6611
rect 713 6584 753 6673
rect 1197 6671 1613 6673
rect 1197 6670 1538 6671
rect 854 6639 964 6653
rect 854 6636 897 6639
rect 854 6631 858 6636
rect 436 6549 753 6584
rect 776 6609 858 6631
rect 887 6609 897 6636
rect 925 6612 932 6639
rect 961 6631 964 6639
rect 961 6612 1026 6631
rect 925 6609 1026 6612
rect 776 6607 1026 6609
rect 437 6473 502 6549
rect 776 6528 813 6607
rect 854 6594 964 6607
rect 928 6538 959 6539
rect 776 6508 785 6528
rect 805 6508 813 6528
rect 776 6498 813 6508
rect 872 6528 959 6538
rect 872 6508 881 6528
rect 901 6508 959 6528
rect 872 6499 959 6508
rect 872 6498 909 6499
rect 437 6455 459 6473
rect 477 6455 502 6473
rect 437 6434 502 6455
rect 650 6453 715 6462
rect 650 6416 660 6453
rect 700 6445 715 6453
rect 928 6446 959 6499
rect 989 6528 1026 6607
rect 1141 6538 1172 6539
rect 989 6508 998 6528
rect 1018 6508 1026 6528
rect 989 6498 1026 6508
rect 1085 6531 1172 6538
rect 1085 6528 1146 6531
rect 1085 6508 1094 6528
rect 1114 6511 1146 6528
rect 1167 6511 1172 6531
rect 1114 6508 1172 6511
rect 1085 6501 1172 6508
rect 1197 6528 1234 6670
rect 1500 6669 1537 6670
rect 1349 6538 1385 6539
rect 1197 6508 1206 6528
rect 1226 6508 1234 6528
rect 1085 6499 1141 6501
rect 1085 6498 1122 6499
rect 1197 6498 1234 6508
rect 1293 6528 1441 6538
rect 1541 6535 1637 6537
rect 1293 6508 1302 6528
rect 1322 6508 1412 6528
rect 1432 6508 1441 6528
rect 1293 6502 1441 6508
rect 1293 6499 1357 6502
rect 1293 6498 1330 6499
rect 1349 6472 1357 6499
rect 1378 6499 1441 6502
rect 1499 6528 1637 6535
rect 1499 6508 1508 6528
rect 1528 6508 1637 6528
rect 1499 6499 1637 6508
rect 1378 6472 1385 6499
rect 1404 6498 1441 6499
rect 1500 6498 1537 6499
rect 1349 6447 1385 6472
rect 820 6445 861 6446
rect 700 6438 861 6445
rect 700 6418 830 6438
rect 850 6418 861 6438
rect 700 6416 861 6418
rect 650 6410 861 6416
rect 928 6442 1287 6446
rect 928 6437 1250 6442
rect 928 6413 1041 6437
rect 1065 6418 1250 6437
rect 1274 6418 1287 6442
rect 1065 6413 1287 6418
rect 928 6410 1287 6413
rect 1349 6410 1384 6447
rect 1452 6444 1552 6447
rect 1452 6440 1519 6444
rect 1452 6414 1464 6440
rect 1490 6418 1519 6440
rect 1545 6418 1552 6444
rect 1490 6414 1552 6418
rect 1452 6410 1552 6414
rect 650 6397 717 6410
rect 442 6374 498 6394
rect 442 6356 461 6374
rect 479 6356 498 6374
rect 442 6243 498 6356
rect 650 6376 664 6397
rect 700 6376 717 6397
rect 928 6389 959 6410
rect 1349 6389 1385 6410
rect 771 6388 808 6389
rect 650 6369 717 6376
rect 770 6379 808 6388
rect 442 6136 497 6243
rect 650 6217 715 6369
rect 770 6359 779 6379
rect 799 6359 808 6379
rect 770 6351 808 6359
rect 874 6383 959 6389
rect 984 6388 1021 6389
rect 874 6363 882 6383
rect 902 6363 959 6383
rect 874 6355 959 6363
rect 983 6379 1021 6388
rect 983 6359 992 6379
rect 1012 6359 1021 6379
rect 874 6354 910 6355
rect 983 6351 1021 6359
rect 1087 6383 1172 6389
rect 1192 6388 1229 6389
rect 1087 6363 1095 6383
rect 1115 6382 1172 6383
rect 1115 6363 1144 6382
rect 1087 6362 1144 6363
rect 1165 6362 1172 6382
rect 1087 6355 1172 6362
rect 1191 6379 1229 6388
rect 1191 6359 1200 6379
rect 1220 6359 1229 6379
rect 1087 6354 1123 6355
rect 1191 6351 1229 6359
rect 1295 6383 1439 6389
rect 1295 6363 1303 6383
rect 1323 6363 1411 6383
rect 1431 6363 1439 6383
rect 1295 6355 1439 6363
rect 1295 6354 1331 6355
rect 1403 6354 1439 6355
rect 1505 6388 1542 6389
rect 1505 6387 1543 6388
rect 1505 6379 1569 6387
rect 1505 6359 1514 6379
rect 1534 6365 1569 6379
rect 1589 6365 1592 6385
rect 1534 6360 1592 6365
rect 1534 6359 1569 6360
rect 771 6322 808 6351
rect 772 6320 808 6322
rect 984 6320 1021 6351
rect 772 6298 1021 6320
rect 853 6292 964 6298
rect 853 6284 894 6292
rect 853 6264 861 6284
rect 880 6264 894 6284
rect 853 6262 894 6264
rect 922 6284 964 6292
rect 922 6264 938 6284
rect 957 6264 964 6284
rect 922 6262 964 6264
rect 853 6247 964 6262
rect 1192 6252 1229 6351
rect 1505 6347 1569 6359
rect 855 6244 959 6247
rect 643 6207 764 6217
rect 643 6205 712 6207
rect 643 6164 656 6205
rect 693 6166 712 6205
rect 749 6166 764 6207
rect 693 6164 764 6166
rect 643 6146 764 6164
rect 435 6102 500 6136
rect 855 6102 959 6104
rect 1190 6102 1231 6252
rect 1609 6244 1636 6499
rect 1698 6489 1778 6500
rect 1698 6463 1715 6489
rect 1755 6463 1778 6489
rect 1698 6436 1778 6463
rect 1698 6410 1719 6436
rect 1759 6410 1778 6436
rect 1698 6391 1778 6410
rect 1698 6365 1722 6391
rect 1762 6365 1778 6391
rect 1698 6314 1778 6365
rect 435 6099 1231 6102
rect 1610 6113 1636 6244
rect 1700 6114 1770 6314
rect 1610 6099 1638 6113
rect 435 6064 1638 6099
rect 1699 6092 1771 6114
rect 435 5907 500 6064
rect 855 6062 959 6064
rect 1190 6062 1231 6064
rect 1699 6044 1713 6092
rect 1759 6044 1771 6092
rect 1699 6027 1771 6044
rect 2801 5994 2873 7833
rect 2979 6066 3071 9370
rect 3465 9353 3496 9374
rect 3886 9353 3922 9374
rect 3308 9352 3345 9353
rect 3307 9343 3345 9352
rect 3307 9323 3316 9343
rect 3336 9323 3345 9343
rect 3307 9315 3345 9323
rect 3411 9347 3496 9353
rect 3521 9352 3558 9353
rect 3411 9327 3419 9347
rect 3439 9327 3496 9347
rect 3411 9319 3496 9327
rect 3520 9343 3558 9352
rect 3520 9323 3529 9343
rect 3549 9323 3558 9343
rect 3411 9318 3447 9319
rect 3520 9315 3558 9323
rect 3624 9347 3709 9353
rect 3729 9352 3766 9353
rect 3624 9327 3632 9347
rect 3652 9346 3709 9347
rect 3652 9327 3681 9346
rect 3624 9326 3681 9327
rect 3702 9326 3709 9346
rect 3624 9319 3709 9326
rect 3728 9343 3766 9352
rect 3728 9323 3737 9343
rect 3757 9323 3766 9343
rect 3624 9318 3660 9319
rect 3728 9315 3766 9323
rect 3832 9347 3976 9353
rect 3832 9327 3840 9347
rect 3860 9327 3948 9347
rect 3968 9327 3976 9347
rect 3832 9319 3976 9327
rect 3832 9318 3868 9319
rect 3940 9318 3976 9319
rect 4042 9352 4079 9353
rect 4042 9351 4080 9352
rect 4042 9343 4106 9351
rect 4042 9323 4051 9343
rect 4071 9329 4106 9343
rect 4126 9329 4129 9349
rect 4071 9324 4129 9329
rect 4071 9323 4106 9324
rect 3308 9286 3345 9315
rect 3309 9284 3345 9286
rect 3521 9284 3558 9315
rect 3309 9262 3558 9284
rect 3390 9256 3501 9262
rect 3390 9248 3431 9256
rect 3390 9228 3398 9248
rect 3417 9228 3431 9248
rect 3390 9226 3431 9228
rect 3459 9248 3501 9256
rect 3459 9228 3475 9248
rect 3494 9228 3501 9248
rect 3459 9226 3501 9228
rect 3390 9211 3501 9226
rect 3729 9194 3766 9315
rect 4042 9311 4106 9323
rect 3847 9194 3876 9198
rect 4146 9196 4173 9463
rect 4005 9194 4173 9196
rect 3729 9168 4173 9194
rect 3688 8900 3733 8909
rect 3688 8862 3698 8900
rect 3723 8862 3733 8900
rect 3688 8851 3733 8862
rect 3691 8843 3733 8851
rect 3691 8138 3734 8843
rect 3847 8229 3876 9168
rect 4005 9167 4173 9168
rect 3845 8208 3882 8229
rect 3845 8171 3856 8208
rect 3873 8171 3882 8208
rect 3845 8161 3882 8171
rect 3691 8118 4085 8138
rect 4105 8118 4108 8138
rect 3692 8113 4108 8118
rect 3692 8112 4033 8113
rect 3349 8081 3459 8095
rect 3349 8078 3392 8081
rect 3349 8073 3353 8078
rect 3271 8051 3353 8073
rect 3382 8051 3392 8078
rect 3420 8054 3427 8081
rect 3456 8073 3459 8081
rect 3456 8054 3521 8073
rect 3420 8051 3521 8054
rect 3271 8049 3521 8051
rect 3271 7970 3308 8049
rect 3349 8036 3459 8049
rect 3423 7980 3454 7981
rect 3271 7950 3280 7970
rect 3300 7950 3308 7970
rect 3271 7940 3308 7950
rect 3367 7970 3454 7980
rect 3367 7950 3376 7970
rect 3396 7950 3454 7970
rect 3367 7941 3454 7950
rect 3367 7940 3404 7941
rect 3423 7888 3454 7941
rect 3484 7970 3521 8049
rect 3636 7980 3667 7981
rect 3484 7950 3493 7970
rect 3513 7950 3521 7970
rect 3484 7940 3521 7950
rect 3580 7973 3667 7980
rect 3580 7970 3641 7973
rect 3580 7950 3589 7970
rect 3609 7953 3641 7970
rect 3662 7953 3667 7973
rect 3609 7950 3667 7953
rect 3580 7943 3667 7950
rect 3692 7970 3729 8112
rect 3995 8111 4032 8112
rect 3844 7980 3880 7981
rect 3692 7950 3701 7970
rect 3721 7950 3729 7970
rect 3580 7941 3636 7943
rect 3580 7940 3617 7941
rect 3692 7940 3729 7950
rect 3788 7970 3936 7980
rect 4036 7977 4132 7979
rect 3788 7950 3797 7970
rect 3817 7950 3907 7970
rect 3927 7950 3936 7970
rect 3788 7944 3936 7950
rect 3788 7941 3852 7944
rect 3788 7940 3825 7941
rect 3844 7914 3852 7941
rect 3873 7941 3936 7944
rect 3994 7970 4132 7977
rect 3994 7950 4003 7970
rect 4023 7950 4132 7970
rect 3994 7941 4132 7950
rect 3873 7914 3880 7941
rect 3899 7940 3936 7941
rect 3995 7940 4032 7941
rect 3844 7889 3880 7914
rect 3315 7887 3356 7888
rect 3235 7882 3356 7887
rect 3186 7880 3356 7882
rect 3186 7869 3325 7880
rect 3186 7846 3209 7869
rect 3235 7860 3325 7869
rect 3345 7860 3356 7880
rect 3235 7852 3356 7860
rect 3423 7884 3782 7888
rect 3423 7879 3745 7884
rect 3423 7855 3536 7879
rect 3560 7860 3745 7879
rect 3769 7860 3782 7884
rect 3560 7855 3782 7860
rect 3423 7852 3782 7855
rect 3844 7852 3879 7889
rect 3947 7886 4047 7889
rect 3947 7882 4014 7886
rect 3947 7856 3959 7882
rect 3985 7860 4014 7882
rect 4040 7860 4047 7886
rect 3985 7856 4047 7860
rect 3947 7852 4047 7856
rect 3235 7846 3243 7852
rect 3186 7838 3243 7846
rect 3423 7831 3454 7852
rect 3844 7831 3880 7852
rect 3266 7830 3303 7831
rect 3265 7821 3303 7830
rect 3265 7801 3274 7821
rect 3294 7801 3303 7821
rect 3265 7793 3303 7801
rect 3369 7825 3454 7831
rect 3479 7830 3516 7831
rect 3369 7805 3377 7825
rect 3397 7805 3454 7825
rect 3369 7797 3454 7805
rect 3478 7821 3516 7830
rect 3478 7801 3487 7821
rect 3507 7801 3516 7821
rect 3369 7796 3405 7797
rect 3478 7793 3516 7801
rect 3582 7825 3667 7831
rect 3687 7830 3724 7831
rect 3582 7805 3590 7825
rect 3610 7824 3667 7825
rect 3610 7805 3639 7824
rect 3582 7804 3639 7805
rect 3660 7804 3667 7824
rect 3582 7797 3667 7804
rect 3686 7821 3724 7830
rect 3686 7801 3695 7821
rect 3715 7801 3724 7821
rect 3582 7796 3618 7797
rect 3686 7793 3724 7801
rect 3790 7825 3934 7831
rect 3790 7805 3798 7825
rect 3818 7805 3906 7825
rect 3926 7805 3934 7825
rect 3790 7797 3934 7805
rect 3790 7796 3826 7797
rect 3898 7796 3934 7797
rect 4000 7830 4037 7831
rect 4000 7829 4038 7830
rect 4000 7821 4064 7829
rect 4000 7801 4009 7821
rect 4029 7807 4064 7821
rect 4084 7807 4087 7827
rect 4029 7802 4087 7807
rect 4029 7801 4064 7802
rect 3266 7764 3303 7793
rect 3267 7762 3303 7764
rect 3479 7762 3516 7793
rect 3267 7740 3516 7762
rect 3348 7734 3459 7740
rect 3348 7726 3389 7734
rect 3348 7706 3356 7726
rect 3375 7706 3389 7726
rect 3348 7704 3389 7706
rect 3417 7726 3459 7734
rect 3417 7706 3433 7726
rect 3452 7706 3459 7726
rect 3417 7704 3459 7706
rect 3348 7689 3459 7704
rect 3687 7678 3724 7793
rect 4000 7789 4064 7801
rect 3680 7672 3727 7678
rect 4104 7674 4131 7941
rect 3963 7672 4131 7674
rect 3680 7646 4131 7672
rect 3680 7511 3727 7646
rect 3963 7645 4131 7646
rect 3678 7462 3737 7511
rect 3678 7434 3696 7462
rect 3724 7434 3737 7462
rect 3678 7424 3737 7434
rect 4793 6687 4871 9727
rect 4793 6667 5193 6687
rect 5213 6667 5216 6687
rect 4793 6665 5216 6667
rect 4800 6662 5216 6665
rect 4800 6661 5141 6662
rect 4457 6630 4567 6644
rect 4457 6627 4500 6630
rect 4457 6622 4461 6627
rect 4379 6600 4461 6622
rect 4490 6600 4500 6627
rect 4528 6603 4535 6630
rect 4564 6622 4567 6630
rect 4564 6603 4629 6622
rect 4528 6600 4629 6603
rect 4379 6598 4629 6600
rect 4379 6519 4416 6598
rect 4457 6585 4567 6598
rect 4531 6529 4562 6530
rect 4379 6499 4388 6519
rect 4408 6499 4416 6519
rect 4379 6489 4416 6499
rect 4475 6519 4562 6529
rect 4475 6499 4484 6519
rect 4504 6499 4562 6519
rect 4475 6490 4562 6499
rect 4475 6489 4512 6490
rect 4249 6436 4360 6439
rect 4531 6437 4562 6490
rect 4592 6519 4629 6598
rect 4744 6529 4775 6530
rect 4592 6499 4601 6519
rect 4621 6499 4629 6519
rect 4592 6489 4629 6499
rect 4688 6522 4775 6529
rect 4688 6519 4749 6522
rect 4688 6499 4697 6519
rect 4717 6502 4749 6519
rect 4770 6502 4775 6522
rect 4717 6499 4775 6502
rect 4688 6492 4775 6499
rect 4800 6519 4837 6661
rect 5103 6660 5140 6661
rect 4952 6529 4988 6530
rect 4800 6499 4809 6519
rect 4829 6499 4837 6519
rect 4688 6490 4744 6492
rect 4688 6489 4725 6490
rect 4800 6489 4837 6499
rect 4896 6519 5044 6529
rect 5144 6526 5240 6528
rect 4896 6499 4905 6519
rect 4925 6499 5015 6519
rect 5035 6499 5044 6519
rect 4896 6493 5044 6499
rect 4896 6490 4960 6493
rect 4896 6489 4933 6490
rect 4952 6463 4960 6490
rect 4981 6490 5044 6493
rect 5102 6519 5240 6526
rect 5102 6499 5111 6519
rect 5131 6499 5240 6519
rect 5102 6490 5240 6499
rect 4981 6463 4988 6490
rect 5007 6489 5044 6490
rect 5103 6489 5140 6490
rect 4952 6438 4988 6463
rect 4423 6436 4464 6437
rect 4249 6429 4464 6436
rect 4249 6428 4314 6429
rect 4249 6404 4257 6428
rect 4281 6405 4314 6428
rect 4338 6409 4433 6429
rect 4453 6409 4464 6429
rect 4338 6405 4464 6409
rect 4281 6404 4464 6405
rect 4249 6401 4464 6404
rect 4531 6433 4890 6437
rect 4531 6428 4853 6433
rect 4531 6404 4644 6428
rect 4668 6409 4853 6428
rect 4877 6409 4890 6433
rect 4668 6404 4890 6409
rect 4531 6401 4890 6404
rect 4952 6401 4987 6438
rect 5055 6435 5155 6438
rect 5055 6431 5122 6435
rect 5055 6405 5067 6431
rect 5093 6409 5122 6431
rect 5148 6409 5155 6435
rect 5093 6405 5155 6409
rect 5055 6401 5155 6405
rect 4249 6397 4360 6401
rect 4531 6380 4562 6401
rect 4952 6380 4988 6401
rect 4374 6379 4411 6380
rect 4373 6370 4411 6379
rect 4373 6350 4382 6370
rect 4402 6350 4411 6370
rect 4373 6342 4411 6350
rect 4477 6374 4562 6380
rect 4587 6379 4624 6380
rect 4477 6354 4485 6374
rect 4505 6354 4562 6374
rect 4477 6346 4562 6354
rect 4586 6370 4624 6379
rect 4586 6350 4595 6370
rect 4615 6350 4624 6370
rect 4477 6345 4513 6346
rect 4586 6342 4624 6350
rect 4690 6374 4775 6380
rect 4795 6379 4832 6380
rect 4690 6354 4698 6374
rect 4718 6373 4775 6374
rect 4718 6354 4747 6373
rect 4690 6353 4747 6354
rect 4768 6353 4775 6373
rect 4690 6346 4775 6353
rect 4794 6370 4832 6379
rect 4794 6350 4803 6370
rect 4823 6350 4832 6370
rect 4690 6345 4726 6346
rect 4794 6342 4832 6350
rect 4898 6374 5042 6380
rect 4898 6354 4906 6374
rect 4926 6354 5014 6374
rect 5034 6354 5042 6374
rect 4898 6346 5042 6354
rect 4898 6345 4934 6346
rect 5006 6345 5042 6346
rect 5108 6379 5145 6380
rect 5108 6378 5146 6379
rect 5108 6370 5172 6378
rect 5108 6350 5117 6370
rect 5137 6356 5172 6370
rect 5192 6356 5195 6376
rect 5137 6351 5195 6356
rect 5137 6350 5172 6351
rect 4374 6313 4411 6342
rect 4375 6311 4411 6313
rect 4587 6311 4624 6342
rect 4375 6289 4624 6311
rect 4456 6283 4567 6289
rect 4456 6275 4497 6283
rect 4456 6255 4464 6275
rect 4483 6255 4497 6275
rect 4456 6253 4497 6255
rect 4525 6275 4567 6283
rect 4525 6255 4541 6275
rect 4560 6255 4567 6275
rect 4525 6253 4567 6255
rect 4456 6238 4567 6253
rect 4795 6227 4832 6342
rect 5108 6338 5172 6350
rect 4791 6221 4846 6227
rect 5212 6223 5239 6490
rect 5071 6221 5239 6223
rect 4791 6196 5239 6221
rect 4791 6162 4800 6196
rect 4829 6195 5239 6196
rect 4829 6162 4846 6195
rect 5071 6194 5239 6195
rect 4791 6136 4846 6162
rect 4791 6102 4799 6136
rect 4828 6102 4846 6136
rect 4791 6090 4846 6102
rect 2987 6045 3071 6066
rect 2987 6017 3015 6045
rect 3059 6017 3071 6045
rect 2801 5966 2875 5994
rect 2801 5918 2824 5966
rect 2861 5918 2875 5966
rect 2987 5988 3071 6017
rect 2987 5960 3012 5988
rect 3056 5960 3071 5988
rect 2987 5935 3071 5960
rect 2801 5909 2875 5918
rect 434 5859 500 5907
rect 2811 5905 2875 5909
rect 3024 5868 3735 5870
rect 2397 5867 3735 5868
rect 1347 5866 1419 5867
rect 434 5785 493 5859
rect 1346 5858 1445 5866
rect 1346 5855 1398 5858
rect 1346 5820 1354 5855
rect 1379 5820 1398 5855
rect 1423 5847 1445 5858
rect 2396 5859 3735 5867
rect 2396 5856 2448 5859
rect 1423 5846 2290 5847
rect 1423 5820 2291 5846
rect 1346 5810 2291 5820
rect 1346 5808 1445 5810
rect 434 5767 456 5785
rect 474 5767 493 5785
rect 434 5745 493 5767
rect 701 5781 1233 5786
rect 701 5761 1587 5781
rect 1607 5761 1610 5781
rect 2246 5777 2291 5810
rect 2396 5821 2404 5856
rect 2429 5821 2448 5856
rect 2473 5821 3735 5859
rect 2396 5812 3735 5821
rect 2396 5809 2485 5812
rect 3024 5810 3735 5812
rect 701 5757 1610 5761
rect 701 5710 744 5757
rect 1194 5756 1610 5757
rect 2242 5757 2635 5777
rect 2655 5757 2658 5777
rect 1194 5755 1535 5756
rect 851 5724 961 5738
rect 851 5721 894 5724
rect 851 5716 855 5721
rect 689 5709 744 5710
rect 433 5686 744 5709
rect 433 5668 458 5686
rect 476 5674 744 5686
rect 773 5694 855 5716
rect 884 5694 894 5721
rect 922 5697 929 5724
rect 958 5716 961 5724
rect 958 5697 1023 5716
rect 922 5694 1023 5697
rect 773 5692 1023 5694
rect 476 5668 498 5674
rect 433 5529 498 5668
rect 773 5613 810 5692
rect 851 5679 961 5692
rect 925 5623 956 5624
rect 773 5593 782 5613
rect 802 5593 810 5613
rect 433 5511 456 5529
rect 474 5511 498 5529
rect 433 5494 498 5511
rect 653 5575 721 5588
rect 773 5583 810 5593
rect 869 5613 956 5623
rect 869 5593 878 5613
rect 898 5593 956 5613
rect 869 5584 956 5593
rect 869 5583 906 5584
rect 653 5533 660 5575
rect 709 5533 721 5575
rect 653 5530 721 5533
rect 925 5531 956 5584
rect 986 5613 1023 5692
rect 1138 5623 1169 5624
rect 986 5593 995 5613
rect 1015 5593 1023 5613
rect 986 5583 1023 5593
rect 1082 5616 1169 5623
rect 1082 5613 1143 5616
rect 1082 5593 1091 5613
rect 1111 5596 1143 5613
rect 1164 5596 1169 5616
rect 1111 5593 1169 5596
rect 1082 5586 1169 5593
rect 1194 5613 1231 5755
rect 1497 5754 1534 5755
rect 2242 5752 2658 5757
rect 2242 5751 2583 5752
rect 1899 5720 2009 5734
rect 1899 5717 1942 5720
rect 1899 5712 1903 5717
rect 1821 5690 1903 5712
rect 1932 5690 1942 5717
rect 1970 5693 1977 5720
rect 2006 5712 2009 5720
rect 2006 5693 2071 5712
rect 1970 5690 2071 5693
rect 1821 5688 2071 5690
rect 1346 5623 1382 5624
rect 1194 5593 1203 5613
rect 1223 5593 1231 5613
rect 1082 5584 1138 5586
rect 1082 5583 1119 5584
rect 1194 5583 1231 5593
rect 1290 5613 1438 5623
rect 1538 5620 1634 5622
rect 1290 5593 1299 5613
rect 1319 5593 1409 5613
rect 1429 5593 1438 5613
rect 1290 5587 1438 5593
rect 1290 5584 1354 5587
rect 1290 5583 1327 5584
rect 1346 5557 1354 5584
rect 1375 5584 1438 5587
rect 1496 5613 1634 5620
rect 1496 5593 1505 5613
rect 1525 5593 1634 5613
rect 1496 5584 1634 5593
rect 1821 5609 1858 5688
rect 1899 5675 2009 5688
rect 1973 5619 2004 5620
rect 1821 5589 1830 5609
rect 1850 5589 1858 5609
rect 1375 5557 1382 5584
rect 1401 5583 1438 5584
rect 1497 5583 1534 5584
rect 1346 5532 1382 5557
rect 817 5530 858 5531
rect 653 5523 858 5530
rect 653 5512 827 5523
rect 653 5479 661 5512
rect 654 5470 661 5479
rect 710 5503 827 5512
rect 847 5503 858 5523
rect 710 5495 858 5503
rect 925 5527 1284 5531
rect 925 5522 1247 5527
rect 925 5498 1038 5522
rect 1062 5503 1247 5522
rect 1271 5503 1284 5527
rect 1062 5498 1284 5503
rect 925 5495 1284 5498
rect 1346 5495 1381 5532
rect 1449 5529 1549 5532
rect 1449 5525 1516 5529
rect 1449 5499 1461 5525
rect 1487 5503 1516 5525
rect 1542 5503 1549 5529
rect 1487 5499 1549 5503
rect 1449 5495 1549 5499
rect 710 5479 721 5495
rect 710 5470 718 5479
rect 925 5474 956 5495
rect 1346 5474 1382 5495
rect 768 5473 805 5474
rect 433 5430 498 5449
rect 433 5412 458 5430
rect 476 5412 498 5430
rect 433 5211 498 5412
rect 654 5286 718 5470
rect 767 5464 805 5473
rect 767 5444 776 5464
rect 796 5444 805 5464
rect 767 5436 805 5444
rect 871 5468 956 5474
rect 981 5473 1018 5474
rect 871 5448 879 5468
rect 899 5448 956 5468
rect 871 5440 956 5448
rect 980 5464 1018 5473
rect 980 5444 989 5464
rect 1009 5444 1018 5464
rect 871 5439 907 5440
rect 980 5436 1018 5444
rect 1084 5468 1169 5474
rect 1189 5473 1226 5474
rect 1084 5448 1092 5468
rect 1112 5467 1169 5468
rect 1112 5448 1141 5467
rect 1084 5447 1141 5448
rect 1162 5447 1169 5467
rect 1084 5440 1169 5447
rect 1188 5464 1226 5473
rect 1188 5444 1197 5464
rect 1217 5444 1226 5464
rect 1084 5439 1120 5440
rect 1188 5436 1226 5444
rect 1292 5468 1436 5474
rect 1292 5448 1300 5468
rect 1320 5448 1408 5468
rect 1428 5448 1436 5468
rect 1292 5440 1436 5448
rect 1292 5439 1328 5440
rect 1400 5439 1436 5440
rect 1502 5473 1539 5474
rect 1502 5472 1540 5473
rect 1502 5464 1566 5472
rect 1502 5444 1511 5464
rect 1531 5450 1566 5464
rect 1586 5450 1589 5470
rect 1531 5445 1589 5450
rect 1531 5444 1566 5445
rect 768 5407 805 5436
rect 769 5405 805 5407
rect 981 5405 1018 5436
rect 769 5383 1018 5405
rect 850 5377 961 5383
rect 850 5369 891 5377
rect 850 5349 858 5369
rect 877 5349 891 5369
rect 850 5347 891 5349
rect 919 5369 961 5377
rect 919 5349 935 5369
rect 954 5349 961 5369
rect 919 5347 961 5349
rect 850 5332 961 5347
rect 654 5276 722 5286
rect 654 5243 671 5276
rect 711 5243 722 5276
rect 654 5231 722 5243
rect 654 5229 718 5231
rect 1189 5212 1226 5436
rect 1502 5432 1566 5444
rect 1606 5214 1633 5584
rect 1821 5579 1858 5589
rect 1917 5609 2004 5619
rect 1917 5589 1926 5609
rect 1946 5589 2004 5609
rect 1917 5580 2004 5589
rect 1917 5579 1954 5580
rect 1697 5566 1767 5571
rect 1692 5560 1767 5566
rect 1692 5527 1700 5560
rect 1753 5527 1767 5560
rect 1973 5527 2004 5580
rect 2034 5609 2071 5688
rect 2186 5619 2217 5620
rect 2034 5589 2043 5609
rect 2063 5589 2071 5609
rect 2034 5579 2071 5589
rect 2130 5612 2217 5619
rect 2130 5609 2191 5612
rect 2130 5589 2139 5609
rect 2159 5592 2191 5609
rect 2212 5592 2217 5612
rect 2159 5589 2217 5592
rect 2130 5582 2217 5589
rect 2242 5609 2279 5751
rect 2545 5750 2582 5751
rect 2394 5619 2430 5620
rect 2242 5589 2251 5609
rect 2271 5589 2279 5609
rect 2130 5580 2186 5582
rect 2130 5579 2167 5580
rect 2242 5579 2279 5589
rect 2338 5609 2486 5619
rect 2586 5616 2682 5618
rect 2338 5589 2347 5609
rect 2367 5589 2457 5609
rect 2477 5589 2486 5609
rect 2338 5583 2486 5589
rect 2338 5580 2402 5583
rect 2338 5579 2375 5580
rect 2394 5553 2402 5580
rect 2423 5580 2486 5583
rect 2544 5609 2682 5616
rect 2544 5589 2553 5609
rect 2573 5589 2682 5609
rect 2544 5580 2682 5589
rect 2423 5553 2430 5580
rect 2449 5579 2486 5580
rect 2545 5579 2582 5580
rect 2394 5528 2430 5553
rect 1692 5526 1775 5527
rect 1865 5526 1906 5527
rect 1692 5519 1906 5526
rect 1692 5502 1875 5519
rect 1692 5469 1705 5502
rect 1758 5499 1875 5502
rect 1895 5499 1906 5519
rect 1758 5491 1906 5499
rect 1973 5523 2332 5527
rect 1973 5518 2295 5523
rect 1973 5494 2086 5518
rect 2110 5499 2295 5518
rect 2319 5499 2332 5523
rect 2110 5494 2332 5499
rect 1973 5491 2332 5494
rect 2394 5491 2429 5528
rect 2497 5525 2597 5528
rect 2497 5521 2564 5525
rect 2497 5495 2509 5521
rect 2535 5499 2564 5521
rect 2590 5499 2597 5525
rect 2535 5495 2597 5499
rect 2497 5491 2597 5495
rect 1758 5469 1775 5491
rect 1973 5470 2004 5491
rect 2394 5470 2430 5491
rect 1816 5469 1853 5470
rect 1692 5455 1775 5469
rect 1465 5212 1633 5214
rect 1189 5211 1633 5212
rect 433 5181 1633 5211
rect 1703 5245 1775 5455
rect 1815 5460 1853 5469
rect 1815 5440 1824 5460
rect 1844 5440 1853 5460
rect 1815 5432 1853 5440
rect 1919 5464 2004 5470
rect 2029 5469 2066 5470
rect 1919 5444 1927 5464
rect 1947 5444 2004 5464
rect 1919 5436 2004 5444
rect 2028 5460 2066 5469
rect 2028 5440 2037 5460
rect 2057 5440 2066 5460
rect 1919 5435 1955 5436
rect 2028 5432 2066 5440
rect 2132 5464 2217 5470
rect 2237 5469 2274 5470
rect 2132 5444 2140 5464
rect 2160 5463 2217 5464
rect 2160 5444 2189 5463
rect 2132 5443 2189 5444
rect 2210 5443 2217 5463
rect 2132 5436 2217 5443
rect 2236 5460 2274 5469
rect 2236 5440 2245 5460
rect 2265 5440 2274 5460
rect 2132 5435 2168 5436
rect 2236 5432 2274 5440
rect 2340 5464 2484 5470
rect 2340 5444 2348 5464
rect 2368 5444 2456 5464
rect 2476 5444 2484 5464
rect 2340 5436 2484 5444
rect 2340 5435 2376 5436
rect 2448 5435 2484 5436
rect 2550 5469 2587 5470
rect 2550 5468 2588 5469
rect 2550 5460 2614 5468
rect 2550 5440 2559 5460
rect 2579 5446 2614 5460
rect 2634 5446 2637 5466
rect 2579 5441 2637 5446
rect 2579 5440 2614 5441
rect 1816 5403 1853 5432
rect 1817 5401 1853 5403
rect 2029 5401 2066 5432
rect 1817 5379 2066 5401
rect 1898 5373 2009 5379
rect 1898 5365 1939 5373
rect 1898 5345 1906 5365
rect 1925 5345 1939 5365
rect 1898 5343 1939 5345
rect 1967 5365 2009 5373
rect 1967 5345 1983 5365
rect 2002 5345 2009 5365
rect 1967 5343 2009 5345
rect 1898 5328 2009 5343
rect 1703 5206 1722 5245
rect 1767 5206 1775 5245
rect 1703 5189 1775 5206
rect 2237 5233 2274 5432
rect 2550 5428 2614 5440
rect 2237 5227 2278 5233
rect 2654 5229 2681 5580
rect 2976 5567 3071 5593
rect 2812 5545 2876 5564
rect 2812 5506 2825 5545
rect 2859 5506 2876 5545
rect 2812 5487 2876 5506
rect 2513 5227 2681 5229
rect 2237 5201 2681 5227
rect 433 5134 498 5181
rect 433 5116 456 5134
rect 474 5116 498 5134
rect 1346 5161 1381 5163
rect 1346 5159 1450 5161
rect 2239 5159 2278 5201
rect 2513 5200 2681 5201
rect 1346 5152 2280 5159
rect 1346 5151 1397 5152
rect 1346 5131 1349 5151
rect 1374 5132 1397 5151
rect 1429 5132 2280 5152
rect 1374 5131 2280 5132
rect 1346 5124 2280 5131
rect 1619 5123 2280 5124
rect 433 5095 498 5116
rect 710 5106 750 5109
rect 710 5102 1613 5106
rect 710 5082 1587 5102
rect 1607 5082 1613 5102
rect 710 5079 1613 5082
rect 434 5035 499 5055
rect 434 5017 458 5035
rect 476 5017 499 5035
rect 434 4990 499 5017
rect 710 4990 750 5079
rect 1194 5077 1610 5079
rect 1194 5076 1535 5077
rect 851 5045 961 5059
rect 851 5042 894 5045
rect 851 5037 855 5042
rect 433 4955 750 4990
rect 773 5015 855 5037
rect 884 5015 894 5042
rect 922 5018 929 5045
rect 958 5037 961 5045
rect 958 5018 1023 5037
rect 922 5015 1023 5018
rect 773 5013 1023 5015
rect 434 4879 499 4955
rect 773 4934 810 5013
rect 851 5000 961 5013
rect 925 4944 956 4945
rect 773 4914 782 4934
rect 802 4914 810 4934
rect 773 4904 810 4914
rect 869 4934 956 4944
rect 869 4914 878 4934
rect 898 4914 956 4934
rect 869 4905 956 4914
rect 869 4904 906 4905
rect 434 4861 456 4879
rect 474 4861 499 4879
rect 434 4840 499 4861
rect 647 4859 712 4868
rect 647 4822 657 4859
rect 697 4851 712 4859
rect 925 4852 956 4905
rect 986 4934 1023 5013
rect 1138 4944 1169 4945
rect 986 4914 995 4934
rect 1015 4914 1023 4934
rect 986 4904 1023 4914
rect 1082 4937 1169 4944
rect 1082 4934 1143 4937
rect 1082 4914 1091 4934
rect 1111 4917 1143 4934
rect 1164 4917 1169 4937
rect 1111 4914 1169 4917
rect 1082 4907 1169 4914
rect 1194 4934 1231 5076
rect 1497 5075 1534 5076
rect 2814 5016 2876 5487
rect 2976 5526 3002 5567
rect 3038 5526 3071 5567
rect 2976 5230 3071 5526
rect 2976 5186 2991 5230
rect 3051 5186 3071 5230
rect 2976 5166 3071 5186
rect 3688 5097 3731 5810
rect 3688 5077 4082 5097
rect 4102 5077 4105 5097
rect 3689 5072 4105 5077
rect 3689 5071 4030 5072
rect 3346 5040 3456 5054
rect 3346 5037 3389 5040
rect 3346 5032 3350 5037
rect 2809 4964 2884 5016
rect 3268 5010 3350 5032
rect 3379 5010 3389 5037
rect 3417 5013 3424 5040
rect 3453 5032 3456 5040
rect 3453 5013 3518 5032
rect 3417 5010 3518 5013
rect 3268 5008 3518 5010
rect 3178 4964 3224 4965
rect 1346 4944 1382 4945
rect 1194 4914 1203 4934
rect 1223 4914 1231 4934
rect 1082 4905 1138 4907
rect 1082 4904 1119 4905
rect 1194 4904 1231 4914
rect 1290 4934 1438 4944
rect 1538 4941 1634 4943
rect 1290 4914 1299 4934
rect 1319 4914 1409 4934
rect 1429 4914 1438 4934
rect 1290 4908 1438 4914
rect 1290 4905 1354 4908
rect 1290 4904 1327 4905
rect 1346 4878 1354 4905
rect 1375 4905 1438 4908
rect 1496 4934 1634 4941
rect 1496 4914 1505 4934
rect 1525 4914 1634 4934
rect 1496 4905 1634 4914
rect 2809 4929 3224 4964
rect 1375 4878 1382 4905
rect 1401 4904 1438 4905
rect 1497 4904 1534 4905
rect 1346 4853 1382 4878
rect 817 4851 858 4852
rect 697 4844 858 4851
rect 697 4824 827 4844
rect 847 4824 858 4844
rect 697 4822 858 4824
rect 647 4816 858 4822
rect 925 4848 1284 4852
rect 925 4843 1247 4848
rect 925 4819 1038 4843
rect 1062 4824 1247 4843
rect 1271 4824 1284 4848
rect 1062 4819 1284 4824
rect 925 4816 1284 4819
rect 1346 4816 1381 4853
rect 1449 4850 1549 4853
rect 1449 4846 1516 4850
rect 1449 4820 1461 4846
rect 1487 4824 1516 4846
rect 1542 4824 1549 4850
rect 1487 4820 1549 4824
rect 1449 4816 1549 4820
rect 647 4803 714 4816
rect 439 4780 495 4800
rect 439 4762 458 4780
rect 476 4762 495 4780
rect 439 4649 495 4762
rect 647 4782 661 4803
rect 697 4782 714 4803
rect 925 4795 956 4816
rect 1346 4795 1382 4816
rect 768 4794 805 4795
rect 647 4775 714 4782
rect 767 4785 805 4794
rect 439 4511 494 4649
rect 647 4623 712 4775
rect 767 4765 776 4785
rect 796 4765 805 4785
rect 767 4757 805 4765
rect 871 4789 956 4795
rect 981 4794 1018 4795
rect 871 4769 879 4789
rect 899 4769 956 4789
rect 871 4761 956 4769
rect 980 4785 1018 4794
rect 980 4765 989 4785
rect 1009 4765 1018 4785
rect 871 4760 907 4761
rect 980 4757 1018 4765
rect 1084 4789 1169 4795
rect 1189 4794 1226 4795
rect 1084 4769 1092 4789
rect 1112 4788 1169 4789
rect 1112 4769 1141 4788
rect 1084 4768 1141 4769
rect 1162 4768 1169 4788
rect 1084 4761 1169 4768
rect 1188 4785 1226 4794
rect 1188 4765 1197 4785
rect 1217 4765 1226 4785
rect 1084 4760 1120 4761
rect 1188 4757 1226 4765
rect 1292 4789 1436 4795
rect 1292 4769 1300 4789
rect 1320 4769 1408 4789
rect 1428 4769 1436 4789
rect 1292 4761 1436 4769
rect 1292 4760 1328 4761
rect 1400 4760 1436 4761
rect 1502 4794 1539 4795
rect 1502 4793 1540 4794
rect 1502 4785 1566 4793
rect 1502 4765 1511 4785
rect 1531 4771 1566 4785
rect 1586 4771 1589 4791
rect 1531 4766 1589 4771
rect 1531 4765 1566 4766
rect 768 4728 805 4757
rect 769 4726 805 4728
rect 981 4726 1018 4757
rect 769 4704 1018 4726
rect 850 4698 961 4704
rect 850 4690 891 4698
rect 850 4670 858 4690
rect 877 4670 891 4690
rect 850 4668 891 4670
rect 919 4690 961 4698
rect 919 4670 935 4690
rect 954 4670 961 4690
rect 919 4668 961 4670
rect 850 4655 961 4668
rect 1189 4658 1226 4757
rect 1502 4753 1566 4765
rect 640 4613 761 4623
rect 640 4611 709 4613
rect 640 4570 653 4611
rect 690 4572 709 4611
rect 746 4572 761 4613
rect 690 4570 761 4572
rect 640 4552 761 4570
rect 432 4508 496 4511
rect 852 4508 956 4514
rect 1187 4508 1228 4658
rect 1606 4650 1633 4905
rect 1695 4895 1775 4906
rect 1695 4869 1712 4895
rect 1752 4869 1775 4895
rect 1695 4842 1775 4869
rect 1695 4816 1716 4842
rect 1756 4816 1775 4842
rect 1695 4797 1775 4816
rect 1695 4771 1719 4797
rect 1759 4771 1775 4797
rect 1695 4720 1775 4771
rect 432 4505 1228 4508
rect 1607 4519 1633 4650
rect 1607 4505 1635 4519
rect 432 4470 1635 4505
rect 1697 4512 1767 4720
rect 2809 4645 2884 4929
rect 3178 4846 3224 4929
rect 3268 4929 3305 5008
rect 3346 4995 3456 5008
rect 3420 4939 3451 4940
rect 3268 4909 3277 4929
rect 3297 4909 3305 4929
rect 3268 4899 3305 4909
rect 3364 4929 3451 4939
rect 3364 4909 3373 4929
rect 3393 4909 3451 4929
rect 3364 4900 3451 4909
rect 3364 4899 3401 4900
rect 3420 4847 3451 4900
rect 3481 4929 3518 5008
rect 3633 4939 3664 4940
rect 3481 4909 3490 4929
rect 3510 4909 3518 4929
rect 3481 4899 3518 4909
rect 3577 4932 3664 4939
rect 3577 4929 3638 4932
rect 3577 4909 3586 4929
rect 3606 4912 3638 4929
rect 3659 4912 3664 4932
rect 3606 4909 3664 4912
rect 3577 4902 3664 4909
rect 3689 4929 3726 5071
rect 3992 5070 4029 5071
rect 3841 4939 3877 4940
rect 3689 4909 3698 4929
rect 3718 4909 3726 4929
rect 3577 4900 3633 4902
rect 3577 4899 3614 4900
rect 3689 4899 3726 4909
rect 3785 4929 3933 4939
rect 4033 4936 4129 4938
rect 3785 4909 3794 4929
rect 3814 4909 3904 4929
rect 3924 4909 3933 4929
rect 3785 4903 3933 4909
rect 3785 4900 3849 4903
rect 3785 4899 3822 4900
rect 3841 4873 3849 4900
rect 3870 4900 3933 4903
rect 3991 4929 4129 4936
rect 3991 4909 4000 4929
rect 4020 4909 4129 4929
rect 3991 4900 4129 4909
rect 3870 4873 3877 4900
rect 3896 4899 3933 4900
rect 3992 4899 4029 4900
rect 3841 4848 3877 4873
rect 3312 4846 3353 4847
rect 3178 4839 3353 4846
rect 2976 4813 3062 4832
rect 2976 4772 2991 4813
rect 3045 4772 3062 4813
rect 3178 4819 3322 4839
rect 3342 4819 3353 4839
rect 3178 4811 3353 4819
rect 3420 4843 3779 4847
rect 3420 4838 3742 4843
rect 3420 4814 3533 4838
rect 3557 4819 3742 4838
rect 3766 4819 3779 4843
rect 3557 4814 3779 4819
rect 3420 4811 3779 4814
rect 3841 4811 3876 4848
rect 3944 4845 4044 4848
rect 3944 4841 4011 4845
rect 3944 4815 3956 4841
rect 3982 4819 4011 4841
rect 4037 4819 4044 4845
rect 3982 4815 4044 4819
rect 3944 4811 4044 4815
rect 3178 4807 3224 4811
rect 3420 4790 3451 4811
rect 3841 4790 3877 4811
rect 3263 4789 3300 4790
rect 2976 4736 3062 4772
rect 3262 4780 3300 4789
rect 3262 4760 3271 4780
rect 3291 4760 3300 4780
rect 3262 4752 3300 4760
rect 3366 4784 3451 4790
rect 3476 4789 3513 4790
rect 3366 4764 3374 4784
rect 3394 4764 3451 4784
rect 3366 4756 3451 4764
rect 3475 4780 3513 4789
rect 3475 4760 3484 4780
rect 3504 4760 3513 4780
rect 3366 4755 3402 4756
rect 3475 4752 3513 4760
rect 3579 4784 3664 4790
rect 3684 4789 3721 4790
rect 3579 4764 3587 4784
rect 3607 4783 3664 4784
rect 3607 4764 3636 4783
rect 3579 4763 3636 4764
rect 3657 4763 3664 4783
rect 3579 4756 3664 4763
rect 3683 4780 3721 4789
rect 3683 4760 3692 4780
rect 3712 4760 3721 4780
rect 3579 4755 3615 4756
rect 3683 4752 3721 4760
rect 3787 4784 3931 4790
rect 3787 4764 3795 4784
rect 3815 4764 3903 4784
rect 3923 4764 3931 4784
rect 3787 4756 3931 4764
rect 3787 4755 3823 4756
rect 432 4409 496 4470
rect 852 4468 956 4470
rect 1187 4468 1228 4470
rect 1697 4467 1718 4512
rect 1698 4446 1718 4467
rect 1748 4467 1767 4512
rect 2804 4603 2884 4645
rect 1748 4446 1765 4467
rect 1698 4427 1765 4446
rect 1347 4419 1419 4420
rect 1346 4411 1445 4419
rect 434 4338 493 4409
rect 1346 4408 1398 4411
rect 1346 4373 1354 4408
rect 1379 4373 1398 4408
rect 1423 4400 1445 4411
rect 1423 4399 2290 4400
rect 1423 4373 2291 4399
rect 1346 4363 2291 4373
rect 1346 4361 1445 4363
rect 434 4320 456 4338
rect 474 4320 493 4338
rect 434 4298 493 4320
rect 701 4334 1233 4339
rect 701 4314 1587 4334
rect 1607 4314 1610 4334
rect 2246 4330 2291 4363
rect 701 4310 1610 4314
rect 701 4263 744 4310
rect 1194 4309 1610 4310
rect 2242 4310 2635 4330
rect 2655 4310 2658 4330
rect 1194 4308 1535 4309
rect 851 4277 961 4291
rect 851 4274 894 4277
rect 851 4269 855 4274
rect 689 4262 744 4263
rect 433 4239 744 4262
rect 433 4221 458 4239
rect 476 4227 744 4239
rect 773 4247 855 4269
rect 884 4247 894 4274
rect 922 4250 929 4277
rect 958 4269 961 4277
rect 958 4250 1023 4269
rect 922 4247 1023 4250
rect 773 4245 1023 4247
rect 476 4221 498 4227
rect 433 4082 498 4221
rect 773 4166 810 4245
rect 851 4232 961 4245
rect 925 4176 956 4177
rect 773 4146 782 4166
rect 802 4146 810 4166
rect 433 4064 456 4082
rect 474 4064 498 4082
rect 433 4047 498 4064
rect 653 4128 721 4141
rect 773 4136 810 4146
rect 869 4166 956 4176
rect 869 4146 878 4166
rect 898 4146 956 4166
rect 869 4137 956 4146
rect 869 4136 906 4137
rect 653 4086 660 4128
rect 709 4086 721 4128
rect 653 4083 721 4086
rect 925 4084 956 4137
rect 986 4166 1023 4245
rect 1138 4176 1169 4177
rect 986 4146 995 4166
rect 1015 4146 1023 4166
rect 986 4136 1023 4146
rect 1082 4169 1169 4176
rect 1082 4166 1143 4169
rect 1082 4146 1091 4166
rect 1111 4149 1143 4166
rect 1164 4149 1169 4169
rect 1111 4146 1169 4149
rect 1082 4139 1169 4146
rect 1194 4166 1231 4308
rect 1497 4307 1534 4308
rect 2242 4305 2658 4310
rect 2242 4304 2583 4305
rect 1899 4273 2009 4287
rect 1899 4270 1942 4273
rect 1899 4265 1903 4270
rect 1821 4243 1903 4265
rect 1932 4243 1942 4270
rect 1970 4246 1977 4273
rect 2006 4265 2009 4273
rect 2006 4246 2071 4265
rect 1970 4243 2071 4246
rect 1821 4241 2071 4243
rect 1346 4176 1382 4177
rect 1194 4146 1203 4166
rect 1223 4146 1231 4166
rect 1082 4137 1138 4139
rect 1082 4136 1119 4137
rect 1194 4136 1231 4146
rect 1290 4166 1438 4176
rect 1538 4173 1634 4175
rect 1290 4146 1299 4166
rect 1319 4146 1409 4166
rect 1429 4146 1438 4166
rect 1290 4140 1438 4146
rect 1290 4137 1354 4140
rect 1290 4136 1327 4137
rect 1346 4110 1354 4137
rect 1375 4137 1438 4140
rect 1496 4166 1634 4173
rect 1496 4146 1505 4166
rect 1525 4146 1634 4166
rect 1496 4137 1634 4146
rect 1821 4162 1858 4241
rect 1899 4228 2009 4241
rect 1973 4172 2004 4173
rect 1821 4142 1830 4162
rect 1850 4142 1858 4162
rect 1375 4110 1382 4137
rect 1401 4136 1438 4137
rect 1497 4136 1534 4137
rect 1346 4085 1382 4110
rect 817 4083 858 4084
rect 653 4076 858 4083
rect 653 4065 827 4076
rect 653 4032 661 4065
rect 654 4023 661 4032
rect 710 4056 827 4065
rect 847 4056 858 4076
rect 710 4048 858 4056
rect 925 4080 1284 4084
rect 925 4075 1247 4080
rect 925 4051 1038 4075
rect 1062 4056 1247 4075
rect 1271 4056 1284 4080
rect 1062 4051 1284 4056
rect 925 4048 1284 4051
rect 1346 4048 1381 4085
rect 1449 4082 1549 4085
rect 1449 4078 1516 4082
rect 1449 4052 1461 4078
rect 1487 4056 1516 4078
rect 1542 4056 1549 4082
rect 1487 4052 1549 4056
rect 1449 4048 1549 4052
rect 710 4032 721 4048
rect 710 4023 718 4032
rect 925 4027 956 4048
rect 1346 4027 1382 4048
rect 768 4026 805 4027
rect 433 3983 498 4002
rect 433 3965 458 3983
rect 476 3965 498 3983
rect 433 3764 498 3965
rect 654 3839 718 4023
rect 767 4017 805 4026
rect 767 3997 776 4017
rect 796 3997 805 4017
rect 767 3989 805 3997
rect 871 4021 956 4027
rect 981 4026 1018 4027
rect 871 4001 879 4021
rect 899 4001 956 4021
rect 871 3993 956 4001
rect 980 4017 1018 4026
rect 980 3997 989 4017
rect 1009 3997 1018 4017
rect 871 3992 907 3993
rect 980 3989 1018 3997
rect 1084 4021 1169 4027
rect 1189 4026 1226 4027
rect 1084 4001 1092 4021
rect 1112 4020 1169 4021
rect 1112 4001 1141 4020
rect 1084 4000 1141 4001
rect 1162 4000 1169 4020
rect 1084 3993 1169 4000
rect 1188 4017 1226 4026
rect 1188 3997 1197 4017
rect 1217 3997 1226 4017
rect 1084 3992 1120 3993
rect 1188 3989 1226 3997
rect 1292 4021 1436 4027
rect 1292 4001 1300 4021
rect 1320 4001 1408 4021
rect 1428 4001 1436 4021
rect 1292 3993 1436 4001
rect 1292 3992 1328 3993
rect 1400 3992 1436 3993
rect 1502 4026 1539 4027
rect 1502 4025 1540 4026
rect 1502 4017 1566 4025
rect 1502 3997 1511 4017
rect 1531 4003 1566 4017
rect 1586 4003 1589 4023
rect 1531 3998 1589 4003
rect 1531 3997 1566 3998
rect 768 3960 805 3989
rect 769 3958 805 3960
rect 981 3958 1018 3989
rect 769 3936 1018 3958
rect 850 3930 961 3936
rect 850 3922 891 3930
rect 850 3902 858 3922
rect 877 3902 891 3922
rect 850 3900 891 3902
rect 919 3922 961 3930
rect 919 3902 935 3922
rect 954 3902 961 3922
rect 919 3900 961 3902
rect 850 3885 961 3900
rect 654 3829 722 3839
rect 654 3796 671 3829
rect 711 3796 722 3829
rect 654 3784 722 3796
rect 654 3782 718 3784
rect 1189 3765 1226 3989
rect 1502 3985 1566 3997
rect 1606 3767 1633 4137
rect 1821 4132 1858 4142
rect 1917 4162 2004 4172
rect 1917 4142 1926 4162
rect 1946 4142 2004 4162
rect 1917 4133 2004 4142
rect 1917 4132 1954 4133
rect 1697 4119 1767 4124
rect 1692 4113 1767 4119
rect 1692 4080 1700 4113
rect 1753 4080 1767 4113
rect 1973 4080 2004 4133
rect 2034 4162 2071 4241
rect 2186 4172 2217 4173
rect 2034 4142 2043 4162
rect 2063 4142 2071 4162
rect 2034 4132 2071 4142
rect 2130 4165 2217 4172
rect 2130 4162 2191 4165
rect 2130 4142 2139 4162
rect 2159 4145 2191 4162
rect 2212 4145 2217 4165
rect 2159 4142 2217 4145
rect 2130 4135 2217 4142
rect 2242 4162 2279 4304
rect 2545 4303 2582 4304
rect 2394 4172 2430 4173
rect 2242 4142 2251 4162
rect 2271 4142 2279 4162
rect 2130 4133 2186 4135
rect 2130 4132 2167 4133
rect 2242 4132 2279 4142
rect 2338 4162 2486 4172
rect 2586 4169 2682 4171
rect 2338 4142 2347 4162
rect 2367 4142 2457 4162
rect 2477 4142 2486 4162
rect 2338 4136 2486 4142
rect 2338 4133 2402 4136
rect 2338 4132 2375 4133
rect 2394 4106 2402 4133
rect 2423 4133 2486 4136
rect 2544 4162 2682 4169
rect 2544 4142 2553 4162
rect 2573 4142 2682 4162
rect 2544 4133 2682 4142
rect 2423 4106 2430 4133
rect 2449 4132 2486 4133
rect 2545 4132 2582 4133
rect 2394 4081 2430 4106
rect 1692 4079 1775 4080
rect 1865 4079 1906 4080
rect 1692 4072 1906 4079
rect 1692 4055 1875 4072
rect 1692 4022 1705 4055
rect 1758 4052 1875 4055
rect 1895 4052 1906 4072
rect 1758 4044 1906 4052
rect 1973 4076 2332 4080
rect 1973 4071 2295 4076
rect 1973 4047 2086 4071
rect 2110 4052 2295 4071
rect 2319 4052 2332 4076
rect 2110 4047 2332 4052
rect 1973 4044 2332 4047
rect 2394 4044 2429 4081
rect 2497 4078 2597 4081
rect 2497 4074 2564 4078
rect 2497 4048 2509 4074
rect 2535 4052 2564 4074
rect 2590 4052 2597 4078
rect 2535 4048 2597 4052
rect 2497 4044 2597 4048
rect 1758 4022 1775 4044
rect 1973 4023 2004 4044
rect 2394 4023 2430 4044
rect 1816 4022 1853 4023
rect 1692 4008 1775 4022
rect 1465 3765 1633 3767
rect 1189 3764 1633 3765
rect 433 3734 1633 3764
rect 1703 3798 1775 4008
rect 1815 4013 1853 4022
rect 1815 3993 1824 4013
rect 1844 3993 1853 4013
rect 1815 3985 1853 3993
rect 1919 4017 2004 4023
rect 2029 4022 2066 4023
rect 1919 3997 1927 4017
rect 1947 3997 2004 4017
rect 1919 3989 2004 3997
rect 2028 4013 2066 4022
rect 2028 3993 2037 4013
rect 2057 3993 2066 4013
rect 1919 3988 1955 3989
rect 2028 3985 2066 3993
rect 2132 4017 2217 4023
rect 2237 4022 2274 4023
rect 2132 3997 2140 4017
rect 2160 4016 2217 4017
rect 2160 3997 2189 4016
rect 2132 3996 2189 3997
rect 2210 3996 2217 4016
rect 2132 3989 2217 3996
rect 2236 4013 2274 4022
rect 2236 3993 2245 4013
rect 2265 3993 2274 4013
rect 2132 3988 2168 3989
rect 2236 3985 2274 3993
rect 2340 4017 2484 4023
rect 2340 3997 2348 4017
rect 2368 3997 2456 4017
rect 2476 3997 2484 4017
rect 2340 3989 2484 3997
rect 2340 3988 2376 3989
rect 2448 3988 2484 3989
rect 2550 4022 2587 4023
rect 2550 4021 2588 4022
rect 2550 4013 2614 4021
rect 2550 3993 2559 4013
rect 2579 3999 2614 4013
rect 2634 3999 2637 4019
rect 2579 3994 2637 3999
rect 2579 3993 2614 3994
rect 1816 3956 1853 3985
rect 1817 3954 1853 3956
rect 2029 3954 2066 3985
rect 1817 3932 2066 3954
rect 1898 3926 2009 3932
rect 1898 3918 1939 3926
rect 1898 3898 1906 3918
rect 1925 3898 1939 3918
rect 1898 3896 1939 3898
rect 1967 3918 2009 3926
rect 1967 3898 1983 3918
rect 2002 3898 2009 3918
rect 1967 3896 2009 3898
rect 1898 3881 2009 3896
rect 1703 3759 1722 3798
rect 1767 3759 1775 3798
rect 1703 3742 1775 3759
rect 2237 3786 2274 3985
rect 2550 3981 2614 3993
rect 2237 3780 2278 3786
rect 2654 3782 2681 4133
rect 2804 4003 2883 4603
rect 2980 4151 3059 4736
rect 3263 4723 3300 4752
rect 3264 4721 3300 4723
rect 3476 4721 3513 4752
rect 3264 4699 3513 4721
rect 3345 4693 3456 4699
rect 3345 4685 3386 4693
rect 3345 4665 3353 4685
rect 3372 4665 3386 4685
rect 3345 4663 3386 4665
rect 3414 4685 3456 4693
rect 3414 4665 3430 4685
rect 3449 4665 3456 4685
rect 3414 4663 3456 4665
rect 3345 4648 3456 4663
rect 3684 4637 3721 4752
rect 3677 4525 3724 4637
rect 3845 4597 3875 4756
rect 3895 4755 3931 4756
rect 3997 4789 4034 4790
rect 3997 4788 4035 4789
rect 3997 4780 4061 4788
rect 3997 4760 4006 4780
rect 4026 4766 4061 4780
rect 4081 4766 4084 4786
rect 4026 4761 4084 4766
rect 4026 4760 4061 4761
rect 3997 4748 4061 4760
rect 3845 4593 3931 4597
rect 3845 4575 3860 4593
rect 3912 4575 3931 4593
rect 3845 4566 3931 4575
rect 4101 4527 4128 4900
rect 3960 4525 4128 4527
rect 3677 4499 4128 4525
rect 3677 4421 3724 4499
rect 3960 4498 4128 4499
rect 3622 4420 3724 4421
rect 3621 4412 3724 4420
rect 3621 4409 3673 4412
rect 3621 4374 3629 4409
rect 3654 4374 3673 4409
rect 3698 4374 3724 4412
rect 3621 4368 3724 4374
rect 3884 4413 3920 4417
rect 3884 4390 3892 4413
rect 3916 4390 3920 4413
rect 3884 4369 3920 4390
rect 3621 4364 3720 4368
rect 3884 4346 3892 4369
rect 3916 4346 3920 4369
rect 2513 3780 2681 3782
rect 2237 3754 2681 3780
rect 433 3687 498 3734
rect 433 3669 456 3687
rect 474 3669 498 3687
rect 1346 3714 1381 3716
rect 1346 3712 1450 3714
rect 2239 3712 2278 3754
rect 2513 3753 2681 3754
rect 1346 3705 2280 3712
rect 1346 3704 1397 3705
rect 1346 3684 1349 3704
rect 1374 3685 1397 3704
rect 1429 3685 2280 3705
rect 1374 3684 2280 3685
rect 1346 3677 2280 3684
rect 1619 3676 2280 3677
rect 433 3648 498 3669
rect 710 3659 750 3662
rect 710 3655 1613 3659
rect 710 3635 1587 3655
rect 1607 3635 1613 3655
rect 710 3632 1613 3635
rect 434 3588 499 3608
rect 434 3570 458 3588
rect 476 3570 499 3588
rect 434 3543 499 3570
rect 710 3543 750 3632
rect 1194 3630 1610 3632
rect 1194 3629 1535 3630
rect 851 3598 961 3612
rect 851 3595 894 3598
rect 851 3590 855 3595
rect 433 3508 750 3543
rect 773 3568 855 3590
rect 884 3568 894 3595
rect 922 3571 929 3598
rect 958 3590 961 3598
rect 958 3571 1023 3590
rect 922 3568 1023 3571
rect 773 3566 1023 3568
rect 434 3432 499 3508
rect 773 3487 810 3566
rect 851 3553 961 3566
rect 925 3497 956 3498
rect 773 3467 782 3487
rect 802 3467 810 3487
rect 773 3457 810 3467
rect 869 3487 956 3497
rect 869 3467 878 3487
rect 898 3467 956 3487
rect 869 3458 956 3467
rect 869 3457 906 3458
rect 434 3414 456 3432
rect 474 3414 499 3432
rect 434 3393 499 3414
rect 647 3412 712 3421
rect 647 3375 657 3412
rect 697 3404 712 3412
rect 925 3405 956 3458
rect 986 3487 1023 3566
rect 1138 3497 1169 3498
rect 986 3467 995 3487
rect 1015 3467 1023 3487
rect 986 3457 1023 3467
rect 1082 3490 1169 3497
rect 1082 3487 1143 3490
rect 1082 3467 1091 3487
rect 1111 3470 1143 3487
rect 1164 3470 1169 3490
rect 1111 3467 1169 3470
rect 1082 3460 1169 3467
rect 1194 3487 1231 3629
rect 1497 3628 1534 3629
rect 1346 3497 1382 3498
rect 1194 3467 1203 3487
rect 1223 3467 1231 3487
rect 1082 3458 1138 3460
rect 1082 3457 1119 3458
rect 1194 3457 1231 3467
rect 1290 3487 1438 3497
rect 1538 3494 1634 3496
rect 1290 3467 1299 3487
rect 1319 3467 1409 3487
rect 1429 3467 1438 3487
rect 1290 3461 1438 3467
rect 1290 3458 1354 3461
rect 1290 3457 1327 3458
rect 1346 3431 1354 3458
rect 1375 3458 1438 3461
rect 1496 3487 1634 3494
rect 1496 3467 1505 3487
rect 1525 3467 1634 3487
rect 1496 3458 1634 3467
rect 1375 3431 1382 3458
rect 1401 3457 1438 3458
rect 1497 3457 1534 3458
rect 1346 3406 1382 3431
rect 817 3404 858 3405
rect 697 3397 858 3404
rect 697 3377 827 3397
rect 847 3377 858 3397
rect 697 3375 858 3377
rect 647 3369 858 3375
rect 925 3401 1284 3405
rect 925 3396 1247 3401
rect 925 3372 1038 3396
rect 1062 3377 1247 3396
rect 1271 3377 1284 3401
rect 1062 3372 1284 3377
rect 925 3369 1284 3372
rect 1346 3369 1381 3406
rect 1449 3403 1549 3406
rect 1449 3399 1516 3403
rect 1449 3373 1461 3399
rect 1487 3377 1516 3399
rect 1542 3377 1549 3403
rect 1487 3373 1549 3377
rect 1449 3369 1549 3373
rect 647 3356 714 3369
rect 439 3333 495 3353
rect 439 3315 458 3333
rect 476 3315 495 3333
rect 439 3202 495 3315
rect 647 3335 661 3356
rect 697 3335 714 3356
rect 925 3348 956 3369
rect 1346 3348 1382 3369
rect 768 3347 805 3348
rect 647 3328 714 3335
rect 767 3338 805 3347
rect 439 3073 494 3202
rect 647 3176 712 3328
rect 767 3318 776 3338
rect 796 3318 805 3338
rect 767 3310 805 3318
rect 871 3342 956 3348
rect 981 3347 1018 3348
rect 871 3322 879 3342
rect 899 3322 956 3342
rect 871 3314 956 3322
rect 980 3338 1018 3347
rect 980 3318 989 3338
rect 1009 3318 1018 3338
rect 871 3313 907 3314
rect 980 3310 1018 3318
rect 1084 3342 1169 3348
rect 1189 3347 1226 3348
rect 1084 3322 1092 3342
rect 1112 3341 1169 3342
rect 1112 3322 1141 3341
rect 1084 3321 1141 3322
rect 1162 3321 1169 3341
rect 1084 3314 1169 3321
rect 1188 3338 1226 3347
rect 1188 3318 1197 3338
rect 1217 3318 1226 3338
rect 1084 3313 1120 3314
rect 1188 3310 1226 3318
rect 1292 3342 1436 3348
rect 1292 3322 1300 3342
rect 1320 3322 1408 3342
rect 1428 3322 1436 3342
rect 1292 3314 1436 3322
rect 1292 3313 1328 3314
rect 1400 3313 1436 3314
rect 1502 3347 1539 3348
rect 1502 3346 1540 3347
rect 1502 3338 1566 3346
rect 1502 3318 1511 3338
rect 1531 3324 1566 3338
rect 1586 3324 1589 3344
rect 1531 3319 1589 3324
rect 1531 3318 1566 3319
rect 768 3281 805 3310
rect 769 3279 805 3281
rect 981 3279 1018 3310
rect 769 3257 1018 3279
rect 850 3251 961 3257
rect 850 3243 891 3251
rect 850 3223 858 3243
rect 877 3223 891 3243
rect 850 3221 891 3223
rect 919 3243 961 3251
rect 919 3223 935 3243
rect 954 3223 961 3243
rect 919 3221 961 3223
rect 850 3206 961 3221
rect 1189 3211 1226 3310
rect 1502 3306 1566 3318
rect 852 3197 956 3206
rect 640 3166 761 3176
rect 640 3164 709 3166
rect 640 3123 653 3164
rect 690 3125 709 3164
rect 746 3125 761 3166
rect 690 3123 761 3125
rect 640 3105 761 3123
rect 433 3061 494 3073
rect 1187 3061 1228 3211
rect 1606 3203 1633 3458
rect 1695 3448 1775 3459
rect 1695 3422 1712 3448
rect 1752 3422 1775 3448
rect 1695 3395 1775 3422
rect 1695 3369 1716 3395
rect 1756 3369 1775 3395
rect 1695 3350 1775 3369
rect 1695 3324 1719 3350
rect 1759 3324 1775 3350
rect 1695 3273 1775 3324
rect 433 3058 1228 3061
rect 1607 3072 1633 3203
rect 1697 3117 1767 3273
rect 1696 3101 1772 3117
rect 1607 3058 1635 3072
rect 433 3023 1635 3058
rect 1696 3064 1711 3101
rect 1755 3064 1772 3101
rect 1696 3044 1772 3064
rect 2810 3094 2880 4003
rect 2979 3402 3060 4151
rect 3884 4046 3920 4346
rect 3808 4017 3921 4046
rect 3808 3652 3839 4017
rect 3732 3632 4125 3652
rect 4145 3632 4148 3652
rect 3732 3627 4148 3632
rect 3732 3626 4073 3627
rect 3389 3595 3499 3609
rect 3389 3592 3432 3595
rect 3389 3587 3393 3592
rect 3311 3565 3393 3587
rect 3422 3565 3432 3592
rect 3460 3568 3467 3595
rect 3496 3587 3499 3595
rect 3496 3568 3561 3587
rect 3460 3565 3561 3568
rect 3311 3563 3561 3565
rect 3311 3484 3348 3563
rect 3389 3550 3499 3563
rect 3463 3494 3494 3495
rect 3311 3464 3320 3484
rect 3340 3464 3348 3484
rect 3311 3454 3348 3464
rect 3407 3484 3494 3494
rect 3407 3464 3416 3484
rect 3436 3464 3494 3484
rect 3407 3455 3494 3464
rect 3407 3454 3444 3455
rect 3463 3402 3494 3455
rect 3524 3484 3561 3563
rect 3676 3494 3707 3495
rect 3524 3464 3533 3484
rect 3553 3464 3561 3484
rect 3524 3454 3561 3464
rect 3620 3487 3707 3494
rect 3620 3484 3681 3487
rect 3620 3464 3629 3484
rect 3649 3467 3681 3484
rect 3702 3467 3707 3487
rect 3649 3464 3707 3467
rect 3620 3457 3707 3464
rect 3732 3484 3769 3626
rect 4035 3625 4072 3626
rect 3884 3494 3920 3495
rect 3732 3464 3741 3484
rect 3761 3464 3769 3484
rect 3620 3455 3676 3457
rect 3620 3454 3657 3455
rect 3732 3454 3769 3464
rect 3828 3484 3976 3494
rect 4076 3491 4172 3493
rect 3828 3464 3837 3484
rect 3857 3464 3947 3484
rect 3967 3464 3976 3484
rect 3828 3458 3976 3464
rect 3828 3455 3892 3458
rect 3828 3454 3865 3455
rect 3884 3428 3892 3455
rect 3913 3455 3976 3458
rect 4034 3484 4172 3491
rect 4034 3464 4043 3484
rect 4063 3464 4172 3484
rect 4034 3455 4172 3464
rect 3913 3428 3920 3455
rect 3939 3454 3976 3455
rect 4035 3454 4072 3455
rect 3884 3403 3920 3428
rect 2979 3401 3313 3402
rect 3355 3401 3396 3402
rect 2979 3394 3396 3401
rect 2979 3374 3365 3394
rect 3385 3374 3396 3394
rect 2979 3366 3396 3374
rect 3463 3398 3822 3402
rect 3463 3393 3785 3398
rect 3463 3369 3576 3393
rect 3600 3374 3785 3393
rect 3809 3374 3822 3398
rect 3600 3369 3822 3374
rect 3463 3366 3822 3369
rect 3884 3366 3919 3403
rect 3987 3400 4087 3403
rect 3987 3396 4054 3400
rect 3987 3370 3999 3396
rect 4025 3374 4054 3396
rect 4080 3374 4087 3400
rect 4025 3370 4087 3374
rect 3987 3366 4087 3370
rect 2979 3362 3313 3366
rect 3463 3345 3494 3366
rect 3884 3345 3920 3366
rect 3306 3344 3343 3345
rect 3305 3335 3343 3344
rect 3305 3315 3314 3335
rect 3334 3315 3343 3335
rect 3305 3307 3343 3315
rect 3409 3339 3494 3345
rect 3519 3344 3556 3345
rect 3409 3319 3417 3339
rect 3437 3319 3494 3339
rect 3409 3311 3494 3319
rect 3518 3335 3556 3344
rect 3518 3315 3527 3335
rect 3547 3315 3556 3335
rect 3409 3310 3445 3311
rect 3518 3307 3556 3315
rect 3622 3339 3707 3345
rect 3727 3344 3764 3345
rect 3622 3319 3630 3339
rect 3650 3338 3707 3339
rect 3650 3319 3679 3338
rect 3622 3318 3679 3319
rect 3700 3318 3707 3338
rect 3622 3311 3707 3318
rect 3726 3335 3764 3344
rect 3726 3315 3735 3335
rect 3755 3315 3764 3335
rect 3622 3310 3658 3311
rect 3726 3307 3764 3315
rect 3830 3339 3974 3345
rect 3830 3319 3838 3339
rect 3858 3319 3946 3339
rect 3966 3319 3974 3339
rect 3830 3311 3974 3319
rect 3830 3310 3866 3311
rect 3938 3310 3974 3311
rect 4040 3344 4077 3345
rect 4040 3343 4078 3344
rect 4040 3335 4104 3343
rect 4040 3315 4049 3335
rect 4069 3321 4104 3335
rect 4124 3321 4127 3341
rect 4069 3316 4127 3321
rect 4069 3315 4104 3316
rect 3306 3278 3343 3307
rect 3307 3276 3343 3278
rect 3519 3276 3556 3307
rect 3307 3254 3556 3276
rect 3388 3248 3499 3254
rect 3388 3240 3429 3248
rect 3388 3220 3396 3240
rect 3415 3220 3429 3240
rect 3388 3218 3429 3220
rect 3457 3240 3499 3248
rect 3457 3220 3473 3240
rect 3492 3220 3499 3240
rect 3457 3218 3499 3220
rect 3388 3203 3499 3218
rect 3727 3186 3764 3307
rect 4040 3303 4104 3315
rect 3845 3186 3874 3190
rect 4144 3188 4171 3455
rect 4003 3186 4171 3188
rect 3727 3160 4171 3186
rect 2810 3044 2882 3094
rect 433 2948 494 3023
rect 852 3021 956 3023
rect 1187 3021 1228 3023
rect 1696 2978 1706 3044
rect 1760 2978 1772 3044
rect 1696 2954 1772 2978
rect 435 2818 494 2948
rect 1348 2899 1420 2900
rect 1347 2891 1446 2899
rect 1347 2888 1399 2891
rect 1347 2853 1355 2888
rect 1380 2853 1399 2888
rect 1424 2880 1446 2891
rect 1424 2879 2291 2880
rect 1424 2853 2292 2879
rect 1347 2843 2292 2853
rect 1347 2841 1446 2843
rect 435 2800 457 2818
rect 475 2800 494 2818
rect 435 2778 494 2800
rect 702 2814 1234 2819
rect 702 2794 1588 2814
rect 1608 2794 1611 2814
rect 2247 2810 2292 2843
rect 702 2790 1611 2794
rect 702 2743 745 2790
rect 1195 2789 1611 2790
rect 2243 2790 2636 2810
rect 2656 2790 2659 2810
rect 1195 2788 1536 2789
rect 852 2757 962 2771
rect 852 2754 895 2757
rect 852 2749 856 2754
rect 690 2742 745 2743
rect 434 2719 745 2742
rect 434 2701 459 2719
rect 477 2707 745 2719
rect 774 2727 856 2749
rect 885 2727 895 2754
rect 923 2730 930 2757
rect 959 2749 962 2757
rect 959 2730 1024 2749
rect 923 2727 1024 2730
rect 774 2725 1024 2727
rect 477 2701 499 2707
rect 434 2562 499 2701
rect 774 2646 811 2725
rect 852 2712 962 2725
rect 926 2656 957 2657
rect 774 2626 783 2646
rect 803 2626 811 2646
rect 434 2544 457 2562
rect 475 2544 499 2562
rect 434 2527 499 2544
rect 654 2608 722 2621
rect 774 2616 811 2626
rect 870 2646 957 2656
rect 870 2626 879 2646
rect 899 2626 957 2646
rect 870 2617 957 2626
rect 870 2616 907 2617
rect 654 2566 661 2608
rect 710 2566 722 2608
rect 654 2563 722 2566
rect 926 2564 957 2617
rect 987 2646 1024 2725
rect 1139 2656 1170 2657
rect 987 2626 996 2646
rect 1016 2626 1024 2646
rect 987 2616 1024 2626
rect 1083 2649 1170 2656
rect 1083 2646 1144 2649
rect 1083 2626 1092 2646
rect 1112 2629 1144 2646
rect 1165 2629 1170 2649
rect 1112 2626 1170 2629
rect 1083 2619 1170 2626
rect 1195 2646 1232 2788
rect 1498 2787 1535 2788
rect 2243 2785 2659 2790
rect 2243 2784 2584 2785
rect 1900 2753 2010 2767
rect 1900 2750 1943 2753
rect 1900 2745 1904 2750
rect 1822 2723 1904 2745
rect 1933 2723 1943 2750
rect 1971 2726 1978 2753
rect 2007 2745 2010 2753
rect 2007 2726 2072 2745
rect 1971 2723 2072 2726
rect 1822 2721 2072 2723
rect 1347 2656 1383 2657
rect 1195 2626 1204 2646
rect 1224 2626 1232 2646
rect 1083 2617 1139 2619
rect 1083 2616 1120 2617
rect 1195 2616 1232 2626
rect 1291 2646 1439 2656
rect 1539 2653 1635 2655
rect 1291 2626 1300 2646
rect 1320 2626 1410 2646
rect 1430 2626 1439 2646
rect 1291 2620 1439 2626
rect 1291 2617 1355 2620
rect 1291 2616 1328 2617
rect 1347 2590 1355 2617
rect 1376 2617 1439 2620
rect 1497 2646 1635 2653
rect 1497 2626 1506 2646
rect 1526 2626 1635 2646
rect 1497 2617 1635 2626
rect 1822 2642 1859 2721
rect 1900 2708 2010 2721
rect 1974 2652 2005 2653
rect 1822 2622 1831 2642
rect 1851 2622 1859 2642
rect 1376 2590 1383 2617
rect 1402 2616 1439 2617
rect 1498 2616 1535 2617
rect 1347 2565 1383 2590
rect 818 2563 859 2564
rect 654 2556 859 2563
rect 654 2545 828 2556
rect 654 2512 662 2545
rect 655 2503 662 2512
rect 711 2536 828 2545
rect 848 2536 859 2556
rect 711 2528 859 2536
rect 926 2560 1285 2564
rect 926 2555 1248 2560
rect 926 2531 1039 2555
rect 1063 2536 1248 2555
rect 1272 2536 1285 2560
rect 1063 2531 1285 2536
rect 926 2528 1285 2531
rect 1347 2528 1382 2565
rect 1450 2562 1550 2565
rect 1450 2558 1517 2562
rect 1450 2532 1462 2558
rect 1488 2536 1517 2558
rect 1543 2536 1550 2562
rect 1488 2532 1550 2536
rect 1450 2528 1550 2532
rect 711 2512 722 2528
rect 711 2503 719 2512
rect 926 2507 957 2528
rect 1347 2507 1383 2528
rect 769 2506 806 2507
rect 434 2463 499 2482
rect 434 2445 459 2463
rect 477 2445 499 2463
rect 434 2244 499 2445
rect 655 2319 719 2503
rect 768 2497 806 2506
rect 768 2477 777 2497
rect 797 2477 806 2497
rect 768 2469 806 2477
rect 872 2501 957 2507
rect 982 2506 1019 2507
rect 872 2481 880 2501
rect 900 2481 957 2501
rect 872 2473 957 2481
rect 981 2497 1019 2506
rect 981 2477 990 2497
rect 1010 2477 1019 2497
rect 872 2472 908 2473
rect 981 2469 1019 2477
rect 1085 2501 1170 2507
rect 1190 2506 1227 2507
rect 1085 2481 1093 2501
rect 1113 2500 1170 2501
rect 1113 2481 1142 2500
rect 1085 2480 1142 2481
rect 1163 2480 1170 2500
rect 1085 2473 1170 2480
rect 1189 2497 1227 2506
rect 1189 2477 1198 2497
rect 1218 2477 1227 2497
rect 1085 2472 1121 2473
rect 1189 2469 1227 2477
rect 1293 2501 1437 2507
rect 1293 2481 1301 2501
rect 1321 2481 1409 2501
rect 1429 2481 1437 2501
rect 1293 2473 1437 2481
rect 1293 2472 1329 2473
rect 1401 2472 1437 2473
rect 1503 2506 1540 2507
rect 1503 2505 1541 2506
rect 1503 2497 1567 2505
rect 1503 2477 1512 2497
rect 1532 2483 1567 2497
rect 1587 2483 1590 2503
rect 1532 2478 1590 2483
rect 1532 2477 1567 2478
rect 769 2440 806 2469
rect 770 2438 806 2440
rect 982 2438 1019 2469
rect 770 2416 1019 2438
rect 851 2410 962 2416
rect 851 2402 892 2410
rect 851 2382 859 2402
rect 878 2382 892 2402
rect 851 2380 892 2382
rect 920 2402 962 2410
rect 920 2382 936 2402
rect 955 2382 962 2402
rect 920 2380 962 2382
rect 851 2365 962 2380
rect 655 2309 723 2319
rect 655 2276 672 2309
rect 712 2276 723 2309
rect 655 2264 723 2276
rect 655 2262 719 2264
rect 1190 2245 1227 2469
rect 1503 2465 1567 2477
rect 1607 2247 1634 2617
rect 1822 2612 1859 2622
rect 1918 2642 2005 2652
rect 1918 2622 1927 2642
rect 1947 2622 2005 2642
rect 1918 2613 2005 2622
rect 1918 2612 1955 2613
rect 1698 2599 1768 2604
rect 1693 2593 1768 2599
rect 1693 2560 1701 2593
rect 1754 2560 1768 2593
rect 1974 2560 2005 2613
rect 2035 2642 2072 2721
rect 2187 2652 2218 2653
rect 2035 2622 2044 2642
rect 2064 2622 2072 2642
rect 2035 2612 2072 2622
rect 2131 2645 2218 2652
rect 2131 2642 2192 2645
rect 2131 2622 2140 2642
rect 2160 2625 2192 2642
rect 2213 2625 2218 2645
rect 2160 2622 2218 2625
rect 2131 2615 2218 2622
rect 2243 2642 2280 2784
rect 2546 2783 2583 2784
rect 2395 2652 2431 2653
rect 2243 2622 2252 2642
rect 2272 2622 2280 2642
rect 2131 2613 2187 2615
rect 2131 2612 2168 2613
rect 2243 2612 2280 2622
rect 2339 2642 2487 2652
rect 2587 2649 2683 2651
rect 2339 2622 2348 2642
rect 2368 2622 2458 2642
rect 2478 2622 2487 2642
rect 2339 2616 2487 2622
rect 2339 2613 2403 2616
rect 2339 2612 2376 2613
rect 2395 2586 2403 2613
rect 2424 2613 2487 2616
rect 2545 2642 2683 2649
rect 2545 2622 2554 2642
rect 2574 2622 2683 2642
rect 2545 2613 2683 2622
rect 2424 2586 2431 2613
rect 2450 2612 2487 2613
rect 2546 2612 2583 2613
rect 2395 2561 2431 2586
rect 1693 2559 1776 2560
rect 1866 2559 1907 2560
rect 1693 2552 1907 2559
rect 1693 2535 1876 2552
rect 1693 2502 1706 2535
rect 1759 2532 1876 2535
rect 1896 2532 1907 2552
rect 1759 2524 1907 2532
rect 1974 2556 2333 2560
rect 1974 2551 2296 2556
rect 1974 2527 2087 2551
rect 2111 2532 2296 2551
rect 2320 2532 2333 2556
rect 2111 2527 2333 2532
rect 1974 2524 2333 2527
rect 2395 2524 2430 2561
rect 2498 2558 2598 2561
rect 2498 2554 2565 2558
rect 2498 2528 2510 2554
rect 2536 2532 2565 2554
rect 2591 2532 2598 2558
rect 2536 2528 2598 2532
rect 2498 2524 2598 2528
rect 1759 2502 1776 2524
rect 1974 2503 2005 2524
rect 2395 2503 2431 2524
rect 1817 2502 1854 2503
rect 1693 2488 1776 2502
rect 1466 2245 1634 2247
rect 1190 2244 1634 2245
rect 434 2214 1634 2244
rect 1704 2278 1776 2488
rect 1816 2493 1854 2502
rect 1816 2473 1825 2493
rect 1845 2473 1854 2493
rect 1816 2465 1854 2473
rect 1920 2497 2005 2503
rect 2030 2502 2067 2503
rect 1920 2477 1928 2497
rect 1948 2477 2005 2497
rect 1920 2469 2005 2477
rect 2029 2493 2067 2502
rect 2029 2473 2038 2493
rect 2058 2473 2067 2493
rect 1920 2468 1956 2469
rect 2029 2465 2067 2473
rect 2133 2497 2218 2503
rect 2238 2502 2275 2503
rect 2133 2477 2141 2497
rect 2161 2496 2218 2497
rect 2161 2477 2190 2496
rect 2133 2476 2190 2477
rect 2211 2476 2218 2496
rect 2133 2469 2218 2476
rect 2237 2493 2275 2502
rect 2237 2473 2246 2493
rect 2266 2473 2275 2493
rect 2133 2468 2169 2469
rect 2237 2465 2275 2473
rect 2341 2497 2485 2503
rect 2341 2477 2349 2497
rect 2369 2477 2457 2497
rect 2477 2477 2485 2497
rect 2341 2469 2485 2477
rect 2341 2468 2377 2469
rect 2449 2468 2485 2469
rect 2551 2502 2588 2503
rect 2551 2501 2589 2502
rect 2551 2493 2615 2501
rect 2551 2473 2560 2493
rect 2580 2479 2615 2493
rect 2635 2479 2638 2499
rect 2580 2474 2638 2479
rect 2580 2473 2615 2474
rect 1817 2436 1854 2465
rect 1818 2434 1854 2436
rect 2030 2434 2067 2465
rect 1818 2412 2067 2434
rect 1899 2406 2010 2412
rect 1899 2398 1940 2406
rect 1899 2378 1907 2398
rect 1926 2378 1940 2398
rect 1899 2376 1940 2378
rect 1968 2398 2010 2406
rect 1968 2378 1984 2398
rect 2003 2378 2010 2398
rect 1968 2376 2010 2378
rect 1899 2361 2010 2376
rect 1704 2239 1723 2278
rect 1768 2239 1776 2278
rect 1704 2222 1776 2239
rect 2238 2266 2275 2465
rect 2551 2461 2615 2473
rect 2238 2260 2279 2266
rect 2655 2262 2682 2613
rect 2811 2565 2882 3044
rect 3686 2892 3731 2901
rect 3686 2854 3696 2892
rect 3721 2854 3731 2892
rect 3686 2843 3731 2854
rect 3689 2835 3731 2843
rect 2811 2481 2880 2565
rect 2514 2260 2682 2262
rect 2238 2234 2682 2260
rect 434 2167 499 2214
rect 434 2149 457 2167
rect 475 2149 499 2167
rect 1347 2194 1382 2196
rect 1347 2192 1451 2194
rect 2240 2192 2279 2234
rect 2514 2233 2682 2234
rect 1347 2185 2281 2192
rect 1347 2184 1398 2185
rect 1347 2164 1350 2184
rect 1375 2165 1398 2184
rect 1430 2165 2281 2185
rect 1375 2164 2281 2165
rect 1347 2157 2281 2164
rect 1620 2156 2281 2157
rect 434 2128 499 2149
rect 711 2139 751 2142
rect 711 2135 1614 2139
rect 711 2115 1588 2135
rect 1608 2115 1614 2135
rect 711 2112 1614 2115
rect 435 2068 500 2088
rect 435 2050 459 2068
rect 477 2050 500 2068
rect 435 2023 500 2050
rect 711 2023 751 2112
rect 1195 2110 1611 2112
rect 1195 2109 1536 2110
rect 852 2078 962 2092
rect 852 2075 895 2078
rect 852 2070 856 2075
rect 434 1988 751 2023
rect 774 2048 856 2070
rect 885 2048 895 2075
rect 923 2051 930 2078
rect 959 2070 962 2078
rect 959 2051 1024 2070
rect 923 2048 1024 2051
rect 774 2046 1024 2048
rect 435 1912 500 1988
rect 774 1967 811 2046
rect 852 2033 962 2046
rect 926 1977 957 1978
rect 774 1947 783 1967
rect 803 1947 811 1967
rect 774 1937 811 1947
rect 870 1967 957 1977
rect 870 1947 879 1967
rect 899 1947 957 1967
rect 870 1938 957 1947
rect 870 1937 907 1938
rect 435 1894 457 1912
rect 475 1894 500 1912
rect 435 1873 500 1894
rect 648 1892 713 1901
rect 648 1855 658 1892
rect 698 1884 713 1892
rect 926 1885 957 1938
rect 987 1967 1024 2046
rect 1139 1977 1170 1978
rect 987 1947 996 1967
rect 1016 1947 1024 1967
rect 987 1937 1024 1947
rect 1083 1970 1170 1977
rect 1083 1967 1144 1970
rect 1083 1947 1092 1967
rect 1112 1950 1144 1967
rect 1165 1950 1170 1970
rect 1112 1947 1170 1950
rect 1083 1940 1170 1947
rect 1195 1967 1232 2109
rect 1498 2108 1535 2109
rect 1347 1977 1383 1978
rect 1195 1947 1204 1967
rect 1224 1947 1232 1967
rect 1083 1938 1139 1940
rect 1083 1937 1120 1938
rect 1195 1937 1232 1947
rect 1291 1967 1439 1977
rect 1539 1974 1635 1976
rect 1291 1947 1300 1967
rect 1320 1947 1410 1967
rect 1430 1947 1439 1967
rect 1291 1941 1439 1947
rect 1291 1938 1355 1941
rect 1291 1937 1328 1938
rect 1347 1911 1355 1938
rect 1376 1938 1439 1941
rect 1497 1967 1635 1974
rect 1497 1947 1506 1967
rect 1526 1947 1635 1967
rect 1497 1938 1635 1947
rect 1376 1911 1383 1938
rect 1402 1937 1439 1938
rect 1498 1937 1535 1938
rect 1347 1886 1383 1911
rect 818 1884 859 1885
rect 698 1877 859 1884
rect 698 1857 828 1877
rect 848 1857 859 1877
rect 698 1855 859 1857
rect 648 1849 859 1855
rect 926 1881 1285 1885
rect 926 1876 1248 1881
rect 926 1852 1039 1876
rect 1063 1857 1248 1876
rect 1272 1857 1285 1881
rect 1063 1852 1285 1857
rect 926 1849 1285 1852
rect 1347 1849 1382 1886
rect 1450 1883 1550 1886
rect 1450 1879 1517 1883
rect 1450 1853 1462 1879
rect 1488 1857 1517 1879
rect 1543 1857 1550 1883
rect 1488 1853 1550 1857
rect 1450 1849 1550 1853
rect 648 1836 715 1849
rect 440 1813 496 1833
rect 440 1795 459 1813
rect 477 1795 496 1813
rect 440 1682 496 1795
rect 648 1815 662 1836
rect 698 1815 715 1836
rect 926 1828 957 1849
rect 1347 1828 1383 1849
rect 769 1827 806 1828
rect 648 1808 715 1815
rect 768 1818 806 1827
rect 440 1544 495 1682
rect 648 1656 713 1808
rect 768 1798 777 1818
rect 797 1798 806 1818
rect 768 1790 806 1798
rect 872 1822 957 1828
rect 982 1827 1019 1828
rect 872 1802 880 1822
rect 900 1802 957 1822
rect 872 1794 957 1802
rect 981 1818 1019 1827
rect 981 1798 990 1818
rect 1010 1798 1019 1818
rect 872 1793 908 1794
rect 981 1790 1019 1798
rect 1085 1822 1170 1828
rect 1190 1827 1227 1828
rect 1085 1802 1093 1822
rect 1113 1821 1170 1822
rect 1113 1802 1142 1821
rect 1085 1801 1142 1802
rect 1163 1801 1170 1821
rect 1085 1794 1170 1801
rect 1189 1818 1227 1827
rect 1189 1798 1198 1818
rect 1218 1798 1227 1818
rect 1085 1793 1121 1794
rect 1189 1790 1227 1798
rect 1293 1822 1437 1828
rect 1293 1802 1301 1822
rect 1321 1802 1409 1822
rect 1429 1802 1437 1822
rect 1293 1794 1437 1802
rect 1293 1793 1329 1794
rect 1401 1793 1437 1794
rect 1503 1827 1540 1828
rect 1503 1826 1541 1827
rect 1503 1818 1567 1826
rect 1503 1798 1512 1818
rect 1532 1804 1567 1818
rect 1587 1804 1590 1824
rect 1532 1799 1590 1804
rect 1532 1798 1567 1799
rect 769 1761 806 1790
rect 770 1759 806 1761
rect 982 1759 1019 1790
rect 770 1737 1019 1759
rect 851 1731 962 1737
rect 851 1723 892 1731
rect 851 1703 859 1723
rect 878 1703 892 1723
rect 851 1701 892 1703
rect 920 1723 962 1731
rect 920 1703 936 1723
rect 955 1703 962 1723
rect 920 1701 962 1703
rect 851 1688 962 1701
rect 1190 1691 1227 1790
rect 1503 1786 1567 1798
rect 641 1646 762 1656
rect 641 1644 710 1646
rect 641 1603 654 1644
rect 691 1605 710 1644
rect 747 1605 762 1646
rect 691 1603 762 1605
rect 641 1585 762 1603
rect 433 1541 497 1544
rect 853 1541 957 1547
rect 1188 1541 1229 1691
rect 1607 1683 1634 1938
rect 1696 1928 1776 1939
rect 2815 1930 2877 2481
rect 3689 2130 3732 2835
rect 3845 2221 3874 3160
rect 4003 3159 4171 3160
rect 3843 2200 3880 2221
rect 3843 2163 3854 2200
rect 3871 2163 3880 2200
rect 3843 2153 3880 2163
rect 3689 2110 4083 2130
rect 4103 2110 4106 2130
rect 3690 2105 4106 2110
rect 3690 2104 4031 2105
rect 3347 2073 3457 2087
rect 3347 2070 3390 2073
rect 3347 2065 3351 2070
rect 3269 2043 3351 2065
rect 3380 2043 3390 2070
rect 3418 2046 3425 2073
rect 3454 2065 3457 2073
rect 3454 2046 3519 2065
rect 3418 2043 3519 2046
rect 3269 2041 3519 2043
rect 3269 1962 3306 2041
rect 3347 2028 3457 2041
rect 3421 1972 3452 1973
rect 3269 1942 3278 1962
rect 3298 1942 3306 1962
rect 3269 1932 3306 1942
rect 3365 1962 3452 1972
rect 3365 1942 3374 1962
rect 3394 1942 3452 1962
rect 3365 1933 3452 1942
rect 3365 1932 3402 1933
rect 1696 1902 1713 1928
rect 1753 1902 1776 1928
rect 1696 1875 1776 1902
rect 1696 1849 1717 1875
rect 1757 1849 1776 1875
rect 1696 1830 1776 1849
rect 1696 1804 1720 1830
rect 1760 1804 1776 1830
rect 2809 1868 2881 1930
rect 3421 1880 3452 1933
rect 3482 1962 3519 2041
rect 3634 1972 3665 1973
rect 3482 1942 3491 1962
rect 3511 1942 3519 1962
rect 3482 1932 3519 1942
rect 3578 1965 3665 1972
rect 3578 1962 3639 1965
rect 3578 1942 3587 1962
rect 3607 1945 3639 1962
rect 3660 1945 3665 1965
rect 3607 1942 3665 1945
rect 3578 1935 3665 1942
rect 3690 1962 3727 2104
rect 3993 2103 4030 2104
rect 3842 1972 3878 1973
rect 3690 1942 3699 1962
rect 3719 1942 3727 1962
rect 3578 1933 3634 1935
rect 3578 1932 3615 1933
rect 3690 1932 3727 1942
rect 3786 1962 3934 1972
rect 4034 1969 4130 1971
rect 3786 1942 3795 1962
rect 3815 1942 3905 1962
rect 3925 1942 3934 1962
rect 3786 1936 3934 1942
rect 3786 1933 3850 1936
rect 3786 1932 3823 1933
rect 3842 1906 3850 1933
rect 3871 1933 3934 1936
rect 3992 1962 4130 1969
rect 3992 1942 4001 1962
rect 4021 1942 4130 1962
rect 3992 1933 4130 1942
rect 3871 1906 3878 1933
rect 3897 1932 3934 1933
rect 3993 1932 4030 1933
rect 3842 1881 3878 1906
rect 3313 1879 3354 1880
rect 3233 1874 3354 1879
rect 2809 1845 2827 1868
rect 2853 1845 2881 1868
rect 2809 1825 2881 1845
rect 3184 1872 3354 1874
rect 3184 1861 3323 1872
rect 3184 1838 3207 1861
rect 3233 1852 3323 1861
rect 3343 1852 3354 1872
rect 3233 1844 3354 1852
rect 3421 1876 3780 1880
rect 3421 1871 3743 1876
rect 3421 1847 3534 1871
rect 3558 1852 3743 1871
rect 3767 1852 3780 1876
rect 3558 1847 3780 1852
rect 3421 1844 3780 1847
rect 3842 1844 3877 1881
rect 3945 1878 4045 1881
rect 3945 1874 4012 1878
rect 3945 1848 3957 1874
rect 3983 1852 4012 1874
rect 4038 1852 4045 1878
rect 3983 1848 4045 1852
rect 3945 1844 4045 1848
rect 3233 1838 3241 1844
rect 3184 1830 3241 1838
rect 3421 1823 3452 1844
rect 3842 1823 3878 1844
rect 3264 1822 3301 1823
rect 1696 1753 1776 1804
rect 3263 1813 3301 1822
rect 3263 1793 3272 1813
rect 3292 1793 3301 1813
rect 3263 1785 3301 1793
rect 3367 1817 3452 1823
rect 3477 1822 3514 1823
rect 3367 1797 3375 1817
rect 3395 1797 3452 1817
rect 3367 1789 3452 1797
rect 3476 1813 3514 1822
rect 3476 1793 3485 1813
rect 3505 1793 3514 1813
rect 3367 1788 3403 1789
rect 3476 1785 3514 1793
rect 3580 1817 3665 1823
rect 3685 1822 3722 1823
rect 3580 1797 3588 1817
rect 3608 1816 3665 1817
rect 3608 1797 3637 1816
rect 3580 1796 3637 1797
rect 3658 1796 3665 1816
rect 3580 1789 3665 1796
rect 3684 1813 3722 1822
rect 3684 1793 3693 1813
rect 3713 1793 3722 1813
rect 3580 1788 3616 1789
rect 3684 1785 3722 1793
rect 3788 1817 3932 1823
rect 3788 1797 3796 1817
rect 3816 1797 3904 1817
rect 3924 1797 3932 1817
rect 3788 1789 3932 1797
rect 3788 1788 3824 1789
rect 3896 1788 3932 1789
rect 3998 1822 4035 1823
rect 3998 1821 4036 1822
rect 3998 1813 4062 1821
rect 3998 1793 4007 1813
rect 4027 1799 4062 1813
rect 4082 1799 4085 1819
rect 4027 1794 4085 1799
rect 4027 1793 4062 1794
rect 3264 1756 3301 1785
rect 3265 1754 3301 1756
rect 3477 1754 3514 1785
rect 433 1538 1229 1541
rect 1608 1552 1634 1683
rect 1608 1538 1636 1552
rect 433 1503 1636 1538
rect 1698 1545 1768 1753
rect 3265 1732 3514 1754
rect 3346 1726 3457 1732
rect 3346 1718 3387 1726
rect 3346 1698 3354 1718
rect 3373 1698 3387 1718
rect 3346 1696 3387 1698
rect 3415 1718 3457 1726
rect 3415 1698 3431 1718
rect 3450 1698 3457 1718
rect 3415 1696 3457 1698
rect 3346 1681 3457 1696
rect 3685 1670 3722 1785
rect 3998 1781 4062 1793
rect 433 1442 497 1503
rect 853 1501 957 1503
rect 1188 1501 1229 1503
rect 1698 1500 1719 1545
rect 1699 1479 1719 1500
rect 1749 1500 1768 1545
rect 3678 1664 3725 1670
rect 4102 1666 4129 1933
rect 3961 1664 4129 1666
rect 3678 1638 4129 1664
rect 3678 1503 3725 1638
rect 3961 1637 4129 1638
rect 1749 1479 1766 1500
rect 1699 1460 1766 1479
rect 3676 1454 3735 1503
rect 1348 1452 1420 1453
rect 1347 1444 1446 1452
rect 435 1371 494 1442
rect 1347 1441 1399 1444
rect 1347 1406 1355 1441
rect 1380 1406 1399 1441
rect 1424 1433 1446 1444
rect 1424 1432 2291 1433
rect 1424 1406 2292 1432
rect 3676 1426 3694 1454
rect 3722 1426 3735 1454
rect 3676 1416 3735 1426
rect 1347 1396 2292 1406
rect 1347 1394 1446 1396
rect 435 1353 457 1371
rect 475 1353 494 1371
rect 435 1331 494 1353
rect 702 1367 1234 1372
rect 702 1347 1588 1367
rect 1608 1347 1611 1367
rect 2247 1363 2292 1396
rect 702 1343 1611 1347
rect 702 1296 745 1343
rect 1195 1342 1611 1343
rect 2243 1343 2636 1363
rect 2656 1343 2659 1363
rect 1195 1341 1536 1342
rect 852 1310 962 1324
rect 852 1307 895 1310
rect 852 1302 856 1307
rect 690 1295 745 1296
rect 434 1272 745 1295
rect 434 1254 459 1272
rect 477 1260 745 1272
rect 774 1280 856 1302
rect 885 1280 895 1307
rect 923 1283 930 1310
rect 959 1302 962 1310
rect 959 1283 1024 1302
rect 923 1280 1024 1283
rect 774 1278 1024 1280
rect 477 1254 499 1260
rect 434 1115 499 1254
rect 774 1199 811 1278
rect 852 1265 962 1278
rect 926 1209 957 1210
rect 774 1179 783 1199
rect 803 1179 811 1199
rect 434 1097 457 1115
rect 475 1097 499 1115
rect 434 1080 499 1097
rect 654 1161 722 1174
rect 774 1169 811 1179
rect 870 1199 957 1209
rect 870 1179 879 1199
rect 899 1179 957 1199
rect 870 1170 957 1179
rect 870 1169 907 1170
rect 654 1119 661 1161
rect 710 1119 722 1161
rect 654 1116 722 1119
rect 926 1117 957 1170
rect 987 1199 1024 1278
rect 1139 1209 1170 1210
rect 987 1179 996 1199
rect 1016 1179 1024 1199
rect 987 1169 1024 1179
rect 1083 1202 1170 1209
rect 1083 1199 1144 1202
rect 1083 1179 1092 1199
rect 1112 1182 1144 1199
rect 1165 1182 1170 1202
rect 1112 1179 1170 1182
rect 1083 1172 1170 1179
rect 1195 1199 1232 1341
rect 1498 1340 1535 1341
rect 2243 1338 2659 1343
rect 2243 1337 2584 1338
rect 1900 1306 2010 1320
rect 1900 1303 1943 1306
rect 1900 1298 1904 1303
rect 1822 1276 1904 1298
rect 1933 1276 1943 1303
rect 1971 1279 1978 1306
rect 2007 1298 2010 1306
rect 2007 1279 2072 1298
rect 1971 1276 2072 1279
rect 1822 1274 2072 1276
rect 1347 1209 1383 1210
rect 1195 1179 1204 1199
rect 1224 1179 1232 1199
rect 1083 1170 1139 1172
rect 1083 1169 1120 1170
rect 1195 1169 1232 1179
rect 1291 1199 1439 1209
rect 1539 1206 1635 1208
rect 1291 1179 1300 1199
rect 1320 1179 1410 1199
rect 1430 1179 1439 1199
rect 1291 1173 1439 1179
rect 1291 1170 1355 1173
rect 1291 1169 1328 1170
rect 1347 1143 1355 1170
rect 1376 1170 1439 1173
rect 1497 1199 1635 1206
rect 1497 1179 1506 1199
rect 1526 1179 1635 1199
rect 1497 1170 1635 1179
rect 1822 1195 1859 1274
rect 1900 1261 2010 1274
rect 1974 1205 2005 1206
rect 1822 1175 1831 1195
rect 1851 1175 1859 1195
rect 1376 1143 1383 1170
rect 1402 1169 1439 1170
rect 1498 1169 1535 1170
rect 1347 1118 1383 1143
rect 818 1116 859 1117
rect 654 1109 859 1116
rect 654 1098 828 1109
rect 654 1065 662 1098
rect 655 1056 662 1065
rect 711 1089 828 1098
rect 848 1089 859 1109
rect 711 1081 859 1089
rect 926 1113 1285 1117
rect 926 1108 1248 1113
rect 926 1084 1039 1108
rect 1063 1089 1248 1108
rect 1272 1089 1285 1113
rect 1063 1084 1285 1089
rect 926 1081 1285 1084
rect 1347 1081 1382 1118
rect 1450 1115 1550 1118
rect 1450 1111 1517 1115
rect 1450 1085 1462 1111
rect 1488 1089 1517 1111
rect 1543 1089 1550 1115
rect 1488 1085 1550 1089
rect 1450 1081 1550 1085
rect 711 1065 722 1081
rect 711 1056 719 1065
rect 926 1060 957 1081
rect 1347 1060 1383 1081
rect 769 1059 806 1060
rect 434 1016 499 1035
rect 434 998 459 1016
rect 477 998 499 1016
rect 434 797 499 998
rect 655 872 719 1056
rect 768 1050 806 1059
rect 768 1030 777 1050
rect 797 1030 806 1050
rect 768 1022 806 1030
rect 872 1054 957 1060
rect 982 1059 1019 1060
rect 872 1034 880 1054
rect 900 1034 957 1054
rect 872 1026 957 1034
rect 981 1050 1019 1059
rect 981 1030 990 1050
rect 1010 1030 1019 1050
rect 872 1025 908 1026
rect 981 1022 1019 1030
rect 1085 1054 1170 1060
rect 1190 1059 1227 1060
rect 1085 1034 1093 1054
rect 1113 1053 1170 1054
rect 1113 1034 1142 1053
rect 1085 1033 1142 1034
rect 1163 1033 1170 1053
rect 1085 1026 1170 1033
rect 1189 1050 1227 1059
rect 1189 1030 1198 1050
rect 1218 1030 1227 1050
rect 1085 1025 1121 1026
rect 1189 1022 1227 1030
rect 1293 1054 1437 1060
rect 1293 1034 1301 1054
rect 1321 1034 1409 1054
rect 1429 1034 1437 1054
rect 1293 1026 1437 1034
rect 1293 1025 1329 1026
rect 1401 1025 1437 1026
rect 1503 1059 1540 1060
rect 1503 1058 1541 1059
rect 1503 1050 1567 1058
rect 1503 1030 1512 1050
rect 1532 1036 1567 1050
rect 1587 1036 1590 1056
rect 1532 1031 1590 1036
rect 1532 1030 1567 1031
rect 769 993 806 1022
rect 770 991 806 993
rect 982 991 1019 1022
rect 770 969 1019 991
rect 851 963 962 969
rect 851 955 892 963
rect 851 935 859 955
rect 878 935 892 955
rect 851 933 892 935
rect 920 955 962 963
rect 920 935 936 955
rect 955 935 962 955
rect 920 933 962 935
rect 851 918 962 933
rect 655 862 723 872
rect 655 829 672 862
rect 712 829 723 862
rect 655 817 723 829
rect 655 815 719 817
rect 1190 798 1227 1022
rect 1503 1018 1567 1030
rect 1607 800 1634 1170
rect 1822 1165 1859 1175
rect 1918 1195 2005 1205
rect 1918 1175 1927 1195
rect 1947 1175 2005 1195
rect 1918 1166 2005 1175
rect 1918 1165 1955 1166
rect 1698 1152 1768 1157
rect 1693 1146 1768 1152
rect 1693 1113 1701 1146
rect 1754 1113 1768 1146
rect 1974 1113 2005 1166
rect 2035 1195 2072 1274
rect 2187 1205 2218 1206
rect 2035 1175 2044 1195
rect 2064 1175 2072 1195
rect 2035 1165 2072 1175
rect 2131 1198 2218 1205
rect 2131 1195 2192 1198
rect 2131 1175 2140 1195
rect 2160 1178 2192 1195
rect 2213 1178 2218 1198
rect 2160 1175 2218 1178
rect 2131 1168 2218 1175
rect 2243 1195 2280 1337
rect 2546 1336 2583 1337
rect 2395 1205 2431 1206
rect 2243 1175 2252 1195
rect 2272 1175 2280 1195
rect 2131 1166 2187 1168
rect 2131 1165 2168 1166
rect 2243 1165 2280 1175
rect 2339 1195 2487 1205
rect 2587 1202 2683 1204
rect 2339 1175 2348 1195
rect 2368 1175 2458 1195
rect 2478 1175 2487 1195
rect 2339 1169 2487 1175
rect 2339 1166 2403 1169
rect 2339 1165 2376 1166
rect 2395 1139 2403 1166
rect 2424 1166 2487 1169
rect 2545 1195 2683 1202
rect 2545 1175 2554 1195
rect 2574 1175 2683 1195
rect 2545 1166 2683 1175
rect 2424 1139 2431 1166
rect 2450 1165 2487 1166
rect 2546 1165 2583 1166
rect 2395 1114 2431 1139
rect 1693 1112 1776 1113
rect 1866 1112 1907 1113
rect 1693 1105 1907 1112
rect 1693 1088 1876 1105
rect 1693 1055 1706 1088
rect 1759 1085 1876 1088
rect 1896 1085 1907 1105
rect 1759 1077 1907 1085
rect 1974 1109 2333 1113
rect 1974 1104 2296 1109
rect 1974 1080 2087 1104
rect 2111 1085 2296 1104
rect 2320 1085 2333 1109
rect 2111 1080 2333 1085
rect 1974 1077 2333 1080
rect 2395 1077 2430 1114
rect 2498 1111 2598 1114
rect 2498 1107 2565 1111
rect 2498 1081 2510 1107
rect 2536 1085 2565 1107
rect 2591 1085 2598 1111
rect 2536 1081 2598 1085
rect 2498 1077 2598 1081
rect 1759 1055 1776 1077
rect 1974 1056 2005 1077
rect 2395 1056 2431 1077
rect 1817 1055 1854 1056
rect 1693 1041 1776 1055
rect 1466 798 1634 800
rect 1190 797 1634 798
rect 434 767 1634 797
rect 1704 831 1776 1041
rect 1816 1046 1854 1055
rect 1816 1026 1825 1046
rect 1845 1026 1854 1046
rect 1816 1018 1854 1026
rect 1920 1050 2005 1056
rect 2030 1055 2067 1056
rect 1920 1030 1928 1050
rect 1948 1030 2005 1050
rect 1920 1022 2005 1030
rect 2029 1046 2067 1055
rect 2029 1026 2038 1046
rect 2058 1026 2067 1046
rect 1920 1021 1956 1022
rect 2029 1018 2067 1026
rect 2133 1050 2218 1056
rect 2238 1055 2275 1056
rect 2133 1030 2141 1050
rect 2161 1049 2218 1050
rect 2161 1030 2190 1049
rect 2133 1029 2190 1030
rect 2211 1029 2218 1049
rect 2133 1022 2218 1029
rect 2237 1046 2275 1055
rect 2237 1026 2246 1046
rect 2266 1026 2275 1046
rect 2133 1021 2169 1022
rect 2237 1018 2275 1026
rect 2341 1050 2485 1056
rect 2341 1030 2349 1050
rect 2369 1030 2457 1050
rect 2477 1030 2485 1050
rect 2341 1022 2485 1030
rect 2341 1021 2377 1022
rect 2449 1021 2485 1022
rect 2551 1055 2588 1056
rect 2551 1054 2589 1055
rect 2551 1046 2615 1054
rect 2551 1026 2560 1046
rect 2580 1032 2615 1046
rect 2635 1032 2638 1052
rect 2580 1027 2638 1032
rect 2580 1026 2615 1027
rect 1817 989 1854 1018
rect 1818 987 1854 989
rect 2030 987 2067 1018
rect 1818 965 2067 987
rect 1899 959 2010 965
rect 1899 951 1940 959
rect 1899 931 1907 951
rect 1926 931 1940 951
rect 1899 929 1940 931
rect 1968 951 2010 959
rect 1968 931 1984 951
rect 2003 931 2010 951
rect 1968 929 2010 931
rect 1899 914 2010 929
rect 1704 792 1723 831
rect 1768 792 1776 831
rect 1704 775 1776 792
rect 2238 819 2275 1018
rect 2551 1014 2615 1026
rect 2238 813 2279 819
rect 2655 815 2682 1166
rect 2514 813 2682 815
rect 2238 787 2682 813
rect 434 720 499 767
rect 434 702 457 720
rect 475 702 499 720
rect 1347 747 1382 749
rect 1347 745 1451 747
rect 2240 745 2279 787
rect 2514 786 2682 787
rect 1347 738 2281 745
rect 1347 737 1398 738
rect 1347 717 1350 737
rect 1375 718 1398 737
rect 1430 718 2281 738
rect 1375 717 2281 718
rect 1347 710 2281 717
rect 1620 709 2281 710
rect 434 681 499 702
rect 711 692 751 695
rect 711 688 1614 692
rect 711 668 1588 688
rect 1608 668 1614 688
rect 711 665 1614 668
rect 435 621 500 641
rect 435 603 459 621
rect 477 603 500 621
rect 435 576 500 603
rect 711 576 751 665
rect 1195 663 1611 665
rect 1195 662 1536 663
rect 852 631 962 645
rect 852 628 895 631
rect 852 623 856 628
rect 434 541 751 576
rect 774 601 856 623
rect 885 601 895 628
rect 923 604 930 631
rect 959 623 962 631
rect 959 604 1024 623
rect 923 601 1024 604
rect 774 599 1024 601
rect 435 465 500 541
rect 774 520 811 599
rect 852 586 962 599
rect 926 530 957 531
rect 774 500 783 520
rect 803 500 811 520
rect 774 490 811 500
rect 870 520 957 530
rect 870 500 879 520
rect 899 500 957 520
rect 870 491 957 500
rect 870 490 907 491
rect 435 447 457 465
rect 475 447 500 465
rect 435 426 500 447
rect 648 445 713 454
rect 648 408 658 445
rect 698 437 713 445
rect 926 438 957 491
rect 987 520 1024 599
rect 1139 530 1170 531
rect 987 500 996 520
rect 1016 500 1024 520
rect 987 490 1024 500
rect 1083 523 1170 530
rect 1083 520 1144 523
rect 1083 500 1092 520
rect 1112 503 1144 520
rect 1165 503 1170 523
rect 1112 500 1170 503
rect 1083 493 1170 500
rect 1195 520 1232 662
rect 1498 661 1535 662
rect 1347 530 1383 531
rect 1195 500 1204 520
rect 1224 500 1232 520
rect 1083 491 1139 493
rect 1083 490 1120 491
rect 1195 490 1232 500
rect 1291 520 1439 530
rect 1539 527 1635 529
rect 1291 500 1300 520
rect 1320 500 1410 520
rect 1430 500 1439 520
rect 1291 494 1439 500
rect 1291 491 1355 494
rect 1291 490 1328 491
rect 1347 464 1355 491
rect 1376 491 1439 494
rect 1497 520 1635 527
rect 1497 500 1506 520
rect 1526 500 1635 520
rect 1497 491 1635 500
rect 1376 464 1383 491
rect 1402 490 1439 491
rect 1498 490 1535 491
rect 1347 439 1383 464
rect 818 437 859 438
rect 698 430 859 437
rect 698 410 828 430
rect 848 410 859 430
rect 698 408 859 410
rect 648 402 859 408
rect 926 434 1285 438
rect 926 429 1248 434
rect 926 405 1039 429
rect 1063 410 1248 429
rect 1272 410 1285 434
rect 1063 405 1285 410
rect 926 402 1285 405
rect 1347 402 1382 439
rect 1450 436 1550 439
rect 1450 432 1517 436
rect 1450 406 1462 432
rect 1488 410 1517 432
rect 1543 410 1550 436
rect 1488 406 1550 410
rect 1450 402 1550 406
rect 648 389 715 402
rect 440 366 496 386
rect 440 348 459 366
rect 477 348 496 366
rect 440 235 496 348
rect 648 368 662 389
rect 698 368 715 389
rect 926 381 957 402
rect 1347 381 1383 402
rect 769 380 806 381
rect 648 361 715 368
rect 768 371 806 380
rect 440 94 495 235
rect 648 209 713 361
rect 768 351 777 371
rect 797 351 806 371
rect 768 343 806 351
rect 872 375 957 381
rect 982 380 1019 381
rect 872 355 880 375
rect 900 355 957 375
rect 872 347 957 355
rect 981 371 1019 380
rect 981 351 990 371
rect 1010 351 1019 371
rect 872 346 908 347
rect 981 343 1019 351
rect 1085 375 1170 381
rect 1190 380 1227 381
rect 1085 355 1093 375
rect 1113 374 1170 375
rect 1113 355 1142 374
rect 1085 354 1142 355
rect 1163 354 1170 374
rect 1085 347 1170 354
rect 1189 371 1227 380
rect 1189 351 1198 371
rect 1218 351 1227 371
rect 1085 346 1121 347
rect 1189 343 1227 351
rect 1293 375 1437 381
rect 1293 355 1301 375
rect 1321 355 1409 375
rect 1429 355 1437 375
rect 1293 347 1437 355
rect 1293 346 1329 347
rect 1401 346 1437 347
rect 1503 380 1540 381
rect 1503 379 1541 380
rect 1503 371 1567 379
rect 1503 351 1512 371
rect 1532 357 1567 371
rect 1587 357 1590 377
rect 1532 352 1590 357
rect 1532 351 1567 352
rect 769 314 806 343
rect 770 312 806 314
rect 982 312 1019 343
rect 770 290 1019 312
rect 851 284 962 290
rect 851 276 892 284
rect 851 256 859 276
rect 878 256 892 276
rect 851 254 892 256
rect 920 276 962 284
rect 920 256 936 276
rect 955 256 962 276
rect 920 254 962 256
rect 851 239 962 254
rect 1190 244 1227 343
rect 1503 339 1567 351
rect 641 199 762 209
rect 641 197 710 199
rect 641 156 654 197
rect 691 158 710 197
rect 747 158 762 199
rect 691 156 762 158
rect 641 138 762 156
rect 853 94 957 239
rect 1188 94 1229 244
rect 1607 236 1634 491
rect 1696 481 1776 492
rect 1696 455 1713 481
rect 1753 455 1776 481
rect 1696 428 1776 455
rect 1696 402 1717 428
rect 1757 402 1776 428
rect 1696 383 1776 402
rect 1696 357 1720 383
rect 1760 357 1776 383
rect 1696 306 1776 357
rect 440 91 1229 94
rect 1608 105 1634 236
rect 1608 91 1636 105
rect 440 58 1636 91
rect 442 56 1636 58
rect 853 54 957 56
rect 1188 54 1229 56
rect 1698 53 1768 306
<< viali >>
rect 2826 11926 2863 11974
rect 1356 11828 1381 11863
rect 1400 11828 1425 11866
rect 1589 11769 1609 11789
rect 2406 11829 2431 11864
rect 2450 11829 2475 11867
rect 2637 11765 2657 11785
rect 857 11702 886 11729
rect 931 11705 960 11732
rect 662 11541 711 11583
rect 1145 11604 1166 11624
rect 1905 11698 1934 11725
rect 1979 11701 2008 11728
rect 1356 11565 1377 11595
rect 663 11478 712 11520
rect 1518 11511 1544 11537
rect 1143 11455 1164 11475
rect 1568 11458 1588 11478
rect 860 11357 879 11377
rect 937 11357 956 11377
rect 673 11251 713 11284
rect 1702 11535 1755 11568
rect 2193 11600 2214 11620
rect 2404 11561 2425 11591
rect 1707 11477 1760 11510
rect 2566 11507 2592 11533
rect 2191 11451 2212 11471
rect 2616 11454 2636 11474
rect 1908 11353 1927 11373
rect 1985 11353 2004 11373
rect 1724 11214 1769 11253
rect 2827 11514 2861 11553
rect 1351 11139 1376 11159
rect 1399 11140 1431 11160
rect 1589 11090 1609 11110
rect 857 11023 886 11050
rect 931 11026 960 11053
rect 659 10830 699 10867
rect 1145 10925 1166 10945
rect 3004 11534 3040 11575
rect 2993 11194 3053 11238
rect 4084 11085 4104 11105
rect 3352 11018 3381 11045
rect 3426 11021 3455 11048
rect 1356 10886 1377 10916
rect 1518 10832 1544 10858
rect 663 10790 699 10811
rect 1143 10776 1164 10796
rect 1568 10779 1588 10799
rect 860 10678 879 10698
rect 937 10678 956 10698
rect 655 10578 692 10619
rect 711 10580 748 10621
rect 1714 10877 1754 10903
rect 1718 10824 1758 10850
rect 1721 10779 1761 10805
rect 3640 10920 3661 10940
rect 3851 10881 3872 10911
rect 2993 10780 3047 10821
rect 4013 10827 4039 10853
rect 3638 10771 3659 10791
rect 1720 10454 1750 10520
rect 1356 10381 1381 10416
rect 1400 10381 1425 10419
rect 1589 10322 1609 10342
rect 2637 10318 2657 10338
rect 857 10255 886 10282
rect 931 10258 960 10285
rect 662 10094 711 10136
rect 1145 10157 1166 10177
rect 1905 10251 1934 10278
rect 1979 10254 2008 10281
rect 1356 10118 1377 10148
rect 663 10031 712 10073
rect 1518 10064 1544 10090
rect 1143 10008 1164 10028
rect 1568 10011 1588 10031
rect 860 9910 879 9930
rect 937 9910 956 9930
rect 673 9804 713 9837
rect 1702 10088 1755 10121
rect 2193 10153 2214 10173
rect 2404 10114 2425 10144
rect 1707 10030 1760 10063
rect 2566 10060 2592 10086
rect 2191 10004 2212 10024
rect 2616 10007 2636 10027
rect 1908 9906 1927 9926
rect 1985 9906 2004 9926
rect 1724 9767 1769 9806
rect 3355 10673 3374 10693
rect 3432 10673 3451 10693
rect 4063 10774 4083 10794
rect 3862 10583 3914 10601
rect 3631 10382 3656 10417
rect 3675 10382 3700 10420
rect 3894 10398 3918 10421
rect 3894 10354 3918 10377
rect 1351 9692 1376 9712
rect 1399 9693 1431 9713
rect 1589 9643 1609 9663
rect 857 9576 886 9603
rect 931 9579 960 9606
rect 659 9383 699 9420
rect 1145 9478 1166 9498
rect 1356 9439 1377 9469
rect 1518 9385 1544 9411
rect 663 9343 699 9364
rect 1143 9329 1164 9349
rect 1568 9332 1588 9352
rect 860 9231 879 9251
rect 937 9231 956 9251
rect 655 9131 692 9172
rect 711 9133 748 9174
rect 1714 9430 1754 9456
rect 1718 9377 1758 9403
rect 1721 9332 1761 9358
rect 1713 9072 1757 9109
rect 3899 9735 3919 9756
rect 3940 9740 3960 9761
rect 4127 9640 4147 9660
rect 3395 9573 3424 9600
rect 3469 9576 3498 9603
rect 3683 9475 3704 9495
rect 3894 9436 3915 9466
rect 4056 9382 4082 9408
rect 1708 8986 1762 9052
rect 1357 8861 1382 8896
rect 1401 8861 1426 8899
rect 1590 8802 1610 8822
rect 2638 8798 2658 8818
rect 858 8735 887 8762
rect 932 8738 961 8765
rect 663 8574 712 8616
rect 1146 8637 1167 8657
rect 1906 8731 1935 8758
rect 1980 8734 2009 8761
rect 1357 8598 1378 8628
rect 664 8511 713 8553
rect 1519 8544 1545 8570
rect 1144 8488 1165 8508
rect 1569 8491 1589 8511
rect 861 8390 880 8410
rect 938 8390 957 8410
rect 674 8284 714 8317
rect 1703 8568 1756 8601
rect 2194 8633 2215 8653
rect 2405 8594 2426 8624
rect 1708 8510 1761 8543
rect 2567 8540 2593 8566
rect 2192 8484 2213 8504
rect 2617 8487 2637 8507
rect 1909 8386 1928 8406
rect 1986 8386 2005 8406
rect 1725 8247 1770 8286
rect 1352 8172 1377 8192
rect 1400 8173 1432 8193
rect 1590 8123 1610 8143
rect 858 8056 887 8083
rect 932 8059 961 8086
rect 660 7863 700 7900
rect 1146 7958 1167 7978
rect 1357 7919 1378 7949
rect 1519 7865 1545 7891
rect 664 7823 700 7844
rect 1144 7809 1165 7829
rect 1569 7812 1589 7832
rect 861 7711 880 7731
rect 938 7711 957 7731
rect 656 7611 693 7652
rect 712 7613 749 7654
rect 1715 7910 1755 7936
rect 1719 7857 1759 7883
rect 1722 7812 1762 7838
rect 2829 7853 2855 7876
rect 1721 7487 1751 7553
rect 1357 7414 1382 7449
rect 1401 7414 1426 7452
rect 1590 7355 1610 7375
rect 2638 7351 2658 7371
rect 858 7288 887 7315
rect 932 7291 961 7318
rect 663 7127 712 7169
rect 1146 7190 1167 7210
rect 1906 7284 1935 7311
rect 1980 7287 2009 7314
rect 1357 7151 1378 7181
rect 664 7064 713 7106
rect 1519 7097 1545 7123
rect 1144 7041 1165 7061
rect 1569 7044 1589 7064
rect 861 6943 880 6963
rect 938 6943 957 6963
rect 674 6837 714 6870
rect 1703 7121 1756 7154
rect 2194 7186 2215 7206
rect 2405 7147 2426 7177
rect 1708 7063 1761 7096
rect 2567 7093 2593 7119
rect 2192 7037 2213 7057
rect 2617 7040 2637 7060
rect 1909 6939 1928 6959
rect 1986 6939 2005 6959
rect 1725 6800 1770 6839
rect 1352 6725 1377 6745
rect 1400 6726 1432 6746
rect 1590 6676 1610 6696
rect 858 6609 887 6636
rect 932 6612 961 6639
rect 660 6416 700 6453
rect 1146 6511 1167 6531
rect 1357 6472 1378 6502
rect 1519 6418 1545 6444
rect 664 6376 700 6397
rect 1144 6362 1165 6382
rect 1569 6365 1589 6385
rect 861 6264 880 6284
rect 938 6264 957 6284
rect 656 6164 693 6205
rect 712 6166 749 6207
rect 1715 6463 1755 6489
rect 1719 6410 1759 6436
rect 1722 6365 1762 6391
rect 1713 6044 1759 6092
rect 3681 9326 3702 9346
rect 4106 9329 4126 9349
rect 3398 9228 3417 9248
rect 3475 9228 3494 9248
rect 3698 8862 3723 8900
rect 3856 8171 3873 8208
rect 4085 8118 4105 8138
rect 3353 8051 3382 8078
rect 3427 8054 3456 8081
rect 3641 7953 3662 7973
rect 3852 7914 3873 7944
rect 3209 7846 3235 7869
rect 4014 7860 4040 7886
rect 3639 7804 3660 7824
rect 4064 7807 4084 7827
rect 3356 7706 3375 7726
rect 3433 7706 3452 7726
rect 3696 7434 3724 7462
rect 5193 6667 5213 6687
rect 4461 6600 4490 6627
rect 4535 6603 4564 6630
rect 4749 6502 4770 6522
rect 4960 6463 4981 6493
rect 4257 6404 4281 6428
rect 4314 6405 4338 6429
rect 5122 6409 5148 6435
rect 4747 6353 4768 6373
rect 5172 6356 5192 6376
rect 4464 6255 4483 6275
rect 4541 6255 4560 6275
rect 4800 6162 4829 6196
rect 4799 6102 4828 6136
rect 3015 6017 3059 6045
rect 2824 5918 2861 5966
rect 3012 5960 3056 5988
rect 1354 5820 1379 5855
rect 1398 5820 1423 5858
rect 1587 5761 1607 5781
rect 2404 5821 2429 5856
rect 2448 5821 2473 5859
rect 2635 5757 2655 5777
rect 855 5694 884 5721
rect 929 5697 958 5724
rect 660 5533 709 5575
rect 1143 5596 1164 5616
rect 1903 5690 1932 5717
rect 1977 5693 2006 5720
rect 1354 5557 1375 5587
rect 661 5470 710 5512
rect 1516 5503 1542 5529
rect 1141 5447 1162 5467
rect 1566 5450 1586 5470
rect 858 5349 877 5369
rect 935 5349 954 5369
rect 671 5243 711 5276
rect 1700 5527 1753 5560
rect 2191 5592 2212 5612
rect 2402 5553 2423 5583
rect 1705 5469 1758 5502
rect 2564 5499 2590 5525
rect 2189 5443 2210 5463
rect 2614 5446 2634 5466
rect 1906 5345 1925 5365
rect 1983 5345 2002 5365
rect 1722 5206 1767 5245
rect 2825 5506 2859 5545
rect 1349 5131 1374 5151
rect 1397 5132 1429 5152
rect 1587 5082 1607 5102
rect 855 5015 884 5042
rect 929 5018 958 5045
rect 657 4822 697 4859
rect 1143 4917 1164 4937
rect 3002 5526 3038 5567
rect 2991 5186 3051 5230
rect 4082 5077 4102 5097
rect 3350 5010 3379 5037
rect 3424 5013 3453 5040
rect 1354 4878 1375 4908
rect 1516 4824 1542 4850
rect 661 4782 697 4803
rect 1141 4768 1162 4788
rect 1566 4771 1586 4791
rect 858 4670 877 4690
rect 935 4670 954 4690
rect 653 4570 690 4611
rect 709 4572 746 4613
rect 1712 4869 1752 4895
rect 1716 4816 1756 4842
rect 1719 4771 1759 4797
rect 3638 4912 3659 4932
rect 3849 4873 3870 4903
rect 2991 4772 3045 4813
rect 4011 4819 4037 4845
rect 3636 4763 3657 4783
rect 1718 4446 1748 4512
rect 1354 4373 1379 4408
rect 1398 4373 1423 4411
rect 1587 4314 1607 4334
rect 2635 4310 2655 4330
rect 855 4247 884 4274
rect 929 4250 958 4277
rect 660 4086 709 4128
rect 1143 4149 1164 4169
rect 1903 4243 1932 4270
rect 1977 4246 2006 4273
rect 1354 4110 1375 4140
rect 661 4023 710 4065
rect 1516 4056 1542 4082
rect 1141 4000 1162 4020
rect 1566 4003 1586 4023
rect 858 3902 877 3922
rect 935 3902 954 3922
rect 671 3796 711 3829
rect 1700 4080 1753 4113
rect 2191 4145 2212 4165
rect 2402 4106 2423 4136
rect 1705 4022 1758 4055
rect 2564 4052 2590 4078
rect 2189 3996 2210 4016
rect 2614 3999 2634 4019
rect 1906 3898 1925 3918
rect 1983 3898 2002 3918
rect 1722 3759 1767 3798
rect 3353 4665 3372 4685
rect 3430 4665 3449 4685
rect 4061 4766 4081 4786
rect 3860 4575 3912 4593
rect 3629 4374 3654 4409
rect 3673 4374 3698 4412
rect 3892 4390 3916 4413
rect 3892 4346 3916 4369
rect 1349 3684 1374 3704
rect 1397 3685 1429 3705
rect 1587 3635 1607 3655
rect 855 3568 884 3595
rect 929 3571 958 3598
rect 657 3375 697 3412
rect 1143 3470 1164 3490
rect 1354 3431 1375 3461
rect 1516 3377 1542 3403
rect 661 3335 697 3356
rect 1141 3321 1162 3341
rect 1566 3324 1586 3344
rect 858 3223 877 3243
rect 935 3223 954 3243
rect 653 3123 690 3164
rect 709 3125 746 3166
rect 1712 3422 1752 3448
rect 1716 3369 1756 3395
rect 1719 3324 1759 3350
rect 1711 3064 1755 3101
rect 4125 3632 4145 3652
rect 3393 3565 3422 3592
rect 3467 3568 3496 3595
rect 3681 3467 3702 3487
rect 3892 3428 3913 3458
rect 4054 3374 4080 3400
rect 3679 3318 3700 3338
rect 4104 3321 4124 3341
rect 3396 3220 3415 3240
rect 3473 3220 3492 3240
rect 1706 2978 1760 3044
rect 1355 2853 1380 2888
rect 1399 2853 1424 2891
rect 1588 2794 1608 2814
rect 2636 2790 2656 2810
rect 856 2727 885 2754
rect 930 2730 959 2757
rect 661 2566 710 2608
rect 1144 2629 1165 2649
rect 1904 2723 1933 2750
rect 1978 2726 2007 2753
rect 1355 2590 1376 2620
rect 662 2503 711 2545
rect 1517 2536 1543 2562
rect 1142 2480 1163 2500
rect 1567 2483 1587 2503
rect 859 2382 878 2402
rect 936 2382 955 2402
rect 672 2276 712 2309
rect 1701 2560 1754 2593
rect 2192 2625 2213 2645
rect 2403 2586 2424 2616
rect 1706 2502 1759 2535
rect 2565 2532 2591 2558
rect 2190 2476 2211 2496
rect 2615 2479 2635 2499
rect 1907 2378 1926 2398
rect 1984 2378 2003 2398
rect 1723 2239 1768 2278
rect 3696 2854 3721 2892
rect 1350 2164 1375 2184
rect 1398 2165 1430 2185
rect 1588 2115 1608 2135
rect 856 2048 885 2075
rect 930 2051 959 2078
rect 658 1855 698 1892
rect 1144 1950 1165 1970
rect 1355 1911 1376 1941
rect 1517 1857 1543 1883
rect 662 1815 698 1836
rect 1142 1801 1163 1821
rect 1567 1804 1587 1824
rect 859 1703 878 1723
rect 936 1703 955 1723
rect 654 1603 691 1644
rect 710 1605 747 1646
rect 3854 2163 3871 2200
rect 4083 2110 4103 2130
rect 3351 2043 3380 2070
rect 3425 2046 3454 2073
rect 1713 1902 1753 1928
rect 1717 1849 1757 1875
rect 1720 1804 1760 1830
rect 3639 1945 3660 1965
rect 3850 1906 3871 1936
rect 2827 1845 2853 1868
rect 3207 1838 3233 1861
rect 4012 1852 4038 1878
rect 3637 1796 3658 1816
rect 4062 1799 4082 1819
rect 3354 1698 3373 1718
rect 3431 1698 3450 1718
rect 1719 1479 1749 1545
rect 1355 1406 1380 1441
rect 1399 1406 1424 1444
rect 3694 1426 3722 1454
rect 1588 1347 1608 1367
rect 2636 1343 2656 1363
rect 856 1280 885 1307
rect 930 1283 959 1310
rect 661 1119 710 1161
rect 1144 1182 1165 1202
rect 1904 1276 1933 1303
rect 1978 1279 2007 1306
rect 1355 1143 1376 1173
rect 662 1056 711 1098
rect 1517 1089 1543 1115
rect 1142 1033 1163 1053
rect 1567 1036 1587 1056
rect 859 935 878 955
rect 936 935 955 955
rect 672 829 712 862
rect 1701 1113 1754 1146
rect 2192 1178 2213 1198
rect 2403 1139 2424 1169
rect 1706 1055 1759 1088
rect 2565 1085 2591 1111
rect 2190 1029 2211 1049
rect 2615 1032 2635 1052
rect 1907 931 1926 951
rect 1984 931 2003 951
rect 1723 792 1768 831
rect 1350 717 1375 737
rect 1398 718 1430 738
rect 1588 668 1608 688
rect 856 601 885 628
rect 930 604 959 631
rect 658 408 698 445
rect 1144 503 1165 523
rect 1355 464 1376 494
rect 1517 410 1543 436
rect 662 368 698 389
rect 1142 354 1163 374
rect 1567 357 1587 377
rect 859 256 878 276
rect 936 256 955 276
rect 654 156 691 197
rect 710 158 747 199
rect 1713 455 1753 481
rect 1717 402 1757 428
rect 1720 357 1760 383
<< metal1 >>
rect 174 11395 281 11992
rect 653 11583 725 11983
rect 1349 11874 1421 11875
rect 1348 11866 1447 11874
rect 1348 11863 1400 11866
rect 1348 11828 1356 11863
rect 1381 11828 1400 11863
rect 1425 11828 1447 11866
rect 1348 11816 1447 11828
rect 1349 11797 1417 11816
rect 1350 11794 1383 11797
rect 1585 11794 1617 11795
rect 760 11733 963 11746
rect 760 11700 784 11733
rect 820 11732 963 11733
rect 820 11729 931 11732
rect 820 11702 857 11729
rect 886 11705 931 11729
rect 960 11705 963 11732
rect 886 11702 963 11705
rect 820 11700 963 11702
rect 760 11687 963 11700
rect 760 11686 861 11687
rect 653 11541 662 11583
rect 711 11541 725 11583
rect 653 11520 725 11541
rect 653 11478 663 11520
rect 712 11478 725 11520
rect 653 11460 725 11478
rect 1138 11624 1170 11631
rect 1138 11604 1145 11624
rect 1166 11604 1170 11624
rect 1138 11539 1170 11604
rect 1350 11595 1381 11794
rect 1582 11789 1617 11794
rect 1582 11769 1589 11789
rect 1609 11769 1617 11789
rect 1582 11761 1617 11769
rect 1350 11565 1356 11595
rect 1377 11565 1381 11595
rect 1350 11557 1381 11565
rect 1508 11539 1548 11540
rect 1138 11537 1550 11539
rect 1138 11511 1518 11537
rect 1544 11511 1550 11537
rect 1138 11503 1550 11511
rect 1138 11475 1170 11503
rect 1583 11483 1617 11761
rect 1699 11574 1769 11984
rect 2813 11974 2878 12009
rect 2813 11970 2826 11974
rect 2814 11926 2826 11970
rect 2863 11970 2878 11974
rect 2863 11926 2876 11970
rect 2399 11875 2471 11876
rect 2398 11867 2487 11875
rect 2398 11864 2450 11867
rect 2398 11829 2406 11864
rect 2431 11829 2450 11864
rect 2475 11829 2487 11867
rect 2398 11817 2487 11829
rect 2398 11816 2467 11817
rect 2398 11798 2434 11816
rect 1808 11729 2011 11742
rect 1808 11696 1832 11729
rect 1868 11728 2011 11729
rect 1868 11725 1979 11728
rect 1868 11698 1905 11725
rect 1934 11701 1979 11725
rect 2008 11701 2011 11728
rect 1934 11698 2011 11701
rect 1868 11696 2011 11698
rect 1808 11683 2011 11696
rect 1808 11682 1909 11683
rect 1138 11455 1143 11475
rect 1164 11455 1170 11475
rect 1138 11448 1170 11455
rect 1561 11478 1617 11483
rect 1561 11458 1568 11478
rect 1588 11458 1617 11478
rect 1694 11568 1769 11574
rect 1694 11535 1702 11568
rect 1755 11535 1769 11568
rect 1694 11510 1769 11535
rect 1694 11477 1707 11510
rect 1760 11477 1769 11510
rect 1694 11468 1769 11477
rect 2186 11620 2218 11627
rect 2186 11600 2193 11620
rect 2214 11600 2218 11620
rect 2186 11535 2218 11600
rect 2398 11591 2429 11798
rect 2633 11790 2665 11791
rect 2630 11785 2665 11790
rect 2630 11765 2637 11785
rect 2657 11765 2665 11785
rect 2630 11757 2665 11765
rect 2398 11561 2404 11591
rect 2425 11561 2429 11591
rect 2398 11553 2429 11561
rect 2556 11535 2596 11536
rect 2186 11533 2598 11535
rect 2186 11507 2566 11533
rect 2592 11507 2598 11533
rect 2186 11499 2598 11507
rect 2186 11471 2218 11499
rect 2631 11479 2665 11757
rect 2814 11572 2876 11926
rect 2983 11575 3065 12004
rect 2814 11553 2878 11572
rect 2814 11514 2827 11553
rect 2861 11514 2878 11553
rect 2814 11495 2878 11514
rect 2983 11534 3004 11575
rect 3040 11534 3065 11575
rect 2983 11505 3065 11534
rect 1694 11463 1752 11468
rect 1561 11451 1617 11458
rect 2186 11451 2191 11471
rect 2212 11451 2218 11471
rect 1561 11450 1596 11451
rect 2186 11444 2218 11451
rect 2609 11474 2665 11479
rect 2609 11454 2616 11474
rect 2636 11454 2665 11474
rect 2609 11447 2665 11454
rect 2609 11446 2644 11447
rect 852 11395 963 11399
rect 2635 11395 3748 11396
rect 174 11377 3748 11395
rect 174 11357 860 11377
rect 879 11357 937 11377
rect 956 11373 3748 11377
rect 956 11357 1908 11373
rect 174 11353 1908 11357
rect 1927 11353 1985 11373
rect 2004 11353 3748 11373
rect 174 11339 3748 11353
rect 174 10716 281 11339
rect 1900 11336 2011 11339
rect 660 11290 724 11294
rect 656 11284 724 11290
rect 656 11251 673 11284
rect 713 11251 724 11284
rect 656 11239 724 11251
rect 1707 11253 1772 11275
rect 656 11237 713 11239
rect 660 10876 711 11237
rect 1707 11214 1724 11253
rect 1769 11214 1772 11253
rect 1348 11169 1383 11171
rect 1348 11160 1452 11169
rect 1348 11159 1399 11160
rect 1348 11139 1351 11159
rect 1376 11140 1399 11159
rect 1431 11140 1452 11160
rect 1376 11139 1452 11140
rect 1348 11132 1452 11139
rect 1348 11120 1383 11132
rect 760 11054 963 11067
rect 760 11021 784 11054
rect 820 11053 963 11054
rect 820 11050 931 11053
rect 820 11023 857 11050
rect 886 11026 931 11050
rect 960 11026 963 11053
rect 886 11023 963 11026
rect 820 11021 963 11023
rect 760 11008 963 11021
rect 760 11007 861 11008
rect 1138 10945 1170 10952
rect 1138 10925 1145 10945
rect 1166 10925 1170 10945
rect 649 10867 714 10876
rect 649 10830 659 10867
rect 699 10833 714 10867
rect 1138 10860 1170 10925
rect 1350 10916 1381 11120
rect 1585 11115 1617 11116
rect 1582 11110 1617 11115
rect 1582 11090 1589 11110
rect 1609 11090 1617 11110
rect 1582 11082 1617 11090
rect 1350 10886 1356 10916
rect 1377 10886 1381 10916
rect 1350 10878 1381 10886
rect 1508 10860 1548 10861
rect 1138 10858 1550 10860
rect 699 10830 716 10833
rect 649 10811 716 10830
rect 649 10790 663 10811
rect 699 10790 716 10811
rect 649 10783 716 10790
rect 1138 10832 1518 10858
rect 1544 10832 1550 10858
rect 1138 10824 1550 10832
rect 1138 10796 1170 10824
rect 1583 10804 1617 11082
rect 1707 10914 1772 11214
rect 2978 11238 3071 11253
rect 2978 11194 2993 11238
rect 3053 11194 3071 11238
rect 1138 10776 1143 10796
rect 1164 10776 1170 10796
rect 1138 10769 1170 10776
rect 1561 10799 1617 10804
rect 1561 10779 1568 10799
rect 1588 10779 1617 10799
rect 1561 10772 1617 10779
rect 1697 10903 1777 10914
rect 1697 10877 1714 10903
rect 1754 10877 1777 10903
rect 1697 10850 1777 10877
rect 1697 10824 1718 10850
rect 1758 10824 1777 10850
rect 1697 10805 1777 10824
rect 1697 10779 1721 10805
rect 1761 10779 1777 10805
rect 1561 10771 1596 10772
rect 1697 10767 1777 10779
rect 2978 10821 3071 11194
rect 3255 11049 3458 11062
rect 3255 11016 3279 11049
rect 3315 11048 3458 11049
rect 3315 11045 3426 11048
rect 3315 11018 3352 11045
rect 3381 11021 3426 11045
rect 3455 11021 3458 11048
rect 3381 11018 3458 11021
rect 3315 11016 3458 11018
rect 3255 11003 3458 11016
rect 3255 11002 3356 11003
rect 2978 10780 2993 10821
rect 3047 10780 3071 10821
rect 2978 10773 3071 10780
rect 3633 10940 3665 10947
rect 3633 10920 3640 10940
rect 3661 10920 3665 10940
rect 3633 10855 3665 10920
rect 3845 10911 3876 11112
rect 4080 11110 4112 11111
rect 4077 11105 4112 11110
rect 4077 11085 4084 11105
rect 4104 11085 4112 11105
rect 4077 11077 4112 11085
rect 3845 10881 3851 10911
rect 3872 10881 3876 10911
rect 3845 10873 3876 10881
rect 4003 10855 4043 10856
rect 3633 10853 4045 10855
rect 3633 10827 4013 10853
rect 4039 10827 4045 10853
rect 3633 10819 4045 10827
rect 3633 10791 3665 10819
rect 4078 10799 4112 11077
rect 3633 10771 3638 10791
rect 3659 10771 3665 10791
rect 3633 10764 3665 10771
rect 4056 10794 4112 10799
rect 4056 10774 4063 10794
rect 4083 10774 4112 10794
rect 4056 10767 4112 10774
rect 4056 10766 4091 10767
rect 852 10716 963 10720
rect 2594 10716 4143 10719
rect 172 10698 4143 10716
rect 172 10678 860 10698
rect 879 10678 937 10698
rect 956 10693 4143 10698
rect 956 10678 3355 10693
rect 172 10673 3355 10678
rect 3374 10673 3432 10693
rect 3451 10673 4143 10693
rect 172 10663 4143 10673
rect 172 10660 797 10663
rect 984 10660 4143 10663
rect 174 10432 281 10660
rect 2594 10659 4143 10660
rect 3347 10656 3458 10659
rect 642 10621 763 10631
rect 642 10619 711 10621
rect 642 10578 655 10619
rect 692 10580 711 10619
rect 748 10580 763 10621
rect 692 10578 763 10580
rect 642 10560 763 10578
rect 3847 10601 3933 10605
rect 3847 10583 3862 10601
rect 3914 10583 3933 10601
rect 3847 10574 3933 10583
rect 648 10458 727 10560
rect 1700 10520 1767 10539
rect 1700 10500 1720 10520
rect 174 10377 282 10432
rect 649 10377 727 10458
rect 1699 10454 1720 10500
rect 1750 10500 1767 10520
rect 1750 10470 1769 10500
rect 1750 10454 1770 10470
rect 1699 10438 1770 10454
rect 1349 10427 1421 10428
rect 1348 10419 1447 10427
rect 1348 10416 1400 10419
rect 1348 10381 1356 10416
rect 1381 10381 1400 10416
rect 1425 10381 1447 10419
rect 174 9948 281 10377
rect 653 10136 725 10377
rect 1348 10369 1447 10381
rect 1349 10350 1417 10369
rect 1350 10347 1383 10350
rect 1585 10347 1617 10348
rect 760 10286 963 10299
rect 760 10253 784 10286
rect 820 10285 963 10286
rect 820 10282 931 10285
rect 820 10255 857 10282
rect 886 10258 931 10282
rect 960 10258 963 10285
rect 886 10255 963 10258
rect 820 10253 963 10255
rect 760 10240 963 10253
rect 760 10239 861 10240
rect 653 10094 662 10136
rect 711 10094 725 10136
rect 653 10073 725 10094
rect 653 10031 663 10073
rect 712 10031 725 10073
rect 653 10013 725 10031
rect 1138 10177 1170 10184
rect 1138 10157 1145 10177
rect 1166 10157 1170 10177
rect 1138 10092 1170 10157
rect 1350 10148 1381 10347
rect 1582 10342 1617 10347
rect 1582 10322 1589 10342
rect 1609 10322 1617 10342
rect 1582 10314 1617 10322
rect 1350 10118 1356 10148
rect 1377 10118 1381 10148
rect 1350 10110 1381 10118
rect 1508 10092 1548 10093
rect 1138 10090 1550 10092
rect 1138 10064 1518 10090
rect 1544 10064 1550 10090
rect 1138 10056 1550 10064
rect 1138 10028 1170 10056
rect 1583 10036 1617 10314
rect 1699 10127 1769 10438
rect 3624 10428 3696 10429
rect 3623 10425 3712 10428
rect 2395 10423 3712 10425
rect 2392 10420 3712 10423
rect 2392 10417 3675 10420
rect 2392 10382 3631 10417
rect 3656 10382 3675 10417
rect 3700 10382 3712 10420
rect 2392 10372 3712 10382
rect 3888 10421 3924 10574
rect 3888 10398 3894 10421
rect 3918 10398 3924 10421
rect 3888 10377 3924 10398
rect 2392 10370 3677 10372
rect 2392 10360 2489 10370
rect 2398 10351 2434 10360
rect 3888 10354 3894 10377
rect 3918 10354 3924 10377
rect 1808 10282 2011 10295
rect 1808 10249 1832 10282
rect 1868 10281 2011 10282
rect 1868 10278 1979 10281
rect 1868 10251 1905 10278
rect 1934 10254 1979 10278
rect 2008 10254 2011 10281
rect 1934 10251 2011 10254
rect 1868 10249 2011 10251
rect 1808 10236 2011 10249
rect 1808 10235 1909 10236
rect 1138 10008 1143 10028
rect 1164 10008 1170 10028
rect 1138 10001 1170 10008
rect 1561 10031 1617 10036
rect 1561 10011 1568 10031
rect 1588 10011 1617 10031
rect 1694 10121 1769 10127
rect 1694 10088 1702 10121
rect 1755 10088 1769 10121
rect 1694 10063 1769 10088
rect 1694 10030 1707 10063
rect 1760 10030 1769 10063
rect 1694 10021 1769 10030
rect 2186 10173 2218 10180
rect 2186 10153 2193 10173
rect 2214 10153 2218 10173
rect 2186 10088 2218 10153
rect 2398 10144 2429 10351
rect 2633 10343 2665 10344
rect 3888 10343 3924 10354
rect 2630 10338 2665 10343
rect 2630 10318 2637 10338
rect 2657 10318 2665 10338
rect 2630 10310 2665 10318
rect 2398 10114 2404 10144
rect 2425 10114 2429 10144
rect 2398 10106 2429 10114
rect 2556 10088 2596 10089
rect 2186 10086 2598 10088
rect 2186 10060 2566 10086
rect 2592 10060 2598 10086
rect 2186 10052 2598 10060
rect 2186 10024 2218 10052
rect 2631 10032 2665 10310
rect 1694 10016 1752 10021
rect 1561 10004 1617 10011
rect 2186 10004 2191 10024
rect 2212 10004 2218 10024
rect 1561 10003 1596 10004
rect 2186 9997 2218 10004
rect 2609 10027 2665 10032
rect 2609 10007 2616 10027
rect 2636 10007 2665 10027
rect 2609 10000 2665 10007
rect 2609 9999 2644 10000
rect 852 9948 963 9952
rect 2727 9948 3968 9949
rect 174 9930 3968 9948
rect 174 9910 860 9930
rect 879 9910 937 9930
rect 956 9926 3968 9930
rect 956 9910 1908 9926
rect 174 9906 1908 9910
rect 1927 9906 1985 9926
rect 2004 9906 3968 9926
rect 174 9892 3968 9906
rect 174 9269 281 9892
rect 1900 9889 2011 9892
rect 660 9843 724 9847
rect 656 9837 724 9843
rect 656 9804 673 9837
rect 713 9804 724 9837
rect 656 9792 724 9804
rect 1707 9806 1772 9828
rect 656 9790 713 9792
rect 660 9429 711 9790
rect 1707 9767 1724 9806
rect 1769 9767 1772 9806
rect 1348 9722 1383 9724
rect 1348 9713 1452 9722
rect 1348 9712 1399 9713
rect 1348 9692 1351 9712
rect 1376 9693 1399 9712
rect 1431 9693 1452 9713
rect 1376 9692 1452 9693
rect 1348 9685 1452 9692
rect 1348 9673 1383 9685
rect 760 9607 963 9620
rect 760 9574 784 9607
rect 820 9606 963 9607
rect 820 9603 931 9606
rect 820 9576 857 9603
rect 886 9579 931 9603
rect 960 9579 963 9606
rect 886 9576 963 9579
rect 820 9574 963 9576
rect 760 9561 963 9574
rect 760 9560 861 9561
rect 1138 9498 1170 9505
rect 1138 9478 1145 9498
rect 1166 9478 1170 9498
rect 649 9420 714 9429
rect 649 9383 659 9420
rect 699 9386 714 9420
rect 1138 9413 1170 9478
rect 1350 9469 1381 9673
rect 1585 9668 1617 9669
rect 1582 9663 1617 9668
rect 1582 9643 1589 9663
rect 1609 9643 1617 9663
rect 1582 9635 1617 9643
rect 1350 9439 1356 9469
rect 1377 9439 1381 9469
rect 1350 9431 1381 9439
rect 1508 9413 1548 9414
rect 1138 9411 1550 9413
rect 699 9383 716 9386
rect 649 9364 716 9383
rect 649 9343 663 9364
rect 699 9343 716 9364
rect 649 9336 716 9343
rect 1138 9385 1518 9411
rect 1544 9385 1550 9411
rect 1138 9377 1550 9385
rect 1138 9349 1170 9377
rect 1583 9357 1617 9635
rect 1707 9467 1772 9767
rect 3886 9761 3991 9770
rect 3886 9756 3940 9761
rect 3886 9735 3899 9756
rect 3919 9740 3940 9756
rect 3960 9740 3991 9761
rect 3919 9735 3991 9740
rect 3886 9704 3991 9735
rect 3889 9687 3924 9704
rect 3888 9669 3924 9687
rect 3298 9604 3501 9617
rect 3298 9571 3322 9604
rect 3358 9603 3501 9604
rect 3358 9600 3469 9603
rect 3358 9573 3395 9600
rect 3424 9576 3469 9600
rect 3498 9576 3501 9603
rect 3424 9573 3501 9576
rect 3358 9571 3501 9573
rect 3298 9558 3501 9571
rect 3298 9557 3399 9558
rect 3676 9495 3708 9502
rect 3676 9475 3683 9495
rect 3704 9475 3708 9495
rect 1138 9329 1143 9349
rect 1164 9329 1170 9349
rect 1138 9322 1170 9329
rect 1561 9352 1617 9357
rect 1561 9332 1568 9352
rect 1588 9332 1617 9352
rect 1561 9325 1617 9332
rect 1697 9456 1777 9467
rect 1697 9430 1714 9456
rect 1754 9430 1777 9456
rect 1697 9403 1777 9430
rect 1697 9377 1718 9403
rect 1758 9377 1777 9403
rect 1697 9358 1777 9377
rect 1697 9332 1721 9358
rect 1761 9332 1777 9358
rect 1561 9324 1596 9325
rect 1697 9320 1777 9332
rect 3676 9410 3708 9475
rect 3888 9466 3919 9669
rect 4123 9665 4155 9666
rect 4120 9660 4155 9665
rect 4120 9640 4127 9660
rect 4147 9640 4155 9660
rect 4120 9632 4155 9640
rect 3888 9436 3894 9466
rect 3915 9436 3919 9466
rect 3888 9428 3919 9436
rect 4046 9410 4086 9411
rect 3676 9408 4088 9410
rect 3676 9382 4056 9408
rect 4082 9382 4088 9408
rect 3676 9374 4088 9382
rect 3676 9346 3708 9374
rect 4121 9354 4155 9632
rect 3676 9326 3681 9346
rect 3702 9326 3708 9346
rect 3676 9319 3708 9326
rect 4099 9349 4155 9354
rect 4099 9329 4106 9349
rect 4126 9329 4155 9349
rect 4099 9322 4155 9329
rect 4099 9321 4134 9322
rect 852 9269 963 9273
rect 2607 9269 2814 9270
rect 3390 9269 3501 9270
rect 172 9251 4192 9269
rect 172 9231 860 9251
rect 879 9231 937 9251
rect 956 9248 4192 9251
rect 956 9231 3398 9248
rect 172 9228 3398 9231
rect 3417 9228 3475 9248
rect 3494 9228 4192 9248
rect 172 9213 4192 9228
rect 174 9025 281 9213
rect 2769 9211 4192 9213
rect 642 9174 763 9184
rect 642 9172 711 9174
rect 642 9131 655 9172
rect 692 9133 711 9172
rect 748 9133 763 9174
rect 692 9131 763 9133
rect 642 9113 763 9131
rect 174 9021 282 9025
rect 648 9021 725 9113
rect 1698 9109 1774 9125
rect 1698 9086 1713 9109
rect 175 8428 282 9021
rect 650 8970 725 9021
rect 1691 9072 1713 9086
rect 1757 9072 1774 9109
rect 1691 9052 1774 9072
rect 1691 8986 1708 9052
rect 1762 8986 1774 9052
rect 650 8927 726 8970
rect 654 8616 726 8927
rect 1691 8962 1774 8986
rect 1691 8942 1767 8962
rect 1691 8923 1770 8942
rect 1350 8907 1422 8908
rect 1349 8899 1448 8907
rect 1349 8896 1401 8899
rect 1349 8861 1357 8896
rect 1382 8861 1401 8896
rect 1426 8861 1448 8899
rect 1349 8849 1448 8861
rect 1350 8830 1418 8849
rect 1351 8827 1384 8830
rect 1586 8827 1618 8828
rect 761 8766 964 8779
rect 761 8733 785 8766
rect 821 8765 964 8766
rect 821 8762 932 8765
rect 821 8735 858 8762
rect 887 8738 932 8762
rect 961 8738 964 8765
rect 887 8735 964 8738
rect 821 8733 964 8735
rect 761 8720 964 8733
rect 761 8719 862 8720
rect 654 8574 663 8616
rect 712 8574 726 8616
rect 654 8553 726 8574
rect 654 8511 664 8553
rect 713 8511 726 8553
rect 654 8493 726 8511
rect 1139 8657 1171 8664
rect 1139 8637 1146 8657
rect 1167 8637 1171 8657
rect 1139 8572 1171 8637
rect 1351 8628 1382 8827
rect 1583 8822 1618 8827
rect 1583 8802 1590 8822
rect 1610 8802 1618 8822
rect 1583 8794 1618 8802
rect 1351 8598 1357 8628
rect 1378 8598 1382 8628
rect 1351 8590 1382 8598
rect 1509 8572 1549 8573
rect 1139 8570 1551 8572
rect 1139 8544 1519 8570
rect 1545 8544 1551 8570
rect 1139 8536 1551 8544
rect 1139 8508 1171 8536
rect 1584 8516 1618 8794
rect 1700 8607 1770 8923
rect 3688 8908 3719 8909
rect 3688 8900 3733 8908
rect 2768 8877 2932 8884
rect 3688 8877 3698 8900
rect 2394 8862 3698 8877
rect 3723 8862 3733 8900
rect 2394 8844 3733 8862
rect 2399 8831 2435 8844
rect 2768 8841 2932 8844
rect 1809 8762 2012 8775
rect 1809 8729 1833 8762
rect 1869 8761 2012 8762
rect 1869 8758 1980 8761
rect 1869 8731 1906 8758
rect 1935 8734 1980 8758
rect 2009 8734 2012 8761
rect 1935 8731 2012 8734
rect 1869 8729 2012 8731
rect 1809 8716 2012 8729
rect 1809 8715 1910 8716
rect 1139 8488 1144 8508
rect 1165 8488 1171 8508
rect 1139 8481 1171 8488
rect 1562 8511 1618 8516
rect 1562 8491 1569 8511
rect 1589 8491 1618 8511
rect 1695 8601 1770 8607
rect 1695 8568 1703 8601
rect 1756 8568 1770 8601
rect 1695 8543 1770 8568
rect 1695 8510 1708 8543
rect 1761 8510 1770 8543
rect 1695 8501 1770 8510
rect 2187 8653 2219 8660
rect 2187 8633 2194 8653
rect 2215 8633 2219 8653
rect 2187 8568 2219 8633
rect 2399 8624 2430 8831
rect 2634 8823 2666 8824
rect 2631 8818 2666 8823
rect 2631 8798 2638 8818
rect 2658 8798 2666 8818
rect 2631 8790 2666 8798
rect 2399 8594 2405 8624
rect 2426 8594 2430 8624
rect 2399 8586 2430 8594
rect 2557 8568 2597 8569
rect 2187 8566 2599 8568
rect 2187 8540 2567 8566
rect 2593 8540 2599 8566
rect 2187 8532 2599 8540
rect 2187 8504 2219 8532
rect 2632 8512 2666 8790
rect 1695 8496 1753 8501
rect 1562 8484 1618 8491
rect 2187 8484 2192 8504
rect 2213 8484 2219 8504
rect 1562 8483 1597 8484
rect 2187 8477 2219 8484
rect 2610 8507 2666 8512
rect 2610 8487 2617 8507
rect 2637 8487 2666 8507
rect 2610 8480 2666 8487
rect 2610 8479 2645 8480
rect 853 8428 964 8432
rect 2636 8428 3936 8429
rect 175 8410 3936 8428
rect 175 8390 861 8410
rect 880 8390 938 8410
rect 957 8406 3936 8410
rect 957 8390 1909 8406
rect 175 8386 1909 8390
rect 1928 8386 1986 8406
rect 2005 8386 3936 8406
rect 175 8372 3936 8386
rect 175 7749 282 8372
rect 1901 8369 2012 8372
rect 661 8323 725 8327
rect 657 8317 725 8323
rect 657 8284 674 8317
rect 714 8284 725 8317
rect 657 8272 725 8284
rect 1708 8286 1773 8308
rect 657 8270 714 8272
rect 661 7909 712 8270
rect 1708 8247 1725 8286
rect 1770 8247 1773 8286
rect 1349 8202 1384 8204
rect 1349 8193 1453 8202
rect 1349 8192 1400 8193
rect 1349 8172 1352 8192
rect 1377 8173 1400 8192
rect 1432 8173 1453 8193
rect 1377 8172 1453 8173
rect 1349 8165 1453 8172
rect 1349 8153 1384 8165
rect 761 8087 964 8100
rect 761 8054 785 8087
rect 821 8086 964 8087
rect 821 8083 932 8086
rect 821 8056 858 8083
rect 887 8059 932 8083
rect 961 8059 964 8086
rect 887 8056 964 8059
rect 821 8054 964 8056
rect 761 8041 964 8054
rect 761 8040 862 8041
rect 1139 7978 1171 7985
rect 1139 7958 1146 7978
rect 1167 7958 1171 7978
rect 650 7900 715 7909
rect 650 7863 660 7900
rect 700 7866 715 7900
rect 1139 7893 1171 7958
rect 1351 7949 1382 8153
rect 1586 8148 1618 8149
rect 1583 8143 1618 8148
rect 1583 8123 1590 8143
rect 1610 8123 1618 8143
rect 1583 8115 1618 8123
rect 1351 7919 1357 7949
rect 1378 7919 1382 7949
rect 1351 7911 1382 7919
rect 1509 7893 1549 7894
rect 1139 7891 1551 7893
rect 700 7863 717 7866
rect 650 7844 717 7863
rect 650 7823 664 7844
rect 700 7823 717 7844
rect 650 7816 717 7823
rect 1139 7865 1519 7891
rect 1545 7865 1551 7891
rect 1139 7857 1551 7865
rect 1139 7829 1171 7857
rect 1584 7837 1618 8115
rect 1708 7947 1773 8247
rect 3845 8208 3882 8229
rect 3845 8171 3856 8208
rect 3873 8184 3882 8208
rect 3873 8171 3883 8184
rect 3845 8161 3883 8171
rect 3846 8157 3883 8161
rect 3846 8151 3879 8157
rect 3256 8082 3459 8095
rect 3256 8049 3280 8082
rect 3316 8081 3459 8082
rect 3316 8078 3427 8081
rect 3316 8051 3353 8078
rect 3382 8054 3427 8078
rect 3456 8054 3459 8081
rect 3382 8051 3459 8054
rect 3316 8049 3459 8051
rect 3256 8036 3459 8049
rect 3256 8035 3357 8036
rect 3634 7973 3666 7980
rect 3634 7953 3641 7973
rect 3662 7953 3666 7973
rect 1139 7809 1144 7829
rect 1165 7809 1171 7829
rect 1139 7802 1171 7809
rect 1562 7832 1618 7837
rect 1562 7812 1569 7832
rect 1589 7812 1618 7832
rect 1562 7805 1618 7812
rect 1698 7936 1778 7947
rect 1698 7910 1715 7936
rect 1755 7910 1778 7936
rect 1698 7883 1778 7910
rect 1698 7857 1719 7883
rect 1759 7857 1778 7883
rect 3634 7888 3666 7953
rect 3846 7944 3877 8151
rect 4081 8143 4113 8144
rect 4078 8138 4113 8143
rect 4078 8118 4085 8138
rect 4105 8118 4113 8138
rect 4078 8110 4113 8118
rect 3846 7914 3852 7944
rect 3873 7914 3877 7944
rect 3846 7906 3877 7914
rect 4004 7888 4044 7889
rect 3634 7886 4046 7888
rect 1698 7838 1778 7857
rect 1698 7812 1722 7838
rect 1762 7812 1778 7838
rect 2811 7876 3248 7882
rect 2811 7853 2829 7876
rect 2855 7869 3248 7876
rect 2855 7853 3209 7869
rect 2811 7846 3209 7853
rect 3235 7846 3248 7869
rect 2811 7833 3248 7846
rect 3634 7860 4014 7886
rect 4040 7860 4046 7886
rect 3634 7852 4046 7860
rect 1562 7804 1597 7805
rect 1698 7800 1778 7812
rect 3634 7824 3666 7852
rect 4079 7832 4113 8110
rect 3634 7804 3639 7824
rect 3660 7804 3666 7824
rect 3634 7797 3666 7804
rect 4057 7827 4113 7832
rect 4057 7807 4064 7827
rect 4084 7807 4113 7827
rect 4057 7800 4113 7807
rect 4057 7799 4092 7800
rect 853 7749 964 7753
rect 2595 7749 4145 7752
rect 173 7731 4145 7749
rect 173 7711 861 7731
rect 880 7711 938 7731
rect 957 7726 4145 7731
rect 957 7711 3356 7726
rect 173 7706 3356 7711
rect 3375 7706 3433 7726
rect 3452 7706 4145 7726
rect 173 7696 4145 7706
rect 173 7693 798 7696
rect 985 7693 4145 7696
rect 175 7465 282 7693
rect 2595 7692 4145 7693
rect 3348 7689 3459 7692
rect 643 7654 764 7664
rect 643 7652 712 7654
rect 643 7611 656 7652
rect 693 7613 712 7652
rect 749 7613 764 7654
rect 693 7611 764 7613
rect 643 7593 764 7611
rect 649 7491 728 7593
rect 1701 7553 1768 7572
rect 1701 7533 1721 7553
rect 175 7410 283 7465
rect 650 7410 728 7491
rect 1700 7487 1721 7533
rect 1751 7533 1768 7553
rect 1751 7503 1770 7533
rect 1751 7487 1771 7503
rect 1700 7471 1771 7487
rect 1350 7460 1422 7461
rect 1349 7452 1448 7460
rect 1349 7449 1401 7452
rect 1349 7414 1357 7449
rect 1382 7414 1401 7449
rect 1426 7414 1448 7452
rect 175 6981 282 7410
rect 654 7169 726 7410
rect 1349 7402 1448 7414
rect 1350 7383 1418 7402
rect 1351 7380 1384 7383
rect 1586 7380 1618 7381
rect 761 7319 964 7332
rect 761 7286 785 7319
rect 821 7318 964 7319
rect 821 7315 932 7318
rect 821 7288 858 7315
rect 887 7291 932 7315
rect 961 7291 964 7318
rect 887 7288 964 7291
rect 821 7286 964 7288
rect 761 7273 964 7286
rect 761 7272 862 7273
rect 654 7127 663 7169
rect 712 7127 726 7169
rect 654 7106 726 7127
rect 654 7064 664 7106
rect 713 7064 726 7106
rect 654 7046 726 7064
rect 1139 7210 1171 7217
rect 1139 7190 1146 7210
rect 1167 7190 1171 7210
rect 1139 7125 1171 7190
rect 1351 7181 1382 7380
rect 1583 7375 1618 7380
rect 1583 7355 1590 7375
rect 1610 7355 1618 7375
rect 1583 7347 1618 7355
rect 1351 7151 1357 7181
rect 1378 7151 1382 7181
rect 1351 7143 1382 7151
rect 1509 7125 1549 7126
rect 1139 7123 1551 7125
rect 1139 7097 1519 7123
rect 1545 7097 1551 7123
rect 1139 7089 1551 7097
rect 1139 7061 1171 7089
rect 1584 7069 1618 7347
rect 1700 7160 1770 7471
rect 2397 7462 3739 7467
rect 2397 7460 3696 7462
rect 2394 7434 3696 7460
rect 3724 7434 3739 7462
rect 2394 7426 3739 7434
rect 2394 7401 2433 7426
rect 2394 7384 2435 7401
rect 2394 7377 2433 7384
rect 1809 7315 2012 7328
rect 1809 7282 1833 7315
rect 1869 7314 2012 7315
rect 1869 7311 1980 7314
rect 1869 7284 1906 7311
rect 1935 7287 1980 7311
rect 2009 7287 2012 7314
rect 1935 7284 2012 7287
rect 1869 7282 2012 7284
rect 1809 7269 2012 7282
rect 1809 7268 1910 7269
rect 1139 7041 1144 7061
rect 1165 7041 1171 7061
rect 1139 7034 1171 7041
rect 1562 7064 1618 7069
rect 1562 7044 1569 7064
rect 1589 7044 1618 7064
rect 1695 7154 1770 7160
rect 1695 7121 1703 7154
rect 1756 7121 1770 7154
rect 1695 7096 1770 7121
rect 1695 7063 1708 7096
rect 1761 7063 1770 7096
rect 1695 7054 1770 7063
rect 2187 7206 2219 7213
rect 2187 7186 2194 7206
rect 2215 7186 2219 7206
rect 2187 7121 2219 7186
rect 2399 7177 2430 7377
rect 2634 7376 2666 7377
rect 2631 7371 2666 7376
rect 2631 7351 2638 7371
rect 2658 7351 2666 7371
rect 2631 7343 2666 7351
rect 2399 7147 2405 7177
rect 2426 7147 2430 7177
rect 2399 7139 2430 7147
rect 2557 7121 2597 7122
rect 2187 7119 2599 7121
rect 2187 7093 2567 7119
rect 2593 7093 2599 7119
rect 2187 7085 2599 7093
rect 2187 7057 2219 7085
rect 2632 7065 2666 7343
rect 1695 7049 1753 7054
rect 1562 7037 1618 7044
rect 2187 7037 2192 7057
rect 2213 7037 2219 7057
rect 1562 7036 1597 7037
rect 2187 7030 2219 7037
rect 2610 7060 2666 7065
rect 2610 7040 2617 7060
rect 2637 7040 2666 7060
rect 2610 7033 2666 7040
rect 2610 7032 2645 7033
rect 853 6981 964 6985
rect 2728 6981 3718 6982
rect 175 6963 3718 6981
rect 175 6943 861 6963
rect 880 6943 938 6963
rect 957 6959 3718 6963
rect 957 6943 1909 6959
rect 175 6939 1909 6943
rect 1928 6939 1986 6959
rect 2005 6939 3718 6959
rect 175 6925 3718 6939
rect 175 6302 282 6925
rect 1901 6922 2012 6925
rect 661 6876 725 6880
rect 657 6870 725 6876
rect 657 6837 674 6870
rect 714 6837 725 6870
rect 657 6825 725 6837
rect 1708 6839 1773 6861
rect 657 6823 714 6825
rect 661 6462 712 6823
rect 1708 6800 1725 6839
rect 1770 6800 1773 6839
rect 1349 6755 1384 6757
rect 1349 6746 1453 6755
rect 1349 6745 1400 6746
rect 1349 6725 1352 6745
rect 1377 6726 1400 6745
rect 1432 6726 1453 6746
rect 1377 6725 1453 6726
rect 1349 6718 1453 6725
rect 1349 6706 1384 6718
rect 761 6640 964 6653
rect 761 6607 785 6640
rect 821 6639 964 6640
rect 821 6636 932 6639
rect 821 6609 858 6636
rect 887 6612 932 6636
rect 961 6612 964 6639
rect 887 6609 964 6612
rect 821 6607 964 6609
rect 761 6594 964 6607
rect 761 6593 862 6594
rect 1139 6531 1171 6538
rect 1139 6511 1146 6531
rect 1167 6511 1171 6531
rect 650 6453 715 6462
rect 650 6416 660 6453
rect 700 6419 715 6453
rect 1139 6446 1171 6511
rect 1351 6502 1382 6706
rect 1586 6701 1618 6702
rect 1583 6696 1618 6701
rect 1583 6676 1590 6696
rect 1610 6676 1618 6696
rect 1583 6668 1618 6676
rect 1351 6472 1357 6502
rect 1378 6472 1382 6502
rect 1351 6464 1382 6472
rect 1509 6446 1549 6447
rect 1139 6444 1551 6446
rect 700 6416 717 6419
rect 650 6397 717 6416
rect 650 6376 664 6397
rect 700 6376 717 6397
rect 650 6369 717 6376
rect 1139 6418 1519 6444
rect 1545 6418 1551 6444
rect 1139 6410 1551 6418
rect 1139 6382 1171 6410
rect 1584 6390 1618 6668
rect 1708 6500 1773 6800
rect 1139 6362 1144 6382
rect 1165 6362 1171 6382
rect 1139 6355 1171 6362
rect 1562 6385 1618 6390
rect 1562 6365 1569 6385
rect 1589 6365 1618 6385
rect 1562 6358 1618 6365
rect 1698 6489 1778 6500
rect 1698 6463 1715 6489
rect 1755 6463 1778 6489
rect 1698 6436 1778 6463
rect 4250 6439 4299 12008
rect 4364 6631 4567 6644
rect 4364 6598 4388 6631
rect 4424 6630 4567 6631
rect 4424 6627 4535 6630
rect 4424 6600 4461 6627
rect 4490 6603 4535 6627
rect 4564 6603 4567 6630
rect 4490 6600 4567 6603
rect 4424 6598 4567 6600
rect 4364 6585 4567 6598
rect 4364 6584 4465 6585
rect 4742 6522 4774 6529
rect 4742 6502 4749 6522
rect 4770 6502 4774 6522
rect 1698 6410 1719 6436
rect 1759 6410 1778 6436
rect 1698 6391 1778 6410
rect 4249 6429 4360 6439
rect 4249 6428 4314 6429
rect 4249 6404 4257 6428
rect 4281 6405 4314 6428
rect 4338 6405 4360 6429
rect 4281 6404 4360 6405
rect 4249 6397 4360 6404
rect 4742 6437 4774 6502
rect 4954 6493 4985 6719
rect 5189 6692 5221 6693
rect 5186 6687 5221 6692
rect 5186 6667 5193 6687
rect 5213 6667 5221 6687
rect 5186 6659 5221 6667
rect 4954 6463 4960 6493
rect 4981 6463 4985 6493
rect 4954 6455 4985 6463
rect 5112 6437 5152 6438
rect 4742 6435 5154 6437
rect 4742 6409 5122 6435
rect 5148 6409 5154 6435
rect 4742 6401 5154 6409
rect 1698 6365 1722 6391
rect 1762 6365 1778 6391
rect 1562 6357 1597 6358
rect 1698 6353 1778 6365
rect 4742 6373 4774 6401
rect 5187 6381 5221 6659
rect 4742 6353 4747 6373
rect 4768 6353 4774 6373
rect 4742 6346 4774 6353
rect 5165 6376 5221 6381
rect 5165 6356 5172 6376
rect 5192 6356 5221 6376
rect 5165 6349 5221 6356
rect 5165 6348 5200 6349
rect 853 6302 964 6306
rect 2608 6302 2815 6303
rect 173 6297 4248 6302
rect 173 6284 4567 6297
rect 173 6264 861 6284
rect 880 6264 938 6284
rect 957 6275 4567 6284
rect 957 6264 4464 6275
rect 173 6255 4464 6264
rect 4483 6255 4541 6275
rect 4560 6255 4567 6275
rect 173 6246 4567 6255
rect 175 6073 282 6246
rect 2770 6244 4567 6246
rect 4456 6238 4567 6244
rect 643 6207 764 6217
rect 643 6205 712 6207
rect 643 6164 656 6205
rect 693 6166 712 6205
rect 749 6166 764 6207
rect 693 6164 764 6166
rect 643 6146 764 6164
rect 4791 6196 4843 6227
rect 4791 6162 4800 6196
rect 4829 6162 4843 6196
rect 166 6046 282 6073
rect 649 6054 714 6146
rect 4791 6136 4843 6162
rect 166 5907 277 6046
rect 647 6008 714 6054
rect 1699 6092 1771 6114
rect 1699 6044 1713 6092
rect 1759 6087 1771 6092
rect 4791 6102 4799 6136
rect 4828 6102 4843 6136
rect 1759 6044 1776 6087
rect 647 5907 712 6008
rect 166 5847 279 5907
rect 647 5869 723 5907
rect 172 5387 279 5847
rect 651 5575 723 5869
rect 1347 5866 1419 5867
rect 1346 5858 1445 5866
rect 1699 5861 1776 6044
rect 2987 6045 3071 6056
rect 2987 6017 3015 6045
rect 3059 6017 3071 6045
rect 2801 5966 2875 5994
rect 2801 5918 2824 5966
rect 2861 5918 2875 5966
rect 2987 5988 3071 6017
rect 2987 5960 3012 5988
rect 3056 5960 3071 5988
rect 2987 5927 3071 5960
rect 2801 5909 2875 5918
rect 2397 5867 2469 5868
rect 1346 5855 1398 5858
rect 1346 5820 1354 5855
rect 1379 5820 1398 5855
rect 1423 5820 1445 5858
rect 1346 5808 1445 5820
rect 1697 5832 1776 5861
rect 2396 5859 2485 5867
rect 2396 5856 2448 5859
rect 1347 5789 1415 5808
rect 1348 5786 1381 5789
rect 1583 5786 1615 5787
rect 758 5725 961 5738
rect 758 5692 782 5725
rect 818 5724 961 5725
rect 818 5721 929 5724
rect 818 5694 855 5721
rect 884 5697 929 5721
rect 958 5697 961 5724
rect 884 5694 961 5697
rect 818 5692 961 5694
rect 758 5679 961 5692
rect 758 5678 859 5679
rect 651 5533 660 5575
rect 709 5533 723 5575
rect 651 5512 723 5533
rect 651 5470 661 5512
rect 710 5470 723 5512
rect 651 5452 723 5470
rect 1136 5616 1168 5623
rect 1136 5596 1143 5616
rect 1164 5596 1168 5616
rect 1136 5531 1168 5596
rect 1348 5587 1379 5786
rect 1580 5781 1615 5786
rect 1580 5761 1587 5781
rect 1607 5761 1615 5781
rect 1580 5753 1615 5761
rect 1348 5557 1354 5587
rect 1375 5557 1379 5587
rect 1348 5549 1379 5557
rect 1506 5531 1546 5532
rect 1136 5529 1548 5531
rect 1136 5503 1516 5529
rect 1542 5503 1548 5529
rect 1136 5495 1548 5503
rect 1136 5467 1168 5495
rect 1581 5475 1615 5753
rect 1697 5566 1767 5832
rect 2396 5821 2404 5856
rect 2429 5821 2448 5856
rect 2473 5821 2485 5859
rect 2396 5809 2485 5821
rect 2396 5808 2465 5809
rect 2396 5790 2432 5808
rect 1806 5721 2009 5734
rect 1806 5688 1830 5721
rect 1866 5720 2009 5721
rect 1866 5717 1977 5720
rect 1866 5690 1903 5717
rect 1932 5693 1977 5717
rect 2006 5693 2009 5720
rect 1932 5690 2009 5693
rect 1866 5688 2009 5690
rect 1806 5675 2009 5688
rect 1806 5674 1907 5675
rect 1136 5447 1141 5467
rect 1162 5447 1168 5467
rect 1136 5440 1168 5447
rect 1559 5470 1615 5475
rect 1559 5450 1566 5470
rect 1586 5450 1615 5470
rect 1692 5560 1767 5566
rect 1692 5527 1700 5560
rect 1753 5527 1767 5560
rect 1692 5502 1767 5527
rect 1692 5469 1705 5502
rect 1758 5469 1767 5502
rect 1692 5460 1767 5469
rect 2184 5612 2216 5619
rect 2184 5592 2191 5612
rect 2212 5592 2216 5612
rect 2184 5527 2216 5592
rect 2396 5583 2427 5790
rect 2631 5782 2663 5783
rect 2628 5777 2663 5782
rect 2628 5757 2635 5777
rect 2655 5757 2663 5777
rect 2628 5749 2663 5757
rect 2396 5553 2402 5583
rect 2423 5553 2427 5583
rect 2396 5545 2427 5553
rect 2554 5527 2594 5528
rect 2184 5525 2596 5527
rect 2184 5499 2564 5525
rect 2590 5499 2596 5525
rect 2184 5491 2596 5499
rect 2184 5463 2216 5491
rect 2629 5471 2663 5749
rect 2812 5564 2874 5909
rect 2981 5882 3071 5927
rect 2981 5567 3063 5882
rect 2812 5545 2876 5564
rect 2812 5506 2825 5545
rect 2859 5506 2876 5545
rect 2812 5487 2876 5506
rect 2981 5526 3002 5567
rect 3038 5526 3063 5567
rect 2981 5497 3063 5526
rect 1692 5455 1750 5460
rect 1559 5443 1615 5450
rect 2184 5443 2189 5463
rect 2210 5443 2216 5463
rect 1559 5442 1594 5443
rect 2184 5436 2216 5443
rect 2607 5466 2663 5471
rect 2607 5446 2614 5466
rect 2634 5446 2663 5466
rect 2607 5439 2663 5446
rect 2607 5438 2642 5439
rect 850 5387 961 5391
rect 2633 5387 4203 5388
rect 172 5369 4203 5387
rect 172 5349 858 5369
rect 877 5349 935 5369
rect 954 5365 4203 5369
rect 954 5349 1906 5365
rect 172 5345 1906 5349
rect 1925 5345 1983 5365
rect 2002 5345 4203 5365
rect 172 5331 4203 5345
rect 172 4708 279 5331
rect 1898 5328 2009 5331
rect 658 5282 722 5286
rect 654 5276 722 5282
rect 654 5243 671 5276
rect 711 5243 722 5276
rect 654 5231 722 5243
rect 1705 5245 1770 5267
rect 654 5229 711 5231
rect 658 4868 709 5229
rect 1705 5206 1722 5245
rect 1767 5206 1770 5245
rect 1346 5161 1381 5163
rect 1346 5152 1450 5161
rect 1346 5151 1397 5152
rect 1346 5131 1349 5151
rect 1374 5132 1397 5151
rect 1429 5132 1450 5152
rect 1374 5131 1450 5132
rect 1346 5124 1450 5131
rect 1346 5112 1381 5124
rect 758 5046 961 5059
rect 758 5013 782 5046
rect 818 5045 961 5046
rect 818 5042 929 5045
rect 818 5015 855 5042
rect 884 5018 929 5042
rect 958 5018 961 5045
rect 884 5015 961 5018
rect 818 5013 961 5015
rect 758 5000 961 5013
rect 758 4999 859 5000
rect 1136 4937 1168 4944
rect 1136 4917 1143 4937
rect 1164 4917 1168 4937
rect 647 4859 712 4868
rect 647 4822 657 4859
rect 697 4825 712 4859
rect 1136 4852 1168 4917
rect 1348 4908 1379 5112
rect 1583 5107 1615 5108
rect 1580 5102 1615 5107
rect 1580 5082 1587 5102
rect 1607 5082 1615 5102
rect 1580 5074 1615 5082
rect 1348 4878 1354 4908
rect 1375 4878 1379 4908
rect 1348 4870 1379 4878
rect 1506 4852 1546 4853
rect 1136 4850 1548 4852
rect 697 4822 714 4825
rect 647 4803 714 4822
rect 647 4782 661 4803
rect 697 4782 714 4803
rect 647 4775 714 4782
rect 1136 4824 1516 4850
rect 1542 4824 1548 4850
rect 1136 4816 1548 4824
rect 1136 4788 1168 4816
rect 1581 4796 1615 5074
rect 1705 4906 1770 5206
rect 2976 5230 3069 5245
rect 2976 5186 2991 5230
rect 3051 5186 3069 5230
rect 1136 4768 1141 4788
rect 1162 4768 1168 4788
rect 1136 4761 1168 4768
rect 1559 4791 1615 4796
rect 1559 4771 1566 4791
rect 1586 4771 1615 4791
rect 1559 4764 1615 4771
rect 1695 4895 1775 4906
rect 1695 4869 1712 4895
rect 1752 4869 1775 4895
rect 1695 4842 1775 4869
rect 1695 4816 1716 4842
rect 1756 4816 1775 4842
rect 1695 4797 1775 4816
rect 1695 4771 1719 4797
rect 1759 4771 1775 4797
rect 1559 4763 1594 4764
rect 1695 4759 1775 4771
rect 2976 4813 3069 5186
rect 3253 5041 3456 5054
rect 3253 5008 3277 5041
rect 3313 5040 3456 5041
rect 3313 5037 3424 5040
rect 3313 5010 3350 5037
rect 3379 5013 3424 5037
rect 3453 5013 3456 5040
rect 3379 5010 3456 5013
rect 3313 5008 3456 5010
rect 3253 4995 3456 5008
rect 3253 4994 3354 4995
rect 2976 4772 2991 4813
rect 3045 4772 3069 4813
rect 2976 4765 3069 4772
rect 3631 4932 3663 4939
rect 3631 4912 3638 4932
rect 3659 4912 3663 4932
rect 3631 4847 3663 4912
rect 3843 4903 3874 5104
rect 4078 5102 4110 5103
rect 4075 5097 4110 5102
rect 4075 5077 4082 5097
rect 4102 5077 4110 5097
rect 4075 5069 4110 5077
rect 3843 4873 3849 4903
rect 3870 4873 3874 4903
rect 3843 4865 3874 4873
rect 4001 4847 4041 4848
rect 3631 4845 4043 4847
rect 3631 4819 4011 4845
rect 4037 4819 4043 4845
rect 3631 4811 4043 4819
rect 3631 4783 3663 4811
rect 4076 4791 4110 5069
rect 3631 4763 3636 4783
rect 3657 4763 3663 4783
rect 3631 4756 3663 4763
rect 4054 4786 4110 4791
rect 4054 4766 4061 4786
rect 4081 4766 4110 4786
rect 4054 4759 4110 4766
rect 4054 4758 4089 4759
rect 850 4708 961 4712
rect 2592 4708 4236 4711
rect 170 4690 4236 4708
rect 170 4670 858 4690
rect 877 4670 935 4690
rect 954 4685 4236 4690
rect 954 4670 3353 4685
rect 170 4665 3353 4670
rect 3372 4665 3430 4685
rect 3449 4665 4236 4685
rect 170 4655 4236 4665
rect 170 4652 795 4655
rect 982 4652 4236 4655
rect 172 4424 279 4652
rect 2592 4651 4236 4652
rect 3345 4648 3456 4651
rect 640 4613 761 4623
rect 640 4611 709 4613
rect 640 4570 653 4611
rect 690 4572 709 4611
rect 746 4572 761 4613
rect 690 4570 761 4572
rect 640 4552 761 4570
rect 3845 4593 3931 4597
rect 3845 4575 3860 4593
rect 3912 4575 3931 4593
rect 3845 4566 3931 4575
rect 646 4450 725 4552
rect 1698 4512 1765 4531
rect 1698 4492 1718 4512
rect 172 4369 280 4424
rect 647 4369 725 4450
rect 1697 4446 1718 4492
rect 1748 4492 1765 4512
rect 1748 4462 1767 4492
rect 1748 4446 1768 4462
rect 1697 4430 1768 4446
rect 1347 4419 1419 4420
rect 1346 4411 1445 4419
rect 1346 4408 1398 4411
rect 1346 4373 1354 4408
rect 1379 4373 1398 4408
rect 1423 4373 1445 4411
rect 172 3940 279 4369
rect 651 4128 723 4369
rect 1346 4361 1445 4373
rect 1347 4342 1415 4361
rect 1348 4339 1381 4342
rect 1583 4339 1615 4340
rect 758 4278 961 4291
rect 758 4245 782 4278
rect 818 4277 961 4278
rect 818 4274 929 4277
rect 818 4247 855 4274
rect 884 4250 929 4274
rect 958 4250 961 4277
rect 884 4247 961 4250
rect 818 4245 961 4247
rect 758 4232 961 4245
rect 758 4231 859 4232
rect 651 4086 660 4128
rect 709 4086 723 4128
rect 651 4065 723 4086
rect 651 4023 661 4065
rect 710 4023 723 4065
rect 651 4005 723 4023
rect 1136 4169 1168 4176
rect 1136 4149 1143 4169
rect 1164 4149 1168 4169
rect 1136 4084 1168 4149
rect 1348 4140 1379 4339
rect 1580 4334 1615 4339
rect 1580 4314 1587 4334
rect 1607 4314 1615 4334
rect 1580 4306 1615 4314
rect 1348 4110 1354 4140
rect 1375 4110 1379 4140
rect 1348 4102 1379 4110
rect 1506 4084 1546 4085
rect 1136 4082 1548 4084
rect 1136 4056 1516 4082
rect 1542 4056 1548 4082
rect 1136 4048 1548 4056
rect 1136 4020 1168 4048
rect 1581 4028 1615 4306
rect 1697 4119 1767 4430
rect 3622 4420 3694 4421
rect 3621 4417 3710 4420
rect 2393 4415 3710 4417
rect 2390 4412 3710 4415
rect 2390 4409 3673 4412
rect 2390 4374 3629 4409
rect 3654 4374 3673 4409
rect 3698 4374 3710 4412
rect 2390 4364 3710 4374
rect 3886 4413 3922 4566
rect 3886 4390 3892 4413
rect 3916 4390 3922 4413
rect 3886 4369 3922 4390
rect 2390 4362 3675 4364
rect 2390 4352 2487 4362
rect 2396 4343 2432 4352
rect 3886 4346 3892 4369
rect 3916 4346 3922 4369
rect 1806 4274 2009 4287
rect 1806 4241 1830 4274
rect 1866 4273 2009 4274
rect 1866 4270 1977 4273
rect 1866 4243 1903 4270
rect 1932 4246 1977 4270
rect 2006 4246 2009 4273
rect 1932 4243 2009 4246
rect 1866 4241 2009 4243
rect 1806 4228 2009 4241
rect 1806 4227 1907 4228
rect 1136 4000 1141 4020
rect 1162 4000 1168 4020
rect 1136 3993 1168 4000
rect 1559 4023 1615 4028
rect 1559 4003 1566 4023
rect 1586 4003 1615 4023
rect 1692 4113 1767 4119
rect 1692 4080 1700 4113
rect 1753 4080 1767 4113
rect 1692 4055 1767 4080
rect 1692 4022 1705 4055
rect 1758 4022 1767 4055
rect 1692 4013 1767 4022
rect 2184 4165 2216 4172
rect 2184 4145 2191 4165
rect 2212 4145 2216 4165
rect 2184 4080 2216 4145
rect 2396 4136 2427 4343
rect 2631 4335 2663 4336
rect 3886 4335 3922 4346
rect 2628 4330 2663 4335
rect 2628 4310 2635 4330
rect 2655 4310 2663 4330
rect 2628 4302 2663 4310
rect 2396 4106 2402 4136
rect 2423 4106 2427 4136
rect 2396 4098 2427 4106
rect 2554 4080 2594 4081
rect 2184 4078 2596 4080
rect 2184 4052 2564 4078
rect 2590 4052 2596 4078
rect 2184 4044 2596 4052
rect 2184 4016 2216 4044
rect 2629 4024 2663 4302
rect 1692 4008 1750 4013
rect 1559 3996 1615 4003
rect 2184 3996 2189 4016
rect 2210 3996 2216 4016
rect 1559 3995 1594 3996
rect 2184 3989 2216 3996
rect 2607 4019 2663 4024
rect 2607 3999 2614 4019
rect 2634 3999 2663 4019
rect 2607 3992 2663 3999
rect 2607 3991 2642 3992
rect 850 3940 961 3944
rect 2725 3940 3884 3941
rect 172 3922 3884 3940
rect 172 3902 858 3922
rect 877 3902 935 3922
rect 954 3918 3884 3922
rect 954 3902 1906 3918
rect 172 3898 1906 3902
rect 1925 3898 1983 3918
rect 2002 3898 3884 3918
rect 172 3884 3884 3898
rect 172 3261 279 3884
rect 1898 3881 2009 3884
rect 658 3835 722 3839
rect 654 3829 722 3835
rect 654 3796 671 3829
rect 711 3796 722 3829
rect 654 3784 722 3796
rect 1705 3798 1770 3820
rect 654 3782 711 3784
rect 658 3421 709 3782
rect 1705 3759 1722 3798
rect 1767 3759 1770 3798
rect 4791 3796 4843 6102
rect 4246 3792 4843 3796
rect 1346 3714 1381 3716
rect 1346 3705 1450 3714
rect 1346 3704 1397 3705
rect 1346 3684 1349 3704
rect 1374 3685 1397 3704
rect 1429 3685 1450 3705
rect 1374 3684 1450 3685
rect 1346 3677 1450 3684
rect 1346 3665 1381 3677
rect 758 3599 961 3612
rect 758 3566 782 3599
rect 818 3598 961 3599
rect 818 3595 929 3598
rect 818 3568 855 3595
rect 884 3571 929 3595
rect 958 3571 961 3598
rect 884 3568 961 3571
rect 818 3566 961 3568
rect 758 3553 961 3566
rect 758 3552 859 3553
rect 1136 3490 1168 3497
rect 1136 3470 1143 3490
rect 1164 3470 1168 3490
rect 647 3412 712 3421
rect 647 3375 657 3412
rect 697 3378 712 3412
rect 1136 3405 1168 3470
rect 1348 3461 1379 3665
rect 1583 3660 1615 3661
rect 1580 3655 1615 3660
rect 1580 3635 1587 3655
rect 1607 3635 1615 3655
rect 1580 3627 1615 3635
rect 1348 3431 1354 3461
rect 1375 3431 1379 3461
rect 1348 3423 1379 3431
rect 1506 3405 1546 3406
rect 1136 3403 1548 3405
rect 697 3375 714 3378
rect 647 3356 714 3375
rect 647 3335 661 3356
rect 697 3335 714 3356
rect 647 3328 714 3335
rect 1136 3377 1516 3403
rect 1542 3377 1548 3403
rect 1136 3369 1548 3377
rect 1136 3341 1168 3369
rect 1581 3349 1615 3627
rect 1705 3459 1770 3759
rect 3883 3747 4843 3792
rect 3883 3743 4296 3747
rect 3883 3654 3917 3743
rect 4121 3657 4153 3658
rect 3296 3596 3499 3609
rect 3296 3563 3320 3596
rect 3356 3595 3499 3596
rect 3356 3592 3467 3595
rect 3356 3565 3393 3592
rect 3422 3568 3467 3592
rect 3496 3568 3499 3595
rect 3422 3565 3499 3568
rect 3356 3563 3499 3565
rect 3296 3550 3499 3563
rect 3296 3549 3397 3550
rect 3674 3487 3706 3494
rect 3674 3467 3681 3487
rect 3702 3467 3706 3487
rect 1136 3321 1141 3341
rect 1162 3321 1168 3341
rect 1136 3314 1168 3321
rect 1559 3344 1615 3349
rect 1559 3324 1566 3344
rect 1586 3324 1615 3344
rect 1559 3317 1615 3324
rect 1695 3448 1775 3459
rect 1695 3422 1712 3448
rect 1752 3422 1775 3448
rect 1695 3395 1775 3422
rect 1695 3369 1716 3395
rect 1756 3369 1775 3395
rect 1695 3350 1775 3369
rect 1695 3324 1719 3350
rect 1759 3324 1775 3350
rect 1559 3316 1594 3317
rect 1695 3312 1775 3324
rect 3674 3402 3706 3467
rect 3886 3458 3917 3654
rect 4118 3652 4153 3657
rect 4118 3632 4125 3652
rect 4145 3632 4153 3652
rect 4118 3624 4153 3632
rect 3886 3428 3892 3458
rect 3913 3428 3917 3458
rect 3886 3420 3917 3428
rect 4044 3402 4084 3403
rect 3674 3400 4086 3402
rect 3674 3374 4054 3400
rect 4080 3374 4086 3400
rect 3674 3366 4086 3374
rect 3674 3338 3706 3366
rect 4119 3346 4153 3624
rect 3674 3318 3679 3338
rect 3700 3318 3706 3338
rect 3674 3311 3706 3318
rect 4097 3341 4153 3346
rect 4097 3321 4104 3341
rect 4124 3321 4153 3341
rect 4097 3314 4153 3321
rect 4097 3313 4132 3314
rect 850 3261 961 3265
rect 2605 3261 2812 3262
rect 3388 3261 3499 3262
rect 170 3243 4236 3261
rect 170 3223 858 3243
rect 877 3223 935 3243
rect 954 3240 4236 3243
rect 954 3223 3396 3240
rect 170 3220 3396 3223
rect 3415 3220 3473 3240
rect 3492 3220 4236 3240
rect 170 3205 4236 3220
rect 172 3017 279 3205
rect 2767 3203 4236 3205
rect 640 3166 761 3176
rect 640 3164 709 3166
rect 640 3123 653 3164
rect 690 3125 709 3164
rect 746 3125 761 3166
rect 690 3123 761 3125
rect 640 3105 761 3123
rect 172 3013 280 3017
rect 646 3013 723 3105
rect 1696 3101 1772 3117
rect 1696 3078 1711 3101
rect 173 2420 280 3013
rect 648 2962 723 3013
rect 1689 3064 1711 3078
rect 1755 3064 1772 3101
rect 1689 3044 1772 3064
rect 1689 2978 1706 3044
rect 1760 2978 1772 3044
rect 648 2919 724 2962
rect 652 2608 724 2919
rect 1689 2954 1772 2978
rect 1689 2934 1765 2954
rect 1689 2915 1768 2934
rect 1348 2899 1420 2900
rect 1347 2891 1446 2899
rect 1347 2888 1399 2891
rect 1347 2853 1355 2888
rect 1380 2853 1399 2888
rect 1424 2853 1446 2891
rect 1347 2841 1446 2853
rect 1348 2822 1416 2841
rect 1349 2819 1382 2822
rect 1584 2819 1616 2820
rect 759 2758 962 2771
rect 759 2725 783 2758
rect 819 2757 962 2758
rect 819 2754 930 2757
rect 819 2727 856 2754
rect 885 2730 930 2754
rect 959 2730 962 2757
rect 885 2727 962 2730
rect 819 2725 962 2727
rect 759 2712 962 2725
rect 759 2711 860 2712
rect 652 2566 661 2608
rect 710 2566 724 2608
rect 652 2545 724 2566
rect 652 2503 662 2545
rect 711 2503 724 2545
rect 652 2485 724 2503
rect 1137 2649 1169 2656
rect 1137 2629 1144 2649
rect 1165 2629 1169 2649
rect 1137 2564 1169 2629
rect 1349 2620 1380 2819
rect 1581 2814 1616 2819
rect 1581 2794 1588 2814
rect 1608 2794 1616 2814
rect 1581 2786 1616 2794
rect 1349 2590 1355 2620
rect 1376 2590 1380 2620
rect 1349 2582 1380 2590
rect 1507 2564 1547 2565
rect 1137 2562 1549 2564
rect 1137 2536 1517 2562
rect 1543 2536 1549 2562
rect 1137 2528 1549 2536
rect 1137 2500 1169 2528
rect 1582 2508 1616 2786
rect 1698 2599 1768 2915
rect 3686 2900 3717 2901
rect 3686 2892 3731 2900
rect 2766 2869 2930 2876
rect 3686 2869 3696 2892
rect 2392 2854 3696 2869
rect 3721 2854 3731 2892
rect 2392 2836 3731 2854
rect 2397 2823 2433 2836
rect 2766 2833 2930 2836
rect 1807 2754 2010 2767
rect 1807 2721 1831 2754
rect 1867 2753 2010 2754
rect 1867 2750 1978 2753
rect 1867 2723 1904 2750
rect 1933 2726 1978 2750
rect 2007 2726 2010 2753
rect 1933 2723 2010 2726
rect 1867 2721 2010 2723
rect 1807 2708 2010 2721
rect 1807 2707 1908 2708
rect 1137 2480 1142 2500
rect 1163 2480 1169 2500
rect 1137 2473 1169 2480
rect 1560 2503 1616 2508
rect 1560 2483 1567 2503
rect 1587 2483 1616 2503
rect 1693 2593 1768 2599
rect 1693 2560 1701 2593
rect 1754 2560 1768 2593
rect 1693 2535 1768 2560
rect 1693 2502 1706 2535
rect 1759 2502 1768 2535
rect 1693 2493 1768 2502
rect 2185 2645 2217 2652
rect 2185 2625 2192 2645
rect 2213 2625 2217 2645
rect 2185 2560 2217 2625
rect 2397 2616 2428 2823
rect 2632 2815 2664 2816
rect 2629 2810 2664 2815
rect 2629 2790 2636 2810
rect 2656 2790 2664 2810
rect 2629 2782 2664 2790
rect 2397 2586 2403 2616
rect 2424 2586 2428 2616
rect 2397 2578 2428 2586
rect 2555 2560 2595 2561
rect 2185 2558 2597 2560
rect 2185 2532 2565 2558
rect 2591 2532 2597 2558
rect 2185 2524 2597 2532
rect 2185 2496 2217 2524
rect 2630 2504 2664 2782
rect 1693 2488 1751 2493
rect 1560 2476 1616 2483
rect 2185 2476 2190 2496
rect 2211 2476 2217 2496
rect 1560 2475 1595 2476
rect 2185 2469 2217 2476
rect 2608 2499 2664 2504
rect 2608 2479 2615 2499
rect 2635 2479 2664 2499
rect 2608 2472 2664 2479
rect 2608 2471 2643 2472
rect 851 2420 962 2424
rect 2634 2420 4204 2421
rect 173 2402 4204 2420
rect 173 2382 859 2402
rect 878 2382 936 2402
rect 955 2398 4204 2402
rect 955 2382 1907 2398
rect 173 2378 1907 2382
rect 1926 2378 1984 2398
rect 2003 2378 4204 2398
rect 173 2364 4204 2378
rect 173 1741 280 2364
rect 1899 2361 2010 2364
rect 659 2315 723 2319
rect 655 2309 723 2315
rect 655 2276 672 2309
rect 712 2276 723 2309
rect 655 2264 723 2276
rect 1706 2278 1771 2300
rect 655 2262 712 2264
rect 659 1901 710 2262
rect 1706 2239 1723 2278
rect 1768 2239 1771 2278
rect 1347 2194 1382 2196
rect 1347 2185 1451 2194
rect 1347 2184 1398 2185
rect 1347 2164 1350 2184
rect 1375 2165 1398 2184
rect 1430 2165 1451 2185
rect 1375 2164 1451 2165
rect 1347 2157 1451 2164
rect 1347 2145 1382 2157
rect 759 2079 962 2092
rect 759 2046 783 2079
rect 819 2078 962 2079
rect 819 2075 930 2078
rect 819 2048 856 2075
rect 885 2051 930 2075
rect 959 2051 962 2078
rect 885 2048 962 2051
rect 819 2046 962 2048
rect 759 2033 962 2046
rect 759 2032 860 2033
rect 1137 1970 1169 1977
rect 1137 1950 1144 1970
rect 1165 1950 1169 1970
rect 648 1892 713 1901
rect 648 1855 658 1892
rect 698 1858 713 1892
rect 1137 1885 1169 1950
rect 1349 1941 1380 2145
rect 1584 2140 1616 2141
rect 1581 2135 1616 2140
rect 1581 2115 1588 2135
rect 1608 2115 1616 2135
rect 1581 2107 1616 2115
rect 1349 1911 1355 1941
rect 1376 1911 1380 1941
rect 1349 1903 1380 1911
rect 1507 1885 1547 1886
rect 1137 1883 1549 1885
rect 698 1855 715 1858
rect 648 1836 715 1855
rect 648 1815 662 1836
rect 698 1815 715 1836
rect 648 1808 715 1815
rect 1137 1857 1517 1883
rect 1543 1857 1549 1883
rect 1137 1849 1549 1857
rect 1137 1821 1169 1849
rect 1582 1829 1616 2107
rect 1706 1939 1771 2239
rect 3843 2200 3880 2221
rect 3843 2163 3854 2200
rect 3871 2176 3880 2200
rect 3871 2163 3881 2176
rect 3843 2153 3881 2163
rect 3844 2149 3881 2153
rect 3844 2143 3877 2149
rect 3254 2074 3457 2087
rect 3254 2041 3278 2074
rect 3314 2073 3457 2074
rect 3314 2070 3425 2073
rect 3314 2043 3351 2070
rect 3380 2046 3425 2070
rect 3454 2046 3457 2073
rect 3380 2043 3457 2046
rect 3314 2041 3457 2043
rect 3254 2028 3457 2041
rect 3254 2027 3355 2028
rect 3632 1965 3664 1972
rect 3632 1945 3639 1965
rect 3660 1945 3664 1965
rect 1137 1801 1142 1821
rect 1163 1801 1169 1821
rect 1137 1794 1169 1801
rect 1560 1824 1616 1829
rect 1560 1804 1567 1824
rect 1587 1804 1616 1824
rect 1560 1797 1616 1804
rect 1696 1928 1776 1939
rect 1696 1902 1713 1928
rect 1753 1902 1776 1928
rect 1696 1875 1776 1902
rect 1696 1849 1717 1875
rect 1757 1849 1776 1875
rect 3632 1880 3664 1945
rect 3844 1936 3875 2143
rect 4079 2135 4111 2136
rect 4076 2130 4111 2135
rect 4076 2110 4083 2130
rect 4103 2110 4111 2130
rect 4076 2102 4111 2110
rect 3844 1906 3850 1936
rect 3871 1906 3875 1936
rect 3844 1898 3875 1906
rect 4002 1880 4042 1881
rect 3632 1878 4044 1880
rect 1696 1830 1776 1849
rect 1696 1804 1720 1830
rect 1760 1804 1776 1830
rect 2809 1868 3246 1874
rect 2809 1845 2827 1868
rect 2853 1861 3246 1868
rect 2853 1845 3207 1861
rect 2809 1838 3207 1845
rect 3233 1838 3246 1861
rect 2809 1825 3246 1838
rect 3632 1852 4012 1878
rect 4038 1852 4044 1878
rect 3632 1844 4044 1852
rect 1560 1796 1595 1797
rect 1696 1792 1776 1804
rect 3632 1816 3664 1844
rect 4077 1824 4111 2102
rect 3632 1796 3637 1816
rect 3658 1796 3664 1816
rect 3632 1789 3664 1796
rect 4055 1819 4111 1824
rect 4055 1799 4062 1819
rect 4082 1799 4111 1819
rect 4055 1792 4111 1799
rect 4055 1791 4090 1792
rect 851 1741 962 1745
rect 2593 1741 4246 1744
rect 171 1723 4246 1741
rect 171 1703 859 1723
rect 878 1703 936 1723
rect 955 1718 4246 1723
rect 955 1703 3354 1718
rect 171 1698 3354 1703
rect 3373 1698 3431 1718
rect 3450 1698 4246 1718
rect 171 1688 4246 1698
rect 171 1685 796 1688
rect 983 1685 4246 1688
rect 173 1457 280 1685
rect 2593 1684 4246 1685
rect 3346 1681 3457 1684
rect 641 1646 762 1656
rect 641 1644 710 1646
rect 641 1603 654 1644
rect 691 1605 710 1644
rect 747 1605 762 1646
rect 691 1603 762 1605
rect 641 1585 762 1603
rect 647 1483 726 1585
rect 1699 1545 1766 1564
rect 1699 1525 1719 1545
rect 173 1402 281 1457
rect 648 1402 726 1483
rect 1698 1479 1719 1525
rect 1749 1525 1766 1545
rect 1749 1495 1768 1525
rect 1749 1479 1769 1495
rect 1698 1463 1769 1479
rect 1348 1452 1420 1453
rect 1347 1444 1446 1452
rect 1347 1441 1399 1444
rect 1347 1406 1355 1441
rect 1380 1406 1399 1441
rect 1424 1406 1446 1444
rect 173 973 280 1402
rect 652 1161 724 1402
rect 1347 1394 1446 1406
rect 1348 1375 1416 1394
rect 1349 1372 1382 1375
rect 1584 1372 1616 1373
rect 759 1311 962 1324
rect 759 1278 783 1311
rect 819 1310 962 1311
rect 819 1307 930 1310
rect 819 1280 856 1307
rect 885 1283 930 1307
rect 959 1283 962 1310
rect 885 1280 962 1283
rect 819 1278 962 1280
rect 759 1265 962 1278
rect 759 1264 860 1265
rect 652 1119 661 1161
rect 710 1119 724 1161
rect 652 1098 724 1119
rect 652 1056 662 1098
rect 711 1056 724 1098
rect 652 1038 724 1056
rect 1137 1202 1169 1209
rect 1137 1182 1144 1202
rect 1165 1182 1169 1202
rect 1137 1117 1169 1182
rect 1349 1173 1380 1372
rect 1581 1367 1616 1372
rect 1581 1347 1588 1367
rect 1608 1347 1616 1367
rect 1581 1339 1616 1347
rect 1349 1143 1355 1173
rect 1376 1143 1380 1173
rect 1349 1135 1380 1143
rect 1507 1117 1547 1118
rect 1137 1115 1549 1117
rect 1137 1089 1517 1115
rect 1543 1089 1549 1115
rect 1137 1081 1549 1089
rect 1137 1053 1169 1081
rect 1582 1061 1616 1339
rect 1698 1152 1768 1463
rect 2395 1454 3737 1459
rect 2395 1452 3694 1454
rect 2392 1426 3694 1452
rect 3722 1426 3737 1454
rect 2392 1418 3737 1426
rect 2392 1393 2431 1418
rect 2392 1376 2433 1393
rect 2392 1369 2431 1376
rect 1807 1307 2010 1320
rect 1807 1274 1831 1307
rect 1867 1306 2010 1307
rect 1867 1303 1978 1306
rect 1867 1276 1904 1303
rect 1933 1279 1978 1303
rect 2007 1279 2010 1306
rect 1933 1276 2010 1279
rect 1867 1274 2010 1276
rect 1807 1261 2010 1274
rect 1807 1260 1908 1261
rect 1137 1033 1142 1053
rect 1163 1033 1169 1053
rect 1137 1026 1169 1033
rect 1560 1056 1616 1061
rect 1560 1036 1567 1056
rect 1587 1036 1616 1056
rect 1693 1146 1768 1152
rect 1693 1113 1701 1146
rect 1754 1113 1768 1146
rect 1693 1088 1768 1113
rect 1693 1055 1706 1088
rect 1759 1055 1768 1088
rect 1693 1046 1768 1055
rect 2185 1198 2217 1205
rect 2185 1178 2192 1198
rect 2213 1178 2217 1198
rect 2185 1113 2217 1178
rect 2397 1169 2428 1369
rect 2632 1368 2664 1369
rect 2629 1363 2664 1368
rect 2629 1343 2636 1363
rect 2656 1343 2664 1363
rect 2629 1335 2664 1343
rect 2397 1139 2403 1169
rect 2424 1139 2428 1169
rect 2397 1131 2428 1139
rect 2555 1113 2595 1114
rect 2185 1111 2597 1113
rect 2185 1085 2565 1111
rect 2591 1085 2597 1111
rect 2185 1077 2597 1085
rect 2185 1049 2217 1077
rect 2630 1057 2664 1335
rect 1693 1041 1751 1046
rect 1560 1029 1616 1036
rect 2185 1029 2190 1049
rect 2211 1029 2217 1049
rect 1560 1028 1595 1029
rect 2185 1022 2217 1029
rect 2608 1052 2664 1057
rect 2608 1032 2615 1052
rect 2635 1032 2664 1052
rect 2608 1025 2664 1032
rect 2608 1024 2643 1025
rect 851 973 962 977
rect 2726 973 4246 974
rect 173 955 4246 973
rect 173 935 859 955
rect 878 935 936 955
rect 955 951 4246 955
rect 955 935 1907 951
rect 173 931 1907 935
rect 1926 931 1984 951
rect 2003 931 4246 951
rect 173 917 4246 931
rect 173 294 280 917
rect 1899 914 2010 917
rect 659 868 723 872
rect 655 862 723 868
rect 655 829 672 862
rect 712 829 723 862
rect 655 817 723 829
rect 1706 831 1771 853
rect 655 815 712 817
rect 659 454 710 815
rect 1706 792 1723 831
rect 1768 792 1771 831
rect 1347 747 1382 749
rect 1347 738 1451 747
rect 1347 737 1398 738
rect 1347 717 1350 737
rect 1375 718 1398 737
rect 1430 718 1451 738
rect 1375 717 1451 718
rect 1347 710 1451 717
rect 1347 698 1382 710
rect 759 632 962 645
rect 759 599 783 632
rect 819 631 962 632
rect 819 628 930 631
rect 819 601 856 628
rect 885 604 930 628
rect 959 604 962 631
rect 885 601 962 604
rect 819 599 962 601
rect 759 586 962 599
rect 759 585 860 586
rect 1137 523 1169 530
rect 1137 503 1144 523
rect 1165 503 1169 523
rect 648 445 713 454
rect 648 408 658 445
rect 698 411 713 445
rect 1137 438 1169 503
rect 1349 494 1380 698
rect 1584 693 1616 694
rect 1581 688 1616 693
rect 1581 668 1588 688
rect 1608 668 1616 688
rect 1581 660 1616 668
rect 1349 464 1355 494
rect 1376 464 1380 494
rect 1349 456 1380 464
rect 1507 438 1547 439
rect 1137 436 1549 438
rect 698 408 715 411
rect 648 389 715 408
rect 648 368 662 389
rect 698 368 715 389
rect 648 361 715 368
rect 1137 410 1517 436
rect 1543 410 1549 436
rect 1137 402 1549 410
rect 1137 374 1169 402
rect 1582 382 1616 660
rect 1706 492 1771 792
rect 1137 354 1142 374
rect 1163 354 1169 374
rect 1137 347 1169 354
rect 1560 377 1616 382
rect 1560 357 1567 377
rect 1587 357 1616 377
rect 1560 350 1616 357
rect 1696 481 1776 492
rect 1696 455 1713 481
rect 1753 455 1776 481
rect 1696 428 1776 455
rect 1696 402 1717 428
rect 1757 402 1776 428
rect 1696 383 1776 402
rect 1696 357 1720 383
rect 1760 357 1776 383
rect 1560 349 1595 350
rect 1696 345 1776 357
rect 851 294 962 298
rect 2606 294 2813 295
rect 171 276 4246 294
rect 171 256 859 276
rect 878 256 936 276
rect 955 256 4246 276
rect 171 238 4246 256
rect 173 38 280 238
rect 2768 236 4246 238
rect 641 199 762 209
rect 641 197 710 199
rect 641 156 654 197
rect 691 158 710 197
rect 747 158 762 199
rect 691 156 762 158
rect 641 138 762 156
rect 647 0 712 138
<< via1 >>
rect 784 11700 820 11733
rect 1832 11696 1868 11729
rect 784 11021 820 11054
rect 3279 11016 3315 11049
rect 784 10253 820 10286
rect 1832 10249 1868 10282
rect 784 9574 820 9607
rect 3322 9571 3358 9604
rect 785 8733 821 8766
rect 1833 8729 1869 8762
rect 785 8054 821 8087
rect 3280 8049 3316 8082
rect 785 7286 821 7319
rect 1833 7282 1869 7315
rect 785 6607 821 6640
rect 4388 6598 4424 6631
rect 782 5692 818 5725
rect 1830 5688 1866 5721
rect 782 5013 818 5046
rect 3277 5008 3313 5041
rect 782 4245 818 4278
rect 1830 4241 1866 4274
rect 782 3566 818 3599
rect 3320 3563 3356 3596
rect 783 2725 819 2758
rect 1831 2721 1867 2754
rect 783 2046 819 2079
rect 3278 2041 3314 2074
rect 783 1278 819 1311
rect 1831 1274 1867 1307
rect 783 599 819 632
<< metal2 >>
rect 3 11748 110 11989
rect 3 11733 3748 11748
rect 3 11700 784 11733
rect 820 11729 3748 11733
rect 820 11700 1832 11729
rect 3 11696 1832 11700
rect 1868 11696 3748 11729
rect 3 11679 3748 11696
rect 3 11073 110 11679
rect 2610 11677 3748 11679
rect 3 11054 4143 11073
rect 3 11021 784 11054
rect 820 11049 4143 11054
rect 820 11021 3279 11049
rect 3 11016 3279 11021
rect 3315 11016 4143 11049
rect 3 11004 4143 11016
rect 3 10301 110 11004
rect 2531 11003 4143 11004
rect 2760 10304 3003 10309
rect 2708 10301 3968 10304
rect 3 10286 3968 10301
rect 3 10253 784 10286
rect 820 10282 3968 10286
rect 820 10253 1832 10282
rect 3 10249 1832 10253
rect 1868 10249 3968 10282
rect 3 10232 3968 10249
rect 3 9626 110 10232
rect 2760 10223 3003 10232
rect 2742 9626 4192 9628
rect 3 9607 4192 9626
rect 3 9574 784 9607
rect 820 9604 4192 9607
rect 820 9574 3322 9604
rect 3 9571 3322 9574
rect 3358 9571 4192 9604
rect 3 9557 4192 9571
rect 3 9022 110 9557
rect 2742 9556 4192 9557
rect 3 9021 111 9022
rect 4 8998 111 9021
rect 2 8954 111 8998
rect 4 8781 111 8954
rect 2752 8781 2940 8783
rect 4 8766 3936 8781
rect 4 8733 785 8766
rect 821 8762 3936 8766
rect 821 8733 1833 8762
rect 4 8729 1833 8733
rect 1869 8729 3936 8762
rect 4 8712 3936 8729
rect 4 8106 111 8712
rect 2611 8710 3936 8712
rect 4 8087 4145 8106
rect 4 8054 785 8087
rect 821 8082 4145 8087
rect 821 8054 3280 8082
rect 4 8049 3280 8054
rect 3316 8049 4145 8082
rect 4 8037 4145 8049
rect 4 7334 111 8037
rect 2532 8036 4145 8037
rect 2709 7334 3718 7337
rect 4 7319 3718 7334
rect 4 7286 785 7319
rect 821 7315 3718 7319
rect 821 7286 1833 7315
rect 4 7282 1833 7286
rect 1869 7282 3718 7315
rect 4 7265 3718 7282
rect 4 6659 111 7265
rect 2743 6660 4248 6661
rect 2743 6659 4448 6660
rect 4 6644 4448 6659
rect 4 6640 4451 6644
rect 4 6607 785 6640
rect 821 6631 4451 6640
rect 821 6607 4388 6631
rect 4 6598 4388 6607
rect 4424 6598 4451 6631
rect 4 6590 4451 6598
rect 4 6073 111 6590
rect 2743 6589 4451 6590
rect 4213 6586 4451 6589
rect -3 5881 113 6073
rect 1 5740 108 5881
rect 1 5725 4180 5740
rect 1 5692 782 5725
rect 818 5721 4180 5725
rect 818 5692 1830 5721
rect 1 5688 1830 5692
rect 1866 5688 4180 5721
rect 1 5671 4180 5688
rect 1 5065 108 5671
rect 2608 5669 4180 5671
rect 1 5046 4236 5065
rect 1 5013 782 5046
rect 818 5041 4236 5046
rect 818 5013 3277 5041
rect 1 5008 3277 5013
rect 3313 5008 4236 5041
rect 1 4996 4236 5008
rect 1 4293 108 4996
rect 2529 4995 4236 4996
rect 2758 4296 3001 4301
rect 2706 4293 4236 4296
rect 1 4278 4236 4293
rect 1 4245 782 4278
rect 818 4274 4236 4278
rect 818 4245 1830 4274
rect 1 4241 1830 4245
rect 1866 4241 4236 4274
rect 1 4224 4236 4241
rect 1 3618 108 4224
rect 2758 4215 3001 4224
rect 2740 3618 4236 3620
rect 1 3599 4236 3618
rect 1 3566 782 3599
rect 818 3596 4236 3599
rect 818 3566 3320 3596
rect 1 3563 3320 3566
rect 3356 3563 4236 3596
rect 1 3549 4236 3563
rect 1 3014 108 3549
rect 2740 3548 4236 3549
rect 1 3013 109 3014
rect 2 2990 109 3013
rect 0 2946 109 2990
rect 2 2773 109 2946
rect 2750 2773 2938 2775
rect 2 2758 4181 2773
rect 2 2725 783 2758
rect 819 2754 4181 2758
rect 819 2725 1831 2754
rect 2 2721 1831 2725
rect 1867 2721 4181 2754
rect 2 2704 4181 2721
rect 2 2098 109 2704
rect 2609 2702 4181 2704
rect 2 2079 4245 2098
rect 2 2046 783 2079
rect 819 2074 4245 2079
rect 819 2046 3278 2074
rect 2 2041 3278 2046
rect 3314 2041 4245 2074
rect 2 2029 4245 2041
rect 2 1326 109 2029
rect 2530 2028 4245 2029
rect 2707 1326 4246 1329
rect 2 1311 4246 1326
rect 2 1278 783 1311
rect 819 1307 4246 1311
rect 819 1278 1831 1307
rect 2 1274 1831 1278
rect 1867 1274 4246 1307
rect 2 1257 4246 1274
rect 2 651 109 1257
rect 2741 651 4246 653
rect 2 632 4246 651
rect 2 599 783 632
rect 819 599 4246 632
rect 2 582 4246 599
rect 2 36 109 582
rect 2741 581 4246 582
<< labels >>
rlabel locali 446 11940 490 11962 1 vref
rlabel metal1 182 11929 278 11962 1 gnd
rlabel metal2 6 11929 102 11962 1 vdd
rlabel metal1 661 11944 723 11971 1 d0
rlabel metal1 1707 11926 1760 11948 1 d1
rlabel metal1 2817 11989 2867 12002 1 d2
rlabel metal1 2993 11972 3045 11991 1 d3
rlabel metal1 4255 11981 4290 11995 1 d4
rlabel metal1 4958 6698 4983 6713 1 vout
<< end >>
