* SPICE3 file created from 6bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 a_1726_3204# a_1513_3204# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X1 a_852_7898# a_431_7898# a_116_8103# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X2 a_116_8333# a_645_8452# a_853_8452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3 gnd d0 a_4079_1330# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X4 a_648_177# a_435_177# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5 gnd d0 a_4080_227# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X6 a_2004_n382# a_2823_4353# a_2774_4543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X7 a_3821_4829# a_4078_4639# a_2883_5073# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X8 gnd d1 a_3138_8192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X9 gnd a_3000_3269# a_2792_3269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X10 a_2746_5488# a_2931_5986# a_2882_6176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X11 a_2889_484# a_3142_471# a_2744_1253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X12 gnd d1 a_3142_471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X13 a_1511_7616# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X14 a_3826_2446# a_3822_2623# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X15 vdd d0 a_4079_1330# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X16 a_3827_3000# a_4080_2987# a_2888_2690# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X17 a_2004_n382# a_2823_4353# a_2778_4366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X18 a_1513_3204# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X19 a_2887_4896# a_3871_5193# a_3822_5383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X20 a_2885_661# a_3142_471# a_2744_1253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X21 vdd d1 a_3142_471# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X22 a_116_8562# a_116_8333# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X23 a_647_5143# a_434_5143# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X24 gnd a_3138_8192# a_2930_8192# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X25 a_3826_2446# a_4079_2433# a_2884_2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X26 a_3820_7035# a_4077_6845# a_2882_7279# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X27 a_119_3234# a_119_3047# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X28 a_119_3047# a_648_2937# a_856_2937# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X29 a_117_6127# a_646_6246# a_854_6246# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X30 a_3822_2623# a_4079_2433# a_2884_2867# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X31 a_1586_2693# a_1373_2693# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X32 a_1694_4326# a_1481_4326# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X33 a_434_5143# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X34 a_2886_7102# a_3870_7399# a_3821_7589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X35 a_118_3691# a_119_3234# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X36 a_117_5897# a_645_5692# a_853_5692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X37 a_2776_6578# a_2790_7681# a_2741_7871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X38 a_2888_2690# a_3872_2987# a_3823_3177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X39 a_646_7349# a_433_7349# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X40 a_3826_1343# a_3822_1520# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X41 a_2884_2867# a_3141_2677# a_2743_3459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X42 a_119_1485# a_647_1280# a_855_1280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X43 a_853_5692# a_1584_6002# a_1792_6002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X44 gnd a_3031_4353# a_2823_4353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X45 a_3825_4652# a_4078_4639# a_2883_5073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X46 a_2776_6578# a_2790_7681# a_2745_7694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X47 a_2741_7871# a_2931_7089# a_2886_7102# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X48 a_855_1280# a_434_1280# a_119_1485# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X49 gnd a_3139_5986# a_2931_5986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X50 a_1373_2693# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X51 a_2778_2166# a_2792_3269# a_2747_3282# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X52 a_1481_4326# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X53 vdd a_3031_4353# a_2823_4353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X54 a_2882_7279# a_3869_6845# a_3824_6858# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X55 gnd a_4079_5193# a_3871_5193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X56 a_118_3921# a_647_4040# a_855_4040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X57 a_433_7349# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X58 a_116_8103# a_644_7898# a_852_7898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X59 gnd d0 a_4078_7399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X60 a_856_1834# a_435_1834# a_119_1944# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X61 a_1727_998# a_1514_998# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X62 a_118_3691# a_646_3486# a_854_3486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X63 a_2883_5073# a_3140_4883# a_2742_5665# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X64 vout a_1682_n382# a_1902_4326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X65 a_2772_6755# a_2791_5475# a_2742_5665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X66 a_857_731# a_436_731# a_120_841# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X67 a_2774_2343# a_2793_1063# a_2744_1253# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X68 a_2743_3459# a_2933_2677# a_2888_2690# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X69 a_2772_6755# a_2791_5475# a_2746_5488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X70 a_117_7000# a_117_6543# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X71 a_3824_6858# a_3820_7035# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X72 a_853_6795# a_432_6795# a_117_7000# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X73 gnd a_4078_7399# a_3870_7399# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X74 a_1792_7105# a_1371_7105# a_853_6795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X75 a_2774_2343# a_2793_1063# a_2748_1076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X76 a_2778_2166# a_3031_2153# a_2774_4543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X77 a_3826_4103# a_3822_4280# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X78 a_3819_8138# a_4076_7948# a_2881_8382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X79 a_3825_4652# a_3821_4829# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X80 a_855_2383# a_434_2383# a_119_2588# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X81 a_3827_1897# a_3823_2074# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X82 gnd a_4080_2987# a_3872_2987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X83 a_120_612# a_649_731# a_857_731# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X84 a_2888_2690# a_3141_2677# a_2743_3459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X85 a_2774_2343# a_3031_2153# a_2774_4543# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X86 vdd a_3139_7089# a_2931_7089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X87 a_3827_1897# a_4080_1884# a_2888_1587# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X88 a_2889_484# a_3873_781# a_3824_971# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X89 a_2778_2166# a_2792_3269# a_2743_3459# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X90 a_2742_5665# a_2932_4883# a_2887_4896# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X91 a_2887_3793# a_3871_4090# a_3822_4280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X92 a_645_8452# a_432_8452# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X93 a_1895_n382# a_1682_n382# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X94 a_649_731# a_436_731# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X95 a_1724_7616# a_1511_7616# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X96 a_3824_5755# a_4077_5742# a_2882_6176# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X97 a_647_4040# a_434_4040# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X98 a_2889_484# a_3873_781# a_3828_794# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X99 a_1794_2693# a_1373_2693# a_855_2383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X100 a_2778_4366# a_2821_6565# a_2772_6755# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X101 a_3826_1343# a_4079_1330# a_2884_1764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X102 a_1726_3204# a_1513_3204# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X103 a_854_4589# a_433_4589# a_118_4794# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X104 a_3822_5383# a_3825_4652# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X105 a_3820_5932# a_4077_5742# a_2882_6176# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X106 a_2774_4543# a_2823_2153# a_2774_2343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X107 a_2881_8382# a_3868_7948# a_3823_7961# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X108 a_119_1944# a_648_1834# a_856_1834# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X109 a_119_3047# a_119_2818# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X110 a_117_5897# a_118_5440# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X111 a_2745_7694# a_2998_7681# a_2776_6578# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X112 a_2778_4366# a_2821_6565# a_2776_6578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X113 a_3822_1520# a_4079_1330# a_2884_1764# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X114 a_432_8452# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X115 a_1682_n382# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X116 vdd a_3141_2677# a_2933_2677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X117 a_2743_3459# a_2933_2677# a_2884_2867# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X118 gnd d0 a_4077_8502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X119 a_1511_7616# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X120 a_2774_4543# a_2823_2153# a_2778_2166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X121 a_3825_7412# a_3821_7589# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X122 a_2886_5999# a_3870_6296# a_3821_6486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X123 a_118_3921# a_118_3691# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X124 a_434_4040# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X125 a_2741_7871# a_2998_7681# a_2776_6578# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X126 a_1513_3204# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X127 a_2885_661# a_3872_227# a_3827_240# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X128 a_2888_1587# a_3872_1884# a_3823_2074# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X129 a_646_6246# a_433_6246# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X130 a_1793_4899# a_1372_4899# a_854_4589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X131 a_3825_3549# a_4078_3536# a_2883_3970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X132 a_1725_5410# a_1512_5410# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X133 a_647_5143# a_434_5143# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X134 a_2882_6176# a_3869_5742# a_3820_5932# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X135 a_1727_998# a_1514_998# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X136 gnd a_4077_8502# a_3869_8502# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X137 a_3823_3177# a_4080_2987# a_2888_2690# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X138 a_3821_3726# a_4078_3536# a_2883_3970# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X139 a_1808_6645# a_1694_6526# a_1808_4445# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X140 a_1585_3796# a_1372_3796# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X141 vdd a_3140_4883# a_2932_4883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X142 a_2882_6176# a_3869_5742# a_3824_5755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X143 gnd a_4079_4090# a_3871_4090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X144 a_2887_3793# a_3140_3780# a_2747_3282# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X145 a_2746_5488# a_2999_5475# a_2772_6755# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X146 a_433_6246# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X147 a_1810_2233# a_1696_2114# a_1803_4326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X148 a_118_4150# a_118_3921# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X149 gnd d0 a_4078_6296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X150 a_1512_5410# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X151 a_434_5143# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X152 a_119_1944# a_119_1715# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X153 gnd a_3029_6565# a_2821_6565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X154 a_2883_3970# a_3140_3780# a_2747_3282# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X155 a_2742_5665# a_2999_5475# a_2772_6755# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X156 a_1514_998# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X157 a_646_7349# a_433_7349# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X158 a_117_7646# a_644_7898# a_852_7898# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X159 gnd a_3031_2153# a_2823_2153# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X160 a_2745_7694# a_2930_8192# a_2885_8205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X161 a_3825_6309# a_3821_6486# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X162 a_855_2383# a_1586_2693# a_1794_2693# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X163 a_1372_3796# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X164 vdd a_3029_6565# a_2821_6565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X165 a_648_2937# a_435_2937# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X166 gnd a_3141_2677# a_2933_2677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X167 a_120_841# a_120_612# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X168 vdd a_3031_2153# a_2823_2153# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X169 a_853_5692# a_432_5692# a_117_5897# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X170 a_2886_7102# a_3870_7399# a_3825_7412# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X171 a_645_6795# a_432_6795# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X172 gnd a_4078_6296# a_3870_6296# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X173 gnd d0 a_4077_6845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X174 a_1792_6002# a_1371_6002# a_853_5692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X175 a_435_177# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X176 a_2885_661# a_3872_227# a_3823_417# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X177 a_1586_1590# a_1373_1590# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X178 gnd a_4080_1884# a_3872_1884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X179 a_647_2383# a_434_2383# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X180 a_2888_2690# a_3872_2987# a_3827_3000# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X181 a_433_7349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X182 a_1808_4445# a_1481_6526# a_1803_6526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X183 a_2888_1587# a_3141_1574# a_2748_1076# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X184 a_2747_3282# a_2932_3780# a_2883_3970# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X185 a_1803_4326# a_1483_2114# a_1805_2114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X186 a_435_2937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X187 a_2884_1764# a_3141_1574# a_2748_1076# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X188 a_432_6795# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X189 a_2747_3282# a_2932_3780# a_2887_3793# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X190 vdd d1 a_3138_8192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X191 gnd a_4077_6845# a_3869_6845# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X192 a_117_7459# a_117_7230# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X193 gnd d0 a_4079_5193# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X194 a_1373_1590# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X195 a_434_2383# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X196 gnd a_4081_781# a_3873_781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X197 a_1791_8208# a_1370_8208# a_852_7898# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X198 a_1794_1590# a_1373_1590# a_855_1280# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X199 a_3823_7961# a_3819_8138# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X200 vdd d0 a_4078_7399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X201 a_854_3486# a_433_3486# a_118_3691# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X202 a_2887_4896# a_3871_5193# a_3826_5206# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X203 a_1792_7105# a_1371_7105# a_854_7349# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X204 a_3824_971# a_3827_240# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X205 a_646_4589# a_433_4589# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X206 vdd a_4081_781# a_3873_781# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X207 vout a_1682_n382# a_2004_n382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X208 a_2886_7102# a_3139_7089# a_2741_7871# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X209 vdd a_3138_8192# a_2930_8192# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X210 a_2748_1076# a_2933_1574# a_2884_1764# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X211 a_3820_5932# a_3826_5206# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X212 a_2746_5488# a_2931_5986# a_2886_5999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X213 gnd d1 a_3140_4883# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X214 vdd a_4078_7399# a_3870_7399# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X215 a_120_1028# a_647_1280# a_855_1280# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X216 a_119_2588# a_119_2131# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X217 a_2748_1076# a_2933_1574# a_2888_1587# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X218 a_645_8452# a_432_8452# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X219 a_433_4589# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X220 vdd a_4080_2987# a_3872_2987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X221 gnd d0 a_4080_2987# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X222 a_1793_3796# a_1372_3796# a_854_3486# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X223 vdd a_4080_227# a_3872_227# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X224 gnd a_3140_3780# a_2932_3780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X225 a_117_6356# a_117_6127# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X226 a_1793_4899# a_1372_4899# a_855_5143# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X227 a_119_1715# a_648_1834# a_856_1834# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X228 vdd d2 a_3000_3269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X229 a_1895_n382# a_1682_n382# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X230 vdd a_3140_3780# a_2932_3780# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X231 a_432_8452# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X232 gnd d1 a_3139_7089# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X233 a_3828_794# a_4081_781# a_2889_484# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X234 vdd a_4079_5193# a_3871_5193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X235 a_117_6543# a_645_6795# a_853_6795# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X236 a_648_2937# a_435_2937# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X237 a_855_5143# a_434_5143# a_118_5024# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X238 a_646_6246# a_433_6246# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X239 gnd d2 a_2999_5475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X240 a_857_731# a_1587_487# a_1795_487# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X241 a_1682_n382# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X242 a_119_2131# a_647_2383# a_855_2383# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X243 a_3824_971# a_4081_781# a_2889_484# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X244 a_119_1485# a_120_1028# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X245 gnd d2 a_3001_1063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X246 gnd a_3141_1574# a_2933_1574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X247 vdd a_3139_5986# a_2931_5986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X248 a_1795_487# a_1374_487# a_857_731# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X249 a_3822_4280# a_3825_3549# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X250 a_1808_4445# a_1694_4326# a_1902_4326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X251 vdd d2 a_2999_5475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X252 a_1374_487# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X253 a_645_5692# a_432_5692# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X254 a_3827_3000# a_3823_3177# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X255 a_2885_8205# a_3138_8192# a_2745_7694# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X256 a_1803_6526# a_1694_6526# a_1808_4445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X257 vdd d2 a_3001_1063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X258 vdd a_3141_1574# a_2933_1574# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X259 a_647_1280# a_434_1280# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X260 a_116_8103# a_117_7646# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X261 a_435_2937# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X262 a_433_6246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X263 a_120_382# a_122_283# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X264 a_1805_2114# a_1696_2114# a_1803_4326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X265 gnd a_4080_227# a_3872_227# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X266 a_854_7349# a_433_7349# a_117_7230# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X267 a_853_8452# a_1583_8208# a_1791_8208# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X268 a_854_3486# a_1585_3796# a_1793_3796# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X269 a_436_731# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X270 a_3823_417# a_4080_227# a_2885_661# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X271 a_647_4040# a_434_4040# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X272 a_118_4337# a_646_4589# a_854_4589# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X273 a_432_5692# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X274 gnd d2 a_3000_3269# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X275 gnd d0 a_4079_4090# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X276 a_434_1280# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X277 a_644_7898# a_431_7898# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X278 gnd d0 a_4076_7948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X279 a_3819_8138# a_3825_7412# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X280 a_1792_6002# a_1371_6002# a_854_6246# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X281 a_1587_487# a_1374_487# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X282 a_646_3486# a_433_3486# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X283 a_2887_3793# a_3871_4090# a_3826_4103# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X284 a_435_177# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X285 a_1902_4326# a_1481_4326# a_1803_4326# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X286 a_2886_5999# a_3139_5986# a_2746_5488# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X287 a_1808_4445# a_1481_6526# a_1808_6645# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X288 gnd a_3142_471# a_2934_471# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X289 a_434_4040# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X290 a_118_4794# a_118_4337# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X291 a_1803_4326# a_1483_2114# a_1810_2233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X292 a_3826_5206# a_4079_5193# a_2887_4896# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X293 a_431_7898# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X294 a_119_2818# a_119_2588# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X295 gnd a_4076_7948# a_3868_7948# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X296 vdd a_3142_471# a_2934_471# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X297 a_855_1280# a_1586_1590# a_1794_1590# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X298 a_1792_6002# a_1725_5410# a_1803_6526# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X299 a_3823_2074# a_4080_1884# a_2888_1587# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X300 a_3822_2623# a_3827_1897# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X301 a_433_3486# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X302 gnd d0 a_4080_1884# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X303 vdd d0 a_4077_8502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X304 a_2886_5999# a_3870_6296# a_3825_6309# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X305 a_1791_8208# a_1370_8208# a_853_8452# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X306 a_3827_240# a_4080_227# a_2885_661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X307 gnd d4 a_3031_4353# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X308 a_3825_7412# a_4078_7399# a_2886_7102# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X309 a_1584_7105# a_1371_7105# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X310 gnd d1 a_3139_5986# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X311 vdd a_4077_8502# a_3869_8502# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X312 a_1791_8208# a_1724_7616# a_1808_6645# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X313 a_2883_5073# a_3870_4639# a_3825_4652# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X314 vref a_116_8562# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X315 a_853_8452# a_432_8452# a_116_8333# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X316 a_3820_8692# a_3823_7961# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X317 a_1793_3796# a_1726_3204# a_1810_2233# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X318 vdd d4 a_3031_4353# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X319 vdd a_4079_4090# a_3871_4090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X320 a_648_1834# a_435_1834# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X321 a_1803_6526# a_1512_5410# a_1793_4899# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X322 a_855_4040# a_434_4040# a_118_3921# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X323 a_118_5440# a_645_5692# a_853_5692# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X324 a_2882_7279# a_3139_7089# a_2741_7871# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X325 a_2888_1587# a_3872_1884# a_3827_1897# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X326 vdd d0 a_4078_6296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X327 a_119_1715# a_119_1485# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X328 a_3826_5206# a_3822_5383# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X329 a_1371_7105# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X330 a_3822_1520# a_3828_794# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X331 a_2884_2867# a_3871_2433# a_3822_2623# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X332 a_1586_2693# a_1373_2693# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X333 a_435_1834# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X334 a_120_612# a_120_382# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X335 vdd d0 a_4080_2987# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X336 vdd d0 a_4078_4639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X337 a_1805_2114# a_1514_998# a_1795_487# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X338 a_2884_2867# a_3871_2433# a_3826_2446# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X339 vdd a_4078_6296# a_3870_6296# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X340 a_1514_998# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X341 a_1808_6645# a_1511_7616# a_1792_7105# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X342 a_854_6246# a_433_6246# a_117_6127# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X343 a_3823_417# a_122_283# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X344 a_1810_2233# a_1513_3204# a_1794_2693# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X345 a_119_3234# a_646_3486# a_854_3486# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X346 a_855_5143# a_434_5143# a_118_5253# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X347 a_1373_2693# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X348 vdd d1 a_3139_7089# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X349 vdd a_4078_4639# a_3870_4639# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X350 a_2883_5073# a_3870_4639# a_3821_4829# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X351 a_1803_4326# a_1694_4326# a_1902_4326# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X352 a_1585_4899# a_1372_4899# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X353 a_117_7230# a_117_7000# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X354 vdd d0 a_4079_5193# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X355 vdd d0 a_4077_6845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X356 a_644_7898# a_431_7898# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X357 a_118_5024# a_118_4794# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X358 vdd a_4080_1884# a_3872_1884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X359 gnd a_4077_8502# a_2885_8205# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X360 a_3827_240# a_3823_417# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X361 a_119_2131# a_119_1944# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X362 a_3821_4829# a_3826_4103# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X363 a_854_7349# a_433_7349# a_117_7459# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X364 a_3826_4103# a_4079_4090# a_2887_3793# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X365 a_852_7898# a_1583_8208# a_1791_8208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X366 a_436_731# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X367 gnd a_4079_2433# a_3871_2433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X368 a_856_2937# a_435_2937# a_119_3047# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X369 a_1372_4899# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X370 vdd a_4077_6845# a_3869_6845# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X371 vdd d1 a_3141_2677# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X372 a_431_7898# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X373 a_2776_6578# a_3029_6565# a_2778_4366# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X374 a_853_6795# a_432_6795# a_117_6543# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X375 gnd d0 a_4078_4639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X376 vdd a_4079_2433# a_3871_2433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X377 a_855_2383# a_434_2383# a_119_2131# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X378 a_1794_2693# a_1373_2693# a_856_2937# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X379 a_2772_6755# a_3029_6565# a_2778_4366# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X380 a_118_5253# a_118_5024# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X381 a_1902_4326# a_1481_4326# a_1808_4445# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X382 a_3825_6309# a_4078_6296# a_2886_5999# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X383 a_118_5253# a_647_5143# a_855_5143# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X384 a_117_6127# a_117_5897# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X385 a_1584_6002# a_1371_6002# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X386 a_2885_8205# a_3869_8502# a_3820_8692# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X387 gnd a_4078_4639# a_3870_4639# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X388 a_1694_6526# a_1481_6526# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X389 vdd d1 a_3140_4883# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X390 a_3821_3726# a_3827_3000# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X391 a_1696_2114# a_1483_2114# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X392 a_118_5440# a_118_5253# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X393 a_3828_794# a_3824_971# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X394 a_854_4589# a_433_4589# a_118_4337# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X395 a_3824_6858# a_4077_6845# a_2882_7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X396 gnd d3 a_3029_6565# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X397 a_1371_6002# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X398 a_647_1280# a_434_1280# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X399 a_3823_3177# a_3826_2446# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X400 a_2884_1764# a_3871_1330# a_3822_1520# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X401 gnd d3 a_3031_2153# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X402 a_1583_8208# a_1370_8208# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X403 vdd d0 a_4076_7948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X404 a_117_7459# a_646_7349# a_854_7349# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X405 a_1481_6526# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X406 a_1586_1590# a_1373_1590# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X407 vdd d3 a_3029_6565# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X408 a_2004_n382# a_1895_n382# vout vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X409 a_1584_7105# a_1371_7105# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X410 a_1483_2114# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X411 gnd d1 a_3141_2677# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X412 a_3825_3549# a_3821_3726# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X413 a_1792_7105# a_1724_7616# a_1808_6645# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X414 a_2884_1764# a_3871_1330# a_3826_1343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X415 vdd d3 a_3031_2153# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X416 a_853_8452# a_432_8452# a_116_8562# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X417 a_2881_8382# a_3138_8192# a_2745_7694# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X418 a_1794_2693# a_1726_3204# a_1810_2233# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X419 a_434_1280# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X420 a_648_1834# a_435_1834# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X421 a_854_7349# a_1584_7105# a_1792_7105# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X422 a_1370_8208# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X423 vdd a_4076_7948# a_3868_7948# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X424 a_1373_1590# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X425 a_3821_7589# a_4078_7399# a_2886_7102# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X426 gnd d0 a_4077_5742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X427 a_1371_7105# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X428 a_2883_3970# a_3870_3536# a_3821_3726# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X429 a_2882_7279# a_3869_6845# a_3820_7035# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X430 a_3820_7035# a_3825_6309# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X431 a_1585_3796# a_1372_3796# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X432 a_118_4337# a_118_4150# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X433 a_645_6795# a_432_6795# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X434 a_856_177# a_435_177# a_122_283# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X435 vdd d0 a_4079_4090# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X436 vdd d0 a_4077_5742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X437 a_2883_3970# a_3870_3536# a_3825_3549# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X438 a_435_1834# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X439 a_647_2383# a_434_2383# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X440 a_3823_2074# a_3826_1343# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X441 a_1585_4899# a_1372_4899# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X442 a_2744_1253# a_2934_471# a_2885_661# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X443 a_2887_4896# a_3140_4883# a_2742_5665# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X444 a_1793_4899# a_1725_5410# a_1803_6526# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X445 a_856_2937# a_435_2937# a_119_2818# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X446 a_1808_6645# a_1511_7616# a_1791_8208# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X447 a_854_6246# a_433_6246# a_117_6356# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X448 gnd a_4077_5742# a_3869_5742# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X449 a_1795_487# a_1727_998# a_1805_2114# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X450 a_856_2937# a_1586_2693# a_1794_2693# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X451 gnd a_4079_1330# a_3871_1330# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X452 a_2744_1253# a_2934_471# a_2889_484# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X453 a_120_382# a_648_177# a_856_177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X454 a_1810_2233# a_1513_3204# a_1793_3796# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X455 a_1372_3796# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X456 a_120_1028# a_120_841# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X457 a_432_6795# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X458 vdd a_4077_5742# a_3869_5742# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X459 a_3822_5383# a_4079_5193# a_2887_4896# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X460 gnd d0 a_4078_3536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X461 a_853_5692# a_432_5692# a_118_5440# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X462 a_434_2383# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X463 vdd a_4079_1330# a_3871_1330# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X464 a_1372_4899# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X465 a_116_8333# a_116_8103# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X466 a_855_1280# a_434_1280# a_120_1028# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X467 a_2743_3459# a_3000_3269# a_2778_2166# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X468 a_646_4589# a_433_4589# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X469 a_116_8562# a_645_8452# a_853_8452# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X470 vdd d0 a_4078_3536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X471 a_648_177# a_435_177# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X472 a_2882_6176# a_3139_5986# a_2746_5488# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X473 gnd d1 a_3140_3780# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X474 a_118_4150# a_647_4040# a_855_4040# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X475 a_1794_1590# a_1727_998# a_1805_2114# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X476 a_117_7646# a_117_7459# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X477 a_855_5143# a_1585_4899# a_1793_4899# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X478 gnd a_4078_3536# a_3870_3536# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X479 a_855_4040# a_434_4040# a_118_4150# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X480 a_2742_5665# a_2932_4883# a_2883_5073# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X481 a_1803_6526# a_1512_5410# a_1792_6002# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X482 a_3821_7589# a_3824_6858# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X483 vdd d1 a_3140_3780# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X484 a_1805_2114# a_1514_998# a_1794_1590# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X485 a_852_7898# a_431_7898# a_117_7646# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X486 a_433_4589# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X487 a_2748_1076# a_3001_1063# a_2774_2343# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X488 vdd a_4078_3536# a_3870_3536# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X489 vdd d0 a_4080_1884# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X490 a_854_3486# a_433_3486# a_119_3234# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X491 a_1793_3796# a_1372_3796# a_855_4040# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X492 a_3824_5755# a_3820_5932# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X493 a_2744_1253# a_3001_1063# a_2774_2343# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X494 a_117_6356# a_646_6246# a_854_6246# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X495 gnd d0 a_4079_2433# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X496 a_1584_6002# a_1371_6002# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X497 gnd d1 a_3141_1574# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X498 a_118_5024# a_647_5143# a_855_5143# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X499 a_2741_7871# a_2931_7089# a_2882_7279# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X500 a_1694_4326# a_1481_4326# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X501 vdd d1 a_3139_5986# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X502 a_1694_6526# a_1481_6526# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X503 vdd d0 a_4079_2433# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X504 gnd d0 a_4081_781# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X505 vdd d1 a_3141_1574# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X506 a_2747_3282# a_3000_3269# a_2778_2166# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X507 gnd d2 a_2998_7681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X508 a_1696_2114# a_1483_2114# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X509 a_117_6543# a_117_6356# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X510 a_854_6246# a_1584_6002# a_1792_6002# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X511 a_3823_7961# a_4076_7948# a_2881_8382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X512 vdd d0 a_4081_781# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X513 a_856_177# a_1587_487# a_1795_487# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X514 a_1794_1590# a_1373_1590# a_856_1834# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X515 vdd d2 a_2998_7681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X516 a_1371_6002# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X517 a_3821_6486# a_3824_5755# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X518 a_1481_4326# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X519 gnd a_3140_4883# a_2932_4883# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X520 a_1481_6526# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X521 a_645_5692# a_432_5692# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X522 a_1583_8208# a_1370_8208# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X523 a_117_7230# a_646_7349# a_854_7349# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X524 gnd a_2998_7681# a_2790_7681# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X525 a_1483_2114# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X526 a_119_2818# a_648_2937# a_856_2937# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X527 gnd a_3820_8692# gnd sky130_fd_pr__res_generic_nd w=17 l=81
X528 a_856_1834# a_435_1834# a_119_1715# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X529 a_117_7000# a_645_6795# a_853_6795# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X530 vdd a_2998_7681# a_2790_7681# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X531 a_856_1834# a_1586_1590# a_1794_1590# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X532 a_857_731# a_436_731# a_120_612# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X533 vdd d0 a_4080_227# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X534 a_3820_8692# a_4077_8502# a_2885_8205# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X535 a_119_2588# a_647_2383# a_855_2383# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X536 vdd a_3000_3269# a_2792_3269# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X537 a_853_6795# a_1584_7105# a_1792_7105# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X538 a_432_5692# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X539 a_1370_8208# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X540 a_1902_4326# a_1895_n382# vout gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X541 gnd a_3139_7089# a_2931_7089# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X542 a_3822_4280# a_4079_4090# a_2887_3793# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X543 a_2881_8382# a_3868_7948# a_3819_8138# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X544 a_1374_487# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X545 a_1795_487# a_1374_487# a_856_177# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X546 a_1725_5410# a_1512_5410# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X547 a_1587_487# a_1374_487# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X548 a_856_177# a_435_177# a_120_382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X549 a_646_3486# a_433_3486# vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X550 a_2778_4366# a_3031_4353# a_2004_n382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X551 a_120_841# a_649_731# a_857_731# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X552 gnd a_2999_5475# a_2791_5475# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X553 a_2745_7694# a_2930_8192# a_2881_8382# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X554 gnd a_3001_1063# a_2793_1063# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X555 a_855_4040# a_1585_3796# a_1793_3796# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X556 a_2774_4543# a_3031_4353# a_2004_n382# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X557 a_118_4794# a_646_4589# a_854_4589# gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X558 vdd a_2999_5475# a_2791_5475# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X559 a_1512_5410# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X560 a_3821_6486# a_4078_6296# a_2886_5999# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X561 vdd a_3001_1063# a_2793_1063# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X562 a_122_283# a_648_177# a_856_177# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X563 a_649_731# a_436_731# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X564 a_854_4589# a_1585_4899# a_1793_4899# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X565 a_2885_8205# a_3869_8502# gnd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X566 a_1724_7616# a_1511_7616# gnd gnd sky130_fd_pr__nfet_01v8 w=42 l=50
X567 a_433_3486# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50
C0 a_1902_4326# a_2004_n382# 8.08fF
C1 a_3823_417# gnd 2.22fF
C2 a_122_283# gnd 6.43fF
C3 d0 gnd 11.73fF
C4 a_3827_240# gnd 2.38fF
C5 a_120_382# gnd 2.23fF
C6 a_2885_661# gnd 2.38fF
C7 d1 gnd 5.62fF
C8 a_856_177# gnd 2.52fF
C9 a_120_612# gnd 2.38fF
C10 a_857_731# gnd 2.18fF
C11 a_120_841# gnd 2.28fF
C12 a_2889_484# gnd 2.52fF
C13 a_3824_971# gnd 2.23fF
C14 a_3828_794# gnd 2.49fF
C15 d2 gnd 3.21fF
C16 a_3822_1520# gnd 2.28fF
C17 a_120_1028# gnd 2.49fF
C18 a_3826_1343# gnd 2.38fF
C19 a_119_1485# gnd 2.23fF
C20 a_2884_1764# gnd 2.18fF
C21 a_855_1280# gnd 2.52fF
C22 a_119_1715# gnd 2.38fF
C23 a_856_1834# gnd 2.45fF
C24 a_119_1944# gnd 2.28fF
C25 a_2888_1587# gnd 2.52fF
C26 a_3823_2074# gnd 2.23fF
C27 a_1805_2114# gnd 2.28fF
C28 a_3827_1897# gnd 2.49fF
C29 a_2774_2343# gnd 2.04fF
C30 a_3822_2623# gnd 2.28fF
C31 a_119_2131# gnd 2.49fF
C32 a_3826_2446# gnd 2.38fF
C33 a_119_2588# gnd 2.23fF
C34 a_2884_2867# gnd 2.45fF
C35 a_855_2383# gnd 2.52fF
C36 a_119_2818# gnd 2.38fF
C37 a_856_2937# gnd 2.18fF
C38 a_119_3047# gnd 2.28fF
C39 a_2888_2690# gnd 2.52fF
C40 a_3823_3177# gnd 2.23fF
C41 a_3827_3000# gnd 2.49fF
C42 a_1810_2233# gnd 2.45fF
C43 a_2778_2166# gnd 2.34fF
C44 a_3821_3726# gnd 2.28fF
C45 a_119_3234# gnd 2.49fF
C46 a_3825_3549# gnd 2.38fF
C47 a_118_3691# gnd 2.23fF
C48 a_2883_3970# gnd 2.18fF
C49 a_854_3486# gnd 2.52fF
C50 a_118_3921# gnd 2.38fF
C51 a_855_4040# gnd 2.45fF
C52 a_118_4150# gnd 2.28fF
C53 a_2887_3793# gnd 2.52fF
C54 a_3822_4280# gnd 2.23fF
C55 a_3826_4103# gnd 2.50fF
C56 a_2004_n382# gnd 6.48fF
C57 a_1803_4326# gnd 3.68fF
C58 a_1902_4326# gnd 5.48fF
C59 a_2774_4543# gnd 3.32fF
C60 a_3821_4829# gnd 2.28fF
C61 a_118_4337# gnd 2.50fF
C62 a_3825_4652# gnd 2.38fF
C63 a_118_4794# gnd 2.23fF
C64 a_2883_5073# gnd 2.45fF
C65 a_854_4589# gnd 2.52fF
C66 a_118_5024# gnd 2.38fF
C67 a_855_5143# gnd 2.18fF
C68 a_118_5253# gnd 2.28fF
C69 a_2887_4896# gnd 2.52fF
C70 a_3822_5383# gnd 2.23fF
C71 a_3826_5206# gnd 2.49fF
C72 a_3820_5932# gnd 2.28fF
C73 a_118_5440# gnd 2.49fF
C74 a_3824_5755# gnd 2.38fF
C75 a_117_5897# gnd 2.23fF
C76 a_2882_6176# gnd 2.18fF
C77 a_853_5692# gnd 2.52fF
C78 a_117_6127# gnd 2.38fF
C79 a_854_6246# gnd 2.45fF
C80 a_117_6356# gnd 2.28fF
C81 a_2886_5999# gnd 2.52fF
C82 a_3821_6486# gnd 2.23fF
C83 a_1803_6526# gnd 2.34fF
C84 a_1808_4445# gnd 3.32fF
C85 a_3825_6309# gnd 2.49fF
C86 a_2778_4366# gnd 3.68fF
C87 a_2772_6755# gnd 2.45fF
C88 a_3820_7035# gnd 2.28fF
C89 a_117_6543# gnd 2.49fF
C90 a_3824_6858# gnd 2.38fF
C91 a_117_7000# gnd 2.23fF
C92 a_2882_7279# gnd 2.45fF
C93 a_853_6795# gnd 2.52fF
C94 a_117_7230# gnd 2.38fF
C95 a_854_7349# gnd 2.18fF
C96 a_117_7459# gnd 2.28fF
C97 a_2886_7102# gnd 2.52fF
C98 a_3821_7589# gnd 2.23fF
C99 a_3825_7412# gnd 2.49fF
C100 a_1808_6645# gnd 2.04fF
C101 a_2776_6578# gnd 2.28fF
C102 a_3819_8138# gnd 2.28fF
C103 a_117_7646# gnd 2.49fF
C104 a_3823_7961# gnd 2.38fF
C105 a_116_8103# gnd 2.23fF
C106 a_2881_8382# gnd 2.18fF
C107 a_852_7898# gnd 2.52fF
C108 a_116_8333# gnd 2.38fF
C109 a_853_8452# gnd 2.38fF
C110 a_116_8562# gnd 2.22fF
C111 a_2885_8205# gnd 2.79fF
C112 a_3820_8692# gnd 2.75fF
C113 vdd gnd 110.57fF
