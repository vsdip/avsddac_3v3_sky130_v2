magic
tech sky130A
timestamp 1633147515
<< nwell >>
rect 41 785 852 1009
rect 1089 781 1900 1005
rect 41 106 852 330
<< nmos >>
rect 105 684 155 726
rect 318 684 368 726
rect 526 684 576 726
rect 734 684 784 726
rect 1153 680 1203 722
rect 1366 680 1416 722
rect 1574 680 1624 722
rect 1782 680 1832 722
rect 105 5 155 47
rect 318 5 368 47
rect 526 5 576 47
rect 734 5 784 47
<< pmos >>
rect 105 803 155 903
rect 318 803 368 903
rect 526 803 576 903
rect 734 803 784 903
rect 1153 799 1203 899
rect 1366 799 1416 899
rect 1574 799 1624 899
rect 1782 799 1832 899
rect 105 124 155 224
rect 318 124 368 224
rect 526 124 576 224
rect 734 124 784 224
<< ndiff >>
rect 56 716 105 726
rect 56 696 67 716
rect 87 696 105 716
rect 56 684 105 696
rect 155 720 199 726
rect 155 700 170 720
rect 190 700 199 720
rect 155 684 199 700
rect 269 716 318 726
rect 269 696 280 716
rect 300 696 318 716
rect 269 684 318 696
rect 368 720 412 726
rect 368 700 383 720
rect 403 700 412 720
rect 368 684 412 700
rect 477 716 526 726
rect 477 696 488 716
rect 508 696 526 716
rect 477 684 526 696
rect 576 720 620 726
rect 576 700 591 720
rect 611 700 620 720
rect 576 684 620 700
rect 690 720 734 726
rect 690 700 699 720
rect 719 700 734 720
rect 690 684 734 700
rect 784 716 833 726
rect 784 696 802 716
rect 822 696 833 716
rect 784 684 833 696
rect 1104 712 1153 722
rect 1104 692 1115 712
rect 1135 692 1153 712
rect 1104 680 1153 692
rect 1203 716 1247 722
rect 1203 696 1218 716
rect 1238 696 1247 716
rect 1203 680 1247 696
rect 1317 712 1366 722
rect 1317 692 1328 712
rect 1348 692 1366 712
rect 1317 680 1366 692
rect 1416 716 1460 722
rect 1416 696 1431 716
rect 1451 696 1460 716
rect 1416 680 1460 696
rect 1525 712 1574 722
rect 1525 692 1536 712
rect 1556 692 1574 712
rect 1525 680 1574 692
rect 1624 716 1668 722
rect 1624 696 1639 716
rect 1659 696 1668 716
rect 1624 680 1668 696
rect 1738 716 1782 722
rect 1738 696 1747 716
rect 1767 696 1782 716
rect 1738 680 1782 696
rect 1832 712 1881 722
rect 1832 692 1850 712
rect 1870 692 1881 712
rect 1832 680 1881 692
rect 56 37 105 47
rect 56 17 67 37
rect 87 17 105 37
rect 56 5 105 17
rect 155 41 199 47
rect 155 21 170 41
rect 190 21 199 41
rect 155 5 199 21
rect 269 37 318 47
rect 269 17 280 37
rect 300 17 318 37
rect 269 5 318 17
rect 368 41 412 47
rect 368 21 383 41
rect 403 21 412 41
rect 368 5 412 21
rect 477 37 526 47
rect 477 17 488 37
rect 508 17 526 37
rect 477 5 526 17
rect 576 41 620 47
rect 576 21 591 41
rect 611 21 620 41
rect 576 5 620 21
rect 690 41 734 47
rect 690 21 699 41
rect 719 21 734 41
rect 690 5 734 21
rect 784 37 833 47
rect 784 17 802 37
rect 822 17 833 37
rect 784 5 833 17
<< pdiff >>
rect 61 865 105 903
rect 61 845 73 865
rect 93 845 105 865
rect 61 803 105 845
rect 155 865 197 903
rect 155 845 169 865
rect 189 845 197 865
rect 155 803 197 845
rect 274 865 318 903
rect 274 845 286 865
rect 306 845 318 865
rect 274 803 318 845
rect 368 865 410 903
rect 368 845 382 865
rect 402 845 410 865
rect 368 803 410 845
rect 482 865 526 903
rect 482 845 494 865
rect 514 845 526 865
rect 482 803 526 845
rect 576 865 618 903
rect 576 845 590 865
rect 610 845 618 865
rect 576 803 618 845
rect 692 865 734 903
rect 692 845 700 865
rect 720 845 734 865
rect 692 803 734 845
rect 784 872 829 903
rect 784 865 828 872
rect 784 845 796 865
rect 816 845 828 865
rect 784 803 828 845
rect 1109 861 1153 899
rect 1109 841 1121 861
rect 1141 841 1153 861
rect 1109 799 1153 841
rect 1203 861 1245 899
rect 1203 841 1217 861
rect 1237 841 1245 861
rect 1203 799 1245 841
rect 1322 861 1366 899
rect 1322 841 1334 861
rect 1354 841 1366 861
rect 1322 799 1366 841
rect 1416 861 1458 899
rect 1416 841 1430 861
rect 1450 841 1458 861
rect 1416 799 1458 841
rect 1530 861 1574 899
rect 1530 841 1542 861
rect 1562 841 1574 861
rect 1530 799 1574 841
rect 1624 861 1666 899
rect 1624 841 1638 861
rect 1658 841 1666 861
rect 1624 799 1666 841
rect 1740 861 1782 899
rect 1740 841 1748 861
rect 1768 841 1782 861
rect 1740 799 1782 841
rect 1832 868 1877 899
rect 1832 861 1876 868
rect 1832 841 1844 861
rect 1864 841 1876 861
rect 1832 799 1876 841
rect 61 186 105 224
rect 61 166 73 186
rect 93 166 105 186
rect 61 124 105 166
rect 155 186 197 224
rect 155 166 169 186
rect 189 166 197 186
rect 155 124 197 166
rect 274 186 318 224
rect 274 166 286 186
rect 306 166 318 186
rect 274 124 318 166
rect 368 186 410 224
rect 368 166 382 186
rect 402 166 410 186
rect 368 124 410 166
rect 482 186 526 224
rect 482 166 494 186
rect 514 166 526 186
rect 482 124 526 166
rect 576 186 618 224
rect 576 166 590 186
rect 610 166 618 186
rect 576 124 618 166
rect 692 186 734 224
rect 692 166 700 186
rect 720 166 734 186
rect 692 124 734 166
rect 784 193 829 224
rect 784 186 828 193
rect 784 166 796 186
rect 816 166 828 186
rect 784 124 828 166
<< ndiffc >>
rect -253 1019 -235 1037
rect -251 920 -233 938
rect -253 763 -235 781
rect 67 696 87 716
rect 170 700 190 720
rect 280 696 300 716
rect 383 700 403 720
rect 488 696 508 716
rect 591 700 611 720
rect 699 700 719 720
rect 802 696 822 716
rect 1115 692 1135 712
rect -251 664 -233 682
rect 1218 696 1238 716
rect 1328 692 1348 712
rect 1431 696 1451 716
rect 1536 692 1556 712
rect 1639 696 1659 716
rect 1747 696 1767 716
rect 1850 692 1870 712
rect -253 368 -235 386
rect -251 269 -233 287
rect -253 113 -235 131
rect -251 14 -233 32
rect 67 17 87 37
rect 170 21 190 41
rect 280 17 300 37
rect 383 21 403 41
rect 488 17 508 37
rect 591 21 611 41
rect 699 21 719 41
rect 802 17 822 37
<< pdiffc >>
rect 73 845 93 865
rect 169 845 189 865
rect 286 845 306 865
rect 382 845 402 865
rect 494 845 514 865
rect 590 845 610 865
rect 700 845 720 865
rect 796 845 816 865
rect 1121 841 1141 861
rect 1217 841 1237 861
rect 1334 841 1354 861
rect 1430 841 1450 861
rect 1542 841 1562 861
rect 1638 841 1658 861
rect 1748 841 1768 861
rect 1844 841 1864 861
rect 73 166 93 186
rect 169 166 189 186
rect 286 166 306 186
rect 382 166 402 186
rect 494 166 514 186
rect 590 166 610 186
rect 700 166 720 186
rect 796 166 816 186
<< psubdiff >>
rect 141 629 252 643
rect 141 599 182 629
rect 210 599 252 629
rect 141 584 252 599
rect 1189 625 1300 639
rect 1189 595 1230 625
rect 1258 595 1300 625
rect 1189 580 1300 595
rect 141 -50 252 -36
rect 141 -80 182 -50
rect 210 -80 252 -50
rect 141 -95 252 -80
<< nsubdiff >>
rect 142 976 252 990
rect 142 946 185 976
rect 213 946 252 976
rect 142 931 252 946
rect 1190 972 1300 986
rect 1190 942 1233 972
rect 1261 942 1300 972
rect 1190 927 1300 942
rect 142 297 252 311
rect 142 267 185 297
rect 213 267 252 297
rect 142 252 252 267
<< psubdiffcont >>
rect 182 599 210 629
rect 1230 595 1258 625
rect 182 -80 210 -50
<< nsubdiffcont >>
rect 185 946 213 976
rect 1233 942 1261 972
rect 185 267 213 297
<< poly >>
rect 105 903 155 916
rect 318 903 368 916
rect 526 903 576 916
rect 734 903 784 916
rect 1153 899 1203 912
rect 1366 899 1416 912
rect 1574 899 1624 912
rect 1782 899 1832 912
rect 105 775 155 803
rect 105 755 118 775
rect 138 755 155 775
rect 105 726 155 755
rect 318 774 368 803
rect 318 750 329 774
rect 353 750 368 774
rect 318 726 368 750
rect 526 779 576 803
rect 526 755 538 779
rect 562 755 576 779
rect 526 726 576 755
rect 734 777 784 803
rect 734 751 752 777
rect 778 751 784 777
rect 734 726 784 751
rect 1153 771 1203 799
rect 1153 751 1166 771
rect 1186 751 1203 771
rect 1153 722 1203 751
rect 1366 770 1416 799
rect 1366 746 1377 770
rect 1401 746 1416 770
rect 1366 722 1416 746
rect 1574 775 1624 799
rect 1574 751 1586 775
rect 1610 751 1624 775
rect 1574 722 1624 751
rect 1782 773 1832 799
rect 1782 747 1800 773
rect 1826 747 1832 773
rect 1782 722 1832 747
rect 105 668 155 684
rect 318 668 368 684
rect 526 668 576 684
rect 734 668 784 684
rect 1153 664 1203 680
rect 1366 664 1416 680
rect 1574 664 1624 680
rect 1782 664 1832 680
rect 105 224 155 237
rect 318 224 368 237
rect 526 224 576 237
rect 734 224 784 237
rect 105 96 155 124
rect 105 76 118 96
rect 138 76 155 96
rect 105 47 155 76
rect 318 95 368 124
rect 318 71 329 95
rect 353 71 368 95
rect 318 47 368 71
rect 526 100 576 124
rect 526 76 538 100
rect 562 76 576 100
rect 526 47 576 76
rect 734 98 784 124
rect 734 72 752 98
rect 778 72 784 98
rect 734 47 784 72
rect 105 -11 155 5
rect 318 -11 368 5
rect 526 -11 576 5
rect 734 -11 784 5
<< polycont >>
rect 118 755 138 775
rect 329 750 353 774
rect 538 755 562 779
rect 752 751 778 777
rect 1166 751 1186 771
rect 1377 746 1401 770
rect 1586 751 1610 775
rect 1800 747 1826 773
rect 118 76 138 96
rect 329 71 353 95
rect 538 76 562 100
rect 752 72 778 98
<< ndiffres >>
rect -274 1037 -217 1056
rect -274 1034 -253 1037
rect -368 1019 -253 1034
rect -235 1019 -217 1037
rect -368 996 -217 1019
rect -368 960 -326 996
rect -369 959 -269 960
rect -369 938 -213 959
rect -369 920 -251 938
rect -233 920 -213 938
rect -369 916 -213 920
rect -274 900 -213 916
rect -274 781 -217 800
rect -274 778 -253 781
rect -368 763 -253 778
rect -235 763 -217 781
rect -368 740 -217 763
rect -368 704 -326 740
rect -369 703 -269 704
rect -369 682 -213 703
rect -369 664 -251 682
rect -233 664 -213 682
rect -369 660 -213 664
rect -274 644 -213 660
rect -274 386 -217 405
rect -274 383 -253 386
rect -368 368 -253 383
rect -235 368 -217 386
rect -368 345 -217 368
rect -368 309 -326 345
rect -369 308 -269 309
rect -369 287 -213 308
rect -369 269 -251 287
rect -233 269 -213 287
rect -369 265 -213 269
rect -274 249 -213 265
rect -274 131 -217 150
rect -274 128 -253 131
rect -368 113 -253 128
rect -235 113 -217 131
rect -368 90 -217 113
rect -368 54 -326 90
rect -369 53 -269 54
rect -369 32 -213 53
rect -369 14 -251 32
rect -233 14 -213 32
rect -369 10 -213 14
rect -274 -6 -213 10
<< locali >>
rect -275 1037 -216 1143
rect 1688 1119 1760 1120
rect 638 1118 710 1119
rect 637 1110 736 1118
rect 637 1107 689 1110
rect 637 1072 645 1107
rect 670 1072 689 1107
rect 714 1099 736 1110
rect 1687 1111 1786 1119
rect 1687 1108 1739 1111
rect 714 1098 1581 1099
rect 714 1072 1582 1098
rect 637 1062 1582 1072
rect 637 1060 736 1062
rect -275 1019 -253 1037
rect -235 1019 -216 1037
rect -275 997 -216 1019
rect -8 1033 524 1038
rect -8 1013 878 1033
rect 898 1013 901 1033
rect 1537 1029 1582 1062
rect 1687 1073 1695 1108
rect 1720 1073 1739 1108
rect 1764 1073 1786 1111
rect 1687 1061 1786 1073
rect -8 1009 901 1013
rect -8 962 35 1009
rect 485 1008 901 1009
rect 1533 1009 1926 1029
rect 1946 1009 1949 1029
rect 485 1007 826 1008
rect 142 976 252 990
rect 142 973 185 976
rect 142 968 146 973
rect -20 961 35 962
rect -276 938 35 961
rect -276 920 -251 938
rect -233 926 35 938
rect 64 946 146 968
rect 175 946 185 973
rect 213 949 220 976
rect 249 968 252 976
rect 249 949 314 968
rect 213 946 314 949
rect 64 944 314 946
rect -233 920 -211 926
rect -276 781 -211 920
rect 64 865 101 944
rect 142 931 252 944
rect 216 875 247 876
rect 64 845 73 865
rect 93 845 101 865
rect -276 763 -253 781
rect -235 763 -211 781
rect -276 746 -211 763
rect -56 827 12 840
rect 64 835 101 845
rect 160 865 247 875
rect 160 845 169 865
rect 189 845 247 865
rect 160 836 247 845
rect 160 835 197 836
rect -56 785 -49 827
rect 0 785 12 827
rect -56 782 12 785
rect 216 783 247 836
rect 277 865 314 944
rect 429 875 460 876
rect 277 845 286 865
rect 306 845 314 865
rect 277 835 314 845
rect 373 868 460 875
rect 373 865 434 868
rect 373 845 382 865
rect 402 848 434 865
rect 455 848 460 868
rect 402 845 460 848
rect 373 838 460 845
rect 485 865 522 1007
rect 788 1006 825 1007
rect 1533 1004 1949 1009
rect 1533 1003 1874 1004
rect 1190 972 1300 986
rect 1190 969 1233 972
rect 1190 964 1194 969
rect 1112 942 1194 964
rect 1223 942 1233 969
rect 1261 945 1268 972
rect 1297 964 1300 972
rect 1297 945 1362 964
rect 1261 942 1362 945
rect 1112 940 1362 942
rect 637 875 673 876
rect 485 845 494 865
rect 514 845 522 865
rect 373 836 429 838
rect 373 835 410 836
rect 485 835 522 845
rect 581 865 729 875
rect 829 872 925 874
rect 581 845 590 865
rect 610 845 700 865
rect 720 845 729 865
rect 581 839 729 845
rect 581 836 645 839
rect 581 835 618 836
rect 637 809 645 836
rect 666 836 729 839
rect 787 865 925 872
rect 787 845 796 865
rect 816 845 925 865
rect 787 836 925 845
rect 1112 861 1149 940
rect 1190 927 1300 940
rect 1264 871 1295 872
rect 1112 841 1121 861
rect 1141 841 1149 861
rect 666 809 673 836
rect 692 835 729 836
rect 788 835 825 836
rect 637 784 673 809
rect 108 782 149 783
rect -56 775 149 782
rect -56 764 118 775
rect -56 731 -48 764
rect -55 722 -48 731
rect 1 755 118 764
rect 138 755 149 775
rect 1 747 149 755
rect 216 779 575 783
rect 216 774 538 779
rect 216 750 329 774
rect 353 755 538 774
rect 562 755 575 779
rect 353 750 575 755
rect 216 747 575 750
rect 637 747 672 784
rect 740 781 840 784
rect 740 777 807 781
rect 740 751 752 777
rect 778 755 807 777
rect 833 755 840 781
rect 778 751 840 755
rect 740 747 840 751
rect 1 731 12 747
rect 1 722 9 731
rect 216 726 247 747
rect 637 726 673 747
rect 59 725 96 726
rect -276 682 -211 701
rect -276 664 -251 682
rect -233 664 -211 682
rect -276 463 -211 664
rect -55 538 9 722
rect 58 716 96 725
rect 58 696 67 716
rect 87 696 96 716
rect 58 688 96 696
rect 162 720 247 726
rect 272 725 309 726
rect 162 700 170 720
rect 190 700 247 720
rect 162 692 247 700
rect 271 716 309 725
rect 271 696 280 716
rect 300 696 309 716
rect 162 691 198 692
rect 271 688 309 696
rect 375 720 460 726
rect 480 725 517 726
rect 375 700 383 720
rect 403 719 460 720
rect 403 700 432 719
rect 375 699 432 700
rect 453 699 460 719
rect 375 692 460 699
rect 479 716 517 725
rect 479 696 488 716
rect 508 696 517 716
rect 375 691 411 692
rect 479 688 517 696
rect 583 720 727 726
rect 583 700 591 720
rect 611 700 699 720
rect 719 700 727 720
rect 583 692 727 700
rect 583 691 619 692
rect 691 691 727 692
rect 793 725 830 726
rect 793 724 831 725
rect 793 716 857 724
rect 793 696 802 716
rect 822 702 857 716
rect 877 702 880 722
rect 822 697 880 702
rect 822 696 857 697
rect 59 659 96 688
rect 60 657 96 659
rect 272 657 309 688
rect 60 635 309 657
rect 141 629 252 635
rect 141 621 182 629
rect 141 601 149 621
rect 168 601 182 621
rect 141 599 182 601
rect 210 621 252 629
rect 210 601 226 621
rect 245 601 252 621
rect 210 599 252 601
rect 141 584 252 599
rect -55 528 13 538
rect -55 495 -38 528
rect 2 495 13 528
rect -55 483 13 495
rect -55 481 9 483
rect 480 464 517 688
rect 793 684 857 696
rect 897 466 924 836
rect 1112 831 1149 841
rect 1208 861 1295 871
rect 1208 841 1217 861
rect 1237 841 1295 861
rect 1208 832 1295 841
rect 1208 831 1245 832
rect 988 818 1058 823
rect 983 812 1058 818
rect 983 779 991 812
rect 1044 779 1058 812
rect 1264 779 1295 832
rect 1325 861 1362 940
rect 1477 871 1508 872
rect 1325 841 1334 861
rect 1354 841 1362 861
rect 1325 831 1362 841
rect 1421 864 1508 871
rect 1421 861 1482 864
rect 1421 841 1430 861
rect 1450 844 1482 861
rect 1503 844 1508 864
rect 1450 841 1508 844
rect 1421 834 1508 841
rect 1533 861 1570 1003
rect 1836 1002 1873 1003
rect 1685 871 1721 872
rect 1533 841 1542 861
rect 1562 841 1570 861
rect 1421 832 1477 834
rect 1421 831 1458 832
rect 1533 831 1570 841
rect 1629 861 1777 871
rect 1877 868 1973 870
rect 1629 841 1638 861
rect 1658 841 1748 861
rect 1768 841 1777 861
rect 1629 835 1777 841
rect 1629 832 1693 835
rect 1629 831 1666 832
rect 1685 805 1693 832
rect 1714 832 1777 835
rect 1835 861 1973 868
rect 1835 841 1844 861
rect 1864 841 1973 861
rect 1835 832 1973 841
rect 1714 805 1721 832
rect 1740 831 1777 832
rect 1836 831 1873 832
rect 1685 780 1721 805
rect 983 778 1066 779
rect 1156 778 1197 779
rect 983 771 1197 778
rect 983 754 1166 771
rect 983 721 996 754
rect 1049 751 1166 754
rect 1186 751 1197 771
rect 1049 743 1197 751
rect 1264 775 1623 779
rect 1264 770 1586 775
rect 1264 746 1377 770
rect 1401 751 1586 770
rect 1610 751 1623 775
rect 1401 746 1623 751
rect 1264 743 1623 746
rect 1685 743 1720 780
rect 1788 777 1888 780
rect 1788 773 1855 777
rect 1788 747 1800 773
rect 1826 751 1855 773
rect 1881 751 1888 777
rect 1826 747 1888 751
rect 1788 743 1888 747
rect 1049 721 1066 743
rect 1264 722 1295 743
rect 1685 722 1721 743
rect 1107 721 1144 722
rect 983 707 1066 721
rect 756 464 924 466
rect 480 463 924 464
rect -276 433 924 463
rect 994 497 1066 707
rect 1106 712 1144 721
rect 1106 692 1115 712
rect 1135 692 1144 712
rect 1106 684 1144 692
rect 1210 716 1295 722
rect 1320 721 1357 722
rect 1210 696 1218 716
rect 1238 696 1295 716
rect 1210 688 1295 696
rect 1319 712 1357 721
rect 1319 692 1328 712
rect 1348 692 1357 712
rect 1210 687 1246 688
rect 1319 684 1357 692
rect 1423 716 1508 722
rect 1528 721 1565 722
rect 1423 696 1431 716
rect 1451 715 1508 716
rect 1451 696 1480 715
rect 1423 695 1480 696
rect 1501 695 1508 715
rect 1423 688 1508 695
rect 1527 712 1565 721
rect 1527 692 1536 712
rect 1556 692 1565 712
rect 1423 687 1459 688
rect 1527 684 1565 692
rect 1631 716 1775 722
rect 1631 696 1639 716
rect 1659 696 1747 716
rect 1767 696 1775 716
rect 1631 688 1775 696
rect 1631 687 1667 688
rect 1739 687 1775 688
rect 1841 721 1878 722
rect 1841 720 1879 721
rect 1841 712 1905 720
rect 1841 692 1850 712
rect 1870 698 1905 712
rect 1925 698 1928 718
rect 1870 693 1928 698
rect 1870 692 1905 693
rect 1107 655 1144 684
rect 1108 653 1144 655
rect 1320 653 1357 684
rect 1108 631 1357 653
rect 1189 625 1300 631
rect 1189 617 1230 625
rect 1189 597 1197 617
rect 1216 597 1230 617
rect 1189 595 1230 597
rect 1258 617 1300 625
rect 1258 597 1274 617
rect 1293 597 1300 617
rect 1258 595 1300 597
rect 1189 580 1300 595
rect 994 458 1013 497
rect 1058 458 1066 497
rect 994 441 1066 458
rect 1528 485 1565 684
rect 1841 680 1905 692
rect 1528 479 1569 485
rect 1945 481 1972 832
rect 1804 479 1972 481
rect 1528 453 1972 479
rect -276 386 -211 433
rect -276 368 -253 386
rect -235 368 -211 386
rect 637 413 672 415
rect 637 411 741 413
rect 1530 411 1569 453
rect 1804 452 1972 453
rect 637 404 1571 411
rect 637 403 688 404
rect 637 383 640 403
rect 665 384 688 403
rect 720 384 1571 404
rect 665 383 1571 384
rect 637 376 1571 383
rect 910 375 1571 376
rect -276 347 -211 368
rect 1 358 41 361
rect 1 354 904 358
rect 1 334 878 354
rect 898 334 904 354
rect 1 331 904 334
rect -275 287 -210 307
rect -275 269 -251 287
rect -233 269 -210 287
rect -275 242 -210 269
rect 1 242 41 331
rect 485 329 901 331
rect 485 328 826 329
rect 142 297 252 311
rect 142 294 185 297
rect 142 289 146 294
rect -276 207 41 242
rect 64 267 146 289
rect 175 267 185 294
rect 213 270 220 297
rect 249 289 252 297
rect 249 270 314 289
rect 213 267 314 270
rect 64 265 314 267
rect -275 131 -210 207
rect 64 186 101 265
rect 142 252 252 265
rect 216 196 247 197
rect 64 166 73 186
rect 93 166 101 186
rect 64 156 101 166
rect 160 186 247 196
rect 160 166 169 186
rect 189 166 247 186
rect 160 157 247 166
rect 160 156 197 157
rect -275 113 -253 131
rect -235 113 -210 131
rect -275 92 -210 113
rect -62 111 3 120
rect -62 74 -52 111
rect -12 103 3 111
rect 216 104 247 157
rect 277 186 314 265
rect 429 196 460 197
rect 277 166 286 186
rect 306 166 314 186
rect 277 156 314 166
rect 373 189 460 196
rect 373 186 434 189
rect 373 166 382 186
rect 402 169 434 186
rect 455 169 460 189
rect 402 166 460 169
rect 373 159 460 166
rect 485 186 522 328
rect 788 327 825 328
rect 637 196 673 197
rect 485 166 494 186
rect 514 166 522 186
rect 373 157 429 159
rect 373 156 410 157
rect 485 156 522 166
rect 581 186 729 196
rect 829 193 925 195
rect 581 166 590 186
rect 610 166 700 186
rect 720 166 729 186
rect 581 160 729 166
rect 581 157 645 160
rect 581 156 618 157
rect 637 130 645 157
rect 666 157 729 160
rect 787 186 925 193
rect 787 166 796 186
rect 816 166 925 186
rect 787 157 925 166
rect 666 130 673 157
rect 692 156 729 157
rect 788 156 825 157
rect 637 105 673 130
rect 108 103 149 104
rect -12 96 149 103
rect -12 76 118 96
rect 138 76 149 96
rect -12 74 149 76
rect -62 68 149 74
rect 216 100 575 104
rect 216 95 538 100
rect 216 71 329 95
rect 353 76 538 95
rect 562 76 575 100
rect 353 71 575 76
rect 216 68 575 71
rect 637 68 672 105
rect 740 102 840 105
rect 740 98 807 102
rect 740 72 752 98
rect 778 76 807 98
rect 833 76 840 102
rect 778 72 840 76
rect 740 68 840 72
rect -62 55 5 68
rect -270 32 -214 52
rect -270 14 -251 32
rect -233 14 -214 32
rect -270 -99 -214 14
rect -62 34 -48 55
rect -12 34 5 55
rect 216 47 247 68
rect 637 47 673 68
rect 59 46 96 47
rect -62 27 5 34
rect 58 37 96 46
rect -270 -240 -215 -99
rect -62 -125 3 27
rect 58 17 67 37
rect 87 17 96 37
rect 58 9 96 17
rect 162 41 247 47
rect 272 46 309 47
rect 162 21 170 41
rect 190 21 247 41
rect 162 13 247 21
rect 271 37 309 46
rect 271 17 280 37
rect 300 17 309 37
rect 162 12 198 13
rect 271 9 309 17
rect 375 41 460 47
rect 480 46 517 47
rect 375 21 383 41
rect 403 40 460 41
rect 403 21 432 40
rect 375 20 432 21
rect 453 20 460 40
rect 375 13 460 20
rect 479 37 517 46
rect 479 17 488 37
rect 508 17 517 37
rect 375 12 411 13
rect 479 9 517 17
rect 583 41 727 47
rect 583 21 591 41
rect 611 21 699 41
rect 719 21 727 41
rect 583 13 727 21
rect 583 12 619 13
rect 691 12 727 13
rect 793 46 830 47
rect 793 45 831 46
rect 793 37 857 45
rect 793 17 802 37
rect 822 23 857 37
rect 877 23 880 43
rect 822 18 880 23
rect 822 17 857 18
rect 59 -20 96 9
rect 60 -22 96 -20
rect 272 -22 309 9
rect 60 -44 309 -22
rect 141 -50 252 -44
rect 141 -58 182 -50
rect 141 -78 149 -58
rect 168 -78 182 -58
rect 141 -80 182 -78
rect 210 -58 252 -50
rect 210 -78 226 -58
rect 245 -78 252 -58
rect 210 -80 252 -78
rect 141 -95 252 -80
rect 480 -90 517 9
rect 793 5 857 17
rect -69 -135 52 -125
rect -69 -137 0 -135
rect -69 -178 -56 -137
rect -19 -176 0 -137
rect 37 -176 52 -135
rect -19 -178 52 -176
rect -69 -196 52 -178
rect 143 -240 247 -95
rect 478 -240 519 -90
rect 897 -98 924 157
rect 986 147 1066 158
rect 986 121 1003 147
rect 1043 121 1066 147
rect 986 94 1066 121
rect 986 68 1007 94
rect 1047 68 1066 94
rect 986 49 1066 68
rect 986 23 1010 49
rect 1050 23 1066 49
rect 986 -28 1066 23
rect -270 -243 519 -240
rect 898 -229 924 -98
rect 898 -243 926 -229
rect -270 -276 926 -243
rect -268 -278 926 -276
rect 143 -280 247 -278
rect 478 -280 519 -278
rect 988 -281 1058 -28
<< viali >>
rect 645 1072 670 1107
rect 689 1072 714 1110
rect 878 1013 898 1033
rect 1695 1073 1720 1108
rect 1739 1073 1764 1111
rect 1926 1009 1946 1029
rect 146 946 175 973
rect 220 949 249 976
rect -49 785 0 827
rect 434 848 455 868
rect 1194 942 1223 969
rect 1268 945 1297 972
rect 645 809 666 839
rect -48 722 1 764
rect 807 755 833 781
rect 432 699 453 719
rect 857 702 877 722
rect 149 601 168 621
rect 226 601 245 621
rect -38 495 2 528
rect 991 779 1044 812
rect 1482 844 1503 864
rect 1693 805 1714 835
rect 996 721 1049 754
rect 1855 751 1881 777
rect 1480 695 1501 715
rect 1905 698 1925 718
rect 1197 597 1216 617
rect 1274 597 1293 617
rect 1013 458 1058 497
rect 640 383 665 403
rect 688 384 720 404
rect 878 334 898 354
rect 146 267 175 294
rect 220 270 249 297
rect -52 74 -12 111
rect 434 169 455 189
rect 645 130 666 160
rect 807 76 833 102
rect -48 34 -12 55
rect 432 20 453 40
rect 857 23 877 43
rect 149 -78 168 -58
rect 226 -78 245 -58
rect -56 -178 -19 -137
rect 0 -176 37 -135
rect 1003 121 1043 147
rect 1007 68 1047 94
rect 1010 23 1050 49
<< metal1 >>
rect -537 639 -430 1152
rect -58 827 14 1143
rect 638 1118 710 1119
rect 637 1110 736 1118
rect 637 1107 689 1110
rect 637 1072 645 1107
rect 670 1072 689 1107
rect 714 1072 736 1110
rect 637 1060 736 1072
rect 638 1041 706 1060
rect 639 1038 672 1041
rect 874 1038 906 1039
rect 49 977 252 990
rect 49 944 73 977
rect 109 976 252 977
rect 109 973 220 976
rect 109 946 146 973
rect 175 949 220 973
rect 249 949 252 976
rect 175 946 252 949
rect 109 944 252 946
rect 49 931 252 944
rect 49 930 150 931
rect -58 785 -49 827
rect 0 785 14 827
rect -58 764 14 785
rect -58 722 -48 764
rect 1 722 14 764
rect -58 704 14 722
rect 427 868 459 875
rect 427 848 434 868
rect 455 848 459 868
rect 427 783 459 848
rect 639 839 670 1038
rect 871 1033 906 1038
rect 871 1013 878 1033
rect 898 1013 906 1033
rect 871 1005 906 1013
rect 639 809 645 839
rect 666 809 670 839
rect 639 801 670 809
rect 797 783 837 784
rect 427 781 839 783
rect 427 755 807 781
rect 833 755 839 781
rect 427 747 839 755
rect 427 719 459 747
rect 872 727 906 1005
rect 988 818 1058 1191
rect 1688 1119 1760 1120
rect 1687 1111 1786 1119
rect 1687 1108 1739 1111
rect 1687 1073 1695 1108
rect 1720 1073 1739 1108
rect 1764 1073 1786 1111
rect 1687 1061 1786 1073
rect 1687 1060 1756 1061
rect 1687 1042 1723 1060
rect 1097 973 1300 986
rect 1097 940 1121 973
rect 1157 972 1300 973
rect 1157 969 1268 972
rect 1157 942 1194 969
rect 1223 945 1268 969
rect 1297 945 1300 972
rect 1223 942 1300 945
rect 1157 940 1300 942
rect 1097 927 1300 940
rect 1097 926 1198 927
rect 427 699 432 719
rect 453 699 459 719
rect 427 692 459 699
rect 850 722 906 727
rect 850 702 857 722
rect 877 702 906 722
rect 983 812 1058 818
rect 983 779 991 812
rect 1044 779 1058 812
rect 983 754 1058 779
rect 983 721 996 754
rect 1049 721 1058 754
rect 983 712 1058 721
rect 1475 864 1507 871
rect 1475 844 1482 864
rect 1503 844 1507 864
rect 1475 779 1507 844
rect 1687 835 1718 1042
rect 1922 1034 1954 1035
rect 1919 1029 1954 1034
rect 1919 1009 1926 1029
rect 1946 1009 1954 1029
rect 1919 1001 1954 1009
rect 1687 805 1693 835
rect 1714 805 1718 835
rect 1687 797 1718 805
rect 1845 779 1885 780
rect 1475 777 1887 779
rect 1475 751 1855 777
rect 1881 751 1887 777
rect 1475 743 1887 751
rect 1475 715 1507 743
rect 1920 723 1954 1001
rect 983 707 1041 712
rect 850 695 906 702
rect 1475 695 1480 715
rect 1501 695 1507 715
rect 850 694 885 695
rect 1475 688 1507 695
rect 1898 718 1954 723
rect 1898 698 1905 718
rect 1925 698 1954 718
rect 1898 691 1954 698
rect 1898 690 1933 691
rect 141 639 252 643
rect -537 621 2139 639
rect -537 601 149 621
rect 168 601 226 621
rect 245 617 2139 621
rect 245 601 1197 617
rect -537 597 1197 601
rect 1216 597 1274 617
rect 1293 597 2139 617
rect -537 583 2139 597
rect -537 -40 -430 583
rect 1189 580 1300 583
rect -51 534 13 538
rect -55 528 13 534
rect -55 495 -38 528
rect 2 495 13 528
rect -55 483 13 495
rect 996 497 1061 519
rect -55 481 2 483
rect -51 120 0 481
rect 996 458 1013 497
rect 1058 458 1061 497
rect 637 413 672 415
rect 637 404 741 413
rect 637 403 688 404
rect 637 383 640 403
rect 665 384 688 403
rect 720 384 741 404
rect 665 383 741 384
rect 637 376 741 383
rect 637 364 672 376
rect 49 298 252 311
rect 49 265 73 298
rect 109 297 252 298
rect 109 294 220 297
rect 109 267 146 294
rect 175 270 220 294
rect 249 270 252 297
rect 175 267 252 270
rect 109 265 252 267
rect 49 252 252 265
rect 49 251 150 252
rect 427 189 459 196
rect 427 169 434 189
rect 455 169 459 189
rect -62 111 3 120
rect -62 74 -52 111
rect -12 77 3 111
rect 427 104 459 169
rect 639 160 670 364
rect 874 359 906 360
rect 871 354 906 359
rect 871 334 878 354
rect 898 334 906 354
rect 871 326 906 334
rect 639 130 645 160
rect 666 130 670 160
rect 639 122 670 130
rect 797 104 837 105
rect 427 102 839 104
rect -12 74 5 77
rect -62 55 5 74
rect -62 34 -48 55
rect -12 34 5 55
rect -62 27 5 34
rect 427 76 807 102
rect 833 76 839 102
rect 427 68 839 76
rect 427 40 459 68
rect 872 48 906 326
rect 996 158 1061 458
rect 427 20 432 40
rect 453 20 459 40
rect 427 13 459 20
rect 850 43 906 48
rect 850 23 857 43
rect 877 23 906 43
rect 850 16 906 23
rect 986 147 1066 158
rect 986 121 1003 147
rect 1043 121 1066 147
rect 986 94 1066 121
rect 986 68 1007 94
rect 1047 68 1066 94
rect 986 49 1066 68
rect 986 23 1010 49
rect 1050 23 1066 49
rect 850 15 885 16
rect 986 11 1066 23
rect 141 -40 252 -36
rect 1896 -40 2131 -39
rect -539 -58 2131 -40
rect -539 -78 149 -58
rect 168 -78 226 -58
rect 245 -78 2131 -58
rect -539 -96 2131 -78
rect -537 -296 -430 -96
rect -69 -135 52 -125
rect -69 -137 0 -135
rect -69 -178 -56 -137
rect -19 -176 0 -137
rect 37 -176 52 -135
rect -19 -178 52 -176
rect -69 -196 52 -178
rect -63 -334 2 -196
<< via1 >>
rect 73 944 109 977
rect 1121 940 1157 973
rect 73 265 109 298
<< metal2 >>
rect -708 992 -601 1149
rect -708 977 2171 992
rect -708 944 73 977
rect 109 973 2171 977
rect 109 944 1121 973
rect -708 940 1121 944
rect 1157 940 2171 973
rect -708 923 2171 940
rect -708 317 -601 923
rect -708 298 2179 317
rect -708 265 73 298
rect 109 265 2179 298
rect -708 248 2179 265
rect -708 -298 -601 248
<< labels >>
rlabel metal1 1778 1070 1786 1110 1 vout
rlabel locali -265 1100 -221 1122 1 vref
rlabel metal1 -529 1089 -433 1122 1 gnd
rlabel metal2 -705 1089 -609 1122 1 vdd
rlabel metal1 -50 1104 12 1131 1 d0
rlabel metal1 996 1133 1049 1155 1 d1
<< end >>
