* SPICE3 file created from resfinal.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a b SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81


V1 a 0 dc 1.8
V2 b 0 0 

.tran 0.1n 10ns

.control
*op line 0 3.3
run
plot V(a)/V1#branch

.endc

.end

