magic
tech sky130A
timestamp 1616159323
<< nwell >>
rect 278 3552 1089 3702
rect 1290 3371 2101 3521
rect 277 3137 1088 3287
rect 1345 2810 2156 2960
rect 283 2571 1094 2721
rect 1295 2390 2106 2540
rect 282 2156 1093 2306
rect 1510 1878 2321 2028
rect 290 1592 1101 1742
rect 1302 1411 2113 1561
rect 289 1177 1100 1327
rect 1357 850 2168 1000
rect 295 611 1106 761
rect 1307 430 2118 580
rect 294 196 1105 346
rect 1605 -114 2416 36
rect 298 -365 1109 -215
rect 1310 -546 2121 -396
rect 297 -780 1108 -630
rect 1365 -1107 2176 -957
rect 303 -1346 1114 -1196
rect 1315 -1527 2126 -1377
rect 302 -1761 1113 -1611
rect 1530 -2039 2341 -1889
rect 310 -2325 1121 -2175
rect 1322 -2506 2133 -2356
rect 309 -2740 1120 -2590
rect 1377 -3067 2188 -2917
rect 315 -3306 1126 -3156
rect 1327 -3487 2138 -3337
rect 314 -3721 1125 -3571
<< nmos >>
rect 342 3451 392 3493
rect 555 3451 605 3493
rect 763 3451 813 3493
rect 971 3451 1021 3493
rect 1354 3270 1404 3312
rect 1567 3270 1617 3312
rect 1775 3270 1825 3312
rect 1983 3270 2033 3312
rect 341 3036 391 3078
rect 554 3036 604 3078
rect 762 3036 812 3078
rect 970 3036 1020 3078
rect 1409 2709 1459 2751
rect 1622 2709 1672 2751
rect 1830 2709 1880 2751
rect 2038 2709 2088 2751
rect 347 2470 397 2512
rect 560 2470 610 2512
rect 768 2470 818 2512
rect 976 2470 1026 2512
rect 1359 2289 1409 2331
rect 1572 2289 1622 2331
rect 1780 2289 1830 2331
rect 1988 2289 2038 2331
rect 346 2055 396 2097
rect 559 2055 609 2097
rect 767 2055 817 2097
rect 975 2055 1025 2097
rect 1574 1777 1624 1819
rect 1787 1777 1837 1819
rect 1995 1777 2045 1819
rect 2203 1777 2253 1819
rect 354 1491 404 1533
rect 567 1491 617 1533
rect 775 1491 825 1533
rect 983 1491 1033 1533
rect 1366 1310 1416 1352
rect 1579 1310 1629 1352
rect 1787 1310 1837 1352
rect 1995 1310 2045 1352
rect 353 1076 403 1118
rect 566 1076 616 1118
rect 774 1076 824 1118
rect 982 1076 1032 1118
rect 1421 749 1471 791
rect 1634 749 1684 791
rect 1842 749 1892 791
rect 2050 749 2100 791
rect 359 510 409 552
rect 572 510 622 552
rect 780 510 830 552
rect 988 510 1038 552
rect 1371 329 1421 371
rect 1584 329 1634 371
rect 1792 329 1842 371
rect 2000 329 2050 371
rect 358 95 408 137
rect 571 95 621 137
rect 779 95 829 137
rect 987 95 1037 137
rect 1669 -215 1719 -173
rect 1882 -215 1932 -173
rect 2090 -215 2140 -173
rect 2298 -215 2348 -173
rect 362 -466 412 -424
rect 575 -466 625 -424
rect 783 -466 833 -424
rect 991 -466 1041 -424
rect 1374 -647 1424 -605
rect 1587 -647 1637 -605
rect 1795 -647 1845 -605
rect 2003 -647 2053 -605
rect 361 -881 411 -839
rect 574 -881 624 -839
rect 782 -881 832 -839
rect 990 -881 1040 -839
rect 1429 -1208 1479 -1166
rect 1642 -1208 1692 -1166
rect 1850 -1208 1900 -1166
rect 2058 -1208 2108 -1166
rect 367 -1447 417 -1405
rect 580 -1447 630 -1405
rect 788 -1447 838 -1405
rect 996 -1447 1046 -1405
rect 1379 -1628 1429 -1586
rect 1592 -1628 1642 -1586
rect 1800 -1628 1850 -1586
rect 2008 -1628 2058 -1586
rect 366 -1862 416 -1820
rect 579 -1862 629 -1820
rect 787 -1862 837 -1820
rect 995 -1862 1045 -1820
rect 1594 -2140 1644 -2098
rect 1807 -2140 1857 -2098
rect 2015 -2140 2065 -2098
rect 2223 -2140 2273 -2098
rect 374 -2426 424 -2384
rect 587 -2426 637 -2384
rect 795 -2426 845 -2384
rect 1003 -2426 1053 -2384
rect 1386 -2607 1436 -2565
rect 1599 -2607 1649 -2565
rect 1807 -2607 1857 -2565
rect 2015 -2607 2065 -2565
rect 373 -2841 423 -2799
rect 586 -2841 636 -2799
rect 794 -2841 844 -2799
rect 1002 -2841 1052 -2799
rect 1441 -3168 1491 -3126
rect 1654 -3168 1704 -3126
rect 1862 -3168 1912 -3126
rect 2070 -3168 2120 -3126
rect 379 -3407 429 -3365
rect 592 -3407 642 -3365
rect 800 -3407 850 -3365
rect 1008 -3407 1058 -3365
rect 1391 -3588 1441 -3546
rect 1604 -3588 1654 -3546
rect 1812 -3588 1862 -3546
rect 2020 -3588 2070 -3546
rect 378 -3822 428 -3780
rect 591 -3822 641 -3780
rect 799 -3822 849 -3780
rect 1007 -3822 1057 -3780
<< pmos >>
rect 342 3570 392 3670
rect 555 3570 605 3670
rect 763 3570 813 3670
rect 971 3570 1021 3670
rect 1354 3389 1404 3489
rect 1567 3389 1617 3489
rect 1775 3389 1825 3489
rect 1983 3389 2033 3489
rect 341 3155 391 3255
rect 554 3155 604 3255
rect 762 3155 812 3255
rect 970 3155 1020 3255
rect 1409 2828 1459 2928
rect 1622 2828 1672 2928
rect 1830 2828 1880 2928
rect 2038 2828 2088 2928
rect 347 2589 397 2689
rect 560 2589 610 2689
rect 768 2589 818 2689
rect 976 2589 1026 2689
rect 1359 2408 1409 2508
rect 1572 2408 1622 2508
rect 1780 2408 1830 2508
rect 1988 2408 2038 2508
rect 346 2174 396 2274
rect 559 2174 609 2274
rect 767 2174 817 2274
rect 975 2174 1025 2274
rect 1574 1896 1624 1996
rect 1787 1896 1837 1996
rect 1995 1896 2045 1996
rect 2203 1896 2253 1996
rect 354 1610 404 1710
rect 567 1610 617 1710
rect 775 1610 825 1710
rect 983 1610 1033 1710
rect 1366 1429 1416 1529
rect 1579 1429 1629 1529
rect 1787 1429 1837 1529
rect 1995 1429 2045 1529
rect 353 1195 403 1295
rect 566 1195 616 1295
rect 774 1195 824 1295
rect 982 1195 1032 1295
rect 1421 868 1471 968
rect 1634 868 1684 968
rect 1842 868 1892 968
rect 2050 868 2100 968
rect 359 629 409 729
rect 572 629 622 729
rect 780 629 830 729
rect 988 629 1038 729
rect 1371 448 1421 548
rect 1584 448 1634 548
rect 1792 448 1842 548
rect 2000 448 2050 548
rect 358 214 408 314
rect 571 214 621 314
rect 779 214 829 314
rect 987 214 1037 314
rect 1669 -96 1719 4
rect 1882 -96 1932 4
rect 2090 -96 2140 4
rect 2298 -96 2348 4
rect 362 -347 412 -247
rect 575 -347 625 -247
rect 783 -347 833 -247
rect 991 -347 1041 -247
rect 1374 -528 1424 -428
rect 1587 -528 1637 -428
rect 1795 -528 1845 -428
rect 2003 -528 2053 -428
rect 361 -762 411 -662
rect 574 -762 624 -662
rect 782 -762 832 -662
rect 990 -762 1040 -662
rect 1429 -1089 1479 -989
rect 1642 -1089 1692 -989
rect 1850 -1089 1900 -989
rect 2058 -1089 2108 -989
rect 367 -1328 417 -1228
rect 580 -1328 630 -1228
rect 788 -1328 838 -1228
rect 996 -1328 1046 -1228
rect 1379 -1509 1429 -1409
rect 1592 -1509 1642 -1409
rect 1800 -1509 1850 -1409
rect 2008 -1509 2058 -1409
rect 366 -1743 416 -1643
rect 579 -1743 629 -1643
rect 787 -1743 837 -1643
rect 995 -1743 1045 -1643
rect 1594 -2021 1644 -1921
rect 1807 -2021 1857 -1921
rect 2015 -2021 2065 -1921
rect 2223 -2021 2273 -1921
rect 374 -2307 424 -2207
rect 587 -2307 637 -2207
rect 795 -2307 845 -2207
rect 1003 -2307 1053 -2207
rect 1386 -2488 1436 -2388
rect 1599 -2488 1649 -2388
rect 1807 -2488 1857 -2388
rect 2015 -2488 2065 -2388
rect 373 -2722 423 -2622
rect 586 -2722 636 -2622
rect 794 -2722 844 -2622
rect 1002 -2722 1052 -2622
rect 1441 -3049 1491 -2949
rect 1654 -3049 1704 -2949
rect 1862 -3049 1912 -2949
rect 2070 -3049 2120 -2949
rect 379 -3288 429 -3188
rect 592 -3288 642 -3188
rect 800 -3288 850 -3188
rect 1008 -3288 1058 -3188
rect 1391 -3469 1441 -3369
rect 1604 -3469 1654 -3369
rect 1812 -3469 1862 -3369
rect 2020 -3469 2070 -3369
rect 378 -3703 428 -3603
rect 591 -3703 641 -3603
rect 799 -3703 849 -3603
rect 1007 -3703 1057 -3603
<< ndiff >>
rect 293 3483 342 3493
rect 293 3463 304 3483
rect 324 3463 342 3483
rect 293 3451 342 3463
rect 392 3487 436 3493
rect 392 3467 407 3487
rect 427 3467 436 3487
rect 392 3451 436 3467
rect 506 3483 555 3493
rect 506 3463 517 3483
rect 537 3463 555 3483
rect 506 3451 555 3463
rect 605 3487 649 3493
rect 605 3467 620 3487
rect 640 3467 649 3487
rect 605 3451 649 3467
rect 714 3483 763 3493
rect 714 3463 725 3483
rect 745 3463 763 3483
rect 714 3451 763 3463
rect 813 3487 857 3493
rect 813 3467 828 3487
rect 848 3467 857 3487
rect 813 3451 857 3467
rect 927 3487 971 3493
rect 927 3467 936 3487
rect 956 3467 971 3487
rect 927 3451 971 3467
rect 1021 3483 1070 3493
rect 1021 3463 1039 3483
rect 1059 3463 1070 3483
rect 1021 3451 1070 3463
rect 1305 3302 1354 3312
rect 1305 3282 1316 3302
rect 1336 3282 1354 3302
rect 1305 3270 1354 3282
rect 1404 3306 1448 3312
rect 1404 3286 1419 3306
rect 1439 3286 1448 3306
rect 1404 3270 1448 3286
rect 1518 3302 1567 3312
rect 1518 3282 1529 3302
rect 1549 3282 1567 3302
rect 1518 3270 1567 3282
rect 1617 3306 1661 3312
rect 1617 3286 1632 3306
rect 1652 3286 1661 3306
rect 1617 3270 1661 3286
rect 1726 3302 1775 3312
rect 1726 3282 1737 3302
rect 1757 3282 1775 3302
rect 1726 3270 1775 3282
rect 1825 3306 1869 3312
rect 1825 3286 1840 3306
rect 1860 3286 1869 3306
rect 1825 3270 1869 3286
rect 1939 3306 1983 3312
rect 1939 3286 1948 3306
rect 1968 3286 1983 3306
rect 1939 3270 1983 3286
rect 2033 3302 2082 3312
rect 2033 3282 2051 3302
rect 2071 3282 2082 3302
rect 2033 3270 2082 3282
rect 292 3068 341 3078
rect 292 3048 303 3068
rect 323 3048 341 3068
rect 292 3036 341 3048
rect 391 3072 435 3078
rect 391 3052 406 3072
rect 426 3052 435 3072
rect 391 3036 435 3052
rect 505 3068 554 3078
rect 505 3048 516 3068
rect 536 3048 554 3068
rect 505 3036 554 3048
rect 604 3072 648 3078
rect 604 3052 619 3072
rect 639 3052 648 3072
rect 604 3036 648 3052
rect 713 3068 762 3078
rect 713 3048 724 3068
rect 744 3048 762 3068
rect 713 3036 762 3048
rect 812 3072 856 3078
rect 812 3052 827 3072
rect 847 3052 856 3072
rect 812 3036 856 3052
rect 926 3072 970 3078
rect 926 3052 935 3072
rect 955 3052 970 3072
rect 926 3036 970 3052
rect 1020 3068 1069 3078
rect 1020 3048 1038 3068
rect 1058 3048 1069 3068
rect 1020 3036 1069 3048
rect 1360 2741 1409 2751
rect 1360 2721 1371 2741
rect 1391 2721 1409 2741
rect 1360 2709 1409 2721
rect 1459 2745 1503 2751
rect 1459 2725 1474 2745
rect 1494 2725 1503 2745
rect 1459 2709 1503 2725
rect 1573 2741 1622 2751
rect 1573 2721 1584 2741
rect 1604 2721 1622 2741
rect 1573 2709 1622 2721
rect 1672 2745 1716 2751
rect 1672 2725 1687 2745
rect 1707 2725 1716 2745
rect 1672 2709 1716 2725
rect 1781 2741 1830 2751
rect 1781 2721 1792 2741
rect 1812 2721 1830 2741
rect 1781 2709 1830 2721
rect 1880 2745 1924 2751
rect 1880 2725 1895 2745
rect 1915 2725 1924 2745
rect 1880 2709 1924 2725
rect 1994 2745 2038 2751
rect 1994 2725 2003 2745
rect 2023 2725 2038 2745
rect 1994 2709 2038 2725
rect 2088 2741 2137 2751
rect 2088 2721 2106 2741
rect 2126 2721 2137 2741
rect 2088 2709 2137 2721
rect 298 2502 347 2512
rect 298 2482 309 2502
rect 329 2482 347 2502
rect 298 2470 347 2482
rect 397 2506 441 2512
rect 397 2486 412 2506
rect 432 2486 441 2506
rect 397 2470 441 2486
rect 511 2502 560 2512
rect 511 2482 522 2502
rect 542 2482 560 2502
rect 511 2470 560 2482
rect 610 2506 654 2512
rect 610 2486 625 2506
rect 645 2486 654 2506
rect 610 2470 654 2486
rect 719 2502 768 2512
rect 719 2482 730 2502
rect 750 2482 768 2502
rect 719 2470 768 2482
rect 818 2506 862 2512
rect 818 2486 833 2506
rect 853 2486 862 2506
rect 818 2470 862 2486
rect 932 2506 976 2512
rect 932 2486 941 2506
rect 961 2486 976 2506
rect 932 2470 976 2486
rect 1026 2502 1075 2512
rect 1026 2482 1044 2502
rect 1064 2482 1075 2502
rect 1026 2470 1075 2482
rect 1310 2321 1359 2331
rect 1310 2301 1321 2321
rect 1341 2301 1359 2321
rect 1310 2289 1359 2301
rect 1409 2325 1453 2331
rect 1409 2305 1424 2325
rect 1444 2305 1453 2325
rect 1409 2289 1453 2305
rect 1523 2321 1572 2331
rect 1523 2301 1534 2321
rect 1554 2301 1572 2321
rect 1523 2289 1572 2301
rect 1622 2325 1666 2331
rect 1622 2305 1637 2325
rect 1657 2305 1666 2325
rect 1622 2289 1666 2305
rect 1731 2321 1780 2331
rect 1731 2301 1742 2321
rect 1762 2301 1780 2321
rect 1731 2289 1780 2301
rect 1830 2325 1874 2331
rect 1830 2305 1845 2325
rect 1865 2305 1874 2325
rect 1830 2289 1874 2305
rect 1944 2325 1988 2331
rect 1944 2305 1953 2325
rect 1973 2305 1988 2325
rect 1944 2289 1988 2305
rect 2038 2321 2087 2331
rect 2038 2301 2056 2321
rect 2076 2301 2087 2321
rect 2038 2289 2087 2301
rect 297 2087 346 2097
rect 297 2067 308 2087
rect 328 2067 346 2087
rect 297 2055 346 2067
rect 396 2091 440 2097
rect 396 2071 411 2091
rect 431 2071 440 2091
rect 396 2055 440 2071
rect 510 2087 559 2097
rect 510 2067 521 2087
rect 541 2067 559 2087
rect 510 2055 559 2067
rect 609 2091 653 2097
rect 609 2071 624 2091
rect 644 2071 653 2091
rect 609 2055 653 2071
rect 718 2087 767 2097
rect 718 2067 729 2087
rect 749 2067 767 2087
rect 718 2055 767 2067
rect 817 2091 861 2097
rect 817 2071 832 2091
rect 852 2071 861 2091
rect 817 2055 861 2071
rect 931 2091 975 2097
rect 931 2071 940 2091
rect 960 2071 975 2091
rect 931 2055 975 2071
rect 1025 2087 1074 2097
rect 1025 2067 1043 2087
rect 1063 2067 1074 2087
rect 1025 2055 1074 2067
rect 1525 1809 1574 1819
rect 1525 1789 1536 1809
rect 1556 1789 1574 1809
rect 1525 1777 1574 1789
rect 1624 1813 1668 1819
rect 1624 1793 1639 1813
rect 1659 1793 1668 1813
rect 1624 1777 1668 1793
rect 1738 1809 1787 1819
rect 1738 1789 1749 1809
rect 1769 1789 1787 1809
rect 1738 1777 1787 1789
rect 1837 1813 1881 1819
rect 1837 1793 1852 1813
rect 1872 1793 1881 1813
rect 1837 1777 1881 1793
rect 1946 1809 1995 1819
rect 1946 1789 1957 1809
rect 1977 1789 1995 1809
rect 1946 1777 1995 1789
rect 2045 1813 2089 1819
rect 2045 1793 2060 1813
rect 2080 1793 2089 1813
rect 2045 1777 2089 1793
rect 2159 1813 2203 1819
rect 2159 1793 2168 1813
rect 2188 1793 2203 1813
rect 2159 1777 2203 1793
rect 2253 1809 2302 1819
rect 2253 1789 2271 1809
rect 2291 1789 2302 1809
rect 2253 1777 2302 1789
rect 305 1523 354 1533
rect 305 1503 316 1523
rect 336 1503 354 1523
rect 305 1491 354 1503
rect 404 1527 448 1533
rect 404 1507 419 1527
rect 439 1507 448 1527
rect 404 1491 448 1507
rect 518 1523 567 1533
rect 518 1503 529 1523
rect 549 1503 567 1523
rect 518 1491 567 1503
rect 617 1527 661 1533
rect 617 1507 632 1527
rect 652 1507 661 1527
rect 617 1491 661 1507
rect 726 1523 775 1533
rect 726 1503 737 1523
rect 757 1503 775 1523
rect 726 1491 775 1503
rect 825 1527 869 1533
rect 825 1507 840 1527
rect 860 1507 869 1527
rect 825 1491 869 1507
rect 939 1527 983 1533
rect 939 1507 948 1527
rect 968 1507 983 1527
rect 939 1491 983 1507
rect 1033 1523 1082 1533
rect 1033 1503 1051 1523
rect 1071 1503 1082 1523
rect 1033 1491 1082 1503
rect 1317 1342 1366 1352
rect 1317 1322 1328 1342
rect 1348 1322 1366 1342
rect 1317 1310 1366 1322
rect 1416 1346 1460 1352
rect 1416 1326 1431 1346
rect 1451 1326 1460 1346
rect 1416 1310 1460 1326
rect 1530 1342 1579 1352
rect 1530 1322 1541 1342
rect 1561 1322 1579 1342
rect 1530 1310 1579 1322
rect 1629 1346 1673 1352
rect 1629 1326 1644 1346
rect 1664 1326 1673 1346
rect 1629 1310 1673 1326
rect 1738 1342 1787 1352
rect 1738 1322 1749 1342
rect 1769 1322 1787 1342
rect 1738 1310 1787 1322
rect 1837 1346 1881 1352
rect 1837 1326 1852 1346
rect 1872 1326 1881 1346
rect 1837 1310 1881 1326
rect 1951 1346 1995 1352
rect 1951 1326 1960 1346
rect 1980 1326 1995 1346
rect 1951 1310 1995 1326
rect 2045 1342 2094 1352
rect 2045 1322 2063 1342
rect 2083 1322 2094 1342
rect 2045 1310 2094 1322
rect 304 1108 353 1118
rect 304 1088 315 1108
rect 335 1088 353 1108
rect 304 1076 353 1088
rect 403 1112 447 1118
rect 403 1092 418 1112
rect 438 1092 447 1112
rect 403 1076 447 1092
rect 517 1108 566 1118
rect 517 1088 528 1108
rect 548 1088 566 1108
rect 517 1076 566 1088
rect 616 1112 660 1118
rect 616 1092 631 1112
rect 651 1092 660 1112
rect 616 1076 660 1092
rect 725 1108 774 1118
rect 725 1088 736 1108
rect 756 1088 774 1108
rect 725 1076 774 1088
rect 824 1112 868 1118
rect 824 1092 839 1112
rect 859 1092 868 1112
rect 824 1076 868 1092
rect 938 1112 982 1118
rect 938 1092 947 1112
rect 967 1092 982 1112
rect 938 1076 982 1092
rect 1032 1108 1081 1118
rect 1032 1088 1050 1108
rect 1070 1088 1081 1108
rect 1032 1076 1081 1088
rect 1372 781 1421 791
rect 1372 761 1383 781
rect 1403 761 1421 781
rect 1372 749 1421 761
rect 1471 785 1515 791
rect 1471 765 1486 785
rect 1506 765 1515 785
rect 1471 749 1515 765
rect 1585 781 1634 791
rect 1585 761 1596 781
rect 1616 761 1634 781
rect 1585 749 1634 761
rect 1684 785 1728 791
rect 1684 765 1699 785
rect 1719 765 1728 785
rect 1684 749 1728 765
rect 1793 781 1842 791
rect 1793 761 1804 781
rect 1824 761 1842 781
rect 1793 749 1842 761
rect 1892 785 1936 791
rect 1892 765 1907 785
rect 1927 765 1936 785
rect 1892 749 1936 765
rect 2006 785 2050 791
rect 2006 765 2015 785
rect 2035 765 2050 785
rect 2006 749 2050 765
rect 2100 781 2149 791
rect 2100 761 2118 781
rect 2138 761 2149 781
rect 2100 749 2149 761
rect 310 542 359 552
rect 310 522 321 542
rect 341 522 359 542
rect 310 510 359 522
rect 409 546 453 552
rect 409 526 424 546
rect 444 526 453 546
rect 409 510 453 526
rect 523 542 572 552
rect 523 522 534 542
rect 554 522 572 542
rect 523 510 572 522
rect 622 546 666 552
rect 622 526 637 546
rect 657 526 666 546
rect 622 510 666 526
rect 731 542 780 552
rect 731 522 742 542
rect 762 522 780 542
rect 731 510 780 522
rect 830 546 874 552
rect 830 526 845 546
rect 865 526 874 546
rect 830 510 874 526
rect 944 546 988 552
rect 944 526 953 546
rect 973 526 988 546
rect 944 510 988 526
rect 1038 542 1087 552
rect 1038 522 1056 542
rect 1076 522 1087 542
rect 1038 510 1087 522
rect 1322 361 1371 371
rect 1322 341 1333 361
rect 1353 341 1371 361
rect 1322 329 1371 341
rect 1421 365 1465 371
rect 1421 345 1436 365
rect 1456 345 1465 365
rect 1421 329 1465 345
rect 1535 361 1584 371
rect 1535 341 1546 361
rect 1566 341 1584 361
rect 1535 329 1584 341
rect 1634 365 1678 371
rect 1634 345 1649 365
rect 1669 345 1678 365
rect 1634 329 1678 345
rect 1743 361 1792 371
rect 1743 341 1754 361
rect 1774 341 1792 361
rect 1743 329 1792 341
rect 1842 365 1886 371
rect 1842 345 1857 365
rect 1877 345 1886 365
rect 1842 329 1886 345
rect 1956 365 2000 371
rect 1956 345 1965 365
rect 1985 345 2000 365
rect 1956 329 2000 345
rect 2050 361 2099 371
rect 2050 341 2068 361
rect 2088 341 2099 361
rect 2050 329 2099 341
rect 309 127 358 137
rect 309 107 320 127
rect 340 107 358 127
rect 309 95 358 107
rect 408 131 452 137
rect 408 111 423 131
rect 443 111 452 131
rect 408 95 452 111
rect 522 127 571 137
rect 522 107 533 127
rect 553 107 571 127
rect 522 95 571 107
rect 621 131 665 137
rect 621 111 636 131
rect 656 111 665 131
rect 621 95 665 111
rect 730 127 779 137
rect 730 107 741 127
rect 761 107 779 127
rect 730 95 779 107
rect 829 131 873 137
rect 829 111 844 131
rect 864 111 873 131
rect 829 95 873 111
rect 943 131 987 137
rect 943 111 952 131
rect 972 111 987 131
rect 943 95 987 111
rect 1037 127 1086 137
rect 1037 107 1055 127
rect 1075 107 1086 127
rect 1037 95 1086 107
rect 1620 -183 1669 -173
rect 1620 -203 1631 -183
rect 1651 -203 1669 -183
rect 1620 -215 1669 -203
rect 1719 -179 1763 -173
rect 1719 -199 1734 -179
rect 1754 -199 1763 -179
rect 1719 -215 1763 -199
rect 1833 -183 1882 -173
rect 1833 -203 1844 -183
rect 1864 -203 1882 -183
rect 1833 -215 1882 -203
rect 1932 -179 1976 -173
rect 1932 -199 1947 -179
rect 1967 -199 1976 -179
rect 1932 -215 1976 -199
rect 2041 -183 2090 -173
rect 2041 -203 2052 -183
rect 2072 -203 2090 -183
rect 2041 -215 2090 -203
rect 2140 -179 2184 -173
rect 2140 -199 2155 -179
rect 2175 -199 2184 -179
rect 2140 -215 2184 -199
rect 2254 -179 2298 -173
rect 2254 -199 2263 -179
rect 2283 -199 2298 -179
rect 2254 -215 2298 -199
rect 2348 -183 2397 -173
rect 2348 -203 2366 -183
rect 2386 -203 2397 -183
rect 2348 -215 2397 -203
rect 313 -434 362 -424
rect 313 -454 324 -434
rect 344 -454 362 -434
rect 313 -466 362 -454
rect 412 -430 456 -424
rect 412 -450 427 -430
rect 447 -450 456 -430
rect 412 -466 456 -450
rect 526 -434 575 -424
rect 526 -454 537 -434
rect 557 -454 575 -434
rect 526 -466 575 -454
rect 625 -430 669 -424
rect 625 -450 640 -430
rect 660 -450 669 -430
rect 625 -466 669 -450
rect 734 -434 783 -424
rect 734 -454 745 -434
rect 765 -454 783 -434
rect 734 -466 783 -454
rect 833 -430 877 -424
rect 833 -450 848 -430
rect 868 -450 877 -430
rect 833 -466 877 -450
rect 947 -430 991 -424
rect 947 -450 956 -430
rect 976 -450 991 -430
rect 947 -466 991 -450
rect 1041 -434 1090 -424
rect 1041 -454 1059 -434
rect 1079 -454 1090 -434
rect 1041 -466 1090 -454
rect 1325 -615 1374 -605
rect 1325 -635 1336 -615
rect 1356 -635 1374 -615
rect 1325 -647 1374 -635
rect 1424 -611 1468 -605
rect 1424 -631 1439 -611
rect 1459 -631 1468 -611
rect 1424 -647 1468 -631
rect 1538 -615 1587 -605
rect 1538 -635 1549 -615
rect 1569 -635 1587 -615
rect 1538 -647 1587 -635
rect 1637 -611 1681 -605
rect 1637 -631 1652 -611
rect 1672 -631 1681 -611
rect 1637 -647 1681 -631
rect 1746 -615 1795 -605
rect 1746 -635 1757 -615
rect 1777 -635 1795 -615
rect 1746 -647 1795 -635
rect 1845 -611 1889 -605
rect 1845 -631 1860 -611
rect 1880 -631 1889 -611
rect 1845 -647 1889 -631
rect 1959 -611 2003 -605
rect 1959 -631 1968 -611
rect 1988 -631 2003 -611
rect 1959 -647 2003 -631
rect 2053 -615 2102 -605
rect 2053 -635 2071 -615
rect 2091 -635 2102 -615
rect 2053 -647 2102 -635
rect 312 -849 361 -839
rect 312 -869 323 -849
rect 343 -869 361 -849
rect 312 -881 361 -869
rect 411 -845 455 -839
rect 411 -865 426 -845
rect 446 -865 455 -845
rect 411 -881 455 -865
rect 525 -849 574 -839
rect 525 -869 536 -849
rect 556 -869 574 -849
rect 525 -881 574 -869
rect 624 -845 668 -839
rect 624 -865 639 -845
rect 659 -865 668 -845
rect 624 -881 668 -865
rect 733 -849 782 -839
rect 733 -869 744 -849
rect 764 -869 782 -849
rect 733 -881 782 -869
rect 832 -845 876 -839
rect 832 -865 847 -845
rect 867 -865 876 -845
rect 832 -881 876 -865
rect 946 -845 990 -839
rect 946 -865 955 -845
rect 975 -865 990 -845
rect 946 -881 990 -865
rect 1040 -849 1089 -839
rect 1040 -869 1058 -849
rect 1078 -869 1089 -849
rect 1040 -881 1089 -869
rect 1380 -1176 1429 -1166
rect 1380 -1196 1391 -1176
rect 1411 -1196 1429 -1176
rect 1380 -1208 1429 -1196
rect 1479 -1172 1523 -1166
rect 1479 -1192 1494 -1172
rect 1514 -1192 1523 -1172
rect 1479 -1208 1523 -1192
rect 1593 -1176 1642 -1166
rect 1593 -1196 1604 -1176
rect 1624 -1196 1642 -1176
rect 1593 -1208 1642 -1196
rect 1692 -1172 1736 -1166
rect 1692 -1192 1707 -1172
rect 1727 -1192 1736 -1172
rect 1692 -1208 1736 -1192
rect 1801 -1176 1850 -1166
rect 1801 -1196 1812 -1176
rect 1832 -1196 1850 -1176
rect 1801 -1208 1850 -1196
rect 1900 -1172 1944 -1166
rect 1900 -1192 1915 -1172
rect 1935 -1192 1944 -1172
rect 1900 -1208 1944 -1192
rect 2014 -1172 2058 -1166
rect 2014 -1192 2023 -1172
rect 2043 -1192 2058 -1172
rect 2014 -1208 2058 -1192
rect 2108 -1176 2157 -1166
rect 2108 -1196 2126 -1176
rect 2146 -1196 2157 -1176
rect 2108 -1208 2157 -1196
rect 318 -1415 367 -1405
rect 318 -1435 329 -1415
rect 349 -1435 367 -1415
rect 318 -1447 367 -1435
rect 417 -1411 461 -1405
rect 417 -1431 432 -1411
rect 452 -1431 461 -1411
rect 417 -1447 461 -1431
rect 531 -1415 580 -1405
rect 531 -1435 542 -1415
rect 562 -1435 580 -1415
rect 531 -1447 580 -1435
rect 630 -1411 674 -1405
rect 630 -1431 645 -1411
rect 665 -1431 674 -1411
rect 630 -1447 674 -1431
rect 739 -1415 788 -1405
rect 739 -1435 750 -1415
rect 770 -1435 788 -1415
rect 739 -1447 788 -1435
rect 838 -1411 882 -1405
rect 838 -1431 853 -1411
rect 873 -1431 882 -1411
rect 838 -1447 882 -1431
rect 952 -1411 996 -1405
rect 952 -1431 961 -1411
rect 981 -1431 996 -1411
rect 952 -1447 996 -1431
rect 1046 -1415 1095 -1405
rect 1046 -1435 1064 -1415
rect 1084 -1435 1095 -1415
rect 1046 -1447 1095 -1435
rect 1330 -1596 1379 -1586
rect 1330 -1616 1341 -1596
rect 1361 -1616 1379 -1596
rect 1330 -1628 1379 -1616
rect 1429 -1592 1473 -1586
rect 1429 -1612 1444 -1592
rect 1464 -1612 1473 -1592
rect 1429 -1628 1473 -1612
rect 1543 -1596 1592 -1586
rect 1543 -1616 1554 -1596
rect 1574 -1616 1592 -1596
rect 1543 -1628 1592 -1616
rect 1642 -1592 1686 -1586
rect 1642 -1612 1657 -1592
rect 1677 -1612 1686 -1592
rect 1642 -1628 1686 -1612
rect 1751 -1596 1800 -1586
rect 1751 -1616 1762 -1596
rect 1782 -1616 1800 -1596
rect 1751 -1628 1800 -1616
rect 1850 -1592 1894 -1586
rect 1850 -1612 1865 -1592
rect 1885 -1612 1894 -1592
rect 1850 -1628 1894 -1612
rect 1964 -1592 2008 -1586
rect 1964 -1612 1973 -1592
rect 1993 -1612 2008 -1592
rect 1964 -1628 2008 -1612
rect 2058 -1596 2107 -1586
rect 2058 -1616 2076 -1596
rect 2096 -1616 2107 -1596
rect 2058 -1628 2107 -1616
rect 317 -1830 366 -1820
rect 317 -1850 328 -1830
rect 348 -1850 366 -1830
rect 317 -1862 366 -1850
rect 416 -1826 460 -1820
rect 416 -1846 431 -1826
rect 451 -1846 460 -1826
rect 416 -1862 460 -1846
rect 530 -1830 579 -1820
rect 530 -1850 541 -1830
rect 561 -1850 579 -1830
rect 530 -1862 579 -1850
rect 629 -1826 673 -1820
rect 629 -1846 644 -1826
rect 664 -1846 673 -1826
rect 629 -1862 673 -1846
rect 738 -1830 787 -1820
rect 738 -1850 749 -1830
rect 769 -1850 787 -1830
rect 738 -1862 787 -1850
rect 837 -1826 881 -1820
rect 837 -1846 852 -1826
rect 872 -1846 881 -1826
rect 837 -1862 881 -1846
rect 951 -1826 995 -1820
rect 951 -1846 960 -1826
rect 980 -1846 995 -1826
rect 951 -1862 995 -1846
rect 1045 -1830 1094 -1820
rect 1045 -1850 1063 -1830
rect 1083 -1850 1094 -1830
rect 1045 -1862 1094 -1850
rect 1545 -2108 1594 -2098
rect 1545 -2128 1556 -2108
rect 1576 -2128 1594 -2108
rect 1545 -2140 1594 -2128
rect 1644 -2104 1688 -2098
rect 1644 -2124 1659 -2104
rect 1679 -2124 1688 -2104
rect 1644 -2140 1688 -2124
rect 1758 -2108 1807 -2098
rect 1758 -2128 1769 -2108
rect 1789 -2128 1807 -2108
rect 1758 -2140 1807 -2128
rect 1857 -2104 1901 -2098
rect 1857 -2124 1872 -2104
rect 1892 -2124 1901 -2104
rect 1857 -2140 1901 -2124
rect 1966 -2108 2015 -2098
rect 1966 -2128 1977 -2108
rect 1997 -2128 2015 -2108
rect 1966 -2140 2015 -2128
rect 2065 -2104 2109 -2098
rect 2065 -2124 2080 -2104
rect 2100 -2124 2109 -2104
rect 2065 -2140 2109 -2124
rect 2179 -2104 2223 -2098
rect 2179 -2124 2188 -2104
rect 2208 -2124 2223 -2104
rect 2179 -2140 2223 -2124
rect 2273 -2108 2322 -2098
rect 2273 -2128 2291 -2108
rect 2311 -2128 2322 -2108
rect 2273 -2140 2322 -2128
rect 325 -2394 374 -2384
rect 325 -2414 336 -2394
rect 356 -2414 374 -2394
rect 325 -2426 374 -2414
rect 424 -2390 468 -2384
rect 424 -2410 439 -2390
rect 459 -2410 468 -2390
rect 424 -2426 468 -2410
rect 538 -2394 587 -2384
rect 538 -2414 549 -2394
rect 569 -2414 587 -2394
rect 538 -2426 587 -2414
rect 637 -2390 681 -2384
rect 637 -2410 652 -2390
rect 672 -2410 681 -2390
rect 637 -2426 681 -2410
rect 746 -2394 795 -2384
rect 746 -2414 757 -2394
rect 777 -2414 795 -2394
rect 746 -2426 795 -2414
rect 845 -2390 889 -2384
rect 845 -2410 860 -2390
rect 880 -2410 889 -2390
rect 845 -2426 889 -2410
rect 959 -2390 1003 -2384
rect 959 -2410 968 -2390
rect 988 -2410 1003 -2390
rect 959 -2426 1003 -2410
rect 1053 -2394 1102 -2384
rect 1053 -2414 1071 -2394
rect 1091 -2414 1102 -2394
rect 1053 -2426 1102 -2414
rect 1337 -2575 1386 -2565
rect 1337 -2595 1348 -2575
rect 1368 -2595 1386 -2575
rect 1337 -2607 1386 -2595
rect 1436 -2571 1480 -2565
rect 1436 -2591 1451 -2571
rect 1471 -2591 1480 -2571
rect 1436 -2607 1480 -2591
rect 1550 -2575 1599 -2565
rect 1550 -2595 1561 -2575
rect 1581 -2595 1599 -2575
rect 1550 -2607 1599 -2595
rect 1649 -2571 1693 -2565
rect 1649 -2591 1664 -2571
rect 1684 -2591 1693 -2571
rect 1649 -2607 1693 -2591
rect 1758 -2575 1807 -2565
rect 1758 -2595 1769 -2575
rect 1789 -2595 1807 -2575
rect 1758 -2607 1807 -2595
rect 1857 -2571 1901 -2565
rect 1857 -2591 1872 -2571
rect 1892 -2591 1901 -2571
rect 1857 -2607 1901 -2591
rect 1971 -2571 2015 -2565
rect 1971 -2591 1980 -2571
rect 2000 -2591 2015 -2571
rect 1971 -2607 2015 -2591
rect 2065 -2575 2114 -2565
rect 2065 -2595 2083 -2575
rect 2103 -2595 2114 -2575
rect 2065 -2607 2114 -2595
rect 324 -2809 373 -2799
rect 324 -2829 335 -2809
rect 355 -2829 373 -2809
rect 324 -2841 373 -2829
rect 423 -2805 467 -2799
rect 423 -2825 438 -2805
rect 458 -2825 467 -2805
rect 423 -2841 467 -2825
rect 537 -2809 586 -2799
rect 537 -2829 548 -2809
rect 568 -2829 586 -2809
rect 537 -2841 586 -2829
rect 636 -2805 680 -2799
rect 636 -2825 651 -2805
rect 671 -2825 680 -2805
rect 636 -2841 680 -2825
rect 745 -2809 794 -2799
rect 745 -2829 756 -2809
rect 776 -2829 794 -2809
rect 745 -2841 794 -2829
rect 844 -2805 888 -2799
rect 844 -2825 859 -2805
rect 879 -2825 888 -2805
rect 844 -2841 888 -2825
rect 958 -2805 1002 -2799
rect 958 -2825 967 -2805
rect 987 -2825 1002 -2805
rect 958 -2841 1002 -2825
rect 1052 -2809 1101 -2799
rect 1052 -2829 1070 -2809
rect 1090 -2829 1101 -2809
rect 1052 -2841 1101 -2829
rect 1392 -3136 1441 -3126
rect 1392 -3156 1403 -3136
rect 1423 -3156 1441 -3136
rect 1392 -3168 1441 -3156
rect 1491 -3132 1535 -3126
rect 1491 -3152 1506 -3132
rect 1526 -3152 1535 -3132
rect 1491 -3168 1535 -3152
rect 1605 -3136 1654 -3126
rect 1605 -3156 1616 -3136
rect 1636 -3156 1654 -3136
rect 1605 -3168 1654 -3156
rect 1704 -3132 1748 -3126
rect 1704 -3152 1719 -3132
rect 1739 -3152 1748 -3132
rect 1704 -3168 1748 -3152
rect 1813 -3136 1862 -3126
rect 1813 -3156 1824 -3136
rect 1844 -3156 1862 -3136
rect 1813 -3168 1862 -3156
rect 1912 -3132 1956 -3126
rect 1912 -3152 1927 -3132
rect 1947 -3152 1956 -3132
rect 1912 -3168 1956 -3152
rect 2026 -3132 2070 -3126
rect 2026 -3152 2035 -3132
rect 2055 -3152 2070 -3132
rect 2026 -3168 2070 -3152
rect 2120 -3136 2169 -3126
rect 2120 -3156 2138 -3136
rect 2158 -3156 2169 -3136
rect 2120 -3168 2169 -3156
rect 330 -3375 379 -3365
rect 330 -3395 341 -3375
rect 361 -3395 379 -3375
rect 330 -3407 379 -3395
rect 429 -3371 473 -3365
rect 429 -3391 444 -3371
rect 464 -3391 473 -3371
rect 429 -3407 473 -3391
rect 543 -3375 592 -3365
rect 543 -3395 554 -3375
rect 574 -3395 592 -3375
rect 543 -3407 592 -3395
rect 642 -3371 686 -3365
rect 642 -3391 657 -3371
rect 677 -3391 686 -3371
rect 642 -3407 686 -3391
rect 751 -3375 800 -3365
rect 751 -3395 762 -3375
rect 782 -3395 800 -3375
rect 751 -3407 800 -3395
rect 850 -3371 894 -3365
rect 850 -3391 865 -3371
rect 885 -3391 894 -3371
rect 850 -3407 894 -3391
rect 964 -3371 1008 -3365
rect 964 -3391 973 -3371
rect 993 -3391 1008 -3371
rect 964 -3407 1008 -3391
rect 1058 -3375 1107 -3365
rect 1058 -3395 1076 -3375
rect 1096 -3395 1107 -3375
rect 1058 -3407 1107 -3395
rect 1342 -3556 1391 -3546
rect 1342 -3576 1353 -3556
rect 1373 -3576 1391 -3556
rect 1342 -3588 1391 -3576
rect 1441 -3552 1485 -3546
rect 1441 -3572 1456 -3552
rect 1476 -3572 1485 -3552
rect 1441 -3588 1485 -3572
rect 1555 -3556 1604 -3546
rect 1555 -3576 1566 -3556
rect 1586 -3576 1604 -3556
rect 1555 -3588 1604 -3576
rect 1654 -3552 1698 -3546
rect 1654 -3572 1669 -3552
rect 1689 -3572 1698 -3552
rect 1654 -3588 1698 -3572
rect 1763 -3556 1812 -3546
rect 1763 -3576 1774 -3556
rect 1794 -3576 1812 -3556
rect 1763 -3588 1812 -3576
rect 1862 -3552 1906 -3546
rect 1862 -3572 1877 -3552
rect 1897 -3572 1906 -3552
rect 1862 -3588 1906 -3572
rect 1976 -3552 2020 -3546
rect 1976 -3572 1985 -3552
rect 2005 -3572 2020 -3552
rect 1976 -3588 2020 -3572
rect 2070 -3556 2119 -3546
rect 2070 -3576 2088 -3556
rect 2108 -3576 2119 -3556
rect 2070 -3588 2119 -3576
rect 329 -3790 378 -3780
rect 329 -3810 340 -3790
rect 360 -3810 378 -3790
rect 329 -3822 378 -3810
rect 428 -3786 472 -3780
rect 428 -3806 443 -3786
rect 463 -3806 472 -3786
rect 428 -3822 472 -3806
rect 542 -3790 591 -3780
rect 542 -3810 553 -3790
rect 573 -3810 591 -3790
rect 542 -3822 591 -3810
rect 641 -3786 685 -3780
rect 641 -3806 656 -3786
rect 676 -3806 685 -3786
rect 641 -3822 685 -3806
rect 750 -3790 799 -3780
rect 750 -3810 761 -3790
rect 781 -3810 799 -3790
rect 750 -3822 799 -3810
rect 849 -3786 893 -3780
rect 849 -3806 864 -3786
rect 884 -3806 893 -3786
rect 849 -3822 893 -3806
rect 963 -3786 1007 -3780
rect 963 -3806 972 -3786
rect 992 -3806 1007 -3786
rect 963 -3822 1007 -3806
rect 1057 -3790 1106 -3780
rect 1057 -3810 1075 -3790
rect 1095 -3810 1106 -3790
rect 1057 -3822 1106 -3810
<< pdiff >>
rect 298 3632 342 3670
rect 298 3612 310 3632
rect 330 3612 342 3632
rect 298 3570 342 3612
rect 392 3632 434 3670
rect 392 3612 406 3632
rect 426 3612 434 3632
rect 392 3570 434 3612
rect 511 3632 555 3670
rect 511 3612 523 3632
rect 543 3612 555 3632
rect 511 3570 555 3612
rect 605 3632 647 3670
rect 605 3612 619 3632
rect 639 3612 647 3632
rect 605 3570 647 3612
rect 719 3632 763 3670
rect 719 3612 731 3632
rect 751 3612 763 3632
rect 719 3570 763 3612
rect 813 3632 855 3670
rect 813 3612 827 3632
rect 847 3612 855 3632
rect 813 3570 855 3612
rect 929 3632 971 3670
rect 929 3612 937 3632
rect 957 3612 971 3632
rect 929 3570 971 3612
rect 1021 3639 1066 3670
rect 1021 3632 1065 3639
rect 1021 3612 1033 3632
rect 1053 3612 1065 3632
rect 1021 3570 1065 3612
rect 1310 3451 1354 3489
rect 1310 3431 1322 3451
rect 1342 3431 1354 3451
rect 1310 3389 1354 3431
rect 1404 3451 1446 3489
rect 1404 3431 1418 3451
rect 1438 3431 1446 3451
rect 1404 3389 1446 3431
rect 1523 3451 1567 3489
rect 1523 3431 1535 3451
rect 1555 3431 1567 3451
rect 1523 3389 1567 3431
rect 1617 3451 1659 3489
rect 1617 3431 1631 3451
rect 1651 3431 1659 3451
rect 1617 3389 1659 3431
rect 1731 3451 1775 3489
rect 1731 3431 1743 3451
rect 1763 3431 1775 3451
rect 1731 3389 1775 3431
rect 1825 3451 1867 3489
rect 1825 3431 1839 3451
rect 1859 3431 1867 3451
rect 1825 3389 1867 3431
rect 1941 3451 1983 3489
rect 1941 3431 1949 3451
rect 1969 3431 1983 3451
rect 1941 3389 1983 3431
rect 2033 3458 2078 3489
rect 2033 3451 2077 3458
rect 2033 3431 2045 3451
rect 2065 3431 2077 3451
rect 2033 3389 2077 3431
rect 297 3217 341 3255
rect 297 3197 309 3217
rect 329 3197 341 3217
rect 297 3155 341 3197
rect 391 3217 433 3255
rect 391 3197 405 3217
rect 425 3197 433 3217
rect 391 3155 433 3197
rect 510 3217 554 3255
rect 510 3197 522 3217
rect 542 3197 554 3217
rect 510 3155 554 3197
rect 604 3217 646 3255
rect 604 3197 618 3217
rect 638 3197 646 3217
rect 604 3155 646 3197
rect 718 3217 762 3255
rect 718 3197 730 3217
rect 750 3197 762 3217
rect 718 3155 762 3197
rect 812 3217 854 3255
rect 812 3197 826 3217
rect 846 3197 854 3217
rect 812 3155 854 3197
rect 928 3217 970 3255
rect 928 3197 936 3217
rect 956 3197 970 3217
rect 928 3155 970 3197
rect 1020 3224 1065 3255
rect 1020 3217 1064 3224
rect 1020 3197 1032 3217
rect 1052 3197 1064 3217
rect 1020 3155 1064 3197
rect 1365 2890 1409 2928
rect 1365 2870 1377 2890
rect 1397 2870 1409 2890
rect 1365 2828 1409 2870
rect 1459 2890 1501 2928
rect 1459 2870 1473 2890
rect 1493 2870 1501 2890
rect 1459 2828 1501 2870
rect 1578 2890 1622 2928
rect 1578 2870 1590 2890
rect 1610 2870 1622 2890
rect 1578 2828 1622 2870
rect 1672 2890 1714 2928
rect 1672 2870 1686 2890
rect 1706 2870 1714 2890
rect 1672 2828 1714 2870
rect 1786 2890 1830 2928
rect 1786 2870 1798 2890
rect 1818 2870 1830 2890
rect 1786 2828 1830 2870
rect 1880 2890 1922 2928
rect 1880 2870 1894 2890
rect 1914 2870 1922 2890
rect 1880 2828 1922 2870
rect 1996 2890 2038 2928
rect 1996 2870 2004 2890
rect 2024 2870 2038 2890
rect 1996 2828 2038 2870
rect 2088 2897 2133 2928
rect 2088 2890 2132 2897
rect 2088 2870 2100 2890
rect 2120 2870 2132 2890
rect 2088 2828 2132 2870
rect 303 2651 347 2689
rect 303 2631 315 2651
rect 335 2631 347 2651
rect 303 2589 347 2631
rect 397 2651 439 2689
rect 397 2631 411 2651
rect 431 2631 439 2651
rect 397 2589 439 2631
rect 516 2651 560 2689
rect 516 2631 528 2651
rect 548 2631 560 2651
rect 516 2589 560 2631
rect 610 2651 652 2689
rect 610 2631 624 2651
rect 644 2631 652 2651
rect 610 2589 652 2631
rect 724 2651 768 2689
rect 724 2631 736 2651
rect 756 2631 768 2651
rect 724 2589 768 2631
rect 818 2651 860 2689
rect 818 2631 832 2651
rect 852 2631 860 2651
rect 818 2589 860 2631
rect 934 2651 976 2689
rect 934 2631 942 2651
rect 962 2631 976 2651
rect 934 2589 976 2631
rect 1026 2658 1071 2689
rect 1026 2651 1070 2658
rect 1026 2631 1038 2651
rect 1058 2631 1070 2651
rect 1026 2589 1070 2631
rect 1315 2470 1359 2508
rect 1315 2450 1327 2470
rect 1347 2450 1359 2470
rect 1315 2408 1359 2450
rect 1409 2470 1451 2508
rect 1409 2450 1423 2470
rect 1443 2450 1451 2470
rect 1409 2408 1451 2450
rect 1528 2470 1572 2508
rect 1528 2450 1540 2470
rect 1560 2450 1572 2470
rect 1528 2408 1572 2450
rect 1622 2470 1664 2508
rect 1622 2450 1636 2470
rect 1656 2450 1664 2470
rect 1622 2408 1664 2450
rect 1736 2470 1780 2508
rect 1736 2450 1748 2470
rect 1768 2450 1780 2470
rect 1736 2408 1780 2450
rect 1830 2470 1872 2508
rect 1830 2450 1844 2470
rect 1864 2450 1872 2470
rect 1830 2408 1872 2450
rect 1946 2470 1988 2508
rect 1946 2450 1954 2470
rect 1974 2450 1988 2470
rect 1946 2408 1988 2450
rect 2038 2477 2083 2508
rect 2038 2470 2082 2477
rect 2038 2450 2050 2470
rect 2070 2450 2082 2470
rect 2038 2408 2082 2450
rect 302 2236 346 2274
rect 302 2216 314 2236
rect 334 2216 346 2236
rect 302 2174 346 2216
rect 396 2236 438 2274
rect 396 2216 410 2236
rect 430 2216 438 2236
rect 396 2174 438 2216
rect 515 2236 559 2274
rect 515 2216 527 2236
rect 547 2216 559 2236
rect 515 2174 559 2216
rect 609 2236 651 2274
rect 609 2216 623 2236
rect 643 2216 651 2236
rect 609 2174 651 2216
rect 723 2236 767 2274
rect 723 2216 735 2236
rect 755 2216 767 2236
rect 723 2174 767 2216
rect 817 2236 859 2274
rect 817 2216 831 2236
rect 851 2216 859 2236
rect 817 2174 859 2216
rect 933 2236 975 2274
rect 933 2216 941 2236
rect 961 2216 975 2236
rect 933 2174 975 2216
rect 1025 2243 1070 2274
rect 1025 2236 1069 2243
rect 1025 2216 1037 2236
rect 1057 2216 1069 2236
rect 1025 2174 1069 2216
rect 1530 1958 1574 1996
rect 1530 1938 1542 1958
rect 1562 1938 1574 1958
rect 1530 1896 1574 1938
rect 1624 1958 1666 1996
rect 1624 1938 1638 1958
rect 1658 1938 1666 1958
rect 1624 1896 1666 1938
rect 1743 1958 1787 1996
rect 1743 1938 1755 1958
rect 1775 1938 1787 1958
rect 1743 1896 1787 1938
rect 1837 1958 1879 1996
rect 1837 1938 1851 1958
rect 1871 1938 1879 1958
rect 1837 1896 1879 1938
rect 1951 1958 1995 1996
rect 1951 1938 1963 1958
rect 1983 1938 1995 1958
rect 1951 1896 1995 1938
rect 2045 1958 2087 1996
rect 2045 1938 2059 1958
rect 2079 1938 2087 1958
rect 2045 1896 2087 1938
rect 2161 1958 2203 1996
rect 2161 1938 2169 1958
rect 2189 1938 2203 1958
rect 2161 1896 2203 1938
rect 2253 1965 2298 1996
rect 2253 1958 2297 1965
rect 2253 1938 2265 1958
rect 2285 1938 2297 1958
rect 2253 1896 2297 1938
rect 310 1672 354 1710
rect 310 1652 322 1672
rect 342 1652 354 1672
rect 310 1610 354 1652
rect 404 1672 446 1710
rect 404 1652 418 1672
rect 438 1652 446 1672
rect 404 1610 446 1652
rect 523 1672 567 1710
rect 523 1652 535 1672
rect 555 1652 567 1672
rect 523 1610 567 1652
rect 617 1672 659 1710
rect 617 1652 631 1672
rect 651 1652 659 1672
rect 617 1610 659 1652
rect 731 1672 775 1710
rect 731 1652 743 1672
rect 763 1652 775 1672
rect 731 1610 775 1652
rect 825 1672 867 1710
rect 825 1652 839 1672
rect 859 1652 867 1672
rect 825 1610 867 1652
rect 941 1672 983 1710
rect 941 1652 949 1672
rect 969 1652 983 1672
rect 941 1610 983 1652
rect 1033 1679 1078 1710
rect 1033 1672 1077 1679
rect 1033 1652 1045 1672
rect 1065 1652 1077 1672
rect 1033 1610 1077 1652
rect 1322 1491 1366 1529
rect 1322 1471 1334 1491
rect 1354 1471 1366 1491
rect 1322 1429 1366 1471
rect 1416 1491 1458 1529
rect 1416 1471 1430 1491
rect 1450 1471 1458 1491
rect 1416 1429 1458 1471
rect 1535 1491 1579 1529
rect 1535 1471 1547 1491
rect 1567 1471 1579 1491
rect 1535 1429 1579 1471
rect 1629 1491 1671 1529
rect 1629 1471 1643 1491
rect 1663 1471 1671 1491
rect 1629 1429 1671 1471
rect 1743 1491 1787 1529
rect 1743 1471 1755 1491
rect 1775 1471 1787 1491
rect 1743 1429 1787 1471
rect 1837 1491 1879 1529
rect 1837 1471 1851 1491
rect 1871 1471 1879 1491
rect 1837 1429 1879 1471
rect 1953 1491 1995 1529
rect 1953 1471 1961 1491
rect 1981 1471 1995 1491
rect 1953 1429 1995 1471
rect 2045 1498 2090 1529
rect 2045 1491 2089 1498
rect 2045 1471 2057 1491
rect 2077 1471 2089 1491
rect 2045 1429 2089 1471
rect 309 1257 353 1295
rect 309 1237 321 1257
rect 341 1237 353 1257
rect 309 1195 353 1237
rect 403 1257 445 1295
rect 403 1237 417 1257
rect 437 1237 445 1257
rect 403 1195 445 1237
rect 522 1257 566 1295
rect 522 1237 534 1257
rect 554 1237 566 1257
rect 522 1195 566 1237
rect 616 1257 658 1295
rect 616 1237 630 1257
rect 650 1237 658 1257
rect 616 1195 658 1237
rect 730 1257 774 1295
rect 730 1237 742 1257
rect 762 1237 774 1257
rect 730 1195 774 1237
rect 824 1257 866 1295
rect 824 1237 838 1257
rect 858 1237 866 1257
rect 824 1195 866 1237
rect 940 1257 982 1295
rect 940 1237 948 1257
rect 968 1237 982 1257
rect 940 1195 982 1237
rect 1032 1264 1077 1295
rect 1032 1257 1076 1264
rect 1032 1237 1044 1257
rect 1064 1237 1076 1257
rect 1032 1195 1076 1237
rect 1377 930 1421 968
rect 1377 910 1389 930
rect 1409 910 1421 930
rect 1377 868 1421 910
rect 1471 930 1513 968
rect 1471 910 1485 930
rect 1505 910 1513 930
rect 1471 868 1513 910
rect 1590 930 1634 968
rect 1590 910 1602 930
rect 1622 910 1634 930
rect 1590 868 1634 910
rect 1684 930 1726 968
rect 1684 910 1698 930
rect 1718 910 1726 930
rect 1684 868 1726 910
rect 1798 930 1842 968
rect 1798 910 1810 930
rect 1830 910 1842 930
rect 1798 868 1842 910
rect 1892 930 1934 968
rect 1892 910 1906 930
rect 1926 910 1934 930
rect 1892 868 1934 910
rect 2008 930 2050 968
rect 2008 910 2016 930
rect 2036 910 2050 930
rect 2008 868 2050 910
rect 2100 937 2145 968
rect 2100 930 2144 937
rect 2100 910 2112 930
rect 2132 910 2144 930
rect 2100 868 2144 910
rect 315 691 359 729
rect 315 671 327 691
rect 347 671 359 691
rect 315 629 359 671
rect 409 691 451 729
rect 409 671 423 691
rect 443 671 451 691
rect 409 629 451 671
rect 528 691 572 729
rect 528 671 540 691
rect 560 671 572 691
rect 528 629 572 671
rect 622 691 664 729
rect 622 671 636 691
rect 656 671 664 691
rect 622 629 664 671
rect 736 691 780 729
rect 736 671 748 691
rect 768 671 780 691
rect 736 629 780 671
rect 830 691 872 729
rect 830 671 844 691
rect 864 671 872 691
rect 830 629 872 671
rect 946 691 988 729
rect 946 671 954 691
rect 974 671 988 691
rect 946 629 988 671
rect 1038 698 1083 729
rect 1038 691 1082 698
rect 1038 671 1050 691
rect 1070 671 1082 691
rect 1038 629 1082 671
rect 1327 510 1371 548
rect 1327 490 1339 510
rect 1359 490 1371 510
rect 1327 448 1371 490
rect 1421 510 1463 548
rect 1421 490 1435 510
rect 1455 490 1463 510
rect 1421 448 1463 490
rect 1540 510 1584 548
rect 1540 490 1552 510
rect 1572 490 1584 510
rect 1540 448 1584 490
rect 1634 510 1676 548
rect 1634 490 1648 510
rect 1668 490 1676 510
rect 1634 448 1676 490
rect 1748 510 1792 548
rect 1748 490 1760 510
rect 1780 490 1792 510
rect 1748 448 1792 490
rect 1842 510 1884 548
rect 1842 490 1856 510
rect 1876 490 1884 510
rect 1842 448 1884 490
rect 1958 510 2000 548
rect 1958 490 1966 510
rect 1986 490 2000 510
rect 1958 448 2000 490
rect 2050 517 2095 548
rect 2050 510 2094 517
rect 2050 490 2062 510
rect 2082 490 2094 510
rect 2050 448 2094 490
rect 314 276 358 314
rect 314 256 326 276
rect 346 256 358 276
rect 314 214 358 256
rect 408 276 450 314
rect 408 256 422 276
rect 442 256 450 276
rect 408 214 450 256
rect 527 276 571 314
rect 527 256 539 276
rect 559 256 571 276
rect 527 214 571 256
rect 621 276 663 314
rect 621 256 635 276
rect 655 256 663 276
rect 621 214 663 256
rect 735 276 779 314
rect 735 256 747 276
rect 767 256 779 276
rect 735 214 779 256
rect 829 276 871 314
rect 829 256 843 276
rect 863 256 871 276
rect 829 214 871 256
rect 945 276 987 314
rect 945 256 953 276
rect 973 256 987 276
rect 945 214 987 256
rect 1037 283 1082 314
rect 1037 276 1081 283
rect 1037 256 1049 276
rect 1069 256 1081 276
rect 1037 214 1081 256
rect 1625 -34 1669 4
rect 1625 -54 1637 -34
rect 1657 -54 1669 -34
rect 1625 -96 1669 -54
rect 1719 -34 1761 4
rect 1719 -54 1733 -34
rect 1753 -54 1761 -34
rect 1719 -96 1761 -54
rect 1838 -34 1882 4
rect 1838 -54 1850 -34
rect 1870 -54 1882 -34
rect 1838 -96 1882 -54
rect 1932 -34 1974 4
rect 1932 -54 1946 -34
rect 1966 -54 1974 -34
rect 1932 -96 1974 -54
rect 2046 -34 2090 4
rect 2046 -54 2058 -34
rect 2078 -54 2090 -34
rect 2046 -96 2090 -54
rect 2140 -34 2182 4
rect 2140 -54 2154 -34
rect 2174 -54 2182 -34
rect 2140 -96 2182 -54
rect 2256 -34 2298 4
rect 2256 -54 2264 -34
rect 2284 -54 2298 -34
rect 2256 -96 2298 -54
rect 2348 -27 2393 4
rect 2348 -34 2392 -27
rect 2348 -54 2360 -34
rect 2380 -54 2392 -34
rect 2348 -96 2392 -54
rect 318 -285 362 -247
rect 318 -305 330 -285
rect 350 -305 362 -285
rect 318 -347 362 -305
rect 412 -285 454 -247
rect 412 -305 426 -285
rect 446 -305 454 -285
rect 412 -347 454 -305
rect 531 -285 575 -247
rect 531 -305 543 -285
rect 563 -305 575 -285
rect 531 -347 575 -305
rect 625 -285 667 -247
rect 625 -305 639 -285
rect 659 -305 667 -285
rect 625 -347 667 -305
rect 739 -285 783 -247
rect 739 -305 751 -285
rect 771 -305 783 -285
rect 739 -347 783 -305
rect 833 -285 875 -247
rect 833 -305 847 -285
rect 867 -305 875 -285
rect 833 -347 875 -305
rect 949 -285 991 -247
rect 949 -305 957 -285
rect 977 -305 991 -285
rect 949 -347 991 -305
rect 1041 -278 1086 -247
rect 1041 -285 1085 -278
rect 1041 -305 1053 -285
rect 1073 -305 1085 -285
rect 1041 -347 1085 -305
rect 1330 -466 1374 -428
rect 1330 -486 1342 -466
rect 1362 -486 1374 -466
rect 1330 -528 1374 -486
rect 1424 -466 1466 -428
rect 1424 -486 1438 -466
rect 1458 -486 1466 -466
rect 1424 -528 1466 -486
rect 1543 -466 1587 -428
rect 1543 -486 1555 -466
rect 1575 -486 1587 -466
rect 1543 -528 1587 -486
rect 1637 -466 1679 -428
rect 1637 -486 1651 -466
rect 1671 -486 1679 -466
rect 1637 -528 1679 -486
rect 1751 -466 1795 -428
rect 1751 -486 1763 -466
rect 1783 -486 1795 -466
rect 1751 -528 1795 -486
rect 1845 -466 1887 -428
rect 1845 -486 1859 -466
rect 1879 -486 1887 -466
rect 1845 -528 1887 -486
rect 1961 -466 2003 -428
rect 1961 -486 1969 -466
rect 1989 -486 2003 -466
rect 1961 -528 2003 -486
rect 2053 -459 2098 -428
rect 2053 -466 2097 -459
rect 2053 -486 2065 -466
rect 2085 -486 2097 -466
rect 2053 -528 2097 -486
rect 317 -700 361 -662
rect 317 -720 329 -700
rect 349 -720 361 -700
rect 317 -762 361 -720
rect 411 -700 453 -662
rect 411 -720 425 -700
rect 445 -720 453 -700
rect 411 -762 453 -720
rect 530 -700 574 -662
rect 530 -720 542 -700
rect 562 -720 574 -700
rect 530 -762 574 -720
rect 624 -700 666 -662
rect 624 -720 638 -700
rect 658 -720 666 -700
rect 624 -762 666 -720
rect 738 -700 782 -662
rect 738 -720 750 -700
rect 770 -720 782 -700
rect 738 -762 782 -720
rect 832 -700 874 -662
rect 832 -720 846 -700
rect 866 -720 874 -700
rect 832 -762 874 -720
rect 948 -700 990 -662
rect 948 -720 956 -700
rect 976 -720 990 -700
rect 948 -762 990 -720
rect 1040 -693 1085 -662
rect 1040 -700 1084 -693
rect 1040 -720 1052 -700
rect 1072 -720 1084 -700
rect 1040 -762 1084 -720
rect 1385 -1027 1429 -989
rect 1385 -1047 1397 -1027
rect 1417 -1047 1429 -1027
rect 1385 -1089 1429 -1047
rect 1479 -1027 1521 -989
rect 1479 -1047 1493 -1027
rect 1513 -1047 1521 -1027
rect 1479 -1089 1521 -1047
rect 1598 -1027 1642 -989
rect 1598 -1047 1610 -1027
rect 1630 -1047 1642 -1027
rect 1598 -1089 1642 -1047
rect 1692 -1027 1734 -989
rect 1692 -1047 1706 -1027
rect 1726 -1047 1734 -1027
rect 1692 -1089 1734 -1047
rect 1806 -1027 1850 -989
rect 1806 -1047 1818 -1027
rect 1838 -1047 1850 -1027
rect 1806 -1089 1850 -1047
rect 1900 -1027 1942 -989
rect 1900 -1047 1914 -1027
rect 1934 -1047 1942 -1027
rect 1900 -1089 1942 -1047
rect 2016 -1027 2058 -989
rect 2016 -1047 2024 -1027
rect 2044 -1047 2058 -1027
rect 2016 -1089 2058 -1047
rect 2108 -1020 2153 -989
rect 2108 -1027 2152 -1020
rect 2108 -1047 2120 -1027
rect 2140 -1047 2152 -1027
rect 2108 -1089 2152 -1047
rect 323 -1266 367 -1228
rect 323 -1286 335 -1266
rect 355 -1286 367 -1266
rect 323 -1328 367 -1286
rect 417 -1266 459 -1228
rect 417 -1286 431 -1266
rect 451 -1286 459 -1266
rect 417 -1328 459 -1286
rect 536 -1266 580 -1228
rect 536 -1286 548 -1266
rect 568 -1286 580 -1266
rect 536 -1328 580 -1286
rect 630 -1266 672 -1228
rect 630 -1286 644 -1266
rect 664 -1286 672 -1266
rect 630 -1328 672 -1286
rect 744 -1266 788 -1228
rect 744 -1286 756 -1266
rect 776 -1286 788 -1266
rect 744 -1328 788 -1286
rect 838 -1266 880 -1228
rect 838 -1286 852 -1266
rect 872 -1286 880 -1266
rect 838 -1328 880 -1286
rect 954 -1266 996 -1228
rect 954 -1286 962 -1266
rect 982 -1286 996 -1266
rect 954 -1328 996 -1286
rect 1046 -1259 1091 -1228
rect 1046 -1266 1090 -1259
rect 1046 -1286 1058 -1266
rect 1078 -1286 1090 -1266
rect 1046 -1328 1090 -1286
rect 1335 -1447 1379 -1409
rect 1335 -1467 1347 -1447
rect 1367 -1467 1379 -1447
rect 1335 -1509 1379 -1467
rect 1429 -1447 1471 -1409
rect 1429 -1467 1443 -1447
rect 1463 -1467 1471 -1447
rect 1429 -1509 1471 -1467
rect 1548 -1447 1592 -1409
rect 1548 -1467 1560 -1447
rect 1580 -1467 1592 -1447
rect 1548 -1509 1592 -1467
rect 1642 -1447 1684 -1409
rect 1642 -1467 1656 -1447
rect 1676 -1467 1684 -1447
rect 1642 -1509 1684 -1467
rect 1756 -1447 1800 -1409
rect 1756 -1467 1768 -1447
rect 1788 -1467 1800 -1447
rect 1756 -1509 1800 -1467
rect 1850 -1447 1892 -1409
rect 1850 -1467 1864 -1447
rect 1884 -1467 1892 -1447
rect 1850 -1509 1892 -1467
rect 1966 -1447 2008 -1409
rect 1966 -1467 1974 -1447
rect 1994 -1467 2008 -1447
rect 1966 -1509 2008 -1467
rect 2058 -1440 2103 -1409
rect 2058 -1447 2102 -1440
rect 2058 -1467 2070 -1447
rect 2090 -1467 2102 -1447
rect 2058 -1509 2102 -1467
rect 322 -1681 366 -1643
rect 322 -1701 334 -1681
rect 354 -1701 366 -1681
rect 322 -1743 366 -1701
rect 416 -1681 458 -1643
rect 416 -1701 430 -1681
rect 450 -1701 458 -1681
rect 416 -1743 458 -1701
rect 535 -1681 579 -1643
rect 535 -1701 547 -1681
rect 567 -1701 579 -1681
rect 535 -1743 579 -1701
rect 629 -1681 671 -1643
rect 629 -1701 643 -1681
rect 663 -1701 671 -1681
rect 629 -1743 671 -1701
rect 743 -1681 787 -1643
rect 743 -1701 755 -1681
rect 775 -1701 787 -1681
rect 743 -1743 787 -1701
rect 837 -1681 879 -1643
rect 837 -1701 851 -1681
rect 871 -1701 879 -1681
rect 837 -1743 879 -1701
rect 953 -1681 995 -1643
rect 953 -1701 961 -1681
rect 981 -1701 995 -1681
rect 953 -1743 995 -1701
rect 1045 -1674 1090 -1643
rect 1045 -1681 1089 -1674
rect 1045 -1701 1057 -1681
rect 1077 -1701 1089 -1681
rect 1045 -1743 1089 -1701
rect 1550 -1959 1594 -1921
rect 1550 -1979 1562 -1959
rect 1582 -1979 1594 -1959
rect 1550 -2021 1594 -1979
rect 1644 -1959 1686 -1921
rect 1644 -1979 1658 -1959
rect 1678 -1979 1686 -1959
rect 1644 -2021 1686 -1979
rect 1763 -1959 1807 -1921
rect 1763 -1979 1775 -1959
rect 1795 -1979 1807 -1959
rect 1763 -2021 1807 -1979
rect 1857 -1959 1899 -1921
rect 1857 -1979 1871 -1959
rect 1891 -1979 1899 -1959
rect 1857 -2021 1899 -1979
rect 1971 -1959 2015 -1921
rect 1971 -1979 1983 -1959
rect 2003 -1979 2015 -1959
rect 1971 -2021 2015 -1979
rect 2065 -1959 2107 -1921
rect 2065 -1979 2079 -1959
rect 2099 -1979 2107 -1959
rect 2065 -2021 2107 -1979
rect 2181 -1959 2223 -1921
rect 2181 -1979 2189 -1959
rect 2209 -1979 2223 -1959
rect 2181 -2021 2223 -1979
rect 2273 -1952 2318 -1921
rect 2273 -1959 2317 -1952
rect 2273 -1979 2285 -1959
rect 2305 -1979 2317 -1959
rect 2273 -2021 2317 -1979
rect 330 -2245 374 -2207
rect 330 -2265 342 -2245
rect 362 -2265 374 -2245
rect 330 -2307 374 -2265
rect 424 -2245 466 -2207
rect 424 -2265 438 -2245
rect 458 -2265 466 -2245
rect 424 -2307 466 -2265
rect 543 -2245 587 -2207
rect 543 -2265 555 -2245
rect 575 -2265 587 -2245
rect 543 -2307 587 -2265
rect 637 -2245 679 -2207
rect 637 -2265 651 -2245
rect 671 -2265 679 -2245
rect 637 -2307 679 -2265
rect 751 -2245 795 -2207
rect 751 -2265 763 -2245
rect 783 -2265 795 -2245
rect 751 -2307 795 -2265
rect 845 -2245 887 -2207
rect 845 -2265 859 -2245
rect 879 -2265 887 -2245
rect 845 -2307 887 -2265
rect 961 -2245 1003 -2207
rect 961 -2265 969 -2245
rect 989 -2265 1003 -2245
rect 961 -2307 1003 -2265
rect 1053 -2238 1098 -2207
rect 1053 -2245 1097 -2238
rect 1053 -2265 1065 -2245
rect 1085 -2265 1097 -2245
rect 1053 -2307 1097 -2265
rect 1342 -2426 1386 -2388
rect 1342 -2446 1354 -2426
rect 1374 -2446 1386 -2426
rect 1342 -2488 1386 -2446
rect 1436 -2426 1478 -2388
rect 1436 -2446 1450 -2426
rect 1470 -2446 1478 -2426
rect 1436 -2488 1478 -2446
rect 1555 -2426 1599 -2388
rect 1555 -2446 1567 -2426
rect 1587 -2446 1599 -2426
rect 1555 -2488 1599 -2446
rect 1649 -2426 1691 -2388
rect 1649 -2446 1663 -2426
rect 1683 -2446 1691 -2426
rect 1649 -2488 1691 -2446
rect 1763 -2426 1807 -2388
rect 1763 -2446 1775 -2426
rect 1795 -2446 1807 -2426
rect 1763 -2488 1807 -2446
rect 1857 -2426 1899 -2388
rect 1857 -2446 1871 -2426
rect 1891 -2446 1899 -2426
rect 1857 -2488 1899 -2446
rect 1973 -2426 2015 -2388
rect 1973 -2446 1981 -2426
rect 2001 -2446 2015 -2426
rect 1973 -2488 2015 -2446
rect 2065 -2419 2110 -2388
rect 2065 -2426 2109 -2419
rect 2065 -2446 2077 -2426
rect 2097 -2446 2109 -2426
rect 2065 -2488 2109 -2446
rect 329 -2660 373 -2622
rect 329 -2680 341 -2660
rect 361 -2680 373 -2660
rect 329 -2722 373 -2680
rect 423 -2660 465 -2622
rect 423 -2680 437 -2660
rect 457 -2680 465 -2660
rect 423 -2722 465 -2680
rect 542 -2660 586 -2622
rect 542 -2680 554 -2660
rect 574 -2680 586 -2660
rect 542 -2722 586 -2680
rect 636 -2660 678 -2622
rect 636 -2680 650 -2660
rect 670 -2680 678 -2660
rect 636 -2722 678 -2680
rect 750 -2660 794 -2622
rect 750 -2680 762 -2660
rect 782 -2680 794 -2660
rect 750 -2722 794 -2680
rect 844 -2660 886 -2622
rect 844 -2680 858 -2660
rect 878 -2680 886 -2660
rect 844 -2722 886 -2680
rect 960 -2660 1002 -2622
rect 960 -2680 968 -2660
rect 988 -2680 1002 -2660
rect 960 -2722 1002 -2680
rect 1052 -2653 1097 -2622
rect 1052 -2660 1096 -2653
rect 1052 -2680 1064 -2660
rect 1084 -2680 1096 -2660
rect 1052 -2722 1096 -2680
rect 1397 -2987 1441 -2949
rect 1397 -3007 1409 -2987
rect 1429 -3007 1441 -2987
rect 1397 -3049 1441 -3007
rect 1491 -2987 1533 -2949
rect 1491 -3007 1505 -2987
rect 1525 -3007 1533 -2987
rect 1491 -3049 1533 -3007
rect 1610 -2987 1654 -2949
rect 1610 -3007 1622 -2987
rect 1642 -3007 1654 -2987
rect 1610 -3049 1654 -3007
rect 1704 -2987 1746 -2949
rect 1704 -3007 1718 -2987
rect 1738 -3007 1746 -2987
rect 1704 -3049 1746 -3007
rect 1818 -2987 1862 -2949
rect 1818 -3007 1830 -2987
rect 1850 -3007 1862 -2987
rect 1818 -3049 1862 -3007
rect 1912 -2987 1954 -2949
rect 1912 -3007 1926 -2987
rect 1946 -3007 1954 -2987
rect 1912 -3049 1954 -3007
rect 2028 -2987 2070 -2949
rect 2028 -3007 2036 -2987
rect 2056 -3007 2070 -2987
rect 2028 -3049 2070 -3007
rect 2120 -2980 2165 -2949
rect 2120 -2987 2164 -2980
rect 2120 -3007 2132 -2987
rect 2152 -3007 2164 -2987
rect 2120 -3049 2164 -3007
rect 335 -3226 379 -3188
rect 335 -3246 347 -3226
rect 367 -3246 379 -3226
rect 335 -3288 379 -3246
rect 429 -3226 471 -3188
rect 429 -3246 443 -3226
rect 463 -3246 471 -3226
rect 429 -3288 471 -3246
rect 548 -3226 592 -3188
rect 548 -3246 560 -3226
rect 580 -3246 592 -3226
rect 548 -3288 592 -3246
rect 642 -3226 684 -3188
rect 642 -3246 656 -3226
rect 676 -3246 684 -3226
rect 642 -3288 684 -3246
rect 756 -3226 800 -3188
rect 756 -3246 768 -3226
rect 788 -3246 800 -3226
rect 756 -3288 800 -3246
rect 850 -3226 892 -3188
rect 850 -3246 864 -3226
rect 884 -3246 892 -3226
rect 850 -3288 892 -3246
rect 966 -3226 1008 -3188
rect 966 -3246 974 -3226
rect 994 -3246 1008 -3226
rect 966 -3288 1008 -3246
rect 1058 -3219 1103 -3188
rect 1058 -3226 1102 -3219
rect 1058 -3246 1070 -3226
rect 1090 -3246 1102 -3226
rect 1058 -3288 1102 -3246
rect 1347 -3407 1391 -3369
rect 1347 -3427 1359 -3407
rect 1379 -3427 1391 -3407
rect 1347 -3469 1391 -3427
rect 1441 -3407 1483 -3369
rect 1441 -3427 1455 -3407
rect 1475 -3427 1483 -3407
rect 1441 -3469 1483 -3427
rect 1560 -3407 1604 -3369
rect 1560 -3427 1572 -3407
rect 1592 -3427 1604 -3407
rect 1560 -3469 1604 -3427
rect 1654 -3407 1696 -3369
rect 1654 -3427 1668 -3407
rect 1688 -3427 1696 -3407
rect 1654 -3469 1696 -3427
rect 1768 -3407 1812 -3369
rect 1768 -3427 1780 -3407
rect 1800 -3427 1812 -3407
rect 1768 -3469 1812 -3427
rect 1862 -3407 1904 -3369
rect 1862 -3427 1876 -3407
rect 1896 -3427 1904 -3407
rect 1862 -3469 1904 -3427
rect 1978 -3407 2020 -3369
rect 1978 -3427 1986 -3407
rect 2006 -3427 2020 -3407
rect 1978 -3469 2020 -3427
rect 2070 -3400 2115 -3369
rect 2070 -3407 2114 -3400
rect 2070 -3427 2082 -3407
rect 2102 -3427 2114 -3407
rect 2070 -3469 2114 -3427
rect 334 -3641 378 -3603
rect 334 -3661 346 -3641
rect 366 -3661 378 -3641
rect 334 -3703 378 -3661
rect 428 -3641 470 -3603
rect 428 -3661 442 -3641
rect 462 -3661 470 -3641
rect 428 -3703 470 -3661
rect 547 -3641 591 -3603
rect 547 -3661 559 -3641
rect 579 -3661 591 -3641
rect 547 -3703 591 -3661
rect 641 -3641 683 -3603
rect 641 -3661 655 -3641
rect 675 -3661 683 -3641
rect 641 -3703 683 -3661
rect 755 -3641 799 -3603
rect 755 -3661 767 -3641
rect 787 -3661 799 -3641
rect 755 -3703 799 -3661
rect 849 -3641 891 -3603
rect 849 -3661 863 -3641
rect 883 -3661 891 -3641
rect 849 -3703 891 -3661
rect 965 -3641 1007 -3603
rect 965 -3661 973 -3641
rect 993 -3661 1007 -3641
rect 965 -3703 1007 -3661
rect 1057 -3634 1102 -3603
rect 1057 -3641 1101 -3634
rect 1057 -3661 1069 -3641
rect 1089 -3661 1101 -3641
rect 1057 -3703 1101 -3661
<< ndiffc >>
rect 118 3847 136 3865
rect 120 3748 138 3766
rect 116 3633 134 3651
rect 118 3534 136 3552
rect 304 3463 324 3483
rect 407 3467 427 3487
rect 517 3463 537 3483
rect 620 3467 640 3487
rect 725 3463 745 3483
rect 828 3467 848 3487
rect 936 3467 956 3487
rect 1039 3463 1059 3483
rect 116 3351 134 3369
rect 1316 3282 1336 3302
rect 1419 3286 1439 3306
rect 1529 3282 1549 3302
rect 1632 3286 1652 3306
rect 1737 3282 1757 3302
rect 1840 3286 1860 3306
rect 1948 3286 1968 3306
rect 2051 3282 2071 3302
rect 118 3252 136 3270
rect 123 3150 141 3168
rect 125 3051 143 3069
rect 303 3048 323 3068
rect 406 3052 426 3072
rect 516 3048 536 3068
rect 619 3052 639 3072
rect 724 3048 744 3068
rect 827 3052 847 3072
rect 935 3052 955 3072
rect 1038 3048 1058 3068
rect 123 2866 141 2884
rect 125 2767 143 2785
rect 1371 2721 1391 2741
rect 1474 2725 1494 2745
rect 1584 2721 1604 2741
rect 1687 2725 1707 2745
rect 1792 2721 1812 2741
rect 1895 2725 1915 2745
rect 2003 2725 2023 2745
rect 2106 2721 2126 2741
rect 121 2652 139 2670
rect 123 2553 141 2571
rect 309 2482 329 2502
rect 412 2486 432 2506
rect 522 2482 542 2502
rect 625 2486 645 2506
rect 730 2482 750 2502
rect 833 2486 853 2506
rect 941 2486 961 2506
rect 1044 2482 1064 2502
rect 121 2370 139 2388
rect 1321 2301 1341 2321
rect 1424 2305 1444 2325
rect 1534 2301 1554 2321
rect 1637 2305 1657 2325
rect 1742 2301 1762 2321
rect 1845 2305 1865 2325
rect 1953 2305 1973 2325
rect 2056 2301 2076 2321
rect 123 2271 141 2289
rect 128 2169 146 2187
rect 130 2070 148 2088
rect 308 2067 328 2087
rect 411 2071 431 2091
rect 521 2067 541 2087
rect 624 2071 644 2091
rect 729 2067 749 2087
rect 832 2071 852 2091
rect 940 2071 960 2091
rect 1043 2067 1063 2087
rect 130 1887 148 1905
rect 132 1788 150 1806
rect 1536 1789 1556 1809
rect 1639 1793 1659 1813
rect 1749 1789 1769 1809
rect 1852 1793 1872 1813
rect 1957 1789 1977 1809
rect 2060 1793 2080 1813
rect 2168 1793 2188 1813
rect 2271 1789 2291 1809
rect 128 1673 146 1691
rect 130 1574 148 1592
rect 316 1503 336 1523
rect 419 1507 439 1527
rect 529 1503 549 1523
rect 632 1507 652 1527
rect 737 1503 757 1523
rect 840 1507 860 1527
rect 948 1507 968 1527
rect 1051 1503 1071 1523
rect 128 1391 146 1409
rect 1328 1322 1348 1342
rect 1431 1326 1451 1346
rect 1541 1322 1561 1342
rect 1644 1326 1664 1346
rect 1749 1322 1769 1342
rect 1852 1326 1872 1346
rect 1960 1326 1980 1346
rect 2063 1322 2083 1342
rect 130 1292 148 1310
rect 135 1190 153 1208
rect 137 1091 155 1109
rect 315 1088 335 1108
rect 418 1092 438 1112
rect 528 1088 548 1108
rect 631 1092 651 1112
rect 736 1088 756 1108
rect 839 1092 859 1112
rect 947 1092 967 1112
rect 1050 1088 1070 1108
rect 135 906 153 924
rect 137 807 155 825
rect 1383 761 1403 781
rect 1486 765 1506 785
rect 1596 761 1616 781
rect 1699 765 1719 785
rect 1804 761 1824 781
rect 1907 765 1927 785
rect 2015 765 2035 785
rect 2118 761 2138 781
rect 133 692 151 710
rect 135 593 153 611
rect 321 522 341 542
rect 424 526 444 546
rect 534 522 554 542
rect 637 526 657 546
rect 742 522 762 542
rect 845 526 865 546
rect 953 526 973 546
rect 1056 522 1076 542
rect 133 410 151 428
rect 1333 341 1353 361
rect 1436 345 1456 365
rect 1546 341 1566 361
rect 1649 345 1669 365
rect 1754 341 1774 361
rect 1857 345 1877 365
rect 1965 345 1985 365
rect 2068 341 2088 361
rect 135 311 153 329
rect 140 209 158 227
rect 142 110 160 128
rect 320 107 340 127
rect 423 111 443 131
rect 533 107 553 127
rect 636 111 656 131
rect 741 107 761 127
rect 844 111 864 131
rect 952 111 972 131
rect 1055 107 1075 127
rect 138 -70 156 -52
rect 140 -169 158 -151
rect 1631 -203 1651 -183
rect 1734 -199 1754 -179
rect 1844 -203 1864 -183
rect 1947 -199 1967 -179
rect 2052 -203 2072 -183
rect 2155 -199 2175 -179
rect 2263 -199 2283 -179
rect 2366 -203 2386 -183
rect 136 -284 154 -266
rect 138 -383 156 -365
rect 324 -454 344 -434
rect 427 -450 447 -430
rect 537 -454 557 -434
rect 640 -450 660 -430
rect 745 -454 765 -434
rect 848 -450 868 -430
rect 956 -450 976 -430
rect 1059 -454 1079 -434
rect 136 -566 154 -548
rect 1336 -635 1356 -615
rect 1439 -631 1459 -611
rect 1549 -635 1569 -615
rect 1652 -631 1672 -611
rect 1757 -635 1777 -615
rect 1860 -631 1880 -611
rect 1968 -631 1988 -611
rect 2071 -635 2091 -615
rect 138 -665 156 -647
rect 143 -767 161 -749
rect 145 -866 163 -848
rect 323 -869 343 -849
rect 426 -865 446 -845
rect 536 -869 556 -849
rect 639 -865 659 -845
rect 744 -869 764 -849
rect 847 -865 867 -845
rect 955 -865 975 -845
rect 1058 -869 1078 -849
rect 143 -1051 161 -1033
rect 145 -1150 163 -1132
rect 1391 -1196 1411 -1176
rect 1494 -1192 1514 -1172
rect 1604 -1196 1624 -1176
rect 1707 -1192 1727 -1172
rect 1812 -1196 1832 -1176
rect 1915 -1192 1935 -1172
rect 2023 -1192 2043 -1172
rect 2126 -1196 2146 -1176
rect 141 -1265 159 -1247
rect 143 -1364 161 -1346
rect 329 -1435 349 -1415
rect 432 -1431 452 -1411
rect 542 -1435 562 -1415
rect 645 -1431 665 -1411
rect 750 -1435 770 -1415
rect 853 -1431 873 -1411
rect 961 -1431 981 -1411
rect 1064 -1435 1084 -1415
rect 141 -1547 159 -1529
rect 1341 -1616 1361 -1596
rect 1444 -1612 1464 -1592
rect 1554 -1616 1574 -1596
rect 1657 -1612 1677 -1592
rect 1762 -1616 1782 -1596
rect 1865 -1612 1885 -1592
rect 1973 -1612 1993 -1592
rect 2076 -1616 2096 -1596
rect 143 -1646 161 -1628
rect 148 -1748 166 -1730
rect 150 -1847 168 -1829
rect 328 -1850 348 -1830
rect 431 -1846 451 -1826
rect 541 -1850 561 -1830
rect 644 -1846 664 -1826
rect 749 -1850 769 -1830
rect 852 -1846 872 -1826
rect 960 -1846 980 -1826
rect 1063 -1850 1083 -1830
rect 150 -2030 168 -2012
rect 152 -2129 170 -2111
rect 1556 -2128 1576 -2108
rect 1659 -2124 1679 -2104
rect 1769 -2128 1789 -2108
rect 1872 -2124 1892 -2104
rect 1977 -2128 1997 -2108
rect 2080 -2124 2100 -2104
rect 2188 -2124 2208 -2104
rect 2291 -2128 2311 -2108
rect 148 -2244 166 -2226
rect 150 -2343 168 -2325
rect 336 -2414 356 -2394
rect 439 -2410 459 -2390
rect 549 -2414 569 -2394
rect 652 -2410 672 -2390
rect 757 -2414 777 -2394
rect 860 -2410 880 -2390
rect 968 -2410 988 -2390
rect 1071 -2414 1091 -2394
rect 148 -2526 166 -2508
rect 1348 -2595 1368 -2575
rect 1451 -2591 1471 -2571
rect 1561 -2595 1581 -2575
rect 1664 -2591 1684 -2571
rect 1769 -2595 1789 -2575
rect 1872 -2591 1892 -2571
rect 1980 -2591 2000 -2571
rect 2083 -2595 2103 -2575
rect 150 -2625 168 -2607
rect 155 -2727 173 -2709
rect 157 -2826 175 -2808
rect 335 -2829 355 -2809
rect 438 -2825 458 -2805
rect 548 -2829 568 -2809
rect 651 -2825 671 -2805
rect 756 -2829 776 -2809
rect 859 -2825 879 -2805
rect 967 -2825 987 -2805
rect 1070 -2829 1090 -2809
rect 155 -3011 173 -2993
rect 157 -3110 175 -3092
rect 1403 -3156 1423 -3136
rect 1506 -3152 1526 -3132
rect 1616 -3156 1636 -3136
rect 1719 -3152 1739 -3132
rect 1824 -3156 1844 -3136
rect 1927 -3152 1947 -3132
rect 2035 -3152 2055 -3132
rect 2138 -3156 2158 -3136
rect 153 -3225 171 -3207
rect 155 -3324 173 -3306
rect 341 -3395 361 -3375
rect 444 -3391 464 -3371
rect 554 -3395 574 -3375
rect 657 -3391 677 -3371
rect 762 -3395 782 -3375
rect 865 -3391 885 -3371
rect 973 -3391 993 -3371
rect 1076 -3395 1096 -3375
rect 153 -3507 171 -3489
rect 1353 -3576 1373 -3556
rect 1456 -3572 1476 -3552
rect 1566 -3576 1586 -3556
rect 1669 -3572 1689 -3552
rect 1774 -3576 1794 -3556
rect 1877 -3572 1897 -3552
rect 1985 -3572 2005 -3552
rect 2088 -3576 2108 -3556
rect 155 -3606 173 -3588
rect 160 -3708 178 -3690
rect 162 -3807 180 -3789
rect 340 -3810 360 -3790
rect 443 -3806 463 -3786
rect 553 -3810 573 -3790
rect 656 -3806 676 -3786
rect 761 -3810 781 -3790
rect 864 -3806 884 -3786
rect 972 -3806 992 -3786
rect 1075 -3810 1095 -3790
<< pdiffc >>
rect 310 3612 330 3632
rect 406 3612 426 3632
rect 523 3612 543 3632
rect 619 3612 639 3632
rect 731 3612 751 3632
rect 827 3612 847 3632
rect 937 3612 957 3632
rect 1033 3612 1053 3632
rect 1322 3431 1342 3451
rect 1418 3431 1438 3451
rect 1535 3431 1555 3451
rect 1631 3431 1651 3451
rect 1743 3431 1763 3451
rect 1839 3431 1859 3451
rect 1949 3431 1969 3451
rect 2045 3431 2065 3451
rect 309 3197 329 3217
rect 405 3197 425 3217
rect 522 3197 542 3217
rect 618 3197 638 3217
rect 730 3197 750 3217
rect 826 3197 846 3217
rect 936 3197 956 3217
rect 1032 3197 1052 3217
rect 1377 2870 1397 2890
rect 1473 2870 1493 2890
rect 1590 2870 1610 2890
rect 1686 2870 1706 2890
rect 1798 2870 1818 2890
rect 1894 2870 1914 2890
rect 2004 2870 2024 2890
rect 2100 2870 2120 2890
rect 315 2631 335 2651
rect 411 2631 431 2651
rect 528 2631 548 2651
rect 624 2631 644 2651
rect 736 2631 756 2651
rect 832 2631 852 2651
rect 942 2631 962 2651
rect 1038 2631 1058 2651
rect 1327 2450 1347 2470
rect 1423 2450 1443 2470
rect 1540 2450 1560 2470
rect 1636 2450 1656 2470
rect 1748 2450 1768 2470
rect 1844 2450 1864 2470
rect 1954 2450 1974 2470
rect 2050 2450 2070 2470
rect 314 2216 334 2236
rect 410 2216 430 2236
rect 527 2216 547 2236
rect 623 2216 643 2236
rect 735 2216 755 2236
rect 831 2216 851 2236
rect 941 2216 961 2236
rect 1037 2216 1057 2236
rect 1542 1938 1562 1958
rect 1638 1938 1658 1958
rect 1755 1938 1775 1958
rect 1851 1938 1871 1958
rect 1963 1938 1983 1958
rect 2059 1938 2079 1958
rect 2169 1938 2189 1958
rect 2265 1938 2285 1958
rect 322 1652 342 1672
rect 418 1652 438 1672
rect 535 1652 555 1672
rect 631 1652 651 1672
rect 743 1652 763 1672
rect 839 1652 859 1672
rect 949 1652 969 1672
rect 1045 1652 1065 1672
rect 1334 1471 1354 1491
rect 1430 1471 1450 1491
rect 1547 1471 1567 1491
rect 1643 1471 1663 1491
rect 1755 1471 1775 1491
rect 1851 1471 1871 1491
rect 1961 1471 1981 1491
rect 2057 1471 2077 1491
rect 321 1237 341 1257
rect 417 1237 437 1257
rect 534 1237 554 1257
rect 630 1237 650 1257
rect 742 1237 762 1257
rect 838 1237 858 1257
rect 948 1237 968 1257
rect 1044 1237 1064 1257
rect 1389 910 1409 930
rect 1485 910 1505 930
rect 1602 910 1622 930
rect 1698 910 1718 930
rect 1810 910 1830 930
rect 1906 910 1926 930
rect 2016 910 2036 930
rect 2112 910 2132 930
rect 327 671 347 691
rect 423 671 443 691
rect 540 671 560 691
rect 636 671 656 691
rect 748 671 768 691
rect 844 671 864 691
rect 954 671 974 691
rect 1050 671 1070 691
rect 1339 490 1359 510
rect 1435 490 1455 510
rect 1552 490 1572 510
rect 1648 490 1668 510
rect 1760 490 1780 510
rect 1856 490 1876 510
rect 1966 490 1986 510
rect 2062 490 2082 510
rect 326 256 346 276
rect 422 256 442 276
rect 539 256 559 276
rect 635 256 655 276
rect 747 256 767 276
rect 843 256 863 276
rect 953 256 973 276
rect 1049 256 1069 276
rect 1637 -54 1657 -34
rect 1733 -54 1753 -34
rect 1850 -54 1870 -34
rect 1946 -54 1966 -34
rect 2058 -54 2078 -34
rect 2154 -54 2174 -34
rect 2264 -54 2284 -34
rect 2360 -54 2380 -34
rect 330 -305 350 -285
rect 426 -305 446 -285
rect 543 -305 563 -285
rect 639 -305 659 -285
rect 751 -305 771 -285
rect 847 -305 867 -285
rect 957 -305 977 -285
rect 1053 -305 1073 -285
rect 1342 -486 1362 -466
rect 1438 -486 1458 -466
rect 1555 -486 1575 -466
rect 1651 -486 1671 -466
rect 1763 -486 1783 -466
rect 1859 -486 1879 -466
rect 1969 -486 1989 -466
rect 2065 -486 2085 -466
rect 329 -720 349 -700
rect 425 -720 445 -700
rect 542 -720 562 -700
rect 638 -720 658 -700
rect 750 -720 770 -700
rect 846 -720 866 -700
rect 956 -720 976 -700
rect 1052 -720 1072 -700
rect 1397 -1047 1417 -1027
rect 1493 -1047 1513 -1027
rect 1610 -1047 1630 -1027
rect 1706 -1047 1726 -1027
rect 1818 -1047 1838 -1027
rect 1914 -1047 1934 -1027
rect 2024 -1047 2044 -1027
rect 2120 -1047 2140 -1027
rect 335 -1286 355 -1266
rect 431 -1286 451 -1266
rect 548 -1286 568 -1266
rect 644 -1286 664 -1266
rect 756 -1286 776 -1266
rect 852 -1286 872 -1266
rect 962 -1286 982 -1266
rect 1058 -1286 1078 -1266
rect 1347 -1467 1367 -1447
rect 1443 -1467 1463 -1447
rect 1560 -1467 1580 -1447
rect 1656 -1467 1676 -1447
rect 1768 -1467 1788 -1447
rect 1864 -1467 1884 -1447
rect 1974 -1467 1994 -1447
rect 2070 -1467 2090 -1447
rect 334 -1701 354 -1681
rect 430 -1701 450 -1681
rect 547 -1701 567 -1681
rect 643 -1701 663 -1681
rect 755 -1701 775 -1681
rect 851 -1701 871 -1681
rect 961 -1701 981 -1681
rect 1057 -1701 1077 -1681
rect 1562 -1979 1582 -1959
rect 1658 -1979 1678 -1959
rect 1775 -1979 1795 -1959
rect 1871 -1979 1891 -1959
rect 1983 -1979 2003 -1959
rect 2079 -1979 2099 -1959
rect 2189 -1979 2209 -1959
rect 2285 -1979 2305 -1959
rect 342 -2265 362 -2245
rect 438 -2265 458 -2245
rect 555 -2265 575 -2245
rect 651 -2265 671 -2245
rect 763 -2265 783 -2245
rect 859 -2265 879 -2245
rect 969 -2265 989 -2245
rect 1065 -2265 1085 -2245
rect 1354 -2446 1374 -2426
rect 1450 -2446 1470 -2426
rect 1567 -2446 1587 -2426
rect 1663 -2446 1683 -2426
rect 1775 -2446 1795 -2426
rect 1871 -2446 1891 -2426
rect 1981 -2446 2001 -2426
rect 2077 -2446 2097 -2426
rect 341 -2680 361 -2660
rect 437 -2680 457 -2660
rect 554 -2680 574 -2660
rect 650 -2680 670 -2660
rect 762 -2680 782 -2660
rect 858 -2680 878 -2660
rect 968 -2680 988 -2660
rect 1064 -2680 1084 -2660
rect 1409 -3007 1429 -2987
rect 1505 -3007 1525 -2987
rect 1622 -3007 1642 -2987
rect 1718 -3007 1738 -2987
rect 1830 -3007 1850 -2987
rect 1926 -3007 1946 -2987
rect 2036 -3007 2056 -2987
rect 2132 -3007 2152 -2987
rect 347 -3246 367 -3226
rect 443 -3246 463 -3226
rect 560 -3246 580 -3226
rect 656 -3246 676 -3226
rect 768 -3246 788 -3226
rect 864 -3246 884 -3226
rect 974 -3246 994 -3226
rect 1070 -3246 1090 -3226
rect 1359 -3427 1379 -3407
rect 1455 -3427 1475 -3407
rect 1572 -3427 1592 -3407
rect 1668 -3427 1688 -3407
rect 1780 -3427 1800 -3407
rect 1876 -3427 1896 -3407
rect 1986 -3427 2006 -3407
rect 2082 -3427 2102 -3407
rect 346 -3661 366 -3641
rect 442 -3661 462 -3641
rect 559 -3661 579 -3641
rect 655 -3661 675 -3641
rect 767 -3661 787 -3641
rect 863 -3661 883 -3641
rect 973 -3661 993 -3641
rect 1069 -3661 1089 -3641
<< poly >>
rect 342 3670 392 3683
rect 555 3670 605 3683
rect 763 3670 813 3683
rect 971 3670 1021 3683
rect 342 3542 392 3570
rect 342 3522 355 3542
rect 375 3522 392 3542
rect 342 3493 392 3522
rect 555 3541 605 3570
rect 555 3517 566 3541
rect 590 3517 605 3541
rect 555 3493 605 3517
rect 763 3546 813 3570
rect 763 3522 775 3546
rect 799 3522 813 3546
rect 763 3493 813 3522
rect 971 3544 1021 3570
rect 971 3518 989 3544
rect 1015 3518 1021 3544
rect 971 3493 1021 3518
rect 1354 3489 1404 3502
rect 1567 3489 1617 3502
rect 1775 3489 1825 3502
rect 1983 3489 2033 3502
rect 342 3435 392 3451
rect 555 3435 605 3451
rect 763 3435 813 3451
rect 971 3435 1021 3451
rect 1354 3361 1404 3389
rect 1354 3341 1367 3361
rect 1387 3341 1404 3361
rect 1354 3312 1404 3341
rect 1567 3360 1617 3389
rect 1567 3336 1578 3360
rect 1602 3336 1617 3360
rect 1567 3312 1617 3336
rect 1775 3365 1825 3389
rect 1775 3341 1787 3365
rect 1811 3341 1825 3365
rect 1775 3312 1825 3341
rect 1983 3363 2033 3389
rect 1983 3337 2001 3363
rect 2027 3337 2033 3363
rect 1983 3312 2033 3337
rect 341 3255 391 3268
rect 554 3255 604 3268
rect 762 3255 812 3268
rect 970 3255 1020 3268
rect 1354 3254 1404 3270
rect 1567 3254 1617 3270
rect 1775 3254 1825 3270
rect 1983 3254 2033 3270
rect 341 3127 391 3155
rect 341 3107 354 3127
rect 374 3107 391 3127
rect 341 3078 391 3107
rect 554 3126 604 3155
rect 554 3102 565 3126
rect 589 3102 604 3126
rect 554 3078 604 3102
rect 762 3131 812 3155
rect 762 3107 774 3131
rect 798 3107 812 3131
rect 762 3078 812 3107
rect 970 3129 1020 3155
rect 970 3103 988 3129
rect 1014 3103 1020 3129
rect 970 3078 1020 3103
rect 341 3020 391 3036
rect 554 3020 604 3036
rect 762 3020 812 3036
rect 970 3020 1020 3036
rect 1409 2928 1459 2941
rect 1622 2928 1672 2941
rect 1830 2928 1880 2941
rect 2038 2928 2088 2941
rect 1409 2800 1459 2828
rect 1409 2780 1422 2800
rect 1442 2780 1459 2800
rect 1409 2751 1459 2780
rect 1622 2799 1672 2828
rect 1622 2775 1633 2799
rect 1657 2775 1672 2799
rect 1622 2751 1672 2775
rect 1830 2804 1880 2828
rect 1830 2780 1842 2804
rect 1866 2780 1880 2804
rect 1830 2751 1880 2780
rect 2038 2802 2088 2828
rect 2038 2776 2056 2802
rect 2082 2776 2088 2802
rect 2038 2751 2088 2776
rect 347 2689 397 2702
rect 560 2689 610 2702
rect 768 2689 818 2702
rect 976 2689 1026 2702
rect 1409 2693 1459 2709
rect 1622 2693 1672 2709
rect 1830 2693 1880 2709
rect 2038 2693 2088 2709
rect 347 2561 397 2589
rect 347 2541 360 2561
rect 380 2541 397 2561
rect 347 2512 397 2541
rect 560 2560 610 2589
rect 560 2536 571 2560
rect 595 2536 610 2560
rect 560 2512 610 2536
rect 768 2565 818 2589
rect 768 2541 780 2565
rect 804 2541 818 2565
rect 768 2512 818 2541
rect 976 2563 1026 2589
rect 976 2537 994 2563
rect 1020 2537 1026 2563
rect 976 2512 1026 2537
rect 1359 2508 1409 2521
rect 1572 2508 1622 2521
rect 1780 2508 1830 2521
rect 1988 2508 2038 2521
rect 347 2454 397 2470
rect 560 2454 610 2470
rect 768 2454 818 2470
rect 976 2454 1026 2470
rect 1359 2380 1409 2408
rect 1359 2360 1372 2380
rect 1392 2360 1409 2380
rect 1359 2331 1409 2360
rect 1572 2379 1622 2408
rect 1572 2355 1583 2379
rect 1607 2355 1622 2379
rect 1572 2331 1622 2355
rect 1780 2384 1830 2408
rect 1780 2360 1792 2384
rect 1816 2360 1830 2384
rect 1780 2331 1830 2360
rect 1988 2382 2038 2408
rect 1988 2356 2006 2382
rect 2032 2356 2038 2382
rect 1988 2331 2038 2356
rect 346 2274 396 2287
rect 559 2274 609 2287
rect 767 2274 817 2287
rect 975 2274 1025 2287
rect 1359 2273 1409 2289
rect 1572 2273 1622 2289
rect 1780 2273 1830 2289
rect 1988 2273 2038 2289
rect 346 2146 396 2174
rect 346 2126 359 2146
rect 379 2126 396 2146
rect 346 2097 396 2126
rect 559 2145 609 2174
rect 559 2121 570 2145
rect 594 2121 609 2145
rect 559 2097 609 2121
rect 767 2150 817 2174
rect 767 2126 779 2150
rect 803 2126 817 2150
rect 767 2097 817 2126
rect 975 2148 1025 2174
rect 975 2122 993 2148
rect 1019 2122 1025 2148
rect 975 2097 1025 2122
rect 346 2039 396 2055
rect 559 2039 609 2055
rect 767 2039 817 2055
rect 975 2039 1025 2055
rect 1574 1996 1624 2009
rect 1787 1996 1837 2009
rect 1995 1996 2045 2009
rect 2203 1996 2253 2009
rect 1574 1868 1624 1896
rect 1574 1848 1587 1868
rect 1607 1848 1624 1868
rect 1574 1819 1624 1848
rect 1787 1867 1837 1896
rect 1787 1843 1798 1867
rect 1822 1843 1837 1867
rect 1787 1819 1837 1843
rect 1995 1872 2045 1896
rect 1995 1848 2007 1872
rect 2031 1848 2045 1872
rect 1995 1819 2045 1848
rect 2203 1870 2253 1896
rect 2203 1844 2221 1870
rect 2247 1844 2253 1870
rect 2203 1819 2253 1844
rect 1574 1761 1624 1777
rect 1787 1761 1837 1777
rect 1995 1761 2045 1777
rect 2203 1761 2253 1777
rect 354 1710 404 1723
rect 567 1710 617 1723
rect 775 1710 825 1723
rect 983 1710 1033 1723
rect 354 1582 404 1610
rect 354 1562 367 1582
rect 387 1562 404 1582
rect 354 1533 404 1562
rect 567 1581 617 1610
rect 567 1557 578 1581
rect 602 1557 617 1581
rect 567 1533 617 1557
rect 775 1586 825 1610
rect 775 1562 787 1586
rect 811 1562 825 1586
rect 775 1533 825 1562
rect 983 1584 1033 1610
rect 983 1558 1001 1584
rect 1027 1558 1033 1584
rect 983 1533 1033 1558
rect 1366 1529 1416 1542
rect 1579 1529 1629 1542
rect 1787 1529 1837 1542
rect 1995 1529 2045 1542
rect 354 1475 404 1491
rect 567 1475 617 1491
rect 775 1475 825 1491
rect 983 1475 1033 1491
rect 1366 1401 1416 1429
rect 1366 1381 1379 1401
rect 1399 1381 1416 1401
rect 1366 1352 1416 1381
rect 1579 1400 1629 1429
rect 1579 1376 1590 1400
rect 1614 1376 1629 1400
rect 1579 1352 1629 1376
rect 1787 1405 1837 1429
rect 1787 1381 1799 1405
rect 1823 1381 1837 1405
rect 1787 1352 1837 1381
rect 1995 1403 2045 1429
rect 1995 1377 2013 1403
rect 2039 1377 2045 1403
rect 1995 1352 2045 1377
rect 353 1295 403 1308
rect 566 1295 616 1308
rect 774 1295 824 1308
rect 982 1295 1032 1308
rect 1366 1294 1416 1310
rect 1579 1294 1629 1310
rect 1787 1294 1837 1310
rect 1995 1294 2045 1310
rect 353 1167 403 1195
rect 353 1147 366 1167
rect 386 1147 403 1167
rect 353 1118 403 1147
rect 566 1166 616 1195
rect 566 1142 577 1166
rect 601 1142 616 1166
rect 566 1118 616 1142
rect 774 1171 824 1195
rect 774 1147 786 1171
rect 810 1147 824 1171
rect 774 1118 824 1147
rect 982 1169 1032 1195
rect 982 1143 1000 1169
rect 1026 1143 1032 1169
rect 982 1118 1032 1143
rect 353 1060 403 1076
rect 566 1060 616 1076
rect 774 1060 824 1076
rect 982 1060 1032 1076
rect 1421 968 1471 981
rect 1634 968 1684 981
rect 1842 968 1892 981
rect 2050 968 2100 981
rect 1421 840 1471 868
rect 1421 820 1434 840
rect 1454 820 1471 840
rect 1421 791 1471 820
rect 1634 839 1684 868
rect 1634 815 1645 839
rect 1669 815 1684 839
rect 1634 791 1684 815
rect 1842 844 1892 868
rect 1842 820 1854 844
rect 1878 820 1892 844
rect 1842 791 1892 820
rect 2050 842 2100 868
rect 2050 816 2068 842
rect 2094 816 2100 842
rect 2050 791 2100 816
rect 359 729 409 742
rect 572 729 622 742
rect 780 729 830 742
rect 988 729 1038 742
rect 1421 733 1471 749
rect 1634 733 1684 749
rect 1842 733 1892 749
rect 2050 733 2100 749
rect 359 601 409 629
rect 359 581 372 601
rect 392 581 409 601
rect 359 552 409 581
rect 572 600 622 629
rect 572 576 583 600
rect 607 576 622 600
rect 572 552 622 576
rect 780 605 830 629
rect 780 581 792 605
rect 816 581 830 605
rect 780 552 830 581
rect 988 603 1038 629
rect 988 577 1006 603
rect 1032 577 1038 603
rect 988 552 1038 577
rect 1371 548 1421 561
rect 1584 548 1634 561
rect 1792 548 1842 561
rect 2000 548 2050 561
rect 359 494 409 510
rect 572 494 622 510
rect 780 494 830 510
rect 988 494 1038 510
rect 1371 420 1421 448
rect 1371 400 1384 420
rect 1404 400 1421 420
rect 1371 371 1421 400
rect 1584 419 1634 448
rect 1584 395 1595 419
rect 1619 395 1634 419
rect 1584 371 1634 395
rect 1792 424 1842 448
rect 1792 400 1804 424
rect 1828 400 1842 424
rect 1792 371 1842 400
rect 2000 422 2050 448
rect 2000 396 2018 422
rect 2044 396 2050 422
rect 2000 371 2050 396
rect 358 314 408 327
rect 571 314 621 327
rect 779 314 829 327
rect 987 314 1037 327
rect 1371 313 1421 329
rect 1584 313 1634 329
rect 1792 313 1842 329
rect 2000 313 2050 329
rect 358 186 408 214
rect 358 166 371 186
rect 391 166 408 186
rect 358 137 408 166
rect 571 185 621 214
rect 571 161 582 185
rect 606 161 621 185
rect 571 137 621 161
rect 779 190 829 214
rect 779 166 791 190
rect 815 166 829 190
rect 779 137 829 166
rect 987 188 1037 214
rect 987 162 1005 188
rect 1031 162 1037 188
rect 987 137 1037 162
rect 358 79 408 95
rect 571 79 621 95
rect 779 79 829 95
rect 987 79 1037 95
rect 1669 4 1719 17
rect 1882 4 1932 17
rect 2090 4 2140 17
rect 2298 4 2348 17
rect 1669 -124 1719 -96
rect 1669 -144 1682 -124
rect 1702 -144 1719 -124
rect 1669 -173 1719 -144
rect 1882 -125 1932 -96
rect 1882 -149 1893 -125
rect 1917 -149 1932 -125
rect 1882 -173 1932 -149
rect 2090 -120 2140 -96
rect 2090 -144 2102 -120
rect 2126 -144 2140 -120
rect 2090 -173 2140 -144
rect 2298 -122 2348 -96
rect 2298 -148 2316 -122
rect 2342 -148 2348 -122
rect 2298 -173 2348 -148
rect 1669 -231 1719 -215
rect 1882 -231 1932 -215
rect 2090 -231 2140 -215
rect 2298 -231 2348 -215
rect 362 -247 412 -234
rect 575 -247 625 -234
rect 783 -247 833 -234
rect 991 -247 1041 -234
rect 362 -375 412 -347
rect 362 -395 375 -375
rect 395 -395 412 -375
rect 362 -424 412 -395
rect 575 -376 625 -347
rect 575 -400 586 -376
rect 610 -400 625 -376
rect 575 -424 625 -400
rect 783 -371 833 -347
rect 783 -395 795 -371
rect 819 -395 833 -371
rect 783 -424 833 -395
rect 991 -373 1041 -347
rect 991 -399 1009 -373
rect 1035 -399 1041 -373
rect 991 -424 1041 -399
rect 1374 -428 1424 -415
rect 1587 -428 1637 -415
rect 1795 -428 1845 -415
rect 2003 -428 2053 -415
rect 362 -482 412 -466
rect 575 -482 625 -466
rect 783 -482 833 -466
rect 991 -482 1041 -466
rect 1374 -556 1424 -528
rect 1374 -576 1387 -556
rect 1407 -576 1424 -556
rect 1374 -605 1424 -576
rect 1587 -557 1637 -528
rect 1587 -581 1598 -557
rect 1622 -581 1637 -557
rect 1587 -605 1637 -581
rect 1795 -552 1845 -528
rect 1795 -576 1807 -552
rect 1831 -576 1845 -552
rect 1795 -605 1845 -576
rect 2003 -554 2053 -528
rect 2003 -580 2021 -554
rect 2047 -580 2053 -554
rect 2003 -605 2053 -580
rect 361 -662 411 -649
rect 574 -662 624 -649
rect 782 -662 832 -649
rect 990 -662 1040 -649
rect 1374 -663 1424 -647
rect 1587 -663 1637 -647
rect 1795 -663 1845 -647
rect 2003 -663 2053 -647
rect 361 -790 411 -762
rect 361 -810 374 -790
rect 394 -810 411 -790
rect 361 -839 411 -810
rect 574 -791 624 -762
rect 574 -815 585 -791
rect 609 -815 624 -791
rect 574 -839 624 -815
rect 782 -786 832 -762
rect 782 -810 794 -786
rect 818 -810 832 -786
rect 782 -839 832 -810
rect 990 -788 1040 -762
rect 990 -814 1008 -788
rect 1034 -814 1040 -788
rect 990 -839 1040 -814
rect 361 -897 411 -881
rect 574 -897 624 -881
rect 782 -897 832 -881
rect 990 -897 1040 -881
rect 1429 -989 1479 -976
rect 1642 -989 1692 -976
rect 1850 -989 1900 -976
rect 2058 -989 2108 -976
rect 1429 -1117 1479 -1089
rect 1429 -1137 1442 -1117
rect 1462 -1137 1479 -1117
rect 1429 -1166 1479 -1137
rect 1642 -1118 1692 -1089
rect 1642 -1142 1653 -1118
rect 1677 -1142 1692 -1118
rect 1642 -1166 1692 -1142
rect 1850 -1113 1900 -1089
rect 1850 -1137 1862 -1113
rect 1886 -1137 1900 -1113
rect 1850 -1166 1900 -1137
rect 2058 -1115 2108 -1089
rect 2058 -1141 2076 -1115
rect 2102 -1141 2108 -1115
rect 2058 -1166 2108 -1141
rect 367 -1228 417 -1215
rect 580 -1228 630 -1215
rect 788 -1228 838 -1215
rect 996 -1228 1046 -1215
rect 1429 -1224 1479 -1208
rect 1642 -1224 1692 -1208
rect 1850 -1224 1900 -1208
rect 2058 -1224 2108 -1208
rect 367 -1356 417 -1328
rect 367 -1376 380 -1356
rect 400 -1376 417 -1356
rect 367 -1405 417 -1376
rect 580 -1357 630 -1328
rect 580 -1381 591 -1357
rect 615 -1381 630 -1357
rect 580 -1405 630 -1381
rect 788 -1352 838 -1328
rect 788 -1376 800 -1352
rect 824 -1376 838 -1352
rect 788 -1405 838 -1376
rect 996 -1354 1046 -1328
rect 996 -1380 1014 -1354
rect 1040 -1380 1046 -1354
rect 996 -1405 1046 -1380
rect 1379 -1409 1429 -1396
rect 1592 -1409 1642 -1396
rect 1800 -1409 1850 -1396
rect 2008 -1409 2058 -1396
rect 367 -1463 417 -1447
rect 580 -1463 630 -1447
rect 788 -1463 838 -1447
rect 996 -1463 1046 -1447
rect 1379 -1537 1429 -1509
rect 1379 -1557 1392 -1537
rect 1412 -1557 1429 -1537
rect 1379 -1586 1429 -1557
rect 1592 -1538 1642 -1509
rect 1592 -1562 1603 -1538
rect 1627 -1562 1642 -1538
rect 1592 -1586 1642 -1562
rect 1800 -1533 1850 -1509
rect 1800 -1557 1812 -1533
rect 1836 -1557 1850 -1533
rect 1800 -1586 1850 -1557
rect 2008 -1535 2058 -1509
rect 2008 -1561 2026 -1535
rect 2052 -1561 2058 -1535
rect 2008 -1586 2058 -1561
rect 366 -1643 416 -1630
rect 579 -1643 629 -1630
rect 787 -1643 837 -1630
rect 995 -1643 1045 -1630
rect 1379 -1644 1429 -1628
rect 1592 -1644 1642 -1628
rect 1800 -1644 1850 -1628
rect 2008 -1644 2058 -1628
rect 366 -1771 416 -1743
rect 366 -1791 379 -1771
rect 399 -1791 416 -1771
rect 366 -1820 416 -1791
rect 579 -1772 629 -1743
rect 579 -1796 590 -1772
rect 614 -1796 629 -1772
rect 579 -1820 629 -1796
rect 787 -1767 837 -1743
rect 787 -1791 799 -1767
rect 823 -1791 837 -1767
rect 787 -1820 837 -1791
rect 995 -1769 1045 -1743
rect 995 -1795 1013 -1769
rect 1039 -1795 1045 -1769
rect 995 -1820 1045 -1795
rect 366 -1878 416 -1862
rect 579 -1878 629 -1862
rect 787 -1878 837 -1862
rect 995 -1878 1045 -1862
rect 1594 -1921 1644 -1908
rect 1807 -1921 1857 -1908
rect 2015 -1921 2065 -1908
rect 2223 -1921 2273 -1908
rect 1594 -2049 1644 -2021
rect 1594 -2069 1607 -2049
rect 1627 -2069 1644 -2049
rect 1594 -2098 1644 -2069
rect 1807 -2050 1857 -2021
rect 1807 -2074 1818 -2050
rect 1842 -2074 1857 -2050
rect 1807 -2098 1857 -2074
rect 2015 -2045 2065 -2021
rect 2015 -2069 2027 -2045
rect 2051 -2069 2065 -2045
rect 2015 -2098 2065 -2069
rect 2223 -2047 2273 -2021
rect 2223 -2073 2241 -2047
rect 2267 -2073 2273 -2047
rect 2223 -2098 2273 -2073
rect 1594 -2156 1644 -2140
rect 1807 -2156 1857 -2140
rect 2015 -2156 2065 -2140
rect 2223 -2156 2273 -2140
rect 374 -2207 424 -2194
rect 587 -2207 637 -2194
rect 795 -2207 845 -2194
rect 1003 -2207 1053 -2194
rect 374 -2335 424 -2307
rect 374 -2355 387 -2335
rect 407 -2355 424 -2335
rect 374 -2384 424 -2355
rect 587 -2336 637 -2307
rect 587 -2360 598 -2336
rect 622 -2360 637 -2336
rect 587 -2384 637 -2360
rect 795 -2331 845 -2307
rect 795 -2355 807 -2331
rect 831 -2355 845 -2331
rect 795 -2384 845 -2355
rect 1003 -2333 1053 -2307
rect 1003 -2359 1021 -2333
rect 1047 -2359 1053 -2333
rect 1003 -2384 1053 -2359
rect 1386 -2388 1436 -2375
rect 1599 -2388 1649 -2375
rect 1807 -2388 1857 -2375
rect 2015 -2388 2065 -2375
rect 374 -2442 424 -2426
rect 587 -2442 637 -2426
rect 795 -2442 845 -2426
rect 1003 -2442 1053 -2426
rect 1386 -2516 1436 -2488
rect 1386 -2536 1399 -2516
rect 1419 -2536 1436 -2516
rect 1386 -2565 1436 -2536
rect 1599 -2517 1649 -2488
rect 1599 -2541 1610 -2517
rect 1634 -2541 1649 -2517
rect 1599 -2565 1649 -2541
rect 1807 -2512 1857 -2488
rect 1807 -2536 1819 -2512
rect 1843 -2536 1857 -2512
rect 1807 -2565 1857 -2536
rect 2015 -2514 2065 -2488
rect 2015 -2540 2033 -2514
rect 2059 -2540 2065 -2514
rect 2015 -2565 2065 -2540
rect 373 -2622 423 -2609
rect 586 -2622 636 -2609
rect 794 -2622 844 -2609
rect 1002 -2622 1052 -2609
rect 1386 -2623 1436 -2607
rect 1599 -2623 1649 -2607
rect 1807 -2623 1857 -2607
rect 2015 -2623 2065 -2607
rect 373 -2750 423 -2722
rect 373 -2770 386 -2750
rect 406 -2770 423 -2750
rect 373 -2799 423 -2770
rect 586 -2751 636 -2722
rect 586 -2775 597 -2751
rect 621 -2775 636 -2751
rect 586 -2799 636 -2775
rect 794 -2746 844 -2722
rect 794 -2770 806 -2746
rect 830 -2770 844 -2746
rect 794 -2799 844 -2770
rect 1002 -2748 1052 -2722
rect 1002 -2774 1020 -2748
rect 1046 -2774 1052 -2748
rect 1002 -2799 1052 -2774
rect 373 -2857 423 -2841
rect 586 -2857 636 -2841
rect 794 -2857 844 -2841
rect 1002 -2857 1052 -2841
rect 1441 -2949 1491 -2936
rect 1654 -2949 1704 -2936
rect 1862 -2949 1912 -2936
rect 2070 -2949 2120 -2936
rect 1441 -3077 1491 -3049
rect 1441 -3097 1454 -3077
rect 1474 -3097 1491 -3077
rect 1441 -3126 1491 -3097
rect 1654 -3078 1704 -3049
rect 1654 -3102 1665 -3078
rect 1689 -3102 1704 -3078
rect 1654 -3126 1704 -3102
rect 1862 -3073 1912 -3049
rect 1862 -3097 1874 -3073
rect 1898 -3097 1912 -3073
rect 1862 -3126 1912 -3097
rect 2070 -3075 2120 -3049
rect 2070 -3101 2088 -3075
rect 2114 -3101 2120 -3075
rect 2070 -3126 2120 -3101
rect 379 -3188 429 -3175
rect 592 -3188 642 -3175
rect 800 -3188 850 -3175
rect 1008 -3188 1058 -3175
rect 1441 -3184 1491 -3168
rect 1654 -3184 1704 -3168
rect 1862 -3184 1912 -3168
rect 2070 -3184 2120 -3168
rect 379 -3316 429 -3288
rect 379 -3336 392 -3316
rect 412 -3336 429 -3316
rect 379 -3365 429 -3336
rect 592 -3317 642 -3288
rect 592 -3341 603 -3317
rect 627 -3341 642 -3317
rect 592 -3365 642 -3341
rect 800 -3312 850 -3288
rect 800 -3336 812 -3312
rect 836 -3336 850 -3312
rect 800 -3365 850 -3336
rect 1008 -3314 1058 -3288
rect 1008 -3340 1026 -3314
rect 1052 -3340 1058 -3314
rect 1008 -3365 1058 -3340
rect 1391 -3369 1441 -3356
rect 1604 -3369 1654 -3356
rect 1812 -3369 1862 -3356
rect 2020 -3369 2070 -3356
rect 379 -3423 429 -3407
rect 592 -3423 642 -3407
rect 800 -3423 850 -3407
rect 1008 -3423 1058 -3407
rect 1391 -3497 1441 -3469
rect 1391 -3517 1404 -3497
rect 1424 -3517 1441 -3497
rect 1391 -3546 1441 -3517
rect 1604 -3498 1654 -3469
rect 1604 -3522 1615 -3498
rect 1639 -3522 1654 -3498
rect 1604 -3546 1654 -3522
rect 1812 -3493 1862 -3469
rect 1812 -3517 1824 -3493
rect 1848 -3517 1862 -3493
rect 1812 -3546 1862 -3517
rect 2020 -3495 2070 -3469
rect 2020 -3521 2038 -3495
rect 2064 -3521 2070 -3495
rect 2020 -3546 2070 -3521
rect 378 -3603 428 -3590
rect 591 -3603 641 -3590
rect 799 -3603 849 -3590
rect 1007 -3603 1057 -3590
rect 1391 -3604 1441 -3588
rect 1604 -3604 1654 -3588
rect 1812 -3604 1862 -3588
rect 2020 -3604 2070 -3588
rect 378 -3731 428 -3703
rect 378 -3751 391 -3731
rect 411 -3751 428 -3731
rect 378 -3780 428 -3751
rect 591 -3732 641 -3703
rect 591 -3756 602 -3732
rect 626 -3756 641 -3732
rect 591 -3780 641 -3756
rect 799 -3727 849 -3703
rect 799 -3751 811 -3727
rect 835 -3751 849 -3727
rect 799 -3780 849 -3751
rect 1007 -3729 1057 -3703
rect 1007 -3755 1025 -3729
rect 1051 -3755 1057 -3729
rect 1007 -3780 1057 -3755
rect 378 -3838 428 -3822
rect 591 -3838 641 -3822
rect 799 -3838 849 -3822
rect 1007 -3838 1057 -3822
<< polycont >>
rect 355 3522 375 3542
rect 566 3517 590 3541
rect 775 3522 799 3546
rect 989 3518 1015 3544
rect 1367 3341 1387 3361
rect 1578 3336 1602 3360
rect 1787 3341 1811 3365
rect 2001 3337 2027 3363
rect 354 3107 374 3127
rect 565 3102 589 3126
rect 774 3107 798 3131
rect 988 3103 1014 3129
rect 1422 2780 1442 2800
rect 1633 2775 1657 2799
rect 1842 2780 1866 2804
rect 2056 2776 2082 2802
rect 360 2541 380 2561
rect 571 2536 595 2560
rect 780 2541 804 2565
rect 994 2537 1020 2563
rect 1372 2360 1392 2380
rect 1583 2355 1607 2379
rect 1792 2360 1816 2384
rect 2006 2356 2032 2382
rect 359 2126 379 2146
rect 570 2121 594 2145
rect 779 2126 803 2150
rect 993 2122 1019 2148
rect 1587 1848 1607 1868
rect 1798 1843 1822 1867
rect 2007 1848 2031 1872
rect 2221 1844 2247 1870
rect 367 1562 387 1582
rect 578 1557 602 1581
rect 787 1562 811 1586
rect 1001 1558 1027 1584
rect 1379 1381 1399 1401
rect 1590 1376 1614 1400
rect 1799 1381 1823 1405
rect 2013 1377 2039 1403
rect 366 1147 386 1167
rect 577 1142 601 1166
rect 786 1147 810 1171
rect 1000 1143 1026 1169
rect 1434 820 1454 840
rect 1645 815 1669 839
rect 1854 820 1878 844
rect 2068 816 2094 842
rect 372 581 392 601
rect 583 576 607 600
rect 792 581 816 605
rect 1006 577 1032 603
rect 1384 400 1404 420
rect 1595 395 1619 419
rect 1804 400 1828 424
rect 2018 396 2044 422
rect 371 166 391 186
rect 582 161 606 185
rect 791 166 815 190
rect 1005 162 1031 188
rect 1682 -144 1702 -124
rect 1893 -149 1917 -125
rect 2102 -144 2126 -120
rect 2316 -148 2342 -122
rect 375 -395 395 -375
rect 586 -400 610 -376
rect 795 -395 819 -371
rect 1009 -399 1035 -373
rect 1387 -576 1407 -556
rect 1598 -581 1622 -557
rect 1807 -576 1831 -552
rect 2021 -580 2047 -554
rect 374 -810 394 -790
rect 585 -815 609 -791
rect 794 -810 818 -786
rect 1008 -814 1034 -788
rect 1442 -1137 1462 -1117
rect 1653 -1142 1677 -1118
rect 1862 -1137 1886 -1113
rect 2076 -1141 2102 -1115
rect 380 -1376 400 -1356
rect 591 -1381 615 -1357
rect 800 -1376 824 -1352
rect 1014 -1380 1040 -1354
rect 1392 -1557 1412 -1537
rect 1603 -1562 1627 -1538
rect 1812 -1557 1836 -1533
rect 2026 -1561 2052 -1535
rect 379 -1791 399 -1771
rect 590 -1796 614 -1772
rect 799 -1791 823 -1767
rect 1013 -1795 1039 -1769
rect 1607 -2069 1627 -2049
rect 1818 -2074 1842 -2050
rect 2027 -2069 2051 -2045
rect 2241 -2073 2267 -2047
rect 387 -2355 407 -2335
rect 598 -2360 622 -2336
rect 807 -2355 831 -2331
rect 1021 -2359 1047 -2333
rect 1399 -2536 1419 -2516
rect 1610 -2541 1634 -2517
rect 1819 -2536 1843 -2512
rect 2033 -2540 2059 -2514
rect 386 -2770 406 -2750
rect 597 -2775 621 -2751
rect 806 -2770 830 -2746
rect 1020 -2774 1046 -2748
rect 1454 -3097 1474 -3077
rect 1665 -3102 1689 -3078
rect 1874 -3097 1898 -3073
rect 2088 -3101 2114 -3075
rect 392 -3336 412 -3316
rect 603 -3341 627 -3317
rect 812 -3336 836 -3312
rect 1026 -3340 1052 -3314
rect 1404 -3517 1424 -3497
rect 1615 -3522 1639 -3498
rect 1824 -3517 1848 -3493
rect 2038 -3521 2064 -3495
rect 391 -3751 411 -3731
rect 602 -3756 626 -3732
rect 811 -3751 835 -3727
rect 1025 -3755 1051 -3729
<< ndiffres >>
rect 97 3865 154 3884
rect 97 3862 118 3865
rect 3 3847 118 3862
rect 136 3847 154 3865
rect 3 3824 154 3847
rect 3 3788 45 3824
rect 2 3787 102 3788
rect 2 3766 158 3787
rect 2 3748 120 3766
rect 138 3748 158 3766
rect 2 3744 158 3748
rect 97 3728 158 3744
rect 95 3651 152 3670
rect 95 3648 116 3651
rect 1 3633 116 3648
rect 134 3633 152 3651
rect 1 3610 152 3633
rect 1 3574 43 3610
rect 0 3573 100 3574
rect 0 3552 156 3573
rect 0 3534 118 3552
rect 136 3534 156 3552
rect 0 3530 156 3534
rect 95 3514 156 3530
rect 95 3369 152 3388
rect 95 3366 116 3369
rect 1 3351 116 3366
rect 134 3351 152 3369
rect 1 3328 152 3351
rect 1 3292 43 3328
rect 0 3291 100 3292
rect 0 3270 156 3291
rect 0 3252 118 3270
rect 136 3252 156 3270
rect 0 3248 156 3252
rect 95 3232 156 3248
rect 102 3168 159 3187
rect 102 3165 123 3168
rect 8 3150 123 3165
rect 141 3150 159 3168
rect 8 3127 159 3150
rect 8 3091 50 3127
rect 7 3090 107 3091
rect 7 3069 163 3090
rect 7 3051 125 3069
rect 143 3051 163 3069
rect 7 3047 163 3051
rect 102 3031 163 3047
rect 102 2884 159 2903
rect 102 2881 123 2884
rect 8 2866 123 2881
rect 141 2866 159 2884
rect 8 2843 159 2866
rect 8 2807 50 2843
rect 7 2806 107 2807
rect 7 2785 163 2806
rect 7 2767 125 2785
rect 143 2767 163 2785
rect 7 2763 163 2767
rect 102 2747 163 2763
rect 100 2670 157 2689
rect 100 2667 121 2670
rect 6 2652 121 2667
rect 139 2652 157 2670
rect 6 2629 157 2652
rect 6 2593 48 2629
rect 5 2592 105 2593
rect 5 2571 161 2592
rect 5 2553 123 2571
rect 141 2553 161 2571
rect 5 2549 161 2553
rect 100 2533 161 2549
rect 100 2388 157 2407
rect 100 2385 121 2388
rect 6 2370 121 2385
rect 139 2370 157 2388
rect 6 2347 157 2370
rect 6 2311 48 2347
rect 5 2310 105 2311
rect 5 2289 161 2310
rect 5 2271 123 2289
rect 141 2271 161 2289
rect 5 2267 161 2271
rect 100 2251 161 2267
rect 107 2187 164 2206
rect 107 2184 128 2187
rect 13 2169 128 2184
rect 146 2169 164 2187
rect 13 2146 164 2169
rect 13 2110 55 2146
rect 12 2109 112 2110
rect 12 2088 168 2109
rect 12 2070 130 2088
rect 148 2070 168 2088
rect 12 2066 168 2070
rect 107 2050 168 2066
rect 109 1905 166 1924
rect 109 1902 130 1905
rect 15 1887 130 1902
rect 148 1887 166 1905
rect 15 1864 166 1887
rect 15 1828 57 1864
rect 14 1827 114 1828
rect 14 1806 170 1827
rect 14 1788 132 1806
rect 150 1788 170 1806
rect 14 1784 170 1788
rect 109 1768 170 1784
rect 107 1691 164 1710
rect 107 1688 128 1691
rect 13 1673 128 1688
rect 146 1673 164 1691
rect 13 1650 164 1673
rect 13 1614 55 1650
rect 12 1613 112 1614
rect 12 1592 168 1613
rect 12 1574 130 1592
rect 148 1574 168 1592
rect 12 1570 168 1574
rect 107 1554 168 1570
rect 107 1409 164 1428
rect 107 1406 128 1409
rect 13 1391 128 1406
rect 146 1391 164 1409
rect 13 1368 164 1391
rect 13 1332 55 1368
rect 12 1331 112 1332
rect 12 1310 168 1331
rect 12 1292 130 1310
rect 148 1292 168 1310
rect 12 1288 168 1292
rect 107 1272 168 1288
rect 114 1208 171 1227
rect 114 1205 135 1208
rect 20 1190 135 1205
rect 153 1190 171 1208
rect 20 1167 171 1190
rect 20 1131 62 1167
rect 19 1130 119 1131
rect 19 1109 175 1130
rect 19 1091 137 1109
rect 155 1091 175 1109
rect 19 1087 175 1091
rect 114 1071 175 1087
rect 114 924 171 943
rect 114 921 135 924
rect 20 906 135 921
rect 153 906 171 924
rect 20 883 171 906
rect 20 847 62 883
rect 19 846 119 847
rect 19 825 175 846
rect 19 807 137 825
rect 155 807 175 825
rect 19 803 175 807
rect 114 787 175 803
rect 112 710 169 729
rect 112 707 133 710
rect 18 692 133 707
rect 151 692 169 710
rect 18 669 169 692
rect 18 633 60 669
rect 17 632 117 633
rect 17 611 173 632
rect 17 593 135 611
rect 153 593 173 611
rect 17 589 173 593
rect 112 573 173 589
rect 112 428 169 447
rect 112 425 133 428
rect 18 410 133 425
rect 151 410 169 428
rect 18 387 169 410
rect 18 351 60 387
rect 17 350 117 351
rect 17 329 173 350
rect 17 311 135 329
rect 153 311 173 329
rect 17 307 173 311
rect 112 291 173 307
rect 119 227 176 246
rect 119 224 140 227
rect 25 209 140 224
rect 158 209 176 227
rect 25 186 176 209
rect 25 150 67 186
rect 24 149 124 150
rect 24 128 180 149
rect 24 110 142 128
rect 160 110 180 128
rect 24 106 180 110
rect 119 90 180 106
rect 117 -52 174 -33
rect 117 -55 138 -52
rect 23 -70 138 -55
rect 156 -70 174 -52
rect 23 -93 174 -70
rect 23 -129 65 -93
rect 22 -130 122 -129
rect 22 -151 178 -130
rect 22 -169 140 -151
rect 158 -169 178 -151
rect 22 -173 178 -169
rect 117 -189 178 -173
rect 115 -266 172 -247
rect 115 -269 136 -266
rect 21 -284 136 -269
rect 154 -284 172 -266
rect 21 -307 172 -284
rect 21 -343 63 -307
rect 20 -344 120 -343
rect 20 -365 176 -344
rect 20 -383 138 -365
rect 156 -383 176 -365
rect 20 -387 176 -383
rect 115 -403 176 -387
rect 115 -548 172 -529
rect 115 -551 136 -548
rect 21 -566 136 -551
rect 154 -566 172 -548
rect 21 -589 172 -566
rect 21 -625 63 -589
rect 20 -626 120 -625
rect 20 -647 176 -626
rect 20 -665 138 -647
rect 156 -665 176 -647
rect 20 -669 176 -665
rect 115 -685 176 -669
rect 122 -749 179 -730
rect 122 -752 143 -749
rect 28 -767 143 -752
rect 161 -767 179 -749
rect 28 -790 179 -767
rect 28 -826 70 -790
rect 27 -827 127 -826
rect 27 -848 183 -827
rect 27 -866 145 -848
rect 163 -866 183 -848
rect 27 -870 183 -866
rect 122 -886 183 -870
rect 122 -1033 179 -1014
rect 122 -1036 143 -1033
rect 28 -1051 143 -1036
rect 161 -1051 179 -1033
rect 28 -1074 179 -1051
rect 28 -1110 70 -1074
rect 27 -1111 127 -1110
rect 27 -1132 183 -1111
rect 27 -1150 145 -1132
rect 163 -1150 183 -1132
rect 27 -1154 183 -1150
rect 122 -1170 183 -1154
rect 120 -1247 177 -1228
rect 120 -1250 141 -1247
rect 26 -1265 141 -1250
rect 159 -1265 177 -1247
rect 26 -1288 177 -1265
rect 26 -1324 68 -1288
rect 25 -1325 125 -1324
rect 25 -1346 181 -1325
rect 25 -1364 143 -1346
rect 161 -1364 181 -1346
rect 25 -1368 181 -1364
rect 120 -1384 181 -1368
rect 120 -1529 177 -1510
rect 120 -1532 141 -1529
rect 26 -1547 141 -1532
rect 159 -1547 177 -1529
rect 26 -1570 177 -1547
rect 26 -1606 68 -1570
rect 25 -1607 125 -1606
rect 25 -1628 181 -1607
rect 25 -1646 143 -1628
rect 161 -1646 181 -1628
rect 25 -1650 181 -1646
rect 120 -1666 181 -1650
rect 127 -1730 184 -1711
rect 127 -1733 148 -1730
rect 33 -1748 148 -1733
rect 166 -1748 184 -1730
rect 33 -1771 184 -1748
rect 33 -1807 75 -1771
rect 32 -1808 132 -1807
rect 32 -1829 188 -1808
rect 32 -1847 150 -1829
rect 168 -1847 188 -1829
rect 32 -1851 188 -1847
rect 127 -1867 188 -1851
rect 129 -2012 186 -1993
rect 129 -2015 150 -2012
rect 35 -2030 150 -2015
rect 168 -2030 186 -2012
rect 35 -2053 186 -2030
rect 35 -2089 77 -2053
rect 34 -2090 134 -2089
rect 34 -2111 190 -2090
rect 34 -2129 152 -2111
rect 170 -2129 190 -2111
rect 34 -2133 190 -2129
rect 129 -2149 190 -2133
rect 127 -2226 184 -2207
rect 127 -2229 148 -2226
rect 33 -2244 148 -2229
rect 166 -2244 184 -2226
rect 33 -2267 184 -2244
rect 33 -2303 75 -2267
rect 32 -2304 132 -2303
rect 32 -2325 188 -2304
rect 32 -2343 150 -2325
rect 168 -2343 188 -2325
rect 32 -2347 188 -2343
rect 127 -2363 188 -2347
rect 127 -2508 184 -2489
rect 127 -2511 148 -2508
rect 33 -2526 148 -2511
rect 166 -2526 184 -2508
rect 33 -2549 184 -2526
rect 33 -2585 75 -2549
rect 32 -2586 132 -2585
rect 32 -2607 188 -2586
rect 32 -2625 150 -2607
rect 168 -2625 188 -2607
rect 32 -2629 188 -2625
rect 127 -2645 188 -2629
rect 134 -2709 191 -2690
rect 134 -2712 155 -2709
rect 40 -2727 155 -2712
rect 173 -2727 191 -2709
rect 40 -2750 191 -2727
rect 40 -2786 82 -2750
rect 39 -2787 139 -2786
rect 39 -2808 195 -2787
rect 39 -2826 157 -2808
rect 175 -2826 195 -2808
rect 39 -2830 195 -2826
rect 134 -2846 195 -2830
rect 134 -2993 191 -2974
rect 134 -2996 155 -2993
rect 40 -3011 155 -2996
rect 173 -3011 191 -2993
rect 40 -3034 191 -3011
rect 40 -3070 82 -3034
rect 39 -3071 139 -3070
rect 39 -3092 195 -3071
rect 39 -3110 157 -3092
rect 175 -3110 195 -3092
rect 39 -3114 195 -3110
rect 134 -3130 195 -3114
rect 132 -3207 189 -3188
rect 132 -3210 153 -3207
rect 38 -3225 153 -3210
rect 171 -3225 189 -3207
rect 38 -3248 189 -3225
rect 38 -3284 80 -3248
rect 37 -3285 137 -3284
rect 37 -3306 193 -3285
rect 37 -3324 155 -3306
rect 173 -3324 193 -3306
rect 37 -3328 193 -3324
rect 132 -3344 193 -3328
rect 132 -3489 189 -3470
rect 132 -3492 153 -3489
rect 38 -3507 153 -3492
rect 171 -3507 189 -3489
rect 38 -3530 189 -3507
rect 38 -3566 80 -3530
rect 37 -3567 137 -3566
rect 37 -3588 193 -3567
rect 37 -3606 155 -3588
rect 173 -3606 193 -3588
rect 37 -3610 193 -3606
rect 132 -3626 193 -3610
rect 139 -3690 196 -3671
rect 139 -3693 160 -3690
rect 45 -3708 160 -3693
rect 178 -3708 196 -3690
rect 45 -3731 196 -3708
rect 45 -3767 87 -3731
rect 44 -3768 144 -3767
rect 44 -3789 200 -3768
rect 44 -3807 162 -3789
rect 180 -3807 200 -3789
rect 44 -3811 200 -3807
rect 139 -3827 200 -3811
<< locali >>
rect 110 3874 145 3922
rect 108 3865 145 3874
rect 108 3847 118 3865
rect 136 3847 145 3865
rect 108 3837 145 3847
rect 111 3773 148 3775
rect 111 3772 759 3773
rect 110 3766 759 3772
rect 110 3748 120 3766
rect 138 3752 759 3766
rect 138 3748 148 3752
rect 589 3751 759 3752
rect 110 3738 148 3748
rect 110 3660 145 3738
rect 722 3728 759 3751
rect 106 3651 145 3660
rect 106 3633 116 3651
rect 134 3633 145 3651
rect 106 3627 145 3633
rect 301 3703 551 3727
rect 301 3632 338 3703
rect 453 3642 484 3643
rect 106 3623 143 3627
rect 301 3612 310 3632
rect 330 3612 338 3632
rect 301 3602 338 3612
rect 397 3632 484 3642
rect 397 3612 406 3632
rect 426 3612 484 3632
rect 397 3603 484 3612
rect 397 3602 434 3603
rect 109 3552 146 3561
rect 107 3534 118 3552
rect 136 3534 146 3552
rect 453 3550 484 3603
rect 514 3632 551 3703
rect 722 3708 1115 3728
rect 1135 3708 1138 3728
rect 722 3703 1138 3708
rect 722 3702 1063 3703
rect 666 3642 697 3643
rect 514 3612 523 3632
rect 543 3612 551 3632
rect 514 3602 551 3612
rect 610 3635 697 3642
rect 610 3632 671 3635
rect 610 3612 619 3632
rect 639 3615 671 3632
rect 692 3615 697 3635
rect 639 3612 697 3615
rect 610 3605 697 3612
rect 722 3632 759 3702
rect 1025 3701 1062 3702
rect 874 3642 910 3643
rect 722 3612 731 3632
rect 751 3612 759 3632
rect 610 3603 666 3605
rect 610 3602 647 3603
rect 722 3602 759 3612
rect 818 3632 966 3642
rect 1066 3639 1162 3641
rect 818 3612 827 3632
rect 847 3612 937 3632
rect 957 3612 966 3632
rect 818 3603 966 3612
rect 1024 3632 1162 3639
rect 1024 3612 1033 3632
rect 1053 3612 1162 3632
rect 1024 3603 1162 3612
rect 818 3602 855 3603
rect 874 3551 910 3603
rect 929 3602 966 3603
rect 1025 3602 1062 3603
rect 345 3549 386 3550
rect 107 3385 146 3534
rect 237 3542 386 3549
rect 237 3522 355 3542
rect 375 3522 386 3542
rect 237 3514 386 3522
rect 453 3546 812 3550
rect 453 3541 775 3546
rect 453 3517 566 3541
rect 590 3522 775 3541
rect 799 3522 812 3546
rect 590 3517 812 3522
rect 453 3514 812 3517
rect 874 3514 909 3551
rect 977 3548 1077 3551
rect 977 3544 1044 3548
rect 977 3518 989 3544
rect 1015 3522 1044 3544
rect 1070 3522 1077 3548
rect 1015 3518 1077 3522
rect 977 3514 1077 3518
rect 453 3493 484 3514
rect 874 3493 910 3514
rect 296 3492 333 3493
rect 295 3483 333 3492
rect 295 3463 304 3483
rect 324 3463 333 3483
rect 295 3455 333 3463
rect 399 3487 484 3493
rect 509 3492 546 3493
rect 399 3467 407 3487
rect 427 3467 484 3487
rect 399 3459 484 3467
rect 508 3483 546 3492
rect 508 3463 517 3483
rect 537 3463 546 3483
rect 399 3458 435 3459
rect 508 3455 546 3463
rect 612 3487 697 3493
rect 717 3492 754 3493
rect 612 3467 620 3487
rect 640 3486 697 3487
rect 640 3467 669 3486
rect 612 3466 669 3467
rect 690 3466 697 3486
rect 612 3459 697 3466
rect 716 3483 754 3492
rect 716 3463 725 3483
rect 745 3463 754 3483
rect 612 3458 648 3459
rect 716 3455 754 3463
rect 820 3488 964 3493
rect 820 3487 885 3488
rect 820 3467 828 3487
rect 848 3467 885 3487
rect 907 3487 964 3488
rect 907 3467 936 3487
rect 956 3467 964 3487
rect 820 3459 964 3467
rect 820 3458 856 3459
rect 928 3458 964 3459
rect 1030 3492 1067 3493
rect 1030 3491 1068 3492
rect 1030 3483 1094 3491
rect 1030 3463 1039 3483
rect 1059 3469 1094 3483
rect 1114 3469 1117 3489
rect 1059 3464 1117 3469
rect 1059 3463 1094 3464
rect 296 3426 333 3455
rect 297 3424 333 3426
rect 509 3424 546 3455
rect 297 3402 546 3424
rect 717 3423 754 3455
rect 1030 3451 1094 3463
rect 1134 3425 1161 3603
rect 993 3423 1161 3425
rect 717 3397 1161 3423
rect 1313 3522 1563 3546
rect 1313 3451 1350 3522
rect 1465 3461 1496 3462
rect 1313 3431 1322 3451
rect 1342 3431 1350 3451
rect 1313 3421 1350 3431
rect 1409 3451 1496 3461
rect 1409 3431 1418 3451
rect 1438 3431 1496 3451
rect 1409 3422 1496 3431
rect 1409 3421 1446 3422
rect 717 3387 739 3397
rect 993 3396 1161 3397
rect 677 3385 739 3387
rect 107 3378 739 3385
rect 106 3369 739 3378
rect 1465 3369 1496 3422
rect 1526 3451 1563 3522
rect 1734 3527 2127 3547
rect 2147 3527 2150 3547
rect 1734 3522 2150 3527
rect 1734 3521 2075 3522
rect 1678 3461 1709 3462
rect 1526 3431 1535 3451
rect 1555 3431 1563 3451
rect 1526 3421 1563 3431
rect 1622 3454 1709 3461
rect 1622 3451 1683 3454
rect 1622 3431 1631 3451
rect 1651 3434 1683 3451
rect 1704 3434 1709 3454
rect 1651 3431 1709 3434
rect 1622 3424 1709 3431
rect 1734 3451 1771 3521
rect 2037 3520 2074 3521
rect 1886 3461 1922 3462
rect 1734 3431 1743 3451
rect 1763 3431 1771 3451
rect 1622 3422 1678 3424
rect 1622 3421 1659 3422
rect 1734 3421 1771 3431
rect 1830 3451 1978 3461
rect 2078 3458 2174 3460
rect 1830 3431 1839 3451
rect 1859 3431 1949 3451
rect 1969 3431 1978 3451
rect 1830 3422 1978 3431
rect 2036 3451 2174 3458
rect 2036 3431 2045 3451
rect 2065 3431 2174 3451
rect 2036 3422 2174 3431
rect 1830 3421 1867 3422
rect 1886 3370 1922 3422
rect 1941 3421 1978 3422
rect 2037 3421 2074 3422
rect 106 3351 116 3369
rect 134 3368 739 3369
rect 1357 3368 1398 3369
rect 134 3363 155 3368
rect 134 3351 146 3363
rect 1249 3361 1398 3368
rect 106 3343 146 3351
rect 189 3350 215 3351
rect 106 3341 143 3343
rect 189 3332 743 3350
rect 1249 3341 1367 3361
rect 1387 3341 1398 3361
rect 1249 3333 1398 3341
rect 1465 3365 1824 3369
rect 1465 3360 1787 3365
rect 1465 3336 1578 3360
rect 1602 3341 1787 3360
rect 1811 3341 1824 3365
rect 1602 3336 1824 3341
rect 1465 3333 1824 3336
rect 1886 3333 1921 3370
rect 1989 3367 2089 3370
rect 1989 3363 2056 3367
rect 1989 3337 2001 3363
rect 2027 3341 2056 3363
rect 2082 3341 2089 3367
rect 2027 3337 2089 3341
rect 1989 3333 2089 3337
rect 109 3273 146 3279
rect 189 3273 215 3332
rect 722 3313 743 3332
rect 109 3270 215 3273
rect 109 3252 118 3270
rect 136 3256 215 3270
rect 300 3288 550 3312
rect 136 3254 212 3256
rect 136 3252 146 3254
rect 109 3242 146 3252
rect 114 3177 145 3242
rect 300 3217 337 3288
rect 452 3227 483 3228
rect 300 3197 309 3217
rect 329 3197 337 3217
rect 300 3187 337 3197
rect 396 3217 483 3227
rect 396 3197 405 3217
rect 425 3197 483 3217
rect 396 3188 483 3197
rect 396 3187 433 3188
rect 113 3168 150 3177
rect 113 3150 123 3168
rect 141 3150 150 3168
rect 113 3140 150 3150
rect 452 3135 483 3188
rect 513 3217 550 3288
rect 721 3293 1114 3313
rect 1134 3293 1137 3313
rect 1465 3312 1496 3333
rect 1886 3312 1922 3333
rect 1308 3311 1345 3312
rect 721 3288 1137 3293
rect 1307 3302 1345 3311
rect 721 3287 1062 3288
rect 665 3227 696 3228
rect 513 3197 522 3217
rect 542 3197 550 3217
rect 513 3187 550 3197
rect 609 3220 696 3227
rect 609 3217 670 3220
rect 609 3197 618 3217
rect 638 3200 670 3217
rect 691 3200 696 3220
rect 638 3197 696 3200
rect 609 3190 696 3197
rect 721 3217 758 3287
rect 1024 3286 1061 3287
rect 1307 3282 1316 3302
rect 1336 3282 1345 3302
rect 1307 3274 1345 3282
rect 1411 3306 1496 3312
rect 1521 3311 1558 3312
rect 1411 3286 1419 3306
rect 1439 3286 1496 3306
rect 1411 3278 1496 3286
rect 1520 3302 1558 3311
rect 1520 3282 1529 3302
rect 1549 3282 1558 3302
rect 1411 3277 1447 3278
rect 1520 3274 1558 3282
rect 1624 3306 1709 3312
rect 1729 3311 1766 3312
rect 1624 3286 1632 3306
rect 1652 3305 1709 3306
rect 1652 3286 1681 3305
rect 1624 3285 1681 3286
rect 1702 3285 1709 3305
rect 1624 3278 1709 3285
rect 1728 3302 1766 3311
rect 1728 3282 1737 3302
rect 1757 3282 1766 3302
rect 1624 3277 1660 3278
rect 1728 3274 1766 3282
rect 1832 3306 1976 3312
rect 1832 3286 1840 3306
rect 1860 3286 1892 3306
rect 1916 3286 1948 3306
rect 1968 3286 1976 3306
rect 1832 3278 1976 3286
rect 1832 3277 1868 3278
rect 1940 3277 1976 3278
rect 2042 3311 2079 3312
rect 2042 3310 2080 3311
rect 2042 3302 2106 3310
rect 2042 3282 2051 3302
rect 2071 3288 2106 3302
rect 2126 3288 2129 3308
rect 2071 3283 2129 3288
rect 2071 3282 2106 3283
rect 1308 3245 1345 3274
rect 1309 3243 1345 3245
rect 1521 3243 1558 3274
rect 873 3227 909 3228
rect 721 3197 730 3217
rect 750 3197 758 3217
rect 609 3188 665 3190
rect 609 3187 646 3188
rect 721 3187 758 3197
rect 817 3217 965 3227
rect 1065 3224 1161 3226
rect 817 3197 826 3217
rect 846 3197 936 3217
rect 956 3197 965 3217
rect 817 3188 965 3197
rect 1023 3217 1161 3224
rect 1309 3221 1558 3243
rect 1729 3242 1766 3274
rect 2042 3270 2106 3282
rect 2146 3244 2173 3422
rect 2005 3242 2173 3244
rect 1729 3238 2173 3242
rect 1023 3197 1032 3217
rect 1052 3197 1161 3217
rect 1729 3219 1778 3238
rect 1798 3219 2173 3238
rect 1729 3216 2173 3219
rect 2005 3215 2173 3216
rect 1023 3188 1161 3197
rect 817 3187 854 3188
rect 873 3136 909 3188
rect 928 3187 965 3188
rect 1024 3187 1061 3188
rect 344 3134 385 3135
rect 236 3127 385 3134
rect 236 3107 354 3127
rect 374 3107 385 3127
rect 236 3099 385 3107
rect 452 3131 811 3135
rect 452 3126 774 3131
rect 452 3102 565 3126
rect 589 3107 774 3126
rect 798 3107 811 3131
rect 589 3102 811 3107
rect 452 3099 811 3102
rect 873 3099 908 3136
rect 976 3133 1076 3136
rect 976 3129 1043 3133
rect 976 3103 988 3129
rect 1014 3107 1043 3129
rect 1069 3107 1076 3133
rect 1014 3103 1076 3107
rect 976 3099 1076 3103
rect 452 3078 483 3099
rect 873 3078 909 3099
rect 116 3069 153 3078
rect 295 3077 332 3078
rect 116 3051 125 3069
rect 143 3051 153 3069
rect 116 3041 153 3051
rect 117 3006 153 3041
rect 294 3068 332 3077
rect 294 3048 303 3068
rect 323 3048 332 3068
rect 294 3040 332 3048
rect 398 3072 483 3078
rect 508 3077 545 3078
rect 398 3052 406 3072
rect 426 3052 483 3072
rect 398 3044 483 3052
rect 507 3068 545 3077
rect 507 3048 516 3068
rect 536 3048 545 3068
rect 398 3043 434 3044
rect 507 3040 545 3048
rect 611 3072 696 3078
rect 716 3077 753 3078
rect 611 3052 619 3072
rect 639 3071 696 3072
rect 639 3052 668 3071
rect 611 3051 668 3052
rect 689 3051 696 3071
rect 611 3044 696 3051
rect 715 3068 753 3077
rect 715 3048 724 3068
rect 744 3048 753 3068
rect 611 3043 647 3044
rect 715 3040 753 3048
rect 819 3072 963 3078
rect 819 3052 827 3072
rect 847 3071 935 3072
rect 847 3052 875 3071
rect 819 3050 875 3052
rect 897 3052 935 3071
rect 955 3052 963 3072
rect 897 3050 963 3052
rect 819 3044 963 3050
rect 819 3043 855 3044
rect 927 3043 963 3044
rect 1029 3077 1066 3078
rect 1029 3076 1067 3077
rect 1029 3068 1093 3076
rect 1029 3048 1038 3068
rect 1058 3054 1093 3068
rect 1113 3054 1116 3074
rect 1058 3049 1116 3054
rect 1058 3048 1093 3049
rect 295 3011 332 3040
rect 115 2965 153 3006
rect 296 3009 332 3011
rect 508 3009 545 3040
rect 296 2987 545 3009
rect 716 3008 753 3040
rect 1029 3036 1093 3048
rect 1133 3010 1160 3188
rect 992 3008 1160 3010
rect 716 2982 1160 3008
rect 717 2965 741 2982
rect 992 2981 1160 2982
rect 115 2947 742 2965
rect 1368 2961 1618 2985
rect 115 2941 153 2947
rect 115 2917 152 2941
rect 115 2893 150 2917
rect 113 2884 150 2893
rect 113 2866 123 2884
rect 141 2866 150 2884
rect 113 2856 150 2866
rect 1368 2890 1405 2961
rect 1520 2900 1551 2901
rect 1368 2870 1377 2890
rect 1397 2870 1405 2890
rect 1368 2860 1405 2870
rect 1464 2890 1551 2900
rect 1464 2870 1473 2890
rect 1493 2870 1551 2890
rect 1464 2861 1551 2870
rect 1464 2860 1501 2861
rect 1520 2808 1551 2861
rect 1581 2890 1618 2961
rect 1789 2966 2182 2986
rect 2202 2966 2205 2986
rect 1789 2961 2205 2966
rect 1789 2960 2130 2961
rect 1733 2900 1764 2901
rect 1581 2870 1590 2890
rect 1610 2870 1618 2890
rect 1581 2860 1618 2870
rect 1677 2893 1764 2900
rect 1677 2890 1738 2893
rect 1677 2870 1686 2890
rect 1706 2873 1738 2890
rect 1759 2873 1764 2893
rect 1706 2870 1764 2873
rect 1677 2863 1764 2870
rect 1789 2890 1826 2960
rect 2092 2959 2129 2960
rect 1941 2900 1977 2901
rect 1789 2870 1798 2890
rect 1818 2870 1826 2890
rect 1677 2861 1733 2863
rect 1677 2860 1714 2861
rect 1789 2860 1826 2870
rect 1885 2890 2033 2900
rect 2133 2897 2229 2899
rect 1885 2870 1894 2890
rect 1914 2870 2004 2890
rect 2024 2870 2033 2890
rect 1885 2861 2033 2870
rect 2091 2890 2229 2897
rect 2091 2870 2100 2890
rect 2120 2870 2229 2890
rect 2091 2861 2229 2870
rect 1885 2860 1922 2861
rect 1941 2809 1977 2861
rect 1996 2860 2033 2861
rect 2092 2860 2129 2861
rect 1412 2807 1453 2808
rect 1304 2800 1453 2807
rect 116 2792 153 2794
rect 116 2791 764 2792
rect 115 2785 764 2791
rect 115 2767 125 2785
rect 143 2771 764 2785
rect 1304 2780 1422 2800
rect 1442 2780 1453 2800
rect 1304 2772 1453 2780
rect 1520 2804 1879 2808
rect 1520 2799 1842 2804
rect 1520 2775 1633 2799
rect 1657 2780 1842 2799
rect 1866 2780 1879 2804
rect 1657 2775 1879 2780
rect 1520 2772 1879 2775
rect 1941 2772 1976 2809
rect 2044 2806 2144 2809
rect 2044 2802 2111 2806
rect 2044 2776 2056 2802
rect 2082 2780 2111 2802
rect 2137 2780 2144 2806
rect 2082 2776 2144 2780
rect 2044 2772 2144 2776
rect 143 2767 153 2771
rect 594 2770 764 2771
rect 115 2757 153 2767
rect 115 2679 150 2757
rect 727 2747 764 2770
rect 1520 2751 1551 2772
rect 1941 2751 1977 2772
rect 1363 2750 1400 2751
rect 111 2670 150 2679
rect 111 2652 121 2670
rect 139 2652 150 2670
rect 111 2646 150 2652
rect 306 2722 556 2746
rect 306 2651 343 2722
rect 458 2661 489 2662
rect 111 2642 148 2646
rect 306 2631 315 2651
rect 335 2631 343 2651
rect 306 2621 343 2631
rect 402 2651 489 2661
rect 402 2631 411 2651
rect 431 2631 489 2651
rect 402 2622 489 2631
rect 402 2621 439 2622
rect 114 2571 151 2580
rect 112 2553 123 2571
rect 141 2553 151 2571
rect 458 2569 489 2622
rect 519 2651 556 2722
rect 727 2727 1120 2747
rect 1140 2727 1143 2747
rect 727 2722 1143 2727
rect 1362 2741 1400 2750
rect 727 2721 1068 2722
rect 1362 2721 1371 2741
rect 1391 2721 1400 2741
rect 671 2661 702 2662
rect 519 2631 528 2651
rect 548 2631 556 2651
rect 519 2621 556 2631
rect 615 2654 702 2661
rect 615 2651 676 2654
rect 615 2631 624 2651
rect 644 2634 676 2651
rect 697 2634 702 2654
rect 644 2631 702 2634
rect 615 2624 702 2631
rect 727 2651 764 2721
rect 1030 2720 1067 2721
rect 1362 2713 1400 2721
rect 1466 2745 1551 2751
rect 1576 2750 1613 2751
rect 1466 2725 1474 2745
rect 1494 2725 1551 2745
rect 1466 2717 1551 2725
rect 1575 2741 1613 2750
rect 1575 2721 1584 2741
rect 1604 2721 1613 2741
rect 1466 2716 1502 2717
rect 1575 2713 1613 2721
rect 1679 2745 1764 2751
rect 1784 2750 1821 2751
rect 1679 2725 1687 2745
rect 1707 2744 1764 2745
rect 1707 2725 1736 2744
rect 1679 2724 1736 2725
rect 1757 2724 1764 2744
rect 1679 2717 1764 2724
rect 1783 2741 1821 2750
rect 1783 2721 1792 2741
rect 1812 2721 1821 2741
rect 1679 2716 1715 2717
rect 1783 2713 1821 2721
rect 1887 2745 2031 2751
rect 1887 2725 1895 2745
rect 1915 2743 2003 2745
rect 1915 2726 1951 2743
rect 1975 2726 2003 2743
rect 1915 2725 2003 2726
rect 2023 2725 2031 2745
rect 1887 2717 2031 2725
rect 1887 2716 1923 2717
rect 1995 2716 2031 2717
rect 2097 2750 2134 2751
rect 2097 2749 2135 2750
rect 2097 2741 2161 2749
rect 2097 2721 2106 2741
rect 2126 2727 2161 2741
rect 2181 2727 2184 2747
rect 2126 2722 2184 2727
rect 2126 2721 2161 2722
rect 1363 2684 1400 2713
rect 1364 2682 1400 2684
rect 1576 2682 1613 2713
rect 879 2661 915 2662
rect 727 2631 736 2651
rect 756 2631 764 2651
rect 615 2622 671 2624
rect 615 2621 652 2622
rect 727 2621 764 2631
rect 823 2651 971 2661
rect 1364 2660 1613 2682
rect 1784 2681 1821 2713
rect 2097 2709 2161 2721
rect 2201 2683 2228 2861
rect 2060 2681 2228 2683
rect 1784 2670 2228 2681
rect 1071 2658 1167 2660
rect 823 2631 832 2651
rect 852 2631 942 2651
rect 962 2631 971 2651
rect 823 2622 971 2631
rect 1029 2651 1167 2658
rect 1784 2655 2230 2670
rect 2060 2654 2230 2655
rect 1029 2631 1038 2651
rect 1058 2631 1167 2651
rect 1029 2622 1167 2631
rect 823 2621 860 2622
rect 879 2570 915 2622
rect 934 2621 971 2622
rect 1030 2621 1067 2622
rect 350 2568 391 2569
rect 112 2404 151 2553
rect 242 2561 391 2568
rect 242 2541 360 2561
rect 380 2541 391 2561
rect 242 2533 391 2541
rect 458 2565 817 2569
rect 458 2560 780 2565
rect 458 2536 571 2560
rect 595 2541 780 2560
rect 804 2541 817 2565
rect 595 2536 817 2541
rect 458 2533 817 2536
rect 879 2533 914 2570
rect 982 2567 1082 2570
rect 982 2563 1049 2567
rect 982 2537 994 2563
rect 1020 2541 1049 2563
rect 1075 2541 1082 2567
rect 1020 2537 1082 2541
rect 982 2533 1082 2537
rect 458 2512 489 2533
rect 879 2512 915 2533
rect 301 2511 338 2512
rect 300 2502 338 2511
rect 300 2482 309 2502
rect 329 2482 338 2502
rect 300 2474 338 2482
rect 404 2506 489 2512
rect 514 2511 551 2512
rect 404 2486 412 2506
rect 432 2486 489 2506
rect 404 2478 489 2486
rect 513 2502 551 2511
rect 513 2482 522 2502
rect 542 2482 551 2502
rect 404 2477 440 2478
rect 513 2474 551 2482
rect 617 2506 702 2512
rect 722 2511 759 2512
rect 617 2486 625 2506
rect 645 2505 702 2506
rect 645 2486 674 2505
rect 617 2485 674 2486
rect 695 2485 702 2505
rect 617 2478 702 2485
rect 721 2502 759 2511
rect 721 2482 730 2502
rect 750 2482 759 2502
rect 617 2477 653 2478
rect 721 2474 759 2482
rect 825 2507 969 2512
rect 825 2506 890 2507
rect 825 2486 833 2506
rect 853 2486 890 2506
rect 912 2506 969 2507
rect 912 2486 941 2506
rect 961 2486 969 2506
rect 825 2478 969 2486
rect 825 2477 861 2478
rect 933 2477 969 2478
rect 1035 2511 1072 2512
rect 1035 2510 1073 2511
rect 1035 2502 1099 2510
rect 1035 2482 1044 2502
rect 1064 2488 1099 2502
rect 1119 2488 1122 2508
rect 1064 2483 1122 2488
rect 1064 2482 1099 2483
rect 301 2445 338 2474
rect 302 2443 338 2445
rect 514 2443 551 2474
rect 302 2421 551 2443
rect 722 2442 759 2474
rect 1035 2470 1099 2482
rect 1139 2444 1166 2622
rect 998 2442 1166 2444
rect 722 2416 1166 2442
rect 1318 2541 1568 2565
rect 1318 2470 1355 2541
rect 1470 2480 1501 2481
rect 1318 2450 1327 2470
rect 1347 2450 1355 2470
rect 1318 2440 1355 2450
rect 1414 2470 1501 2480
rect 1414 2450 1423 2470
rect 1443 2450 1501 2470
rect 1414 2441 1501 2450
rect 1414 2440 1451 2441
rect 722 2406 744 2416
rect 998 2415 1166 2416
rect 682 2404 744 2406
rect 112 2397 744 2404
rect 111 2388 744 2397
rect 1470 2388 1501 2441
rect 1531 2470 1568 2541
rect 1739 2546 2132 2566
rect 2152 2546 2155 2566
rect 1739 2541 2155 2546
rect 1739 2540 2080 2541
rect 1683 2480 1714 2481
rect 1531 2450 1540 2470
rect 1560 2450 1568 2470
rect 1531 2440 1568 2450
rect 1627 2473 1714 2480
rect 1627 2470 1688 2473
rect 1627 2450 1636 2470
rect 1656 2453 1688 2470
rect 1709 2453 1714 2473
rect 1656 2450 1714 2453
rect 1627 2443 1714 2450
rect 1739 2470 1776 2540
rect 2042 2539 2079 2540
rect 1891 2480 1927 2481
rect 1739 2450 1748 2470
rect 1768 2450 1776 2470
rect 1627 2441 1683 2443
rect 1627 2440 1664 2441
rect 1739 2440 1776 2450
rect 1835 2470 1983 2480
rect 2083 2477 2179 2479
rect 1835 2450 1844 2470
rect 1864 2450 1954 2470
rect 1974 2450 1983 2470
rect 1835 2441 1983 2450
rect 2041 2470 2179 2477
rect 2041 2450 2050 2470
rect 2070 2450 2179 2470
rect 2041 2441 2179 2450
rect 1835 2440 1872 2441
rect 1891 2389 1927 2441
rect 1946 2440 1983 2441
rect 2042 2440 2079 2441
rect 111 2370 121 2388
rect 139 2387 744 2388
rect 1362 2387 1403 2388
rect 139 2382 160 2387
rect 139 2370 151 2382
rect 1254 2380 1403 2387
rect 111 2362 151 2370
rect 194 2369 220 2370
rect 111 2360 148 2362
rect 194 2351 748 2369
rect 1254 2360 1372 2380
rect 1392 2360 1403 2380
rect 1254 2352 1403 2360
rect 1470 2384 1829 2388
rect 1470 2379 1792 2384
rect 1470 2355 1583 2379
rect 1607 2360 1792 2379
rect 1816 2360 1829 2384
rect 1607 2355 1829 2360
rect 1470 2352 1829 2355
rect 1891 2352 1926 2389
rect 1994 2386 2094 2389
rect 1994 2382 2061 2386
rect 1994 2356 2006 2382
rect 2032 2360 2061 2382
rect 2087 2360 2094 2386
rect 2032 2356 2094 2360
rect 1994 2352 2094 2356
rect 114 2292 151 2298
rect 194 2292 220 2351
rect 727 2332 748 2351
rect 114 2289 220 2292
rect 114 2271 123 2289
rect 141 2275 220 2289
rect 305 2307 555 2331
rect 141 2273 217 2275
rect 141 2271 151 2273
rect 114 2261 151 2271
rect 119 2196 150 2261
rect 305 2236 342 2307
rect 457 2246 488 2247
rect 305 2216 314 2236
rect 334 2216 342 2236
rect 305 2206 342 2216
rect 401 2236 488 2246
rect 401 2216 410 2236
rect 430 2216 488 2236
rect 401 2207 488 2216
rect 401 2206 438 2207
rect 118 2187 155 2196
rect 118 2169 128 2187
rect 146 2169 155 2187
rect 118 2159 155 2169
rect 457 2154 488 2207
rect 518 2236 555 2307
rect 726 2312 1119 2332
rect 1139 2312 1142 2332
rect 1470 2331 1501 2352
rect 1891 2331 1927 2352
rect 1313 2330 1350 2331
rect 726 2307 1142 2312
rect 1312 2321 1350 2330
rect 726 2306 1067 2307
rect 670 2246 701 2247
rect 518 2216 527 2236
rect 547 2216 555 2236
rect 518 2206 555 2216
rect 614 2239 701 2246
rect 614 2236 675 2239
rect 614 2216 623 2236
rect 643 2219 675 2236
rect 696 2219 701 2239
rect 643 2216 701 2219
rect 614 2209 701 2216
rect 726 2236 763 2306
rect 1029 2305 1066 2306
rect 1312 2301 1321 2321
rect 1341 2301 1350 2321
rect 1312 2293 1350 2301
rect 1416 2325 1501 2331
rect 1526 2330 1563 2331
rect 1416 2305 1424 2325
rect 1444 2305 1501 2325
rect 1416 2297 1501 2305
rect 1525 2321 1563 2330
rect 1525 2301 1534 2321
rect 1554 2301 1563 2321
rect 1416 2296 1452 2297
rect 1525 2293 1563 2301
rect 1629 2325 1714 2331
rect 1734 2330 1771 2331
rect 1629 2305 1637 2325
rect 1657 2324 1714 2325
rect 1657 2305 1686 2324
rect 1629 2304 1686 2305
rect 1707 2304 1714 2324
rect 1629 2297 1714 2304
rect 1733 2321 1771 2330
rect 1733 2301 1742 2321
rect 1762 2301 1771 2321
rect 1629 2296 1665 2297
rect 1733 2293 1771 2301
rect 1837 2326 1981 2331
rect 1837 2325 1896 2326
rect 1837 2305 1845 2325
rect 1865 2306 1896 2325
rect 1920 2325 1981 2326
rect 1920 2306 1953 2325
rect 1865 2305 1953 2306
rect 1973 2305 1981 2325
rect 1837 2297 1981 2305
rect 1837 2296 1873 2297
rect 1945 2296 1981 2297
rect 2047 2330 2084 2331
rect 2047 2329 2085 2330
rect 2047 2321 2111 2329
rect 2047 2301 2056 2321
rect 2076 2307 2111 2321
rect 2131 2307 2134 2327
rect 2076 2302 2134 2307
rect 2076 2301 2111 2302
rect 1313 2264 1350 2293
rect 1314 2262 1350 2264
rect 1526 2262 1563 2293
rect 878 2246 914 2247
rect 726 2216 735 2236
rect 755 2216 763 2236
rect 614 2207 670 2209
rect 614 2206 651 2207
rect 726 2206 763 2216
rect 822 2236 970 2246
rect 1070 2243 1166 2245
rect 822 2216 831 2236
rect 851 2216 941 2236
rect 961 2216 970 2236
rect 822 2207 970 2216
rect 1028 2236 1166 2243
rect 1314 2240 1563 2262
rect 1734 2261 1771 2293
rect 2047 2289 2111 2301
rect 2151 2263 2178 2441
rect 2010 2261 2178 2263
rect 1734 2257 2178 2261
rect 1028 2216 1037 2236
rect 1057 2216 1166 2236
rect 1734 2238 1783 2257
rect 1803 2238 2178 2257
rect 1734 2235 2178 2238
rect 2010 2234 2178 2235
rect 2199 2260 2230 2654
rect 2199 2234 2204 2260
rect 2223 2234 2230 2260
rect 2199 2231 2230 2234
rect 1028 2207 1166 2216
rect 822 2206 859 2207
rect 878 2155 914 2207
rect 933 2206 970 2207
rect 1029 2206 1066 2207
rect 349 2153 390 2154
rect 241 2146 390 2153
rect 241 2126 359 2146
rect 379 2126 390 2146
rect 241 2118 390 2126
rect 457 2150 816 2154
rect 457 2145 779 2150
rect 457 2121 570 2145
rect 594 2126 779 2145
rect 803 2126 816 2150
rect 594 2121 816 2126
rect 457 2118 816 2121
rect 878 2118 913 2155
rect 981 2152 1081 2155
rect 981 2148 1048 2152
rect 981 2122 993 2148
rect 1019 2126 1048 2148
rect 1074 2126 1081 2152
rect 1019 2122 1081 2126
rect 981 2118 1081 2122
rect 457 2097 488 2118
rect 878 2097 914 2118
rect 121 2088 158 2097
rect 300 2096 337 2097
rect 121 2070 130 2088
rect 148 2070 158 2088
rect 121 2060 158 2070
rect 122 2025 158 2060
rect 299 2087 337 2096
rect 299 2067 308 2087
rect 328 2067 337 2087
rect 299 2059 337 2067
rect 403 2091 488 2097
rect 513 2096 550 2097
rect 403 2071 411 2091
rect 431 2071 488 2091
rect 403 2063 488 2071
rect 512 2087 550 2096
rect 512 2067 521 2087
rect 541 2067 550 2087
rect 403 2062 439 2063
rect 512 2059 550 2067
rect 616 2091 701 2097
rect 721 2096 758 2097
rect 616 2071 624 2091
rect 644 2090 701 2091
rect 644 2071 673 2090
rect 616 2070 673 2071
rect 694 2070 701 2090
rect 616 2063 701 2070
rect 720 2087 758 2096
rect 720 2067 729 2087
rect 749 2067 758 2087
rect 616 2062 652 2063
rect 720 2059 758 2067
rect 824 2091 968 2097
rect 824 2071 832 2091
rect 852 2090 940 2091
rect 852 2071 880 2090
rect 824 2069 880 2071
rect 902 2071 940 2090
rect 960 2071 968 2091
rect 902 2069 968 2071
rect 824 2063 968 2069
rect 824 2062 860 2063
rect 932 2062 968 2063
rect 1034 2096 1071 2097
rect 1034 2095 1072 2096
rect 1034 2087 1098 2095
rect 1034 2067 1043 2087
rect 1063 2073 1098 2087
rect 1118 2073 1121 2093
rect 1063 2068 1121 2073
rect 1063 2067 1098 2068
rect 300 2030 337 2059
rect 120 1984 158 2025
rect 301 2028 337 2030
rect 513 2028 550 2059
rect 301 2006 550 2028
rect 721 2027 758 2059
rect 1034 2055 1098 2067
rect 1138 2029 1165 2207
rect 997 2027 1165 2029
rect 721 2001 1165 2027
rect 722 1984 746 2001
rect 997 2000 1165 2001
rect 1533 2029 1783 2053
rect 120 1966 747 1984
rect 120 1960 158 1966
rect 122 1914 157 1960
rect 1533 1958 1570 2029
rect 1685 1968 1716 1969
rect 1533 1938 1542 1958
rect 1562 1938 1570 1958
rect 1533 1928 1570 1938
rect 1629 1958 1716 1968
rect 1629 1938 1638 1958
rect 1658 1938 1716 1958
rect 1629 1929 1716 1938
rect 1629 1928 1666 1929
rect 120 1905 157 1914
rect 120 1887 130 1905
rect 148 1887 157 1905
rect 120 1877 157 1887
rect 1685 1876 1716 1929
rect 1746 1958 1783 2029
rect 1954 2034 2347 2054
rect 2367 2034 2370 2054
rect 1954 2029 2370 2034
rect 1954 2028 2295 2029
rect 1898 1968 1929 1969
rect 1746 1938 1755 1958
rect 1775 1938 1783 1958
rect 1746 1928 1783 1938
rect 1842 1961 1929 1968
rect 1842 1958 1903 1961
rect 1842 1938 1851 1958
rect 1871 1941 1903 1958
rect 1924 1941 1929 1961
rect 1871 1938 1929 1941
rect 1842 1931 1929 1938
rect 1954 1958 1991 2028
rect 2257 2027 2294 2028
rect 2106 1968 2142 1969
rect 1954 1938 1963 1958
rect 1983 1938 1991 1958
rect 1842 1929 1898 1931
rect 1842 1928 1879 1929
rect 1954 1928 1991 1938
rect 2050 1958 2198 1968
rect 2298 1965 2394 1967
rect 2050 1938 2059 1958
rect 2079 1938 2169 1958
rect 2189 1938 2198 1958
rect 2050 1929 2198 1938
rect 2256 1958 2394 1965
rect 2256 1938 2265 1958
rect 2285 1938 2394 1958
rect 2256 1929 2394 1938
rect 2050 1928 2087 1929
rect 2106 1877 2142 1929
rect 2161 1928 2198 1929
rect 2257 1928 2294 1929
rect 1577 1875 1618 1876
rect 1469 1868 1618 1875
rect 1469 1848 1587 1868
rect 1607 1848 1618 1868
rect 1469 1840 1618 1848
rect 1685 1872 2044 1876
rect 1685 1867 2007 1872
rect 1685 1843 1798 1867
rect 1822 1848 2007 1867
rect 2031 1848 2044 1872
rect 1822 1843 2044 1848
rect 1685 1840 2044 1843
rect 2106 1840 2141 1877
rect 2209 1874 2309 1877
rect 2209 1870 2276 1874
rect 2209 1844 2221 1870
rect 2247 1848 2276 1870
rect 2302 1848 2309 1874
rect 2247 1844 2309 1848
rect 2209 1840 2309 1844
rect 1685 1819 1716 1840
rect 2106 1819 2142 1840
rect 1528 1818 1565 1819
rect 123 1813 160 1815
rect 123 1812 771 1813
rect 122 1806 771 1812
rect 122 1788 132 1806
rect 150 1792 771 1806
rect 150 1788 160 1792
rect 601 1791 771 1792
rect 122 1778 160 1788
rect 122 1700 157 1778
rect 734 1768 771 1791
rect 1527 1809 1565 1818
rect 1527 1789 1536 1809
rect 1556 1789 1565 1809
rect 1527 1781 1565 1789
rect 1631 1813 1716 1819
rect 1741 1818 1778 1819
rect 1631 1793 1639 1813
rect 1659 1793 1716 1813
rect 1631 1785 1716 1793
rect 1740 1809 1778 1818
rect 1740 1789 1749 1809
rect 1769 1789 1778 1809
rect 1631 1784 1667 1785
rect 1740 1781 1778 1789
rect 1844 1813 1929 1819
rect 1949 1818 1986 1819
rect 1844 1793 1852 1813
rect 1872 1812 1929 1813
rect 1872 1793 1901 1812
rect 1844 1792 1901 1793
rect 1922 1792 1929 1812
rect 1844 1785 1929 1792
rect 1948 1809 1986 1818
rect 1948 1789 1957 1809
rect 1977 1789 1986 1809
rect 1844 1784 1880 1785
rect 1948 1781 1986 1789
rect 2052 1817 2196 1819
rect 2052 1813 2110 1817
rect 2052 1793 2060 1813
rect 2080 1793 2110 1813
rect 2052 1791 2110 1793
rect 2135 1813 2196 1817
rect 2135 1793 2168 1813
rect 2188 1793 2196 1813
rect 2135 1791 2196 1793
rect 2052 1785 2196 1791
rect 2052 1784 2088 1785
rect 2160 1784 2196 1785
rect 2262 1818 2299 1819
rect 2262 1817 2300 1818
rect 2262 1809 2326 1817
rect 2262 1789 2271 1809
rect 2291 1795 2326 1809
rect 2346 1795 2349 1815
rect 2291 1790 2349 1795
rect 2291 1789 2326 1790
rect 118 1691 157 1700
rect 118 1673 128 1691
rect 146 1673 157 1691
rect 118 1667 157 1673
rect 313 1743 563 1767
rect 313 1672 350 1743
rect 465 1682 496 1683
rect 118 1663 155 1667
rect 313 1652 322 1672
rect 342 1652 350 1672
rect 313 1642 350 1652
rect 409 1672 496 1682
rect 409 1652 418 1672
rect 438 1652 496 1672
rect 409 1643 496 1652
rect 409 1642 446 1643
rect 121 1592 158 1601
rect 119 1574 130 1592
rect 148 1574 158 1592
rect 465 1590 496 1643
rect 526 1672 563 1743
rect 734 1748 1127 1768
rect 1147 1748 1150 1768
rect 1528 1752 1565 1781
rect 734 1743 1150 1748
rect 1529 1750 1565 1752
rect 1741 1750 1778 1781
rect 734 1742 1075 1743
rect 678 1682 709 1683
rect 526 1652 535 1672
rect 555 1652 563 1672
rect 526 1642 563 1652
rect 622 1675 709 1682
rect 622 1672 683 1675
rect 622 1652 631 1672
rect 651 1655 683 1672
rect 704 1655 709 1675
rect 651 1652 709 1655
rect 622 1645 709 1652
rect 734 1672 771 1742
rect 1037 1741 1074 1742
rect 1529 1728 1778 1750
rect 1949 1749 1986 1781
rect 2262 1777 2326 1789
rect 2366 1751 2393 1929
rect 2225 1749 2393 1751
rect 1949 1723 2393 1749
rect 2225 1722 2393 1723
rect 886 1682 922 1683
rect 734 1652 743 1672
rect 763 1652 771 1672
rect 622 1643 678 1645
rect 622 1642 659 1643
rect 734 1642 771 1652
rect 830 1672 978 1682
rect 1078 1679 1174 1681
rect 830 1652 839 1672
rect 859 1652 949 1672
rect 969 1652 978 1672
rect 830 1643 978 1652
rect 1036 1672 1174 1679
rect 1036 1652 1045 1672
rect 1065 1652 1174 1672
rect 1036 1643 1174 1652
rect 830 1642 867 1643
rect 886 1591 922 1643
rect 941 1642 978 1643
rect 1037 1642 1074 1643
rect 357 1589 398 1590
rect 119 1425 158 1574
rect 249 1582 398 1589
rect 249 1562 367 1582
rect 387 1562 398 1582
rect 249 1554 398 1562
rect 465 1586 824 1590
rect 465 1581 787 1586
rect 465 1557 578 1581
rect 602 1562 787 1581
rect 811 1562 824 1586
rect 602 1557 824 1562
rect 465 1554 824 1557
rect 886 1554 921 1591
rect 989 1588 1089 1591
rect 989 1584 1056 1588
rect 989 1558 1001 1584
rect 1027 1562 1056 1584
rect 1082 1562 1089 1588
rect 1027 1558 1089 1562
rect 989 1554 1089 1558
rect 465 1533 496 1554
rect 886 1533 922 1554
rect 308 1532 345 1533
rect 307 1523 345 1532
rect 307 1503 316 1523
rect 336 1503 345 1523
rect 307 1495 345 1503
rect 411 1527 496 1533
rect 521 1532 558 1533
rect 411 1507 419 1527
rect 439 1507 496 1527
rect 411 1499 496 1507
rect 520 1523 558 1532
rect 520 1503 529 1523
rect 549 1503 558 1523
rect 411 1498 447 1499
rect 520 1495 558 1503
rect 624 1527 709 1533
rect 729 1532 766 1533
rect 624 1507 632 1527
rect 652 1526 709 1527
rect 652 1507 681 1526
rect 624 1506 681 1507
rect 702 1506 709 1526
rect 624 1499 709 1506
rect 728 1523 766 1532
rect 728 1503 737 1523
rect 757 1503 766 1523
rect 624 1498 660 1499
rect 728 1495 766 1503
rect 832 1528 976 1533
rect 832 1527 897 1528
rect 832 1507 840 1527
rect 860 1507 897 1527
rect 919 1527 976 1528
rect 919 1507 948 1527
rect 968 1507 976 1527
rect 832 1499 976 1507
rect 832 1498 868 1499
rect 940 1498 976 1499
rect 1042 1532 1079 1533
rect 1042 1531 1080 1532
rect 1042 1523 1106 1531
rect 1042 1503 1051 1523
rect 1071 1509 1106 1523
rect 1126 1509 1129 1529
rect 1071 1504 1129 1509
rect 1071 1503 1106 1504
rect 308 1466 345 1495
rect 309 1464 345 1466
rect 521 1464 558 1495
rect 309 1442 558 1464
rect 729 1463 766 1495
rect 1042 1491 1106 1503
rect 1146 1465 1173 1643
rect 1005 1463 1173 1465
rect 729 1437 1173 1463
rect 1325 1562 1575 1586
rect 1325 1491 1362 1562
rect 1477 1501 1508 1502
rect 1325 1471 1334 1491
rect 1354 1471 1362 1491
rect 1325 1461 1362 1471
rect 1421 1491 1508 1501
rect 1421 1471 1430 1491
rect 1450 1471 1508 1491
rect 1421 1462 1508 1471
rect 1421 1461 1458 1462
rect 729 1427 751 1437
rect 1005 1436 1173 1437
rect 689 1425 751 1427
rect 119 1418 751 1425
rect 118 1409 751 1418
rect 1477 1409 1508 1462
rect 1538 1491 1575 1562
rect 1746 1567 2139 1587
rect 2159 1567 2162 1587
rect 1746 1562 2162 1567
rect 1746 1561 2087 1562
rect 1690 1501 1721 1502
rect 1538 1471 1547 1491
rect 1567 1471 1575 1491
rect 1538 1461 1575 1471
rect 1634 1494 1721 1501
rect 1634 1491 1695 1494
rect 1634 1471 1643 1491
rect 1663 1474 1695 1491
rect 1716 1474 1721 1494
rect 1663 1471 1721 1474
rect 1634 1464 1721 1471
rect 1746 1491 1783 1561
rect 2049 1560 2086 1561
rect 1898 1501 1934 1502
rect 1746 1471 1755 1491
rect 1775 1471 1783 1491
rect 1634 1462 1690 1464
rect 1634 1461 1671 1462
rect 1746 1461 1783 1471
rect 1842 1491 1990 1501
rect 2090 1498 2186 1500
rect 1842 1471 1851 1491
rect 1871 1471 1961 1491
rect 1981 1471 1990 1491
rect 1842 1462 1990 1471
rect 2048 1491 2186 1498
rect 2048 1471 2057 1491
rect 2077 1471 2186 1491
rect 2048 1462 2186 1471
rect 1842 1461 1879 1462
rect 1898 1410 1934 1462
rect 1953 1461 1990 1462
rect 2049 1461 2086 1462
rect 118 1391 128 1409
rect 146 1408 751 1409
rect 1369 1408 1410 1409
rect 146 1403 167 1408
rect 146 1391 158 1403
rect 1261 1401 1410 1408
rect 118 1383 158 1391
rect 201 1390 227 1391
rect 118 1381 155 1383
rect 201 1372 755 1390
rect 1261 1381 1379 1401
rect 1399 1381 1410 1401
rect 1261 1373 1410 1381
rect 1477 1405 1836 1409
rect 1477 1400 1799 1405
rect 1477 1376 1590 1400
rect 1614 1381 1799 1400
rect 1823 1381 1836 1405
rect 1614 1376 1836 1381
rect 1477 1373 1836 1376
rect 1898 1373 1933 1410
rect 2001 1407 2101 1410
rect 2001 1403 2068 1407
rect 2001 1377 2013 1403
rect 2039 1381 2068 1403
rect 2094 1381 2101 1407
rect 2039 1377 2101 1381
rect 2001 1373 2101 1377
rect 121 1313 158 1319
rect 201 1313 227 1372
rect 734 1353 755 1372
rect 121 1310 227 1313
rect 121 1292 130 1310
rect 148 1296 227 1310
rect 312 1328 562 1352
rect 148 1294 224 1296
rect 148 1292 158 1294
rect 121 1282 158 1292
rect 126 1217 157 1282
rect 312 1257 349 1328
rect 464 1267 495 1268
rect 312 1237 321 1257
rect 341 1237 349 1257
rect 312 1227 349 1237
rect 408 1257 495 1267
rect 408 1237 417 1257
rect 437 1237 495 1257
rect 408 1228 495 1237
rect 408 1227 445 1228
rect 125 1208 162 1217
rect 125 1190 135 1208
rect 153 1190 162 1208
rect 125 1180 162 1190
rect 464 1175 495 1228
rect 525 1257 562 1328
rect 733 1333 1126 1353
rect 1146 1333 1149 1353
rect 1477 1352 1508 1373
rect 1898 1352 1934 1373
rect 1320 1351 1357 1352
rect 733 1328 1149 1333
rect 1319 1342 1357 1351
rect 733 1327 1074 1328
rect 677 1267 708 1268
rect 525 1237 534 1257
rect 554 1237 562 1257
rect 525 1227 562 1237
rect 621 1260 708 1267
rect 621 1257 682 1260
rect 621 1237 630 1257
rect 650 1240 682 1257
rect 703 1240 708 1260
rect 650 1237 708 1240
rect 621 1230 708 1237
rect 733 1257 770 1327
rect 1036 1326 1073 1327
rect 1319 1322 1328 1342
rect 1348 1322 1357 1342
rect 1319 1314 1357 1322
rect 1423 1346 1508 1352
rect 1533 1351 1570 1352
rect 1423 1326 1431 1346
rect 1451 1326 1508 1346
rect 1423 1318 1508 1326
rect 1532 1342 1570 1351
rect 1532 1322 1541 1342
rect 1561 1322 1570 1342
rect 1423 1317 1459 1318
rect 1532 1314 1570 1322
rect 1636 1346 1721 1352
rect 1741 1351 1778 1352
rect 1636 1326 1644 1346
rect 1664 1345 1721 1346
rect 1664 1326 1693 1345
rect 1636 1325 1693 1326
rect 1714 1325 1721 1345
rect 1636 1318 1721 1325
rect 1740 1342 1778 1351
rect 1740 1322 1749 1342
rect 1769 1322 1778 1342
rect 1636 1317 1672 1318
rect 1740 1314 1778 1322
rect 1844 1346 1988 1352
rect 1844 1326 1852 1346
rect 1872 1326 1904 1346
rect 1928 1326 1960 1346
rect 1980 1326 1988 1346
rect 1844 1318 1988 1326
rect 1844 1317 1880 1318
rect 1952 1317 1988 1318
rect 2054 1351 2091 1352
rect 2054 1350 2092 1351
rect 2054 1342 2118 1350
rect 2054 1322 2063 1342
rect 2083 1328 2118 1342
rect 2138 1328 2141 1348
rect 2083 1323 2141 1328
rect 2083 1322 2118 1323
rect 1320 1285 1357 1314
rect 1321 1283 1357 1285
rect 1533 1283 1570 1314
rect 885 1267 921 1268
rect 733 1237 742 1257
rect 762 1237 770 1257
rect 621 1228 677 1230
rect 621 1227 658 1228
rect 733 1227 770 1237
rect 829 1257 977 1267
rect 1077 1264 1173 1266
rect 829 1237 838 1257
rect 858 1237 948 1257
rect 968 1237 977 1257
rect 829 1228 977 1237
rect 1035 1257 1173 1264
rect 1321 1261 1570 1283
rect 1741 1282 1778 1314
rect 2054 1310 2118 1322
rect 2158 1284 2185 1462
rect 2017 1282 2185 1284
rect 1741 1278 2185 1282
rect 1035 1237 1044 1257
rect 1064 1237 1173 1257
rect 1741 1259 1790 1278
rect 1810 1259 2185 1278
rect 1741 1256 2185 1259
rect 2017 1255 2185 1256
rect 1035 1228 1173 1237
rect 829 1227 866 1228
rect 885 1176 921 1228
rect 940 1227 977 1228
rect 1036 1227 1073 1228
rect 356 1174 397 1175
rect 248 1167 397 1174
rect 248 1147 366 1167
rect 386 1147 397 1167
rect 248 1139 397 1147
rect 464 1171 823 1175
rect 464 1166 786 1171
rect 464 1142 577 1166
rect 601 1147 786 1166
rect 810 1147 823 1171
rect 601 1142 823 1147
rect 464 1139 823 1142
rect 885 1139 920 1176
rect 988 1173 1088 1176
rect 988 1169 1055 1173
rect 988 1143 1000 1169
rect 1026 1147 1055 1169
rect 1081 1147 1088 1173
rect 1026 1143 1088 1147
rect 988 1139 1088 1143
rect 464 1118 495 1139
rect 885 1118 921 1139
rect 128 1109 165 1118
rect 307 1117 344 1118
rect 128 1091 137 1109
rect 155 1091 165 1109
rect 128 1081 165 1091
rect 129 1046 165 1081
rect 306 1108 344 1117
rect 306 1088 315 1108
rect 335 1088 344 1108
rect 306 1080 344 1088
rect 410 1112 495 1118
rect 520 1117 557 1118
rect 410 1092 418 1112
rect 438 1092 495 1112
rect 410 1084 495 1092
rect 519 1108 557 1117
rect 519 1088 528 1108
rect 548 1088 557 1108
rect 410 1083 446 1084
rect 519 1080 557 1088
rect 623 1112 708 1118
rect 728 1117 765 1118
rect 623 1092 631 1112
rect 651 1111 708 1112
rect 651 1092 680 1111
rect 623 1091 680 1092
rect 701 1091 708 1111
rect 623 1084 708 1091
rect 727 1108 765 1117
rect 727 1088 736 1108
rect 756 1088 765 1108
rect 623 1083 659 1084
rect 727 1080 765 1088
rect 831 1112 975 1118
rect 831 1092 839 1112
rect 859 1111 947 1112
rect 859 1092 887 1111
rect 831 1090 887 1092
rect 909 1092 947 1111
rect 967 1092 975 1112
rect 909 1090 975 1092
rect 831 1084 975 1090
rect 831 1083 867 1084
rect 939 1083 975 1084
rect 1041 1117 1078 1118
rect 1041 1116 1079 1117
rect 1041 1108 1105 1116
rect 1041 1088 1050 1108
rect 1070 1094 1105 1108
rect 1125 1094 1128 1114
rect 1070 1089 1128 1094
rect 1070 1088 1105 1089
rect 307 1051 344 1080
rect 127 1005 165 1046
rect 308 1049 344 1051
rect 520 1049 557 1080
rect 308 1027 557 1049
rect 728 1048 765 1080
rect 1041 1076 1105 1088
rect 1145 1050 1172 1228
rect 1004 1048 1172 1050
rect 728 1022 1172 1048
rect 729 1005 753 1022
rect 1004 1021 1172 1022
rect 127 987 754 1005
rect 1380 1001 1630 1025
rect 127 981 165 987
rect 127 957 164 981
rect 127 933 162 957
rect 125 924 162 933
rect 125 906 135 924
rect 153 906 162 924
rect 125 896 162 906
rect 1380 930 1417 1001
rect 1532 940 1563 941
rect 1380 910 1389 930
rect 1409 910 1417 930
rect 1380 900 1417 910
rect 1476 930 1563 940
rect 1476 910 1485 930
rect 1505 910 1563 930
rect 1476 901 1563 910
rect 1476 900 1513 901
rect 1532 848 1563 901
rect 1593 930 1630 1001
rect 1801 1006 2194 1026
rect 2214 1006 2217 1026
rect 1801 1001 2217 1006
rect 1801 1000 2142 1001
rect 1745 940 1776 941
rect 1593 910 1602 930
rect 1622 910 1630 930
rect 1593 900 1630 910
rect 1689 933 1776 940
rect 1689 930 1750 933
rect 1689 910 1698 930
rect 1718 913 1750 930
rect 1771 913 1776 933
rect 1718 910 1776 913
rect 1689 903 1776 910
rect 1801 930 1838 1000
rect 2104 999 2141 1000
rect 1953 940 1989 941
rect 1801 910 1810 930
rect 1830 910 1838 930
rect 1689 901 1745 903
rect 1689 900 1726 901
rect 1801 900 1838 910
rect 1897 930 2045 940
rect 2145 937 2241 939
rect 1897 910 1906 930
rect 1926 910 2016 930
rect 2036 910 2045 930
rect 1897 901 2045 910
rect 2103 930 2241 937
rect 2103 910 2112 930
rect 2132 910 2241 930
rect 2103 901 2241 910
rect 1897 900 1934 901
rect 1953 849 1989 901
rect 2008 900 2045 901
rect 2104 900 2141 901
rect 1424 847 1465 848
rect 1316 840 1465 847
rect 128 832 165 834
rect 128 831 776 832
rect 127 825 776 831
rect 127 807 137 825
rect 155 811 776 825
rect 1316 820 1434 840
rect 1454 820 1465 840
rect 1316 812 1465 820
rect 1532 844 1891 848
rect 1532 839 1854 844
rect 1532 815 1645 839
rect 1669 820 1854 839
rect 1878 820 1891 844
rect 1669 815 1891 820
rect 1532 812 1891 815
rect 1953 812 1988 849
rect 2056 846 2156 849
rect 2056 842 2123 846
rect 2056 816 2068 842
rect 2094 820 2123 842
rect 2149 820 2156 846
rect 2094 816 2156 820
rect 2056 812 2156 816
rect 155 807 165 811
rect 606 810 776 811
rect 127 797 165 807
rect 127 719 162 797
rect 739 787 776 810
rect 1532 791 1563 812
rect 1953 791 1989 812
rect 1375 790 1412 791
rect 123 710 162 719
rect 123 692 133 710
rect 151 692 162 710
rect 123 686 162 692
rect 318 762 568 786
rect 318 691 355 762
rect 470 701 501 702
rect 123 682 160 686
rect 318 671 327 691
rect 347 671 355 691
rect 318 661 355 671
rect 414 691 501 701
rect 414 671 423 691
rect 443 671 501 691
rect 414 662 501 671
rect 414 661 451 662
rect 126 611 163 620
rect 124 593 135 611
rect 153 593 163 611
rect 470 609 501 662
rect 531 691 568 762
rect 739 767 1132 787
rect 1152 767 1155 787
rect 739 762 1155 767
rect 1374 781 1412 790
rect 739 761 1080 762
rect 1374 761 1383 781
rect 1403 761 1412 781
rect 683 701 714 702
rect 531 671 540 691
rect 560 671 568 691
rect 531 661 568 671
rect 627 694 714 701
rect 627 691 688 694
rect 627 671 636 691
rect 656 674 688 691
rect 709 674 714 694
rect 656 671 714 674
rect 627 664 714 671
rect 739 691 776 761
rect 1042 760 1079 761
rect 1374 753 1412 761
rect 1478 785 1563 791
rect 1588 790 1625 791
rect 1478 765 1486 785
rect 1506 765 1563 785
rect 1478 757 1563 765
rect 1587 781 1625 790
rect 1587 761 1596 781
rect 1616 761 1625 781
rect 1478 756 1514 757
rect 1587 753 1625 761
rect 1691 785 1776 791
rect 1796 790 1833 791
rect 1691 765 1699 785
rect 1719 784 1776 785
rect 1719 765 1748 784
rect 1691 764 1748 765
rect 1769 764 1776 784
rect 1691 757 1776 764
rect 1795 781 1833 790
rect 1795 761 1804 781
rect 1824 761 1833 781
rect 1691 756 1727 757
rect 1795 753 1833 761
rect 1899 785 2043 791
rect 1899 765 1907 785
rect 1927 784 2015 785
rect 1927 765 1960 784
rect 1983 765 2015 784
rect 2035 765 2043 785
rect 1899 757 2043 765
rect 1899 756 1935 757
rect 2007 756 2043 757
rect 2109 790 2146 791
rect 2109 789 2147 790
rect 2109 781 2173 789
rect 2109 761 2118 781
rect 2138 767 2173 781
rect 2193 767 2196 787
rect 2138 762 2196 767
rect 2138 761 2173 762
rect 1375 724 1412 753
rect 1376 722 1412 724
rect 1588 722 1625 753
rect 891 701 927 702
rect 739 671 748 691
rect 768 671 776 691
rect 627 662 683 664
rect 627 661 664 662
rect 739 661 776 671
rect 835 691 983 701
rect 1376 700 1625 722
rect 1796 721 1833 753
rect 2109 749 2173 761
rect 2213 723 2240 901
rect 2072 721 2240 723
rect 1796 710 2240 721
rect 2303 721 2333 1722
rect 2303 716 2335 721
rect 1083 698 1179 700
rect 835 671 844 691
rect 864 671 954 691
rect 974 671 983 691
rect 835 662 983 671
rect 1041 691 1179 698
rect 1796 695 2242 710
rect 2072 694 2242 695
rect 1041 671 1050 691
rect 1070 671 1179 691
rect 1041 662 1179 671
rect 835 661 872 662
rect 891 610 927 662
rect 946 661 983 662
rect 1042 661 1079 662
rect 362 608 403 609
rect 124 444 163 593
rect 254 601 403 608
rect 254 581 372 601
rect 392 581 403 601
rect 254 573 403 581
rect 470 605 829 609
rect 470 600 792 605
rect 470 576 583 600
rect 607 581 792 600
rect 816 581 829 605
rect 607 576 829 581
rect 470 573 829 576
rect 891 573 926 610
rect 994 607 1094 610
rect 994 603 1061 607
rect 994 577 1006 603
rect 1032 581 1061 603
rect 1087 581 1094 607
rect 1032 577 1094 581
rect 994 573 1094 577
rect 470 552 501 573
rect 891 552 927 573
rect 313 551 350 552
rect 312 542 350 551
rect 312 522 321 542
rect 341 522 350 542
rect 312 514 350 522
rect 416 546 501 552
rect 526 551 563 552
rect 416 526 424 546
rect 444 526 501 546
rect 416 518 501 526
rect 525 542 563 551
rect 525 522 534 542
rect 554 522 563 542
rect 416 517 452 518
rect 525 514 563 522
rect 629 546 714 552
rect 734 551 771 552
rect 629 526 637 546
rect 657 545 714 546
rect 657 526 686 545
rect 629 525 686 526
rect 707 525 714 545
rect 629 518 714 525
rect 733 542 771 551
rect 733 522 742 542
rect 762 522 771 542
rect 629 517 665 518
rect 733 514 771 522
rect 837 547 981 552
rect 837 546 902 547
rect 837 526 845 546
rect 865 526 902 546
rect 924 546 981 547
rect 924 526 953 546
rect 973 526 981 546
rect 837 518 981 526
rect 837 517 873 518
rect 945 517 981 518
rect 1047 551 1084 552
rect 1047 550 1085 551
rect 1047 542 1111 550
rect 1047 522 1056 542
rect 1076 528 1111 542
rect 1131 528 1134 548
rect 1076 523 1134 528
rect 1076 522 1111 523
rect 313 485 350 514
rect 314 483 350 485
rect 526 483 563 514
rect 314 461 563 483
rect 734 482 771 514
rect 1047 510 1111 522
rect 1151 484 1178 662
rect 1010 482 1178 484
rect 734 456 1178 482
rect 1330 581 1580 605
rect 1330 510 1367 581
rect 1482 520 1513 521
rect 1330 490 1339 510
rect 1359 490 1367 510
rect 1330 480 1367 490
rect 1426 510 1513 520
rect 1426 490 1435 510
rect 1455 490 1513 510
rect 1426 481 1513 490
rect 1426 480 1463 481
rect 734 446 756 456
rect 1010 455 1178 456
rect 694 444 756 446
rect 124 437 756 444
rect 123 428 756 437
rect 1482 428 1513 481
rect 1543 510 1580 581
rect 1751 586 2144 606
rect 2164 586 2167 606
rect 1751 581 2167 586
rect 1751 580 2092 581
rect 1695 520 1726 521
rect 1543 490 1552 510
rect 1572 490 1580 510
rect 1543 480 1580 490
rect 1639 513 1726 520
rect 1639 510 1700 513
rect 1639 490 1648 510
rect 1668 493 1700 510
rect 1721 493 1726 513
rect 1668 490 1726 493
rect 1639 483 1726 490
rect 1751 510 1788 580
rect 2054 579 2091 580
rect 1903 520 1939 521
rect 1751 490 1760 510
rect 1780 490 1788 510
rect 1639 481 1695 483
rect 1639 480 1676 481
rect 1751 480 1788 490
rect 1847 510 1995 520
rect 2095 517 2191 519
rect 1847 490 1856 510
rect 1876 490 1966 510
rect 1986 490 1995 510
rect 1847 481 1995 490
rect 2053 510 2191 517
rect 2053 490 2062 510
rect 2082 490 2191 510
rect 2053 481 2191 490
rect 1847 480 1884 481
rect 1903 429 1939 481
rect 1958 480 1995 481
rect 2054 480 2091 481
rect 123 410 133 428
rect 151 427 756 428
rect 1374 427 1415 428
rect 151 422 172 427
rect 151 410 163 422
rect 1266 420 1415 427
rect 123 402 163 410
rect 206 409 232 410
rect 123 400 160 402
rect 206 391 760 409
rect 1266 400 1384 420
rect 1404 400 1415 420
rect 1266 392 1415 400
rect 1482 424 1841 428
rect 1482 419 1804 424
rect 1482 395 1595 419
rect 1619 400 1804 419
rect 1828 400 1841 424
rect 1619 395 1841 400
rect 1482 392 1841 395
rect 1903 392 1938 429
rect 2006 426 2106 429
rect 2006 422 2073 426
rect 2006 396 2018 422
rect 2044 400 2073 422
rect 2099 400 2106 426
rect 2044 396 2106 400
rect 2006 392 2106 396
rect 126 332 163 338
rect 206 332 232 391
rect 739 372 760 391
rect 126 329 232 332
rect 126 311 135 329
rect 153 315 232 329
rect 317 347 567 371
rect 153 313 229 315
rect 153 311 163 313
rect 126 301 163 311
rect 131 236 162 301
rect 317 276 354 347
rect 469 286 500 287
rect 317 256 326 276
rect 346 256 354 276
rect 317 246 354 256
rect 413 276 500 286
rect 413 256 422 276
rect 442 256 500 276
rect 413 247 500 256
rect 413 246 450 247
rect 130 227 167 236
rect 130 209 140 227
rect 158 209 167 227
rect 130 199 167 209
rect 469 194 500 247
rect 530 276 567 347
rect 738 352 1131 372
rect 1151 352 1154 372
rect 1482 371 1513 392
rect 1903 371 1939 392
rect 1325 370 1362 371
rect 738 347 1154 352
rect 1324 361 1362 370
rect 738 346 1079 347
rect 682 286 713 287
rect 530 256 539 276
rect 559 256 567 276
rect 530 246 567 256
rect 626 279 713 286
rect 626 276 687 279
rect 626 256 635 276
rect 655 259 687 276
rect 708 259 713 279
rect 655 256 713 259
rect 626 249 713 256
rect 738 276 775 346
rect 1041 345 1078 346
rect 1324 341 1333 361
rect 1353 341 1362 361
rect 1324 333 1362 341
rect 1428 365 1513 371
rect 1538 370 1575 371
rect 1428 345 1436 365
rect 1456 345 1513 365
rect 1428 337 1513 345
rect 1537 361 1575 370
rect 1537 341 1546 361
rect 1566 341 1575 361
rect 1428 336 1464 337
rect 1537 333 1575 341
rect 1641 365 1726 371
rect 1746 370 1783 371
rect 1641 345 1649 365
rect 1669 364 1726 365
rect 1669 345 1698 364
rect 1641 344 1698 345
rect 1719 344 1726 364
rect 1641 337 1726 344
rect 1745 361 1783 370
rect 1745 341 1754 361
rect 1774 341 1783 361
rect 1641 336 1677 337
rect 1745 333 1783 341
rect 1849 366 1993 371
rect 1849 365 1908 366
rect 1849 345 1857 365
rect 1877 346 1908 365
rect 1932 365 1993 366
rect 1932 346 1965 365
rect 1877 345 1965 346
rect 1985 345 1993 365
rect 1849 337 1993 345
rect 1849 336 1885 337
rect 1957 336 1993 337
rect 2059 370 2096 371
rect 2059 369 2097 370
rect 2059 361 2123 369
rect 2059 341 2068 361
rect 2088 347 2123 361
rect 2143 347 2146 367
rect 2088 342 2146 347
rect 2088 341 2123 342
rect 1325 304 1362 333
rect 1326 302 1362 304
rect 1538 302 1575 333
rect 890 286 926 287
rect 738 256 747 276
rect 767 256 775 276
rect 626 247 682 249
rect 626 246 663 247
rect 738 246 775 256
rect 834 276 982 286
rect 1082 283 1178 285
rect 834 256 843 276
rect 863 256 953 276
rect 973 256 982 276
rect 834 247 982 256
rect 1040 276 1178 283
rect 1326 280 1575 302
rect 1746 301 1783 333
rect 2059 329 2123 341
rect 2163 303 2190 481
rect 2022 301 2190 303
rect 1746 297 2190 301
rect 1040 256 1049 276
rect 1069 256 1178 276
rect 1746 278 1795 297
rect 1815 278 2190 297
rect 1746 275 2190 278
rect 2022 274 2190 275
rect 2211 300 2242 694
rect 2303 698 2308 716
rect 2328 698 2335 716
rect 2303 693 2335 698
rect 2306 691 2335 693
rect 2211 274 2216 300
rect 2235 274 2242 300
rect 2211 271 2242 274
rect 1040 247 1178 256
rect 834 246 871 247
rect 890 195 926 247
rect 945 246 982 247
rect 1041 246 1078 247
rect 361 193 402 194
rect 253 186 402 193
rect 253 166 371 186
rect 391 166 402 186
rect 253 158 402 166
rect 469 190 828 194
rect 469 185 791 190
rect 469 161 582 185
rect 606 166 791 185
rect 815 166 828 190
rect 606 161 828 166
rect 469 158 828 161
rect 890 158 925 195
rect 993 192 1093 195
rect 993 188 1060 192
rect 993 162 1005 188
rect 1031 166 1060 188
rect 1086 166 1093 192
rect 1031 162 1093 166
rect 993 158 1093 162
rect 469 137 500 158
rect 890 137 926 158
rect 133 128 170 137
rect 312 136 349 137
rect 133 110 142 128
rect 160 110 170 128
rect 133 100 170 110
rect 134 65 170 100
rect 311 127 349 136
rect 311 107 320 127
rect 340 107 349 127
rect 311 99 349 107
rect 415 131 500 137
rect 525 136 562 137
rect 415 111 423 131
rect 443 111 500 131
rect 415 103 500 111
rect 524 127 562 136
rect 524 107 533 127
rect 553 107 562 127
rect 415 102 451 103
rect 524 99 562 107
rect 628 131 713 137
rect 733 136 770 137
rect 628 111 636 131
rect 656 130 713 131
rect 656 111 685 130
rect 628 110 685 111
rect 706 110 713 130
rect 628 103 713 110
rect 732 127 770 136
rect 732 107 741 127
rect 761 107 770 127
rect 628 102 664 103
rect 732 99 770 107
rect 836 131 980 137
rect 836 111 844 131
rect 864 130 952 131
rect 864 111 892 130
rect 836 109 892 111
rect 914 111 952 130
rect 972 111 980 131
rect 914 109 980 111
rect 836 103 980 109
rect 836 102 872 103
rect 944 102 980 103
rect 1046 136 1083 137
rect 1046 135 1084 136
rect 1046 127 1110 135
rect 1046 107 1055 127
rect 1075 113 1110 127
rect 1130 113 1133 133
rect 1075 108 1133 113
rect 1075 107 1110 108
rect 312 70 349 99
rect 132 24 170 65
rect 313 68 349 70
rect 525 68 562 99
rect 313 46 562 68
rect 733 67 770 99
rect 1046 95 1110 107
rect 1150 69 1177 247
rect 1009 67 1177 69
rect 733 41 1177 67
rect 734 24 758 41
rect 1009 40 1177 41
rect 1628 37 1878 61
rect 132 6 759 24
rect 132 5 170 6
rect 130 0 170 5
rect 130 -43 165 0
rect 128 -52 165 -43
rect 128 -70 138 -52
rect 156 -70 165 -52
rect 1628 -34 1665 37
rect 1780 -24 1811 -23
rect 1628 -54 1637 -34
rect 1657 -54 1665 -34
rect 1628 -64 1665 -54
rect 1724 -34 1811 -24
rect 1724 -54 1733 -34
rect 1753 -54 1811 -34
rect 1724 -63 1811 -54
rect 1724 -64 1761 -63
rect 128 -80 165 -70
rect 1780 -116 1811 -63
rect 1841 -34 1878 37
rect 2049 42 2442 62
rect 2462 42 2465 62
rect 2049 37 2465 42
rect 2049 36 2390 37
rect 1993 -24 2024 -23
rect 1841 -54 1850 -34
rect 1870 -54 1878 -34
rect 1841 -64 1878 -54
rect 1937 -31 2024 -24
rect 1937 -34 1998 -31
rect 1937 -54 1946 -34
rect 1966 -51 1998 -34
rect 2019 -51 2024 -31
rect 1966 -54 2024 -51
rect 1937 -61 2024 -54
rect 2049 -34 2086 36
rect 2352 35 2389 36
rect 2201 -24 2237 -23
rect 2049 -54 2058 -34
rect 2078 -54 2086 -34
rect 1937 -63 1993 -61
rect 1937 -64 1974 -63
rect 2049 -64 2086 -54
rect 2145 -34 2293 -24
rect 2393 -27 2489 -25
rect 2145 -54 2154 -34
rect 2174 -54 2264 -34
rect 2284 -54 2293 -34
rect 2145 -63 2293 -54
rect 2351 -34 2489 -27
rect 2351 -54 2360 -34
rect 2380 -54 2489 -34
rect 2351 -63 2489 -54
rect 2145 -64 2182 -63
rect 2201 -115 2237 -63
rect 2256 -64 2293 -63
rect 2352 -64 2389 -63
rect 1672 -117 1713 -116
rect 1564 -124 1713 -117
rect 131 -144 168 -142
rect 1564 -144 1682 -124
rect 1702 -144 1713 -124
rect 131 -145 779 -144
rect 130 -151 779 -145
rect 130 -169 140 -151
rect 158 -165 779 -151
rect 1564 -152 1713 -144
rect 1780 -120 2139 -116
rect 1780 -125 2102 -120
rect 1780 -149 1893 -125
rect 1917 -144 2102 -125
rect 2126 -144 2139 -120
rect 1917 -149 2139 -144
rect 1780 -152 2139 -149
rect 2201 -152 2236 -115
rect 2304 -118 2404 -115
rect 2304 -122 2371 -118
rect 2304 -148 2316 -122
rect 2342 -144 2371 -122
rect 2397 -144 2404 -118
rect 2342 -148 2404 -144
rect 2304 -152 2404 -148
rect 158 -169 168 -165
rect 609 -166 779 -165
rect 130 -179 168 -169
rect 130 -257 165 -179
rect 742 -189 779 -166
rect 1780 -173 1811 -152
rect 2201 -173 2237 -152
rect 1623 -174 1660 -173
rect 1622 -183 1660 -174
rect 126 -266 165 -257
rect 126 -284 136 -266
rect 154 -284 165 -266
rect 126 -290 165 -284
rect 321 -214 571 -190
rect 321 -285 358 -214
rect 473 -275 504 -274
rect 126 -294 163 -290
rect 321 -305 330 -285
rect 350 -305 358 -285
rect 321 -315 358 -305
rect 417 -285 504 -275
rect 417 -305 426 -285
rect 446 -305 504 -285
rect 417 -314 504 -305
rect 417 -315 454 -314
rect 129 -365 166 -356
rect 127 -383 138 -365
rect 156 -383 166 -365
rect 473 -367 504 -314
rect 534 -285 571 -214
rect 742 -209 1135 -189
rect 1155 -209 1158 -189
rect 742 -214 1158 -209
rect 1622 -203 1631 -183
rect 1651 -203 1660 -183
rect 1622 -211 1660 -203
rect 1726 -179 1811 -173
rect 1836 -174 1873 -173
rect 1726 -199 1734 -179
rect 1754 -199 1811 -179
rect 1726 -207 1811 -199
rect 1835 -183 1873 -174
rect 1835 -203 1844 -183
rect 1864 -203 1873 -183
rect 1726 -208 1762 -207
rect 1835 -211 1873 -203
rect 1939 -179 2024 -173
rect 2044 -174 2081 -173
rect 1939 -199 1947 -179
rect 1967 -180 2024 -179
rect 1967 -199 1996 -180
rect 1939 -200 1996 -199
rect 2017 -200 2024 -180
rect 1939 -207 2024 -200
rect 2043 -183 2081 -174
rect 2043 -203 2052 -183
rect 2072 -203 2081 -183
rect 1939 -208 1975 -207
rect 2043 -211 2081 -203
rect 2147 -178 2291 -173
rect 2147 -179 2211 -178
rect 2147 -199 2155 -179
rect 2175 -197 2211 -179
rect 2237 -179 2291 -178
rect 2237 -197 2263 -179
rect 2175 -199 2263 -197
rect 2283 -199 2291 -179
rect 2147 -207 2291 -199
rect 2147 -208 2183 -207
rect 2255 -208 2291 -207
rect 2357 -174 2394 -173
rect 2357 -175 2395 -174
rect 2357 -183 2421 -175
rect 2357 -203 2366 -183
rect 2386 -197 2421 -183
rect 2441 -197 2444 -177
rect 2386 -202 2444 -197
rect 2386 -203 2421 -202
rect 742 -215 1083 -214
rect 686 -275 717 -274
rect 534 -305 543 -285
rect 563 -305 571 -285
rect 534 -315 571 -305
rect 630 -282 717 -275
rect 630 -285 691 -282
rect 630 -305 639 -285
rect 659 -302 691 -285
rect 712 -302 717 -282
rect 659 -305 717 -302
rect 630 -312 717 -305
rect 742 -285 779 -215
rect 1045 -216 1082 -215
rect 1623 -240 1660 -211
rect 1624 -242 1660 -240
rect 1836 -242 1873 -211
rect 1624 -264 1873 -242
rect 2044 -243 2081 -211
rect 2357 -215 2421 -203
rect 2461 -238 2488 -63
rect 2441 -241 2488 -238
rect 2320 -243 2488 -241
rect 2044 -269 2488 -243
rect 2320 -270 2488 -269
rect 894 -275 930 -274
rect 742 -305 751 -285
rect 771 -305 779 -285
rect 630 -314 686 -312
rect 630 -315 667 -314
rect 742 -315 779 -305
rect 838 -285 986 -275
rect 1086 -278 1182 -276
rect 838 -305 847 -285
rect 867 -305 957 -285
rect 977 -305 986 -285
rect 838 -314 986 -305
rect 1044 -285 1182 -278
rect 1044 -305 1053 -285
rect 1073 -305 1182 -285
rect 1044 -314 1182 -305
rect 838 -315 875 -314
rect 894 -366 930 -314
rect 949 -315 986 -314
rect 1045 -315 1082 -314
rect 365 -368 406 -367
rect 127 -532 166 -383
rect 257 -375 406 -368
rect 257 -395 375 -375
rect 395 -395 406 -375
rect 257 -403 406 -395
rect 473 -371 832 -367
rect 473 -376 795 -371
rect 473 -400 586 -376
rect 610 -395 795 -376
rect 819 -395 832 -371
rect 610 -400 832 -395
rect 473 -403 832 -400
rect 894 -403 929 -366
rect 997 -369 1097 -366
rect 997 -373 1064 -369
rect 997 -399 1009 -373
rect 1035 -395 1064 -373
rect 1090 -395 1097 -369
rect 1035 -399 1097 -395
rect 997 -403 1097 -399
rect 473 -424 504 -403
rect 894 -424 930 -403
rect 316 -425 353 -424
rect 315 -434 353 -425
rect 315 -454 324 -434
rect 344 -454 353 -434
rect 315 -462 353 -454
rect 419 -430 504 -424
rect 529 -425 566 -424
rect 419 -450 427 -430
rect 447 -450 504 -430
rect 419 -458 504 -450
rect 528 -434 566 -425
rect 528 -454 537 -434
rect 557 -454 566 -434
rect 419 -459 455 -458
rect 528 -462 566 -454
rect 632 -430 717 -424
rect 737 -425 774 -424
rect 632 -450 640 -430
rect 660 -431 717 -430
rect 660 -450 689 -431
rect 632 -451 689 -450
rect 710 -451 717 -431
rect 632 -458 717 -451
rect 736 -434 774 -425
rect 736 -454 745 -434
rect 765 -454 774 -434
rect 632 -459 668 -458
rect 736 -462 774 -454
rect 840 -429 984 -424
rect 840 -430 905 -429
rect 840 -450 848 -430
rect 868 -450 905 -430
rect 927 -430 984 -429
rect 927 -450 956 -430
rect 976 -450 984 -430
rect 840 -458 984 -450
rect 840 -459 876 -458
rect 948 -459 984 -458
rect 1050 -425 1087 -424
rect 1050 -426 1088 -425
rect 1050 -434 1114 -426
rect 1050 -454 1059 -434
rect 1079 -448 1114 -434
rect 1134 -448 1137 -428
rect 1079 -453 1137 -448
rect 1079 -454 1114 -453
rect 316 -491 353 -462
rect 317 -493 353 -491
rect 529 -493 566 -462
rect 317 -515 566 -493
rect 737 -494 774 -462
rect 1050 -466 1114 -454
rect 1154 -492 1181 -314
rect 1013 -494 1181 -492
rect 737 -520 1181 -494
rect 1333 -395 1583 -371
rect 1333 -466 1370 -395
rect 1485 -456 1516 -455
rect 1333 -486 1342 -466
rect 1362 -486 1370 -466
rect 1333 -496 1370 -486
rect 1429 -466 1516 -456
rect 1429 -486 1438 -466
rect 1458 -486 1516 -466
rect 1429 -495 1516 -486
rect 1429 -496 1466 -495
rect 737 -530 759 -520
rect 1013 -521 1181 -520
rect 697 -532 759 -530
rect 127 -539 759 -532
rect 126 -548 759 -539
rect 1485 -548 1516 -495
rect 1546 -466 1583 -395
rect 1754 -390 2147 -370
rect 2167 -390 2170 -370
rect 1754 -395 2170 -390
rect 1754 -396 2095 -395
rect 1698 -456 1729 -455
rect 1546 -486 1555 -466
rect 1575 -486 1583 -466
rect 1546 -496 1583 -486
rect 1642 -463 1729 -456
rect 1642 -466 1703 -463
rect 1642 -486 1651 -466
rect 1671 -483 1703 -466
rect 1724 -483 1729 -463
rect 1671 -486 1729 -483
rect 1642 -493 1729 -486
rect 1754 -466 1791 -396
rect 2057 -397 2094 -396
rect 1906 -456 1942 -455
rect 1754 -486 1763 -466
rect 1783 -486 1791 -466
rect 1642 -495 1698 -493
rect 1642 -496 1679 -495
rect 1754 -496 1791 -486
rect 1850 -466 1998 -456
rect 2098 -459 2194 -457
rect 1850 -486 1859 -466
rect 1879 -486 1969 -466
rect 1989 -486 1998 -466
rect 1850 -495 1998 -486
rect 2056 -466 2194 -459
rect 2056 -486 2065 -466
rect 2085 -486 2194 -466
rect 2056 -495 2194 -486
rect 1850 -496 1887 -495
rect 1906 -547 1942 -495
rect 1961 -496 1998 -495
rect 2057 -496 2094 -495
rect 126 -566 136 -548
rect 154 -549 759 -548
rect 1377 -549 1418 -548
rect 154 -554 175 -549
rect 154 -566 166 -554
rect 1269 -556 1418 -549
rect 126 -574 166 -566
rect 209 -567 235 -566
rect 126 -576 163 -574
rect 209 -585 763 -567
rect 1269 -576 1387 -556
rect 1407 -576 1418 -556
rect 1269 -584 1418 -576
rect 1485 -552 1844 -548
rect 1485 -557 1807 -552
rect 1485 -581 1598 -557
rect 1622 -576 1807 -557
rect 1831 -576 1844 -552
rect 1622 -581 1844 -576
rect 1485 -584 1844 -581
rect 1906 -584 1941 -547
rect 2009 -550 2109 -547
rect 2009 -554 2076 -550
rect 2009 -580 2021 -554
rect 2047 -576 2076 -554
rect 2102 -576 2109 -550
rect 2047 -580 2109 -576
rect 2009 -584 2109 -580
rect 129 -644 166 -638
rect 209 -644 235 -585
rect 742 -604 763 -585
rect 129 -647 235 -644
rect 129 -665 138 -647
rect 156 -661 235 -647
rect 320 -629 570 -605
rect 156 -663 232 -661
rect 156 -665 166 -663
rect 129 -675 166 -665
rect 134 -740 165 -675
rect 320 -700 357 -629
rect 472 -690 503 -689
rect 320 -720 329 -700
rect 349 -720 357 -700
rect 320 -730 357 -720
rect 416 -700 503 -690
rect 416 -720 425 -700
rect 445 -720 503 -700
rect 416 -729 503 -720
rect 416 -730 453 -729
rect 133 -749 170 -740
rect 133 -767 143 -749
rect 161 -767 170 -749
rect 133 -777 170 -767
rect 472 -782 503 -729
rect 533 -700 570 -629
rect 741 -624 1134 -604
rect 1154 -624 1157 -604
rect 1485 -605 1516 -584
rect 1906 -605 1942 -584
rect 1328 -606 1365 -605
rect 741 -629 1157 -624
rect 1327 -615 1365 -606
rect 741 -630 1082 -629
rect 685 -690 716 -689
rect 533 -720 542 -700
rect 562 -720 570 -700
rect 533 -730 570 -720
rect 629 -697 716 -690
rect 629 -700 690 -697
rect 629 -720 638 -700
rect 658 -717 690 -700
rect 711 -717 716 -697
rect 658 -720 716 -717
rect 629 -727 716 -720
rect 741 -700 778 -630
rect 1044 -631 1081 -630
rect 1327 -635 1336 -615
rect 1356 -635 1365 -615
rect 1327 -643 1365 -635
rect 1431 -611 1516 -605
rect 1541 -606 1578 -605
rect 1431 -631 1439 -611
rect 1459 -631 1516 -611
rect 1431 -639 1516 -631
rect 1540 -615 1578 -606
rect 1540 -635 1549 -615
rect 1569 -635 1578 -615
rect 1431 -640 1467 -639
rect 1540 -643 1578 -635
rect 1644 -611 1729 -605
rect 1749 -606 1786 -605
rect 1644 -631 1652 -611
rect 1672 -612 1729 -611
rect 1672 -631 1701 -612
rect 1644 -632 1701 -631
rect 1722 -632 1729 -612
rect 1644 -639 1729 -632
rect 1748 -615 1786 -606
rect 1748 -635 1757 -615
rect 1777 -635 1786 -615
rect 1644 -640 1680 -639
rect 1748 -643 1786 -635
rect 1852 -611 1996 -605
rect 1852 -631 1860 -611
rect 1880 -631 1912 -611
rect 1936 -631 1968 -611
rect 1988 -631 1996 -611
rect 1852 -639 1996 -631
rect 1852 -640 1888 -639
rect 1960 -640 1996 -639
rect 2062 -606 2099 -605
rect 2062 -607 2100 -606
rect 2062 -615 2126 -607
rect 2062 -635 2071 -615
rect 2091 -629 2126 -615
rect 2146 -629 2149 -609
rect 2091 -634 2149 -629
rect 2091 -635 2126 -634
rect 1328 -672 1365 -643
rect 1329 -674 1365 -672
rect 1541 -674 1578 -643
rect 893 -690 929 -689
rect 741 -720 750 -700
rect 770 -720 778 -700
rect 629 -729 685 -727
rect 629 -730 666 -729
rect 741 -730 778 -720
rect 837 -700 985 -690
rect 1085 -693 1181 -691
rect 837 -720 846 -700
rect 866 -720 956 -700
rect 976 -720 985 -700
rect 837 -729 985 -720
rect 1043 -700 1181 -693
rect 1329 -696 1578 -674
rect 1749 -675 1786 -643
rect 2062 -647 2126 -635
rect 2166 -673 2193 -495
rect 2025 -675 2193 -673
rect 1749 -679 2193 -675
rect 1043 -720 1052 -700
rect 1072 -720 1181 -700
rect 1749 -698 1798 -679
rect 1818 -698 2193 -679
rect 1749 -701 2193 -698
rect 2025 -702 2193 -701
rect 1043 -729 1181 -720
rect 837 -730 874 -729
rect 893 -781 929 -729
rect 948 -730 985 -729
rect 1044 -730 1081 -729
rect 364 -783 405 -782
rect 256 -790 405 -783
rect 256 -810 374 -790
rect 394 -810 405 -790
rect 256 -818 405 -810
rect 472 -786 831 -782
rect 472 -791 794 -786
rect 472 -815 585 -791
rect 609 -810 794 -791
rect 818 -810 831 -786
rect 609 -815 831 -810
rect 472 -818 831 -815
rect 893 -818 928 -781
rect 996 -784 1096 -781
rect 996 -788 1063 -784
rect 996 -814 1008 -788
rect 1034 -810 1063 -788
rect 1089 -810 1096 -784
rect 1034 -814 1096 -810
rect 996 -818 1096 -814
rect 472 -839 503 -818
rect 893 -839 929 -818
rect 136 -848 173 -839
rect 315 -840 352 -839
rect 136 -866 145 -848
rect 163 -866 173 -848
rect 136 -876 173 -866
rect 137 -911 173 -876
rect 314 -849 352 -840
rect 314 -869 323 -849
rect 343 -869 352 -849
rect 314 -877 352 -869
rect 418 -845 503 -839
rect 528 -840 565 -839
rect 418 -865 426 -845
rect 446 -865 503 -845
rect 418 -873 503 -865
rect 527 -849 565 -840
rect 527 -869 536 -849
rect 556 -869 565 -849
rect 418 -874 454 -873
rect 527 -877 565 -869
rect 631 -845 716 -839
rect 736 -840 773 -839
rect 631 -865 639 -845
rect 659 -846 716 -845
rect 659 -865 688 -846
rect 631 -866 688 -865
rect 709 -866 716 -846
rect 631 -873 716 -866
rect 735 -849 773 -840
rect 735 -869 744 -849
rect 764 -869 773 -849
rect 631 -874 667 -873
rect 735 -877 773 -869
rect 839 -845 983 -839
rect 839 -865 847 -845
rect 867 -846 955 -845
rect 867 -865 895 -846
rect 839 -867 895 -865
rect 917 -865 955 -846
rect 975 -865 983 -845
rect 917 -867 983 -865
rect 839 -873 983 -867
rect 839 -874 875 -873
rect 947 -874 983 -873
rect 1049 -840 1086 -839
rect 1049 -841 1087 -840
rect 1049 -849 1113 -841
rect 1049 -869 1058 -849
rect 1078 -863 1113 -849
rect 1133 -863 1136 -843
rect 1078 -868 1136 -863
rect 1078 -869 1113 -868
rect 315 -906 352 -877
rect 135 -952 173 -911
rect 316 -908 352 -906
rect 528 -908 565 -877
rect 316 -930 565 -908
rect 736 -909 773 -877
rect 1049 -881 1113 -869
rect 1153 -907 1180 -729
rect 1012 -909 1180 -907
rect 736 -935 1180 -909
rect 737 -952 761 -935
rect 1012 -936 1180 -935
rect 135 -970 762 -952
rect 1388 -956 1638 -932
rect 135 -976 173 -970
rect 135 -1000 172 -976
rect 135 -1024 170 -1000
rect 133 -1033 170 -1024
rect 133 -1051 143 -1033
rect 161 -1051 170 -1033
rect 133 -1061 170 -1051
rect 1388 -1027 1425 -956
rect 1540 -1017 1571 -1016
rect 1388 -1047 1397 -1027
rect 1417 -1047 1425 -1027
rect 1388 -1057 1425 -1047
rect 1484 -1027 1571 -1017
rect 1484 -1047 1493 -1027
rect 1513 -1047 1571 -1027
rect 1484 -1056 1571 -1047
rect 1484 -1057 1521 -1056
rect 1540 -1109 1571 -1056
rect 1601 -1027 1638 -956
rect 1809 -951 2202 -931
rect 2222 -951 2225 -931
rect 1809 -956 2225 -951
rect 1809 -957 2150 -956
rect 1753 -1017 1784 -1016
rect 1601 -1047 1610 -1027
rect 1630 -1047 1638 -1027
rect 1601 -1057 1638 -1047
rect 1697 -1024 1784 -1017
rect 1697 -1027 1758 -1024
rect 1697 -1047 1706 -1027
rect 1726 -1044 1758 -1027
rect 1779 -1044 1784 -1024
rect 1726 -1047 1784 -1044
rect 1697 -1054 1784 -1047
rect 1809 -1027 1846 -957
rect 2112 -958 2149 -957
rect 1961 -1017 1997 -1016
rect 1809 -1047 1818 -1027
rect 1838 -1047 1846 -1027
rect 1697 -1056 1753 -1054
rect 1697 -1057 1734 -1056
rect 1809 -1057 1846 -1047
rect 1905 -1027 2053 -1017
rect 2153 -1020 2249 -1018
rect 1905 -1047 1914 -1027
rect 1934 -1047 2024 -1027
rect 2044 -1047 2053 -1027
rect 1905 -1056 2053 -1047
rect 2111 -1027 2249 -1020
rect 2111 -1047 2120 -1027
rect 2140 -1047 2249 -1027
rect 2111 -1056 2249 -1047
rect 1905 -1057 1942 -1056
rect 1961 -1108 1997 -1056
rect 2016 -1057 2053 -1056
rect 2112 -1057 2149 -1056
rect 1432 -1110 1473 -1109
rect 1324 -1117 1473 -1110
rect 136 -1125 173 -1123
rect 136 -1126 784 -1125
rect 135 -1132 784 -1126
rect 135 -1150 145 -1132
rect 163 -1146 784 -1132
rect 1324 -1137 1442 -1117
rect 1462 -1137 1473 -1117
rect 1324 -1145 1473 -1137
rect 1540 -1113 1899 -1109
rect 1540 -1118 1862 -1113
rect 1540 -1142 1653 -1118
rect 1677 -1137 1862 -1118
rect 1886 -1137 1899 -1113
rect 1677 -1142 1899 -1137
rect 1540 -1145 1899 -1142
rect 1961 -1145 1996 -1108
rect 2064 -1111 2164 -1108
rect 2064 -1115 2131 -1111
rect 2064 -1141 2076 -1115
rect 2102 -1137 2131 -1115
rect 2157 -1137 2164 -1111
rect 2102 -1141 2164 -1137
rect 2064 -1145 2164 -1141
rect 163 -1150 173 -1146
rect 614 -1147 784 -1146
rect 135 -1160 173 -1150
rect 135 -1238 170 -1160
rect 747 -1170 784 -1147
rect 1540 -1166 1571 -1145
rect 1961 -1166 1997 -1145
rect 1383 -1167 1420 -1166
rect 131 -1247 170 -1238
rect 131 -1265 141 -1247
rect 159 -1265 170 -1247
rect 131 -1271 170 -1265
rect 326 -1195 576 -1171
rect 326 -1266 363 -1195
rect 478 -1256 509 -1255
rect 131 -1275 168 -1271
rect 326 -1286 335 -1266
rect 355 -1286 363 -1266
rect 326 -1296 363 -1286
rect 422 -1266 509 -1256
rect 422 -1286 431 -1266
rect 451 -1286 509 -1266
rect 422 -1295 509 -1286
rect 422 -1296 459 -1295
rect 134 -1346 171 -1337
rect 132 -1364 143 -1346
rect 161 -1364 171 -1346
rect 478 -1348 509 -1295
rect 539 -1266 576 -1195
rect 747 -1190 1140 -1170
rect 1160 -1190 1163 -1170
rect 747 -1195 1163 -1190
rect 1382 -1176 1420 -1167
rect 747 -1196 1088 -1195
rect 1382 -1196 1391 -1176
rect 1411 -1196 1420 -1176
rect 691 -1256 722 -1255
rect 539 -1286 548 -1266
rect 568 -1286 576 -1266
rect 539 -1296 576 -1286
rect 635 -1263 722 -1256
rect 635 -1266 696 -1263
rect 635 -1286 644 -1266
rect 664 -1283 696 -1266
rect 717 -1283 722 -1263
rect 664 -1286 722 -1283
rect 635 -1293 722 -1286
rect 747 -1266 784 -1196
rect 1050 -1197 1087 -1196
rect 1382 -1204 1420 -1196
rect 1486 -1172 1571 -1166
rect 1596 -1167 1633 -1166
rect 1486 -1192 1494 -1172
rect 1514 -1192 1571 -1172
rect 1486 -1200 1571 -1192
rect 1595 -1176 1633 -1167
rect 1595 -1196 1604 -1176
rect 1624 -1196 1633 -1176
rect 1486 -1201 1522 -1200
rect 1595 -1204 1633 -1196
rect 1699 -1172 1784 -1166
rect 1804 -1167 1841 -1166
rect 1699 -1192 1707 -1172
rect 1727 -1173 1784 -1172
rect 1727 -1192 1756 -1173
rect 1699 -1193 1756 -1192
rect 1777 -1193 1784 -1173
rect 1699 -1200 1784 -1193
rect 1803 -1176 1841 -1167
rect 1803 -1196 1812 -1176
rect 1832 -1196 1841 -1176
rect 1699 -1201 1735 -1200
rect 1803 -1204 1841 -1196
rect 1907 -1172 2051 -1166
rect 1907 -1192 1915 -1172
rect 1935 -1174 2023 -1172
rect 1935 -1191 1971 -1174
rect 1995 -1191 2023 -1174
rect 1935 -1192 2023 -1191
rect 2043 -1192 2051 -1172
rect 1907 -1200 2051 -1192
rect 1907 -1201 1943 -1200
rect 2015 -1201 2051 -1200
rect 2117 -1167 2154 -1166
rect 2117 -1168 2155 -1167
rect 2117 -1176 2181 -1168
rect 2117 -1196 2126 -1176
rect 2146 -1190 2181 -1176
rect 2201 -1190 2204 -1170
rect 2146 -1195 2204 -1190
rect 2146 -1196 2181 -1195
rect 1383 -1233 1420 -1204
rect 1384 -1235 1420 -1233
rect 1596 -1235 1633 -1204
rect 899 -1256 935 -1255
rect 747 -1286 756 -1266
rect 776 -1286 784 -1266
rect 635 -1295 691 -1293
rect 635 -1296 672 -1295
rect 747 -1296 784 -1286
rect 843 -1266 991 -1256
rect 1384 -1257 1633 -1235
rect 1804 -1236 1841 -1204
rect 2117 -1208 2181 -1196
rect 2221 -1234 2248 -1056
rect 2080 -1236 2248 -1234
rect 1804 -1247 2248 -1236
rect 1091 -1259 1187 -1257
rect 843 -1286 852 -1266
rect 872 -1286 962 -1266
rect 982 -1286 991 -1266
rect 843 -1295 991 -1286
rect 1049 -1266 1187 -1259
rect 1804 -1262 2250 -1247
rect 2080 -1263 2250 -1262
rect 1049 -1286 1058 -1266
rect 1078 -1286 1187 -1266
rect 1049 -1295 1187 -1286
rect 843 -1296 880 -1295
rect 899 -1347 935 -1295
rect 954 -1296 991 -1295
rect 1050 -1296 1087 -1295
rect 370 -1349 411 -1348
rect 132 -1513 171 -1364
rect 262 -1356 411 -1349
rect 262 -1376 380 -1356
rect 400 -1376 411 -1356
rect 262 -1384 411 -1376
rect 478 -1352 837 -1348
rect 478 -1357 800 -1352
rect 478 -1381 591 -1357
rect 615 -1376 800 -1357
rect 824 -1376 837 -1352
rect 615 -1381 837 -1376
rect 478 -1384 837 -1381
rect 899 -1384 934 -1347
rect 1002 -1350 1102 -1347
rect 1002 -1354 1069 -1350
rect 1002 -1380 1014 -1354
rect 1040 -1376 1069 -1354
rect 1095 -1376 1102 -1350
rect 1040 -1380 1102 -1376
rect 1002 -1384 1102 -1380
rect 478 -1405 509 -1384
rect 899 -1405 935 -1384
rect 321 -1406 358 -1405
rect 320 -1415 358 -1406
rect 320 -1435 329 -1415
rect 349 -1435 358 -1415
rect 320 -1443 358 -1435
rect 424 -1411 509 -1405
rect 534 -1406 571 -1405
rect 424 -1431 432 -1411
rect 452 -1431 509 -1411
rect 424 -1439 509 -1431
rect 533 -1415 571 -1406
rect 533 -1435 542 -1415
rect 562 -1435 571 -1415
rect 424 -1440 460 -1439
rect 533 -1443 571 -1435
rect 637 -1411 722 -1405
rect 742 -1406 779 -1405
rect 637 -1431 645 -1411
rect 665 -1412 722 -1411
rect 665 -1431 694 -1412
rect 637 -1432 694 -1431
rect 715 -1432 722 -1412
rect 637 -1439 722 -1432
rect 741 -1415 779 -1406
rect 741 -1435 750 -1415
rect 770 -1435 779 -1415
rect 637 -1440 673 -1439
rect 741 -1443 779 -1435
rect 845 -1410 989 -1405
rect 845 -1411 910 -1410
rect 845 -1431 853 -1411
rect 873 -1431 910 -1411
rect 932 -1411 989 -1410
rect 932 -1431 961 -1411
rect 981 -1431 989 -1411
rect 845 -1439 989 -1431
rect 845 -1440 881 -1439
rect 953 -1440 989 -1439
rect 1055 -1406 1092 -1405
rect 1055 -1407 1093 -1406
rect 1055 -1415 1119 -1407
rect 1055 -1435 1064 -1415
rect 1084 -1429 1119 -1415
rect 1139 -1429 1142 -1409
rect 1084 -1434 1142 -1429
rect 1084 -1435 1119 -1434
rect 321 -1472 358 -1443
rect 322 -1474 358 -1472
rect 534 -1474 571 -1443
rect 322 -1496 571 -1474
rect 742 -1475 779 -1443
rect 1055 -1447 1119 -1435
rect 1159 -1473 1186 -1295
rect 1018 -1475 1186 -1473
rect 742 -1501 1186 -1475
rect 1338 -1376 1588 -1352
rect 1338 -1447 1375 -1376
rect 1490 -1437 1521 -1436
rect 1338 -1467 1347 -1447
rect 1367 -1467 1375 -1447
rect 1338 -1477 1375 -1467
rect 1434 -1447 1521 -1437
rect 1434 -1467 1443 -1447
rect 1463 -1467 1521 -1447
rect 1434 -1476 1521 -1467
rect 1434 -1477 1471 -1476
rect 742 -1511 764 -1501
rect 1018 -1502 1186 -1501
rect 702 -1513 764 -1511
rect 132 -1520 764 -1513
rect 131 -1529 764 -1520
rect 1490 -1529 1521 -1476
rect 1551 -1447 1588 -1376
rect 1759 -1371 2152 -1351
rect 2172 -1371 2175 -1351
rect 1759 -1376 2175 -1371
rect 1759 -1377 2100 -1376
rect 1703 -1437 1734 -1436
rect 1551 -1467 1560 -1447
rect 1580 -1467 1588 -1447
rect 1551 -1477 1588 -1467
rect 1647 -1444 1734 -1437
rect 1647 -1447 1708 -1444
rect 1647 -1467 1656 -1447
rect 1676 -1464 1708 -1447
rect 1729 -1464 1734 -1444
rect 1676 -1467 1734 -1464
rect 1647 -1474 1734 -1467
rect 1759 -1447 1796 -1377
rect 2062 -1378 2099 -1377
rect 1911 -1437 1947 -1436
rect 1759 -1467 1768 -1447
rect 1788 -1467 1796 -1447
rect 1647 -1476 1703 -1474
rect 1647 -1477 1684 -1476
rect 1759 -1477 1796 -1467
rect 1855 -1447 2003 -1437
rect 2103 -1440 2199 -1438
rect 1855 -1467 1864 -1447
rect 1884 -1467 1974 -1447
rect 1994 -1467 2003 -1447
rect 1855 -1476 2003 -1467
rect 2061 -1447 2199 -1440
rect 2061 -1467 2070 -1447
rect 2090 -1467 2199 -1447
rect 2061 -1476 2199 -1467
rect 1855 -1477 1892 -1476
rect 1911 -1528 1947 -1476
rect 1966 -1477 2003 -1476
rect 2062 -1477 2099 -1476
rect 131 -1547 141 -1529
rect 159 -1530 764 -1529
rect 1382 -1530 1423 -1529
rect 159 -1535 180 -1530
rect 159 -1547 171 -1535
rect 1274 -1537 1423 -1530
rect 131 -1555 171 -1547
rect 214 -1548 240 -1547
rect 131 -1557 168 -1555
rect 214 -1566 768 -1548
rect 1274 -1557 1392 -1537
rect 1412 -1557 1423 -1537
rect 1274 -1565 1423 -1557
rect 1490 -1533 1849 -1529
rect 1490 -1538 1812 -1533
rect 1490 -1562 1603 -1538
rect 1627 -1557 1812 -1538
rect 1836 -1557 1849 -1533
rect 1627 -1562 1849 -1557
rect 1490 -1565 1849 -1562
rect 1911 -1565 1946 -1528
rect 2014 -1531 2114 -1528
rect 2014 -1535 2081 -1531
rect 2014 -1561 2026 -1535
rect 2052 -1557 2081 -1535
rect 2107 -1557 2114 -1531
rect 2052 -1561 2114 -1557
rect 2014 -1565 2114 -1561
rect 134 -1625 171 -1619
rect 214 -1625 240 -1566
rect 747 -1585 768 -1566
rect 134 -1628 240 -1625
rect 134 -1646 143 -1628
rect 161 -1642 240 -1628
rect 325 -1610 575 -1586
rect 161 -1644 237 -1642
rect 161 -1646 171 -1644
rect 134 -1656 171 -1646
rect 139 -1721 170 -1656
rect 325 -1681 362 -1610
rect 477 -1671 508 -1670
rect 325 -1701 334 -1681
rect 354 -1701 362 -1681
rect 325 -1711 362 -1701
rect 421 -1681 508 -1671
rect 421 -1701 430 -1681
rect 450 -1701 508 -1681
rect 421 -1710 508 -1701
rect 421 -1711 458 -1710
rect 138 -1730 175 -1721
rect 138 -1748 148 -1730
rect 166 -1748 175 -1730
rect 138 -1758 175 -1748
rect 477 -1763 508 -1710
rect 538 -1681 575 -1610
rect 746 -1605 1139 -1585
rect 1159 -1605 1162 -1585
rect 1490 -1586 1521 -1565
rect 1911 -1586 1947 -1565
rect 1333 -1587 1370 -1586
rect 746 -1610 1162 -1605
rect 1332 -1596 1370 -1587
rect 746 -1611 1087 -1610
rect 690 -1671 721 -1670
rect 538 -1701 547 -1681
rect 567 -1701 575 -1681
rect 538 -1711 575 -1701
rect 634 -1678 721 -1671
rect 634 -1681 695 -1678
rect 634 -1701 643 -1681
rect 663 -1698 695 -1681
rect 716 -1698 721 -1678
rect 663 -1701 721 -1698
rect 634 -1708 721 -1701
rect 746 -1681 783 -1611
rect 1049 -1612 1086 -1611
rect 1332 -1616 1341 -1596
rect 1361 -1616 1370 -1596
rect 1332 -1624 1370 -1616
rect 1436 -1592 1521 -1586
rect 1546 -1587 1583 -1586
rect 1436 -1612 1444 -1592
rect 1464 -1612 1521 -1592
rect 1436 -1620 1521 -1612
rect 1545 -1596 1583 -1587
rect 1545 -1616 1554 -1596
rect 1574 -1616 1583 -1596
rect 1436 -1621 1472 -1620
rect 1545 -1624 1583 -1616
rect 1649 -1592 1734 -1586
rect 1754 -1587 1791 -1586
rect 1649 -1612 1657 -1592
rect 1677 -1593 1734 -1592
rect 1677 -1612 1706 -1593
rect 1649 -1613 1706 -1612
rect 1727 -1613 1734 -1593
rect 1649 -1620 1734 -1613
rect 1753 -1596 1791 -1587
rect 1753 -1616 1762 -1596
rect 1782 -1616 1791 -1596
rect 1649 -1621 1685 -1620
rect 1753 -1624 1791 -1616
rect 1857 -1591 2001 -1586
rect 1857 -1592 1916 -1591
rect 1857 -1612 1865 -1592
rect 1885 -1611 1916 -1592
rect 1940 -1592 2001 -1591
rect 1940 -1611 1973 -1592
rect 1885 -1612 1973 -1611
rect 1993 -1612 2001 -1592
rect 1857 -1620 2001 -1612
rect 1857 -1621 1893 -1620
rect 1965 -1621 2001 -1620
rect 2067 -1587 2104 -1586
rect 2067 -1588 2105 -1587
rect 2067 -1596 2131 -1588
rect 2067 -1616 2076 -1596
rect 2096 -1610 2131 -1596
rect 2151 -1610 2154 -1590
rect 2096 -1615 2154 -1610
rect 2096 -1616 2131 -1615
rect 1333 -1653 1370 -1624
rect 1334 -1655 1370 -1653
rect 1546 -1655 1583 -1624
rect 898 -1671 934 -1670
rect 746 -1701 755 -1681
rect 775 -1701 783 -1681
rect 634 -1710 690 -1708
rect 634 -1711 671 -1710
rect 746 -1711 783 -1701
rect 842 -1681 990 -1671
rect 1090 -1674 1186 -1672
rect 842 -1701 851 -1681
rect 871 -1701 961 -1681
rect 981 -1701 990 -1681
rect 842 -1710 990 -1701
rect 1048 -1681 1186 -1674
rect 1334 -1677 1583 -1655
rect 1754 -1656 1791 -1624
rect 2067 -1628 2131 -1616
rect 2171 -1654 2198 -1476
rect 2030 -1656 2198 -1654
rect 1754 -1660 2198 -1656
rect 1048 -1701 1057 -1681
rect 1077 -1701 1186 -1681
rect 1754 -1679 1803 -1660
rect 1823 -1679 2198 -1660
rect 1754 -1682 2198 -1679
rect 2030 -1683 2198 -1682
rect 2219 -1657 2250 -1263
rect 2219 -1683 2224 -1657
rect 2243 -1683 2250 -1657
rect 2219 -1686 2250 -1683
rect 1048 -1710 1186 -1701
rect 842 -1711 879 -1710
rect 898 -1762 934 -1710
rect 953 -1711 990 -1710
rect 1049 -1711 1086 -1710
rect 369 -1764 410 -1763
rect 261 -1771 410 -1764
rect 261 -1791 379 -1771
rect 399 -1791 410 -1771
rect 261 -1799 410 -1791
rect 477 -1767 836 -1763
rect 477 -1772 799 -1767
rect 477 -1796 590 -1772
rect 614 -1791 799 -1772
rect 823 -1791 836 -1767
rect 614 -1796 836 -1791
rect 477 -1799 836 -1796
rect 898 -1799 933 -1762
rect 1001 -1765 1101 -1762
rect 1001 -1769 1068 -1765
rect 1001 -1795 1013 -1769
rect 1039 -1791 1068 -1769
rect 1094 -1791 1101 -1765
rect 1039 -1795 1101 -1791
rect 1001 -1799 1101 -1795
rect 477 -1820 508 -1799
rect 898 -1820 934 -1799
rect 141 -1829 178 -1820
rect 320 -1821 357 -1820
rect 141 -1847 150 -1829
rect 168 -1847 178 -1829
rect 141 -1857 178 -1847
rect 142 -1892 178 -1857
rect 319 -1830 357 -1821
rect 319 -1850 328 -1830
rect 348 -1850 357 -1830
rect 319 -1858 357 -1850
rect 423 -1826 508 -1820
rect 533 -1821 570 -1820
rect 423 -1846 431 -1826
rect 451 -1846 508 -1826
rect 423 -1854 508 -1846
rect 532 -1830 570 -1821
rect 532 -1850 541 -1830
rect 561 -1850 570 -1830
rect 423 -1855 459 -1854
rect 532 -1858 570 -1850
rect 636 -1826 721 -1820
rect 741 -1821 778 -1820
rect 636 -1846 644 -1826
rect 664 -1827 721 -1826
rect 664 -1846 693 -1827
rect 636 -1847 693 -1846
rect 714 -1847 721 -1827
rect 636 -1854 721 -1847
rect 740 -1830 778 -1821
rect 740 -1850 749 -1830
rect 769 -1850 778 -1830
rect 636 -1855 672 -1854
rect 740 -1858 778 -1850
rect 844 -1826 988 -1820
rect 844 -1846 852 -1826
rect 872 -1827 960 -1826
rect 872 -1846 900 -1827
rect 844 -1848 900 -1846
rect 922 -1846 960 -1827
rect 980 -1846 988 -1826
rect 922 -1848 988 -1846
rect 844 -1854 988 -1848
rect 844 -1855 880 -1854
rect 952 -1855 988 -1854
rect 1054 -1821 1091 -1820
rect 1054 -1822 1092 -1821
rect 1054 -1830 1118 -1822
rect 1054 -1850 1063 -1830
rect 1083 -1844 1118 -1830
rect 1138 -1844 1141 -1824
rect 1083 -1849 1141 -1844
rect 1083 -1850 1118 -1849
rect 320 -1887 357 -1858
rect 140 -1933 178 -1892
rect 321 -1889 357 -1887
rect 533 -1889 570 -1858
rect 321 -1911 570 -1889
rect 741 -1890 778 -1858
rect 1054 -1862 1118 -1850
rect 1158 -1888 1185 -1710
rect 1017 -1890 1185 -1888
rect 741 -1916 1185 -1890
rect 742 -1933 766 -1916
rect 1017 -1917 1185 -1916
rect 1553 -1888 1803 -1864
rect 140 -1951 767 -1933
rect 140 -1957 178 -1951
rect 142 -2003 177 -1957
rect 1553 -1959 1590 -1888
rect 1705 -1949 1736 -1948
rect 1553 -1979 1562 -1959
rect 1582 -1979 1590 -1959
rect 1553 -1989 1590 -1979
rect 1649 -1959 1736 -1949
rect 1649 -1979 1658 -1959
rect 1678 -1979 1736 -1959
rect 1649 -1988 1736 -1979
rect 1649 -1989 1686 -1988
rect 140 -2012 177 -2003
rect 140 -2030 150 -2012
rect 168 -2030 177 -2012
rect 140 -2040 177 -2030
rect 1705 -2041 1736 -1988
rect 1766 -1959 1803 -1888
rect 1974 -1883 2367 -1863
rect 2387 -1883 2390 -1863
rect 1974 -1888 2390 -1883
rect 1974 -1889 2315 -1888
rect 1918 -1949 1949 -1948
rect 1766 -1979 1775 -1959
rect 1795 -1979 1803 -1959
rect 1766 -1989 1803 -1979
rect 1862 -1956 1949 -1949
rect 1862 -1959 1923 -1956
rect 1862 -1979 1871 -1959
rect 1891 -1976 1923 -1959
rect 1944 -1976 1949 -1956
rect 1891 -1979 1949 -1976
rect 1862 -1986 1949 -1979
rect 1974 -1959 2011 -1889
rect 2277 -1890 2314 -1889
rect 2126 -1949 2162 -1948
rect 1974 -1979 1983 -1959
rect 2003 -1979 2011 -1959
rect 1862 -1988 1918 -1986
rect 1862 -1989 1899 -1988
rect 1974 -1989 2011 -1979
rect 2070 -1959 2218 -1949
rect 2318 -1952 2414 -1950
rect 2070 -1979 2079 -1959
rect 2099 -1979 2189 -1959
rect 2209 -1979 2218 -1959
rect 2070 -1988 2218 -1979
rect 2276 -1959 2414 -1952
rect 2276 -1979 2285 -1959
rect 2305 -1979 2414 -1959
rect 2276 -1988 2414 -1979
rect 2070 -1989 2107 -1988
rect 2126 -2040 2162 -1988
rect 2181 -1989 2218 -1988
rect 2277 -1989 2314 -1988
rect 1597 -2042 1638 -2041
rect 1489 -2049 1638 -2042
rect 1489 -2069 1607 -2049
rect 1627 -2069 1638 -2049
rect 1489 -2077 1638 -2069
rect 1705 -2045 2064 -2041
rect 1705 -2050 2027 -2045
rect 1705 -2074 1818 -2050
rect 1842 -2069 2027 -2050
rect 2051 -2069 2064 -2045
rect 1842 -2074 2064 -2069
rect 1705 -2077 2064 -2074
rect 2126 -2077 2161 -2040
rect 2229 -2043 2329 -2040
rect 2229 -2047 2296 -2043
rect 2229 -2073 2241 -2047
rect 2267 -2069 2296 -2047
rect 2322 -2069 2329 -2043
rect 2267 -2073 2329 -2069
rect 2229 -2077 2329 -2073
rect 1705 -2098 1736 -2077
rect 2126 -2098 2162 -2077
rect 1548 -2099 1585 -2098
rect 143 -2104 180 -2102
rect 143 -2105 791 -2104
rect 142 -2111 791 -2105
rect 142 -2129 152 -2111
rect 170 -2125 791 -2111
rect 170 -2129 180 -2125
rect 621 -2126 791 -2125
rect 142 -2139 180 -2129
rect 142 -2217 177 -2139
rect 754 -2149 791 -2126
rect 1547 -2108 1585 -2099
rect 1547 -2128 1556 -2108
rect 1576 -2128 1585 -2108
rect 1547 -2136 1585 -2128
rect 1651 -2104 1736 -2098
rect 1761 -2099 1798 -2098
rect 1651 -2124 1659 -2104
rect 1679 -2124 1736 -2104
rect 1651 -2132 1736 -2124
rect 1760 -2108 1798 -2099
rect 1760 -2128 1769 -2108
rect 1789 -2128 1798 -2108
rect 1651 -2133 1687 -2132
rect 1760 -2136 1798 -2128
rect 1864 -2104 1949 -2098
rect 1969 -2099 2006 -2098
rect 1864 -2124 1872 -2104
rect 1892 -2105 1949 -2104
rect 1892 -2124 1921 -2105
rect 1864 -2125 1921 -2124
rect 1942 -2125 1949 -2105
rect 1864 -2132 1949 -2125
rect 1968 -2108 2006 -2099
rect 1968 -2128 1977 -2108
rect 1997 -2128 2006 -2108
rect 1864 -2133 1900 -2132
rect 1968 -2136 2006 -2128
rect 2072 -2104 2216 -2098
rect 2072 -2124 2080 -2104
rect 2100 -2123 2136 -2104
rect 2159 -2123 2188 -2104
rect 2100 -2124 2188 -2123
rect 2208 -2124 2216 -2104
rect 2072 -2132 2216 -2124
rect 2072 -2133 2108 -2132
rect 2180 -2133 2216 -2132
rect 2282 -2099 2319 -2098
rect 2282 -2100 2320 -2099
rect 2282 -2108 2346 -2100
rect 2282 -2128 2291 -2108
rect 2311 -2122 2346 -2108
rect 2366 -2122 2369 -2102
rect 2311 -2127 2369 -2122
rect 2311 -2128 2346 -2127
rect 138 -2226 177 -2217
rect 138 -2244 148 -2226
rect 166 -2244 177 -2226
rect 138 -2250 177 -2244
rect 333 -2174 583 -2150
rect 333 -2245 370 -2174
rect 485 -2235 516 -2234
rect 138 -2254 175 -2250
rect 333 -2265 342 -2245
rect 362 -2265 370 -2245
rect 333 -2275 370 -2265
rect 429 -2245 516 -2235
rect 429 -2265 438 -2245
rect 458 -2265 516 -2245
rect 429 -2274 516 -2265
rect 429 -2275 466 -2274
rect 141 -2325 178 -2316
rect 139 -2343 150 -2325
rect 168 -2343 178 -2325
rect 485 -2327 516 -2274
rect 546 -2245 583 -2174
rect 754 -2169 1147 -2149
rect 1167 -2169 1170 -2149
rect 1548 -2165 1585 -2136
rect 754 -2174 1170 -2169
rect 1549 -2167 1585 -2165
rect 1761 -2167 1798 -2136
rect 754 -2175 1095 -2174
rect 698 -2235 729 -2234
rect 546 -2265 555 -2245
rect 575 -2265 583 -2245
rect 546 -2275 583 -2265
rect 642 -2242 729 -2235
rect 642 -2245 703 -2242
rect 642 -2265 651 -2245
rect 671 -2262 703 -2245
rect 724 -2262 729 -2242
rect 671 -2265 729 -2262
rect 642 -2272 729 -2265
rect 754 -2245 791 -2175
rect 1057 -2176 1094 -2175
rect 1549 -2189 1798 -2167
rect 1969 -2168 2006 -2136
rect 2282 -2140 2346 -2128
rect 2386 -2166 2413 -1988
rect 2441 -2101 2479 -270
rect 2443 -2161 2476 -2101
rect 2245 -2168 2413 -2166
rect 1969 -2194 2413 -2168
rect 2245 -2195 2413 -2194
rect 2442 -2172 2479 -2161
rect 2442 -2191 2448 -2172
rect 2471 -2191 2479 -2172
rect 906 -2235 942 -2234
rect 754 -2265 763 -2245
rect 783 -2265 791 -2245
rect 642 -2274 698 -2272
rect 642 -2275 679 -2274
rect 754 -2275 791 -2265
rect 850 -2245 998 -2235
rect 1098 -2238 1194 -2236
rect 850 -2265 859 -2245
rect 879 -2265 969 -2245
rect 989 -2265 998 -2245
rect 850 -2274 998 -2265
rect 1056 -2245 1194 -2238
rect 1056 -2265 1065 -2245
rect 1085 -2265 1194 -2245
rect 1056 -2274 1194 -2265
rect 850 -2275 887 -2274
rect 906 -2326 942 -2274
rect 961 -2275 998 -2274
rect 1057 -2275 1094 -2274
rect 377 -2328 418 -2327
rect 139 -2492 178 -2343
rect 269 -2335 418 -2328
rect 269 -2355 387 -2335
rect 407 -2355 418 -2335
rect 269 -2363 418 -2355
rect 485 -2331 844 -2327
rect 485 -2336 807 -2331
rect 485 -2360 598 -2336
rect 622 -2355 807 -2336
rect 831 -2355 844 -2331
rect 622 -2360 844 -2355
rect 485 -2363 844 -2360
rect 906 -2363 941 -2326
rect 1009 -2329 1109 -2326
rect 1009 -2333 1076 -2329
rect 1009 -2359 1021 -2333
rect 1047 -2355 1076 -2333
rect 1102 -2355 1109 -2329
rect 1047 -2359 1109 -2355
rect 1009 -2363 1109 -2359
rect 485 -2384 516 -2363
rect 906 -2384 942 -2363
rect 328 -2385 365 -2384
rect 327 -2394 365 -2385
rect 327 -2414 336 -2394
rect 356 -2414 365 -2394
rect 327 -2422 365 -2414
rect 431 -2390 516 -2384
rect 541 -2385 578 -2384
rect 431 -2410 439 -2390
rect 459 -2410 516 -2390
rect 431 -2418 516 -2410
rect 540 -2394 578 -2385
rect 540 -2414 549 -2394
rect 569 -2414 578 -2394
rect 431 -2419 467 -2418
rect 540 -2422 578 -2414
rect 644 -2390 729 -2384
rect 749 -2385 786 -2384
rect 644 -2410 652 -2390
rect 672 -2391 729 -2390
rect 672 -2410 701 -2391
rect 644 -2411 701 -2410
rect 722 -2411 729 -2391
rect 644 -2418 729 -2411
rect 748 -2394 786 -2385
rect 748 -2414 757 -2394
rect 777 -2414 786 -2394
rect 644 -2419 680 -2418
rect 748 -2422 786 -2414
rect 852 -2389 996 -2384
rect 852 -2390 917 -2389
rect 852 -2410 860 -2390
rect 880 -2410 917 -2390
rect 939 -2390 996 -2389
rect 939 -2410 968 -2390
rect 988 -2410 996 -2390
rect 852 -2418 996 -2410
rect 852 -2419 888 -2418
rect 960 -2419 996 -2418
rect 1062 -2385 1099 -2384
rect 1062 -2386 1100 -2385
rect 1062 -2394 1126 -2386
rect 1062 -2414 1071 -2394
rect 1091 -2408 1126 -2394
rect 1146 -2408 1149 -2388
rect 1091 -2413 1149 -2408
rect 1091 -2414 1126 -2413
rect 328 -2451 365 -2422
rect 329 -2453 365 -2451
rect 541 -2453 578 -2422
rect 329 -2475 578 -2453
rect 749 -2454 786 -2422
rect 1062 -2426 1126 -2414
rect 1166 -2452 1193 -2274
rect 1025 -2454 1193 -2452
rect 749 -2480 1193 -2454
rect 1345 -2355 1595 -2331
rect 1345 -2426 1382 -2355
rect 1497 -2416 1528 -2415
rect 1345 -2446 1354 -2426
rect 1374 -2446 1382 -2426
rect 1345 -2456 1382 -2446
rect 1441 -2426 1528 -2416
rect 1441 -2446 1450 -2426
rect 1470 -2446 1528 -2426
rect 1441 -2455 1528 -2446
rect 1441 -2456 1478 -2455
rect 749 -2490 771 -2480
rect 1025 -2481 1193 -2480
rect 709 -2492 771 -2490
rect 139 -2499 771 -2492
rect 138 -2508 771 -2499
rect 1497 -2508 1528 -2455
rect 1558 -2426 1595 -2355
rect 1766 -2350 2159 -2330
rect 2179 -2350 2182 -2330
rect 1766 -2355 2182 -2350
rect 1766 -2356 2107 -2355
rect 1710 -2416 1741 -2415
rect 1558 -2446 1567 -2426
rect 1587 -2446 1595 -2426
rect 1558 -2456 1595 -2446
rect 1654 -2423 1741 -2416
rect 1654 -2426 1715 -2423
rect 1654 -2446 1663 -2426
rect 1683 -2443 1715 -2426
rect 1736 -2443 1741 -2423
rect 1683 -2446 1741 -2443
rect 1654 -2453 1741 -2446
rect 1766 -2426 1803 -2356
rect 2069 -2357 2106 -2356
rect 1918 -2416 1954 -2415
rect 1766 -2446 1775 -2426
rect 1795 -2446 1803 -2426
rect 1654 -2455 1710 -2453
rect 1654 -2456 1691 -2455
rect 1766 -2456 1803 -2446
rect 1862 -2426 2010 -2416
rect 2110 -2419 2206 -2417
rect 1862 -2446 1871 -2426
rect 1891 -2446 1981 -2426
rect 2001 -2446 2010 -2426
rect 1862 -2455 2010 -2446
rect 2068 -2426 2206 -2419
rect 2068 -2446 2077 -2426
rect 2097 -2446 2206 -2426
rect 2068 -2455 2206 -2446
rect 1862 -2456 1899 -2455
rect 1918 -2507 1954 -2455
rect 1973 -2456 2010 -2455
rect 2069 -2456 2106 -2455
rect 138 -2526 148 -2508
rect 166 -2509 771 -2508
rect 1389 -2509 1430 -2508
rect 166 -2514 187 -2509
rect 166 -2526 178 -2514
rect 1281 -2516 1430 -2509
rect 138 -2534 178 -2526
rect 221 -2527 247 -2526
rect 138 -2536 175 -2534
rect 221 -2545 775 -2527
rect 1281 -2536 1399 -2516
rect 1419 -2536 1430 -2516
rect 1281 -2544 1430 -2536
rect 1497 -2512 1856 -2508
rect 1497 -2517 1819 -2512
rect 1497 -2541 1610 -2517
rect 1634 -2536 1819 -2517
rect 1843 -2536 1856 -2512
rect 1634 -2541 1856 -2536
rect 1497 -2544 1856 -2541
rect 1918 -2544 1953 -2507
rect 2021 -2510 2121 -2507
rect 2021 -2514 2088 -2510
rect 2021 -2540 2033 -2514
rect 2059 -2536 2088 -2514
rect 2114 -2536 2121 -2510
rect 2059 -2540 2121 -2536
rect 2021 -2544 2121 -2540
rect 141 -2604 178 -2598
rect 221 -2604 247 -2545
rect 754 -2564 775 -2545
rect 141 -2607 247 -2604
rect 141 -2625 150 -2607
rect 168 -2621 247 -2607
rect 332 -2589 582 -2565
rect 168 -2623 244 -2621
rect 168 -2625 178 -2623
rect 141 -2635 178 -2625
rect 146 -2700 177 -2635
rect 332 -2660 369 -2589
rect 484 -2650 515 -2649
rect 332 -2680 341 -2660
rect 361 -2680 369 -2660
rect 332 -2690 369 -2680
rect 428 -2660 515 -2650
rect 428 -2680 437 -2660
rect 457 -2680 515 -2660
rect 428 -2689 515 -2680
rect 428 -2690 465 -2689
rect 145 -2709 182 -2700
rect 145 -2727 155 -2709
rect 173 -2727 182 -2709
rect 145 -2737 182 -2727
rect 484 -2742 515 -2689
rect 545 -2660 582 -2589
rect 753 -2584 1146 -2564
rect 1166 -2584 1169 -2564
rect 1497 -2565 1528 -2544
rect 1918 -2565 1954 -2544
rect 1340 -2566 1377 -2565
rect 753 -2589 1169 -2584
rect 1339 -2575 1377 -2566
rect 753 -2590 1094 -2589
rect 697 -2650 728 -2649
rect 545 -2680 554 -2660
rect 574 -2680 582 -2660
rect 545 -2690 582 -2680
rect 641 -2657 728 -2650
rect 641 -2660 702 -2657
rect 641 -2680 650 -2660
rect 670 -2677 702 -2660
rect 723 -2677 728 -2657
rect 670 -2680 728 -2677
rect 641 -2687 728 -2680
rect 753 -2660 790 -2590
rect 1056 -2591 1093 -2590
rect 1339 -2595 1348 -2575
rect 1368 -2595 1377 -2575
rect 1339 -2603 1377 -2595
rect 1443 -2571 1528 -2565
rect 1553 -2566 1590 -2565
rect 1443 -2591 1451 -2571
rect 1471 -2591 1528 -2571
rect 1443 -2599 1528 -2591
rect 1552 -2575 1590 -2566
rect 1552 -2595 1561 -2575
rect 1581 -2595 1590 -2575
rect 1443 -2600 1479 -2599
rect 1552 -2603 1590 -2595
rect 1656 -2571 1741 -2565
rect 1761 -2566 1798 -2565
rect 1656 -2591 1664 -2571
rect 1684 -2572 1741 -2571
rect 1684 -2591 1713 -2572
rect 1656 -2592 1713 -2591
rect 1734 -2592 1741 -2572
rect 1656 -2599 1741 -2592
rect 1760 -2575 1798 -2566
rect 1760 -2595 1769 -2575
rect 1789 -2595 1798 -2575
rect 1656 -2600 1692 -2599
rect 1760 -2603 1798 -2595
rect 1864 -2571 2008 -2565
rect 1864 -2591 1872 -2571
rect 1892 -2591 1924 -2571
rect 1948 -2591 1980 -2571
rect 2000 -2591 2008 -2571
rect 1864 -2599 2008 -2591
rect 1864 -2600 1900 -2599
rect 1972 -2600 2008 -2599
rect 2074 -2566 2111 -2565
rect 2074 -2567 2112 -2566
rect 2074 -2575 2138 -2567
rect 2074 -2595 2083 -2575
rect 2103 -2589 2138 -2575
rect 2158 -2589 2161 -2569
rect 2103 -2594 2161 -2589
rect 2103 -2595 2138 -2594
rect 1340 -2632 1377 -2603
rect 1341 -2634 1377 -2632
rect 1553 -2634 1590 -2603
rect 905 -2650 941 -2649
rect 753 -2680 762 -2660
rect 782 -2680 790 -2660
rect 641 -2689 697 -2687
rect 641 -2690 678 -2689
rect 753 -2690 790 -2680
rect 849 -2660 997 -2650
rect 1097 -2653 1193 -2651
rect 849 -2680 858 -2660
rect 878 -2680 968 -2660
rect 988 -2680 997 -2660
rect 849 -2689 997 -2680
rect 1055 -2660 1193 -2653
rect 1341 -2656 1590 -2634
rect 1761 -2635 1798 -2603
rect 2074 -2607 2138 -2595
rect 2178 -2633 2205 -2455
rect 2037 -2635 2205 -2633
rect 1761 -2639 2205 -2635
rect 1055 -2680 1064 -2660
rect 1084 -2680 1193 -2660
rect 1761 -2658 1810 -2639
rect 1830 -2658 2205 -2639
rect 1761 -2661 2205 -2658
rect 2037 -2662 2205 -2661
rect 1055 -2689 1193 -2680
rect 849 -2690 886 -2689
rect 905 -2741 941 -2689
rect 960 -2690 997 -2689
rect 1056 -2690 1093 -2689
rect 376 -2743 417 -2742
rect 268 -2750 417 -2743
rect 268 -2770 386 -2750
rect 406 -2770 417 -2750
rect 268 -2778 417 -2770
rect 484 -2746 843 -2742
rect 484 -2751 806 -2746
rect 484 -2775 597 -2751
rect 621 -2770 806 -2751
rect 830 -2770 843 -2746
rect 621 -2775 843 -2770
rect 484 -2778 843 -2775
rect 905 -2778 940 -2741
rect 1008 -2744 1108 -2741
rect 1008 -2748 1075 -2744
rect 1008 -2774 1020 -2748
rect 1046 -2770 1075 -2748
rect 1101 -2770 1108 -2744
rect 1046 -2774 1108 -2770
rect 1008 -2778 1108 -2774
rect 484 -2799 515 -2778
rect 905 -2799 941 -2778
rect 148 -2808 185 -2799
rect 327 -2800 364 -2799
rect 148 -2826 157 -2808
rect 175 -2826 185 -2808
rect 148 -2836 185 -2826
rect 149 -2871 185 -2836
rect 326 -2809 364 -2800
rect 326 -2829 335 -2809
rect 355 -2829 364 -2809
rect 326 -2837 364 -2829
rect 430 -2805 515 -2799
rect 540 -2800 577 -2799
rect 430 -2825 438 -2805
rect 458 -2825 515 -2805
rect 430 -2833 515 -2825
rect 539 -2809 577 -2800
rect 539 -2829 548 -2809
rect 568 -2829 577 -2809
rect 430 -2834 466 -2833
rect 539 -2837 577 -2829
rect 643 -2805 728 -2799
rect 748 -2800 785 -2799
rect 643 -2825 651 -2805
rect 671 -2806 728 -2805
rect 671 -2825 700 -2806
rect 643 -2826 700 -2825
rect 721 -2826 728 -2806
rect 643 -2833 728 -2826
rect 747 -2809 785 -2800
rect 747 -2829 756 -2809
rect 776 -2829 785 -2809
rect 643 -2834 679 -2833
rect 747 -2837 785 -2829
rect 851 -2805 995 -2799
rect 851 -2825 859 -2805
rect 879 -2806 967 -2805
rect 879 -2825 907 -2806
rect 851 -2827 907 -2825
rect 929 -2825 967 -2806
rect 987 -2825 995 -2805
rect 929 -2827 995 -2825
rect 851 -2833 995 -2827
rect 851 -2834 887 -2833
rect 959 -2834 995 -2833
rect 1061 -2800 1098 -2799
rect 1061 -2801 1099 -2800
rect 1061 -2809 1125 -2801
rect 1061 -2829 1070 -2809
rect 1090 -2823 1125 -2809
rect 1145 -2823 1148 -2803
rect 1090 -2828 1148 -2823
rect 1090 -2829 1125 -2828
rect 327 -2866 364 -2837
rect 147 -2912 185 -2871
rect 328 -2868 364 -2866
rect 540 -2868 577 -2837
rect 328 -2890 577 -2868
rect 748 -2869 785 -2837
rect 1061 -2841 1125 -2829
rect 1165 -2867 1192 -2689
rect 1024 -2869 1192 -2867
rect 748 -2895 1192 -2869
rect 749 -2912 773 -2895
rect 1024 -2896 1192 -2895
rect 147 -2930 774 -2912
rect 1400 -2916 1650 -2892
rect 147 -2936 185 -2930
rect 147 -2960 184 -2936
rect 147 -2984 182 -2960
rect 145 -2993 182 -2984
rect 145 -3011 155 -2993
rect 173 -3011 182 -2993
rect 145 -3021 182 -3011
rect 1400 -2987 1437 -2916
rect 1552 -2977 1583 -2976
rect 1400 -3007 1409 -2987
rect 1429 -3007 1437 -2987
rect 1400 -3017 1437 -3007
rect 1496 -2987 1583 -2977
rect 1496 -3007 1505 -2987
rect 1525 -3007 1583 -2987
rect 1496 -3016 1583 -3007
rect 1496 -3017 1533 -3016
rect 1552 -3069 1583 -3016
rect 1613 -2987 1650 -2916
rect 1821 -2911 2214 -2891
rect 2234 -2911 2237 -2891
rect 1821 -2916 2237 -2911
rect 1821 -2917 2162 -2916
rect 1765 -2977 1796 -2976
rect 1613 -3007 1622 -2987
rect 1642 -3007 1650 -2987
rect 1613 -3017 1650 -3007
rect 1709 -2984 1796 -2977
rect 1709 -2987 1770 -2984
rect 1709 -3007 1718 -2987
rect 1738 -3004 1770 -2987
rect 1791 -3004 1796 -2984
rect 1738 -3007 1796 -3004
rect 1709 -3014 1796 -3007
rect 1821 -2987 1858 -2917
rect 2124 -2918 2161 -2917
rect 1973 -2977 2009 -2976
rect 1821 -3007 1830 -2987
rect 1850 -3007 1858 -2987
rect 1709 -3016 1765 -3014
rect 1709 -3017 1746 -3016
rect 1821 -3017 1858 -3007
rect 1917 -2987 2065 -2977
rect 2165 -2980 2261 -2978
rect 1917 -3007 1926 -2987
rect 1946 -3007 2036 -2987
rect 2056 -3007 2065 -2987
rect 1917 -3016 2065 -3007
rect 2123 -2987 2261 -2980
rect 2123 -3007 2132 -2987
rect 2152 -3007 2261 -2987
rect 2123 -3016 2261 -3007
rect 1917 -3017 1954 -3016
rect 1973 -3068 2009 -3016
rect 2028 -3017 2065 -3016
rect 2124 -3017 2161 -3016
rect 1444 -3070 1485 -3069
rect 1336 -3077 1485 -3070
rect 148 -3085 185 -3083
rect 148 -3086 796 -3085
rect 147 -3092 796 -3086
rect 147 -3110 157 -3092
rect 175 -3106 796 -3092
rect 1336 -3097 1454 -3077
rect 1474 -3097 1485 -3077
rect 1336 -3105 1485 -3097
rect 1552 -3073 1911 -3069
rect 1552 -3078 1874 -3073
rect 1552 -3102 1665 -3078
rect 1689 -3097 1874 -3078
rect 1898 -3097 1911 -3073
rect 1689 -3102 1911 -3097
rect 1552 -3105 1911 -3102
rect 1973 -3105 2008 -3068
rect 2076 -3071 2176 -3068
rect 2076 -3075 2143 -3071
rect 2076 -3101 2088 -3075
rect 2114 -3097 2143 -3075
rect 2169 -3097 2176 -3071
rect 2114 -3101 2176 -3097
rect 2076 -3105 2176 -3101
rect 175 -3110 185 -3106
rect 626 -3107 796 -3106
rect 147 -3120 185 -3110
rect 147 -3198 182 -3120
rect 759 -3130 796 -3107
rect 1552 -3126 1583 -3105
rect 1973 -3126 2009 -3105
rect 1395 -3127 1432 -3126
rect 143 -3207 182 -3198
rect 143 -3225 153 -3207
rect 171 -3225 182 -3207
rect 143 -3231 182 -3225
rect 338 -3155 588 -3131
rect 338 -3226 375 -3155
rect 490 -3216 521 -3215
rect 143 -3235 180 -3231
rect 338 -3246 347 -3226
rect 367 -3246 375 -3226
rect 338 -3256 375 -3246
rect 434 -3226 521 -3216
rect 434 -3246 443 -3226
rect 463 -3246 521 -3226
rect 434 -3255 521 -3246
rect 434 -3256 471 -3255
rect 146 -3306 183 -3297
rect 144 -3324 155 -3306
rect 173 -3324 183 -3306
rect 490 -3308 521 -3255
rect 551 -3226 588 -3155
rect 759 -3150 1152 -3130
rect 1172 -3150 1175 -3130
rect 759 -3155 1175 -3150
rect 1394 -3136 1432 -3127
rect 759 -3156 1100 -3155
rect 1394 -3156 1403 -3136
rect 1423 -3156 1432 -3136
rect 703 -3216 734 -3215
rect 551 -3246 560 -3226
rect 580 -3246 588 -3226
rect 551 -3256 588 -3246
rect 647 -3223 734 -3216
rect 647 -3226 708 -3223
rect 647 -3246 656 -3226
rect 676 -3243 708 -3226
rect 729 -3243 734 -3223
rect 676 -3246 734 -3243
rect 647 -3253 734 -3246
rect 759 -3226 796 -3156
rect 1062 -3157 1099 -3156
rect 1394 -3164 1432 -3156
rect 1498 -3132 1583 -3126
rect 1608 -3127 1645 -3126
rect 1498 -3152 1506 -3132
rect 1526 -3152 1583 -3132
rect 1498 -3160 1583 -3152
rect 1607 -3136 1645 -3127
rect 1607 -3156 1616 -3136
rect 1636 -3156 1645 -3136
rect 1498 -3161 1534 -3160
rect 1607 -3164 1645 -3156
rect 1711 -3132 1796 -3126
rect 1816 -3127 1853 -3126
rect 1711 -3152 1719 -3132
rect 1739 -3133 1796 -3132
rect 1739 -3152 1768 -3133
rect 1711 -3153 1768 -3152
rect 1789 -3153 1796 -3133
rect 1711 -3160 1796 -3153
rect 1815 -3136 1853 -3127
rect 1815 -3156 1824 -3136
rect 1844 -3156 1853 -3136
rect 1711 -3161 1747 -3160
rect 1815 -3164 1853 -3156
rect 1919 -3132 2063 -3126
rect 1919 -3152 1927 -3132
rect 1947 -3133 2035 -3132
rect 1947 -3152 1980 -3133
rect 2003 -3152 2035 -3133
rect 2055 -3152 2063 -3132
rect 1919 -3160 2063 -3152
rect 1919 -3161 1955 -3160
rect 2027 -3161 2063 -3160
rect 2129 -3127 2166 -3126
rect 2129 -3128 2167 -3127
rect 2129 -3136 2193 -3128
rect 2129 -3156 2138 -3136
rect 2158 -3150 2193 -3136
rect 2213 -3150 2216 -3130
rect 2158 -3155 2216 -3150
rect 2158 -3156 2193 -3155
rect 1395 -3193 1432 -3164
rect 1396 -3195 1432 -3193
rect 1608 -3195 1645 -3164
rect 911 -3216 947 -3215
rect 759 -3246 768 -3226
rect 788 -3246 796 -3226
rect 647 -3255 703 -3253
rect 647 -3256 684 -3255
rect 759 -3256 796 -3246
rect 855 -3226 1003 -3216
rect 1396 -3217 1645 -3195
rect 1816 -3196 1853 -3164
rect 2129 -3168 2193 -3156
rect 2233 -3194 2260 -3016
rect 2092 -3196 2260 -3194
rect 1816 -3207 2260 -3196
rect 2323 -3196 2353 -2195
rect 2442 -2202 2479 -2191
rect 2323 -3201 2355 -3196
rect 1103 -3219 1199 -3217
rect 855 -3246 864 -3226
rect 884 -3246 974 -3226
rect 994 -3246 1003 -3226
rect 855 -3255 1003 -3246
rect 1061 -3226 1199 -3219
rect 1816 -3222 2262 -3207
rect 2092 -3223 2262 -3222
rect 1061 -3246 1070 -3226
rect 1090 -3246 1199 -3226
rect 1061 -3255 1199 -3246
rect 855 -3256 892 -3255
rect 911 -3307 947 -3255
rect 966 -3256 1003 -3255
rect 1062 -3256 1099 -3255
rect 382 -3309 423 -3308
rect 144 -3473 183 -3324
rect 274 -3316 423 -3309
rect 274 -3336 392 -3316
rect 412 -3336 423 -3316
rect 274 -3344 423 -3336
rect 490 -3312 849 -3308
rect 490 -3317 812 -3312
rect 490 -3341 603 -3317
rect 627 -3336 812 -3317
rect 836 -3336 849 -3312
rect 627 -3341 849 -3336
rect 490 -3344 849 -3341
rect 911 -3344 946 -3307
rect 1014 -3310 1114 -3307
rect 1014 -3314 1081 -3310
rect 1014 -3340 1026 -3314
rect 1052 -3336 1081 -3314
rect 1107 -3336 1114 -3310
rect 1052 -3340 1114 -3336
rect 1014 -3344 1114 -3340
rect 490 -3365 521 -3344
rect 911 -3365 947 -3344
rect 333 -3366 370 -3365
rect 332 -3375 370 -3366
rect 332 -3395 341 -3375
rect 361 -3395 370 -3375
rect 332 -3403 370 -3395
rect 436 -3371 521 -3365
rect 546 -3366 583 -3365
rect 436 -3391 444 -3371
rect 464 -3391 521 -3371
rect 436 -3399 521 -3391
rect 545 -3375 583 -3366
rect 545 -3395 554 -3375
rect 574 -3395 583 -3375
rect 436 -3400 472 -3399
rect 545 -3403 583 -3395
rect 649 -3371 734 -3365
rect 754 -3366 791 -3365
rect 649 -3391 657 -3371
rect 677 -3372 734 -3371
rect 677 -3391 706 -3372
rect 649 -3392 706 -3391
rect 727 -3392 734 -3372
rect 649 -3399 734 -3392
rect 753 -3375 791 -3366
rect 753 -3395 762 -3375
rect 782 -3395 791 -3375
rect 649 -3400 685 -3399
rect 753 -3403 791 -3395
rect 857 -3370 1001 -3365
rect 857 -3371 922 -3370
rect 857 -3391 865 -3371
rect 885 -3391 922 -3371
rect 944 -3371 1001 -3370
rect 944 -3391 973 -3371
rect 993 -3391 1001 -3371
rect 857 -3399 1001 -3391
rect 857 -3400 893 -3399
rect 965 -3400 1001 -3399
rect 1067 -3366 1104 -3365
rect 1067 -3367 1105 -3366
rect 1067 -3375 1131 -3367
rect 1067 -3395 1076 -3375
rect 1096 -3389 1131 -3375
rect 1151 -3389 1154 -3369
rect 1096 -3394 1154 -3389
rect 1096 -3395 1131 -3394
rect 333 -3432 370 -3403
rect 334 -3434 370 -3432
rect 546 -3434 583 -3403
rect 334 -3456 583 -3434
rect 754 -3435 791 -3403
rect 1067 -3407 1131 -3395
rect 1171 -3433 1198 -3255
rect 1030 -3435 1198 -3433
rect 754 -3461 1198 -3435
rect 1350 -3336 1600 -3312
rect 1350 -3407 1387 -3336
rect 1502 -3397 1533 -3396
rect 1350 -3427 1359 -3407
rect 1379 -3427 1387 -3407
rect 1350 -3437 1387 -3427
rect 1446 -3407 1533 -3397
rect 1446 -3427 1455 -3407
rect 1475 -3427 1533 -3407
rect 1446 -3436 1533 -3427
rect 1446 -3437 1483 -3436
rect 754 -3471 776 -3461
rect 1030 -3462 1198 -3461
rect 714 -3473 776 -3471
rect 144 -3480 776 -3473
rect 143 -3489 776 -3480
rect 1502 -3489 1533 -3436
rect 1563 -3407 1600 -3336
rect 1771 -3331 2164 -3311
rect 2184 -3331 2187 -3311
rect 1771 -3336 2187 -3331
rect 1771 -3337 2112 -3336
rect 1715 -3397 1746 -3396
rect 1563 -3427 1572 -3407
rect 1592 -3427 1600 -3407
rect 1563 -3437 1600 -3427
rect 1659 -3404 1746 -3397
rect 1659 -3407 1720 -3404
rect 1659 -3427 1668 -3407
rect 1688 -3424 1720 -3407
rect 1741 -3424 1746 -3404
rect 1688 -3427 1746 -3424
rect 1659 -3434 1746 -3427
rect 1771 -3407 1808 -3337
rect 2074 -3338 2111 -3337
rect 1923 -3397 1959 -3396
rect 1771 -3427 1780 -3407
rect 1800 -3427 1808 -3407
rect 1659 -3436 1715 -3434
rect 1659 -3437 1696 -3436
rect 1771 -3437 1808 -3427
rect 1867 -3407 2015 -3397
rect 2115 -3400 2211 -3398
rect 1867 -3427 1876 -3407
rect 1896 -3427 1986 -3407
rect 2006 -3427 2015 -3407
rect 1867 -3436 2015 -3427
rect 2073 -3407 2211 -3400
rect 2073 -3427 2082 -3407
rect 2102 -3427 2211 -3407
rect 2073 -3436 2211 -3427
rect 1867 -3437 1904 -3436
rect 1923 -3488 1959 -3436
rect 1978 -3437 2015 -3436
rect 2074 -3437 2111 -3436
rect 143 -3507 153 -3489
rect 171 -3490 776 -3489
rect 1394 -3490 1435 -3489
rect 171 -3495 192 -3490
rect 171 -3507 183 -3495
rect 1286 -3497 1435 -3490
rect 143 -3515 183 -3507
rect 226 -3508 252 -3507
rect 143 -3517 180 -3515
rect 226 -3526 780 -3508
rect 1286 -3517 1404 -3497
rect 1424 -3517 1435 -3497
rect 1286 -3525 1435 -3517
rect 1502 -3493 1861 -3489
rect 1502 -3498 1824 -3493
rect 1502 -3522 1615 -3498
rect 1639 -3517 1824 -3498
rect 1848 -3517 1861 -3493
rect 1639 -3522 1861 -3517
rect 1502 -3525 1861 -3522
rect 1923 -3525 1958 -3488
rect 2026 -3491 2126 -3488
rect 2026 -3495 2093 -3491
rect 2026 -3521 2038 -3495
rect 2064 -3517 2093 -3495
rect 2119 -3517 2126 -3491
rect 2064 -3521 2126 -3517
rect 2026 -3525 2126 -3521
rect 146 -3585 183 -3579
rect 226 -3585 252 -3526
rect 759 -3545 780 -3526
rect 146 -3588 252 -3585
rect 146 -3606 155 -3588
rect 173 -3602 252 -3588
rect 337 -3570 587 -3546
rect 173 -3604 249 -3602
rect 173 -3606 183 -3604
rect 146 -3616 183 -3606
rect 151 -3681 182 -3616
rect 337 -3641 374 -3570
rect 489 -3631 520 -3630
rect 337 -3661 346 -3641
rect 366 -3661 374 -3641
rect 337 -3671 374 -3661
rect 433 -3641 520 -3631
rect 433 -3661 442 -3641
rect 462 -3661 520 -3641
rect 433 -3670 520 -3661
rect 433 -3671 470 -3670
rect 150 -3690 187 -3681
rect 150 -3708 160 -3690
rect 178 -3708 187 -3690
rect 150 -3718 187 -3708
rect 489 -3723 520 -3670
rect 550 -3641 587 -3570
rect 758 -3565 1151 -3545
rect 1171 -3565 1174 -3545
rect 1502 -3546 1533 -3525
rect 1923 -3546 1959 -3525
rect 1345 -3547 1382 -3546
rect 758 -3570 1174 -3565
rect 1344 -3556 1382 -3547
rect 758 -3571 1099 -3570
rect 702 -3631 733 -3630
rect 550 -3661 559 -3641
rect 579 -3661 587 -3641
rect 550 -3671 587 -3661
rect 646 -3638 733 -3631
rect 646 -3641 707 -3638
rect 646 -3661 655 -3641
rect 675 -3658 707 -3641
rect 728 -3658 733 -3638
rect 675 -3661 733 -3658
rect 646 -3668 733 -3661
rect 758 -3641 795 -3571
rect 1061 -3572 1098 -3571
rect 1344 -3576 1353 -3556
rect 1373 -3576 1382 -3556
rect 1344 -3584 1382 -3576
rect 1448 -3552 1533 -3546
rect 1558 -3547 1595 -3546
rect 1448 -3572 1456 -3552
rect 1476 -3572 1533 -3552
rect 1448 -3580 1533 -3572
rect 1557 -3556 1595 -3547
rect 1557 -3576 1566 -3556
rect 1586 -3576 1595 -3556
rect 1448 -3581 1484 -3580
rect 1557 -3584 1595 -3576
rect 1661 -3552 1746 -3546
rect 1766 -3547 1803 -3546
rect 1661 -3572 1669 -3552
rect 1689 -3553 1746 -3552
rect 1689 -3572 1718 -3553
rect 1661 -3573 1718 -3572
rect 1739 -3573 1746 -3553
rect 1661 -3580 1746 -3573
rect 1765 -3556 1803 -3547
rect 1765 -3576 1774 -3556
rect 1794 -3576 1803 -3556
rect 1661 -3581 1697 -3580
rect 1765 -3584 1803 -3576
rect 1869 -3551 2013 -3546
rect 1869 -3552 1928 -3551
rect 1869 -3572 1877 -3552
rect 1897 -3571 1928 -3552
rect 1952 -3552 2013 -3551
rect 1952 -3571 1985 -3552
rect 1897 -3572 1985 -3571
rect 2005 -3572 2013 -3552
rect 1869 -3580 2013 -3572
rect 1869 -3581 1905 -3580
rect 1977 -3581 2013 -3580
rect 2079 -3547 2116 -3546
rect 2079 -3548 2117 -3547
rect 2079 -3556 2143 -3548
rect 2079 -3576 2088 -3556
rect 2108 -3570 2143 -3556
rect 2163 -3570 2166 -3550
rect 2108 -3575 2166 -3570
rect 2108 -3576 2143 -3575
rect 1345 -3613 1382 -3584
rect 1346 -3615 1382 -3613
rect 1558 -3615 1595 -3584
rect 910 -3631 946 -3630
rect 758 -3661 767 -3641
rect 787 -3661 795 -3641
rect 646 -3670 702 -3668
rect 646 -3671 683 -3670
rect 758 -3671 795 -3661
rect 854 -3641 1002 -3631
rect 1102 -3634 1198 -3632
rect 854 -3661 863 -3641
rect 883 -3661 973 -3641
rect 993 -3661 1002 -3641
rect 854 -3670 1002 -3661
rect 1060 -3641 1198 -3634
rect 1346 -3637 1595 -3615
rect 1766 -3616 1803 -3584
rect 2079 -3588 2143 -3576
rect 2183 -3614 2210 -3436
rect 2042 -3616 2210 -3614
rect 1766 -3620 2210 -3616
rect 1060 -3661 1069 -3641
rect 1089 -3661 1198 -3641
rect 1766 -3639 1815 -3620
rect 1835 -3639 2210 -3620
rect 1766 -3642 2210 -3639
rect 2042 -3643 2210 -3642
rect 2231 -3617 2262 -3223
rect 2323 -3219 2328 -3201
rect 2348 -3219 2355 -3201
rect 2323 -3224 2355 -3219
rect 2326 -3226 2355 -3224
rect 2231 -3643 2236 -3617
rect 2255 -3643 2262 -3617
rect 2231 -3646 2262 -3643
rect 1060 -3670 1198 -3661
rect 854 -3671 891 -3670
rect 910 -3722 946 -3670
rect 965 -3671 1002 -3670
rect 1061 -3671 1098 -3670
rect 381 -3724 422 -3723
rect 273 -3731 422 -3724
rect 273 -3751 391 -3731
rect 411 -3751 422 -3731
rect 273 -3759 422 -3751
rect 489 -3727 848 -3723
rect 489 -3732 811 -3727
rect 489 -3756 602 -3732
rect 626 -3751 811 -3732
rect 835 -3751 848 -3727
rect 626 -3756 848 -3751
rect 489 -3759 848 -3756
rect 910 -3759 945 -3722
rect 1013 -3725 1113 -3722
rect 1013 -3729 1080 -3725
rect 1013 -3755 1025 -3729
rect 1051 -3751 1080 -3729
rect 1106 -3751 1113 -3725
rect 1051 -3755 1113 -3751
rect 1013 -3759 1113 -3755
rect 489 -3780 520 -3759
rect 910 -3780 946 -3759
rect 153 -3789 190 -3780
rect 332 -3781 369 -3780
rect 153 -3807 162 -3789
rect 180 -3807 190 -3789
rect 153 -3817 190 -3807
rect 154 -3852 190 -3817
rect 331 -3790 369 -3781
rect 331 -3810 340 -3790
rect 360 -3810 369 -3790
rect 331 -3818 369 -3810
rect 435 -3786 520 -3780
rect 545 -3781 582 -3780
rect 435 -3806 443 -3786
rect 463 -3806 520 -3786
rect 435 -3814 520 -3806
rect 544 -3790 582 -3781
rect 544 -3810 553 -3790
rect 573 -3810 582 -3790
rect 435 -3815 471 -3814
rect 544 -3818 582 -3810
rect 648 -3786 733 -3780
rect 753 -3781 790 -3780
rect 648 -3806 656 -3786
rect 676 -3787 733 -3786
rect 676 -3806 705 -3787
rect 648 -3807 705 -3806
rect 726 -3807 733 -3787
rect 648 -3814 733 -3807
rect 752 -3790 790 -3781
rect 752 -3810 761 -3790
rect 781 -3810 790 -3790
rect 648 -3815 684 -3814
rect 752 -3818 790 -3810
rect 856 -3786 1000 -3780
rect 856 -3806 864 -3786
rect 884 -3787 972 -3786
rect 884 -3806 912 -3787
rect 856 -3808 912 -3806
rect 934 -3806 972 -3787
rect 992 -3806 1000 -3786
rect 934 -3808 1000 -3806
rect 856 -3814 1000 -3808
rect 856 -3815 892 -3814
rect 964 -3815 1000 -3814
rect 1066 -3781 1103 -3780
rect 1066 -3782 1104 -3781
rect 1066 -3790 1130 -3782
rect 1066 -3810 1075 -3790
rect 1095 -3804 1130 -3790
rect 1150 -3804 1153 -3784
rect 1095 -3809 1153 -3804
rect 1095 -3810 1130 -3809
rect 332 -3847 369 -3818
rect 152 -3893 190 -3852
rect 333 -3849 369 -3847
rect 545 -3849 582 -3818
rect 333 -3871 582 -3849
rect 753 -3850 790 -3818
rect 1066 -3822 1130 -3810
rect 1170 -3848 1197 -3670
rect 1029 -3850 1197 -3848
rect 753 -3876 1197 -3850
rect 754 -3893 778 -3876
rect 1029 -3877 1197 -3876
rect 152 -3911 779 -3893
rect 152 -3917 190 -3911
<< viali >>
rect 1115 3708 1135 3728
rect 671 3615 692 3635
rect 1044 3522 1070 3548
rect 669 3466 690 3486
rect 885 3467 907 3488
rect 1094 3469 1114 3489
rect 2127 3527 2147 3547
rect 1683 3434 1704 3454
rect 2056 3341 2082 3367
rect 1114 3293 1134 3313
rect 670 3200 691 3220
rect 1681 3285 1702 3305
rect 1892 3286 1916 3306
rect 2106 3288 2126 3308
rect 1778 3219 1798 3238
rect 1043 3107 1069 3133
rect 668 3051 689 3071
rect 875 3050 897 3071
rect 1093 3054 1113 3074
rect 2182 2966 2202 2986
rect 1738 2873 1759 2893
rect 2111 2780 2137 2806
rect 1120 2727 1140 2747
rect 676 2634 697 2654
rect 1736 2724 1757 2744
rect 1951 2726 1975 2743
rect 2161 2727 2181 2747
rect 1049 2541 1075 2567
rect 674 2485 695 2505
rect 890 2486 912 2507
rect 1099 2488 1119 2508
rect 2132 2546 2152 2566
rect 1688 2453 1709 2473
rect 2061 2360 2087 2386
rect 1119 2312 1139 2332
rect 675 2219 696 2239
rect 1686 2304 1707 2324
rect 1896 2306 1920 2326
rect 2111 2307 2131 2327
rect 1783 2238 1803 2257
rect 2204 2234 2223 2260
rect 1048 2126 1074 2152
rect 673 2070 694 2090
rect 880 2069 902 2090
rect 1098 2073 1118 2093
rect 2347 2034 2367 2054
rect 1903 1941 1924 1961
rect 2276 1848 2302 1874
rect 1901 1792 1922 1812
rect 2110 1791 2135 1817
rect 2326 1795 2346 1815
rect 1127 1748 1147 1768
rect 683 1655 704 1675
rect 1056 1562 1082 1588
rect 681 1506 702 1526
rect 897 1507 919 1528
rect 1106 1509 1126 1529
rect 2139 1567 2159 1587
rect 1695 1474 1716 1494
rect 2068 1381 2094 1407
rect 1126 1333 1146 1353
rect 682 1240 703 1260
rect 1693 1325 1714 1345
rect 1904 1326 1928 1346
rect 2118 1328 2138 1348
rect 1790 1259 1810 1278
rect 1055 1147 1081 1173
rect 680 1091 701 1111
rect 887 1090 909 1111
rect 1105 1094 1125 1114
rect 2194 1006 2214 1026
rect 1750 913 1771 933
rect 2123 820 2149 846
rect 1132 767 1152 787
rect 688 674 709 694
rect 1748 764 1769 784
rect 1960 765 1983 784
rect 2173 767 2193 787
rect 1061 581 1087 607
rect 686 525 707 545
rect 902 526 924 547
rect 1111 528 1131 548
rect 2144 586 2164 606
rect 1700 493 1721 513
rect 2073 400 2099 426
rect 1131 352 1151 372
rect 687 259 708 279
rect 1698 344 1719 364
rect 1908 346 1932 366
rect 2123 347 2143 367
rect 1795 278 1815 297
rect 2308 698 2328 716
rect 2216 274 2235 300
rect 1060 166 1086 192
rect 685 110 706 130
rect 892 109 914 130
rect 1110 113 1130 133
rect 2442 42 2462 62
rect 1998 -51 2019 -31
rect 2371 -144 2397 -118
rect 1135 -209 1155 -189
rect 1996 -200 2017 -180
rect 2211 -197 2237 -178
rect 2421 -197 2441 -177
rect 691 -302 712 -282
rect 1064 -395 1090 -369
rect 689 -451 710 -431
rect 905 -450 927 -429
rect 1114 -448 1134 -428
rect 2147 -390 2167 -370
rect 1703 -483 1724 -463
rect 2076 -576 2102 -550
rect 1134 -624 1154 -604
rect 690 -717 711 -697
rect 1701 -632 1722 -612
rect 1912 -631 1936 -611
rect 2126 -629 2146 -609
rect 1798 -698 1818 -679
rect 1063 -810 1089 -784
rect 688 -866 709 -846
rect 895 -867 917 -846
rect 1113 -863 1133 -843
rect 2202 -951 2222 -931
rect 1758 -1044 1779 -1024
rect 2131 -1137 2157 -1111
rect 1140 -1190 1160 -1170
rect 696 -1283 717 -1263
rect 1756 -1193 1777 -1173
rect 1971 -1191 1995 -1174
rect 2181 -1190 2201 -1170
rect 1069 -1376 1095 -1350
rect 694 -1432 715 -1412
rect 910 -1431 932 -1410
rect 1119 -1429 1139 -1409
rect 2152 -1371 2172 -1351
rect 1708 -1464 1729 -1444
rect 2081 -1557 2107 -1531
rect 1139 -1605 1159 -1585
rect 695 -1698 716 -1678
rect 1706 -1613 1727 -1593
rect 1916 -1611 1940 -1591
rect 2131 -1610 2151 -1590
rect 1803 -1679 1823 -1660
rect 2224 -1683 2243 -1657
rect 1068 -1791 1094 -1765
rect 693 -1847 714 -1827
rect 900 -1848 922 -1827
rect 1118 -1844 1138 -1824
rect 2367 -1883 2387 -1863
rect 1923 -1976 1944 -1956
rect 2296 -2069 2322 -2043
rect 1921 -2125 1942 -2105
rect 2136 -2123 2159 -2104
rect 2346 -2122 2366 -2102
rect 1147 -2169 1167 -2149
rect 703 -2262 724 -2242
rect 2448 -2191 2471 -2172
rect 1076 -2355 1102 -2329
rect 701 -2411 722 -2391
rect 917 -2410 939 -2389
rect 1126 -2408 1146 -2388
rect 2159 -2350 2179 -2330
rect 1715 -2443 1736 -2423
rect 2088 -2536 2114 -2510
rect 1146 -2584 1166 -2564
rect 702 -2677 723 -2657
rect 1713 -2592 1734 -2572
rect 1924 -2591 1948 -2571
rect 2138 -2589 2158 -2569
rect 1810 -2658 1830 -2639
rect 1075 -2770 1101 -2744
rect 700 -2826 721 -2806
rect 907 -2827 929 -2806
rect 1125 -2823 1145 -2803
rect 2214 -2911 2234 -2891
rect 1770 -3004 1791 -2984
rect 2143 -3097 2169 -3071
rect 1152 -3150 1172 -3130
rect 708 -3243 729 -3223
rect 1768 -3153 1789 -3133
rect 1980 -3152 2003 -3133
rect 2193 -3150 2213 -3130
rect 1081 -3336 1107 -3310
rect 706 -3392 727 -3372
rect 922 -3391 944 -3370
rect 1131 -3389 1151 -3369
rect 2164 -3331 2184 -3311
rect 1720 -3424 1741 -3404
rect 2093 -3517 2119 -3491
rect 1151 -3565 1171 -3545
rect 707 -3658 728 -3638
rect 1718 -3573 1739 -3553
rect 1928 -3571 1952 -3551
rect 2143 -3570 2163 -3550
rect 1815 -3639 1835 -3620
rect 2328 -3219 2348 -3201
rect 2236 -3643 2255 -3617
rect 1080 -3751 1106 -3725
rect 705 -3807 726 -3787
rect 912 -3808 934 -3787
rect 1130 -3804 1150 -3784
<< metal1 >>
rect 1111 3733 1143 3734
rect 1108 3728 1143 3733
rect 1108 3708 1115 3728
rect 1135 3708 1143 3728
rect 1108 3700 1143 3708
rect 664 3635 696 3642
rect 664 3615 671 3635
rect 692 3615 696 3635
rect 664 3550 696 3615
rect 1034 3550 1074 3551
rect 664 3548 1076 3550
rect 664 3522 1044 3548
rect 1070 3522 1076 3548
rect 664 3514 1076 3522
rect 664 3486 696 3514
rect 1109 3494 1143 3700
rect 664 3466 669 3486
rect 690 3466 696 3486
rect 664 3459 696 3466
rect 873 3488 913 3493
rect 873 3467 885 3488
rect 907 3467 913 3488
rect 873 3455 913 3467
rect 1087 3489 1143 3494
rect 1087 3469 1094 3489
rect 1114 3469 1143 3489
rect 1087 3462 1143 3469
rect 1200 3563 2157 3582
rect 1087 3461 1122 3462
rect 879 3423 907 3455
rect 1200 3423 1231 3563
rect 2120 3547 2155 3563
rect 2120 3527 2127 3547
rect 2147 3527 2155 3547
rect 2120 3519 2155 3527
rect 879 3392 1231 3423
rect 1676 3454 1708 3461
rect 1676 3434 1683 3454
rect 1704 3434 1708 3454
rect 1676 3369 1708 3434
rect 2046 3369 2086 3370
rect 1676 3367 2088 3369
rect 1676 3341 2056 3367
rect 2082 3341 2088 3367
rect 1676 3333 2088 3341
rect 1110 3318 1142 3319
rect 1107 3313 1142 3318
rect 1107 3293 1114 3313
rect 1134 3293 1142 3313
rect 1107 3285 1142 3293
rect 663 3220 695 3227
rect 663 3200 670 3220
rect 691 3200 695 3220
rect 663 3135 695 3200
rect 1033 3135 1073 3136
rect 663 3133 1075 3135
rect 663 3107 1043 3133
rect 1069 3107 1075 3133
rect 663 3099 1075 3107
rect 663 3071 695 3099
rect 663 3051 668 3071
rect 689 3051 695 3071
rect 663 3044 695 3051
rect 863 3071 913 3080
rect 1108 3079 1142 3285
rect 1676 3305 1708 3333
rect 1676 3285 1681 3305
rect 1702 3285 1708 3305
rect 1676 3278 1708 3285
rect 1883 3306 1925 3314
rect 2121 3313 2155 3519
rect 1883 3286 1892 3306
rect 1916 3286 1925 3306
rect 1883 3274 1925 3286
rect 2099 3308 2155 3313
rect 2099 3288 2106 3308
rect 2126 3288 2155 3308
rect 2099 3281 2155 3288
rect 2099 3280 2134 3281
rect 1885 3245 1920 3274
rect 1885 3244 2195 3245
rect 1770 3238 1806 3242
rect 1770 3219 1778 3238
rect 1798 3219 1806 3238
rect 1770 3216 1806 3219
rect 1771 3188 1805 3216
rect 1885 3210 2212 3244
rect 863 3050 875 3071
rect 897 3050 913 3071
rect 863 3042 913 3050
rect 1086 3074 1142 3079
rect 1086 3054 1093 3074
rect 1113 3054 1142 3074
rect 1086 3047 1142 3054
rect 1243 3160 1806 3188
rect 1086 3046 1121 3047
rect 868 3009 909 3042
rect 1243 3009 1283 3160
rect 868 2980 1283 3009
rect 2172 2986 2212 3210
rect 868 2979 1277 2980
rect 2172 2966 2182 2986
rect 2202 2966 2212 2986
rect 2172 2956 2212 2966
rect 1731 2893 1763 2900
rect 1731 2873 1738 2893
rect 1759 2873 1763 2893
rect 1731 2808 1763 2873
rect 2101 2808 2141 2809
rect 1731 2806 2143 2808
rect 1731 2780 2111 2806
rect 2137 2780 2143 2806
rect 1731 2772 2143 2780
rect 1116 2752 1148 2753
rect 1113 2747 1148 2752
rect 1113 2727 1120 2747
rect 1140 2727 1148 2747
rect 1113 2719 1148 2727
rect 669 2654 701 2661
rect 669 2634 676 2654
rect 697 2634 701 2654
rect 669 2569 701 2634
rect 1039 2569 1079 2570
rect 669 2567 1081 2569
rect 669 2541 1049 2567
rect 1075 2541 1081 2567
rect 669 2533 1081 2541
rect 669 2505 701 2533
rect 1114 2513 1148 2719
rect 1731 2744 1763 2772
rect 1731 2724 1736 2744
rect 1757 2724 1763 2744
rect 1731 2717 1763 2724
rect 1942 2743 1980 2755
rect 2176 2752 2210 2956
rect 1942 2726 1951 2743
rect 1975 2726 1980 2743
rect 1942 2683 1980 2726
rect 2154 2747 2210 2752
rect 2154 2727 2161 2747
rect 2181 2727 2210 2747
rect 2154 2720 2210 2727
rect 2154 2719 2189 2720
rect 2288 2683 2372 2688
rect 1942 2654 2372 2683
rect 669 2485 674 2505
rect 695 2485 701 2505
rect 669 2478 701 2485
rect 878 2507 918 2512
rect 878 2486 890 2507
rect 912 2486 918 2507
rect 878 2474 918 2486
rect 1092 2508 1148 2513
rect 1092 2488 1099 2508
rect 1119 2488 1148 2508
rect 1092 2481 1148 2488
rect 1205 2582 2162 2601
rect 1092 2480 1127 2481
rect 884 2442 912 2474
rect 1205 2442 1236 2582
rect 2125 2566 2160 2582
rect 2125 2546 2132 2566
rect 2152 2546 2160 2566
rect 2125 2538 2160 2546
rect 884 2411 1236 2442
rect 1681 2473 1713 2480
rect 1681 2453 1688 2473
rect 1709 2453 1713 2473
rect 1681 2388 1713 2453
rect 2051 2388 2091 2389
rect 1681 2386 2093 2388
rect 1681 2360 2061 2386
rect 2087 2360 2093 2386
rect 1681 2352 2093 2360
rect 1115 2337 1147 2338
rect 1112 2332 1147 2337
rect 1112 2312 1119 2332
rect 1139 2312 1147 2332
rect 1112 2304 1147 2312
rect 668 2239 700 2246
rect 668 2219 675 2239
rect 696 2219 700 2239
rect 668 2154 700 2219
rect 1038 2154 1078 2155
rect 668 2152 1080 2154
rect 668 2126 1048 2152
rect 1074 2126 1080 2152
rect 668 2118 1080 2126
rect 668 2090 700 2118
rect 668 2070 673 2090
rect 694 2070 700 2090
rect 668 2063 700 2070
rect 868 2090 918 2099
rect 1113 2098 1147 2304
rect 1681 2324 1713 2352
rect 1681 2304 1686 2324
rect 1707 2304 1713 2324
rect 1886 2326 1928 2335
rect 2126 2332 2160 2538
rect 1886 2312 1896 2326
rect 1681 2297 1713 2304
rect 1885 2306 1896 2312
rect 1920 2306 1928 2326
rect 1885 2295 1928 2306
rect 2104 2327 2160 2332
rect 2104 2307 2111 2327
rect 2131 2307 2160 2327
rect 2104 2300 2160 2307
rect 2104 2299 2139 2300
rect 1885 2265 1925 2295
rect 1775 2257 1811 2261
rect 1775 2238 1783 2257
rect 1803 2238 1811 2257
rect 1775 2235 1811 2238
rect 1885 2260 2232 2265
rect 1776 2207 1810 2235
rect 1885 2234 2204 2260
rect 2223 2234 2232 2260
rect 1885 2230 2232 2234
rect 868 2069 880 2090
rect 902 2069 918 2090
rect 868 2061 918 2069
rect 1091 2093 1147 2098
rect 1091 2073 1098 2093
rect 1118 2073 1147 2093
rect 1091 2066 1147 2073
rect 1248 2179 1811 2207
rect 1091 2065 1126 2066
rect 873 2028 914 2061
rect 1248 2028 1288 2179
rect 2337 2060 2372 2654
rect 2337 2054 2375 2060
rect 2337 2034 2347 2054
rect 2367 2034 2375 2054
rect 2337 2032 2375 2034
rect 873 1999 1288 2028
rect 2340 2026 2375 2032
rect 873 1998 1282 1999
rect 1896 1961 1928 1968
rect 1896 1941 1903 1961
rect 1924 1941 1928 1961
rect 1896 1876 1928 1941
rect 2266 1876 2306 1877
rect 1896 1874 2308 1876
rect 1896 1848 2276 1874
rect 2302 1848 2308 1874
rect 1896 1840 2308 1848
rect 1896 1812 1928 1840
rect 1896 1792 1901 1812
rect 1922 1792 1928 1812
rect 1896 1785 1928 1792
rect 2100 1817 2147 1823
rect 2341 1820 2375 2026
rect 2100 1791 2110 1817
rect 2135 1791 2147 1817
rect 2100 1789 2147 1791
rect 2319 1815 2375 1820
rect 2319 1795 2326 1815
rect 2346 1795 2375 1815
rect 1123 1773 1155 1774
rect 1120 1768 1155 1773
rect 1120 1748 1127 1768
rect 1147 1748 1155 1768
rect 1120 1740 1155 1748
rect 676 1675 708 1682
rect 676 1655 683 1675
rect 704 1655 708 1675
rect 676 1590 708 1655
rect 1046 1590 1086 1591
rect 676 1588 1088 1590
rect 676 1562 1056 1588
rect 1082 1562 1088 1588
rect 676 1554 1088 1562
rect 676 1526 708 1554
rect 1121 1534 1155 1740
rect 2105 1754 2142 1789
rect 2319 1788 2375 1795
rect 2319 1787 2354 1788
rect 2439 1754 2471 1756
rect 2105 1721 2475 1754
rect 676 1506 681 1526
rect 702 1506 708 1526
rect 676 1499 708 1506
rect 885 1528 925 1533
rect 885 1507 897 1528
rect 919 1507 925 1528
rect 885 1495 925 1507
rect 1099 1529 1155 1534
rect 1099 1509 1106 1529
rect 1126 1509 1155 1529
rect 1099 1502 1155 1509
rect 1212 1603 2169 1622
rect 1099 1501 1134 1502
rect 891 1463 919 1495
rect 1212 1463 1243 1603
rect 2132 1587 2167 1603
rect 2132 1567 2139 1587
rect 2159 1567 2167 1587
rect 2132 1559 2167 1567
rect 891 1432 1243 1463
rect 1688 1494 1720 1501
rect 1688 1474 1695 1494
rect 1716 1474 1720 1494
rect 1688 1409 1720 1474
rect 2058 1409 2098 1410
rect 1688 1407 2100 1409
rect 1688 1381 2068 1407
rect 2094 1381 2100 1407
rect 1688 1373 2100 1381
rect 1122 1358 1154 1359
rect 1119 1353 1154 1358
rect 1119 1333 1126 1353
rect 1146 1333 1154 1353
rect 1119 1325 1154 1333
rect 675 1260 707 1267
rect 675 1240 682 1260
rect 703 1240 707 1260
rect 675 1175 707 1240
rect 1045 1175 1085 1176
rect 675 1173 1087 1175
rect 675 1147 1055 1173
rect 1081 1147 1087 1173
rect 675 1139 1087 1147
rect 675 1111 707 1139
rect 675 1091 680 1111
rect 701 1091 707 1111
rect 675 1084 707 1091
rect 875 1111 925 1120
rect 1120 1119 1154 1325
rect 1688 1345 1720 1373
rect 1688 1325 1693 1345
rect 1714 1325 1720 1345
rect 1688 1318 1720 1325
rect 1895 1346 1937 1354
rect 2133 1353 2167 1559
rect 1895 1326 1904 1346
rect 1928 1326 1937 1346
rect 1895 1314 1937 1326
rect 2111 1348 2167 1353
rect 2111 1328 2118 1348
rect 2138 1328 2167 1348
rect 2111 1321 2167 1328
rect 2111 1320 2146 1321
rect 1897 1285 1932 1314
rect 1897 1284 2207 1285
rect 1782 1278 1818 1282
rect 1782 1259 1790 1278
rect 1810 1259 1818 1278
rect 1782 1256 1818 1259
rect 1783 1228 1817 1256
rect 1897 1250 2224 1284
rect 875 1090 887 1111
rect 909 1090 925 1111
rect 875 1082 925 1090
rect 1098 1114 1154 1119
rect 1098 1094 1105 1114
rect 1125 1094 1154 1114
rect 1098 1087 1154 1094
rect 1255 1200 1818 1228
rect 1098 1086 1133 1087
rect 880 1049 921 1082
rect 1255 1049 1295 1200
rect 880 1020 1295 1049
rect 2184 1026 2224 1250
rect 880 1019 1289 1020
rect 2184 1006 2194 1026
rect 2214 1006 2224 1026
rect 2184 996 2224 1006
rect 1743 933 1775 940
rect 1743 913 1750 933
rect 1771 913 1775 933
rect 1743 848 1775 913
rect 2113 848 2153 849
rect 1743 846 2155 848
rect 1743 820 2123 846
rect 2149 820 2155 846
rect 1743 812 2155 820
rect 1128 792 1160 793
rect 1125 787 1160 792
rect 1125 767 1132 787
rect 1152 767 1160 787
rect 1125 759 1160 767
rect 681 694 713 701
rect 681 674 688 694
rect 709 674 713 694
rect 681 609 713 674
rect 1051 609 1091 610
rect 681 607 1093 609
rect 681 581 1061 607
rect 1087 581 1093 607
rect 681 573 1093 581
rect 681 545 713 573
rect 1126 553 1160 759
rect 1743 784 1775 812
rect 2188 792 2222 996
rect 1743 764 1748 784
rect 1769 764 1775 784
rect 1743 757 1775 764
rect 1954 784 1991 790
rect 1954 765 1960 784
rect 1983 765 1991 784
rect 1954 760 1991 765
rect 2166 787 2222 792
rect 2166 767 2173 787
rect 2193 767 2222 787
rect 2166 760 2222 767
rect 1962 723 1986 760
rect 2166 759 2201 760
rect 1962 721 2330 723
rect 1962 716 2335 721
rect 1962 698 2308 716
rect 2328 698 2335 716
rect 1962 693 2335 698
rect 2306 691 2335 693
rect 681 525 686 545
rect 707 525 713 545
rect 681 518 713 525
rect 890 547 930 552
rect 890 526 902 547
rect 924 526 930 547
rect 890 514 930 526
rect 1104 548 1160 553
rect 1104 528 1111 548
rect 1131 528 1160 548
rect 1104 521 1160 528
rect 1217 622 2174 641
rect 1104 520 1139 521
rect 896 482 924 514
rect 1217 482 1248 622
rect 2137 606 2172 622
rect 2137 586 2144 606
rect 2164 586 2172 606
rect 2137 578 2172 586
rect 896 451 1248 482
rect 1693 513 1725 520
rect 1693 493 1700 513
rect 1721 493 1725 513
rect 1693 428 1725 493
rect 2063 428 2103 429
rect 1693 426 2105 428
rect 1693 400 2073 426
rect 2099 400 2105 426
rect 1693 392 2105 400
rect 1127 377 1159 378
rect 1124 372 1159 377
rect 1124 352 1131 372
rect 1151 352 1159 372
rect 1124 344 1159 352
rect 680 279 712 286
rect 680 259 687 279
rect 708 259 712 279
rect 680 194 712 259
rect 1050 194 1090 195
rect 680 192 1092 194
rect 680 166 1060 192
rect 1086 166 1092 192
rect 680 158 1092 166
rect 680 130 712 158
rect 680 110 685 130
rect 706 110 712 130
rect 680 103 712 110
rect 880 130 930 139
rect 1125 138 1159 344
rect 1693 364 1725 392
rect 1693 344 1698 364
rect 1719 344 1725 364
rect 1898 366 1940 375
rect 2138 372 2172 578
rect 1898 352 1908 366
rect 1693 337 1725 344
rect 1897 346 1908 352
rect 1932 346 1940 366
rect 1897 335 1940 346
rect 2116 367 2172 372
rect 2116 347 2123 367
rect 2143 347 2172 367
rect 2116 340 2172 347
rect 2116 339 2151 340
rect 1897 305 1937 335
rect 1787 297 1823 301
rect 1787 278 1795 297
rect 1815 278 1823 297
rect 1787 275 1823 278
rect 1897 300 2244 305
rect 1788 247 1822 275
rect 1897 274 2216 300
rect 2235 274 2244 300
rect 1897 270 2244 274
rect 880 109 892 130
rect 914 109 930 130
rect 880 101 930 109
rect 1103 133 1159 138
rect 1103 113 1110 133
rect 1130 113 1159 133
rect 1103 106 1159 113
rect 1260 219 1823 247
rect 1103 105 1138 106
rect 885 68 926 101
rect 1260 68 1300 219
rect 2439 68 2471 1721
rect 885 39 1300 68
rect 2438 67 2471 68
rect 2435 62 2471 67
rect 2435 42 2442 62
rect 2462 42 2471 62
rect 885 38 1294 39
rect 2435 37 2471 42
rect 2435 34 2470 37
rect 1991 -31 2023 -24
rect 1991 -51 1998 -31
rect 2019 -51 2023 -31
rect 1991 -116 2023 -51
rect 2361 -116 2401 -115
rect 1991 -118 2403 -116
rect 1991 -144 2371 -118
rect 2397 -144 2403 -118
rect 1991 -152 2403 -144
rect 1991 -180 2023 -152
rect 1131 -184 1163 -183
rect 1128 -189 1163 -184
rect 1128 -209 1135 -189
rect 1155 -209 1163 -189
rect 1991 -200 1996 -180
rect 2017 -200 2023 -180
rect 1991 -207 2023 -200
rect 2196 -178 2245 -168
rect 2436 -172 2470 34
rect 2196 -197 2211 -178
rect 2237 -197 2245 -178
rect 2196 -206 2245 -197
rect 2414 -177 2470 -172
rect 2414 -197 2421 -177
rect 2441 -197 2470 -177
rect 2414 -204 2470 -197
rect 2414 -205 2449 -204
rect 1128 -217 1163 -209
rect 684 -282 716 -275
rect 684 -302 691 -282
rect 712 -302 716 -282
rect 684 -367 716 -302
rect 1054 -367 1094 -366
rect 684 -369 1096 -367
rect 684 -395 1064 -369
rect 1090 -395 1096 -369
rect 684 -403 1096 -395
rect 684 -431 716 -403
rect 1129 -423 1163 -217
rect 2205 -244 2240 -206
rect 2205 -274 2529 -244
rect 684 -451 689 -431
rect 710 -451 716 -431
rect 684 -458 716 -451
rect 893 -429 933 -424
rect 893 -450 905 -429
rect 927 -450 933 -429
rect 893 -462 933 -450
rect 1107 -428 1163 -423
rect 1107 -448 1114 -428
rect 1134 -448 1163 -428
rect 1107 -455 1163 -448
rect 1220 -354 2177 -335
rect 1107 -456 1142 -455
rect 899 -494 927 -462
rect 1220 -494 1251 -354
rect 2140 -370 2175 -354
rect 2140 -390 2147 -370
rect 2167 -390 2175 -370
rect 2140 -398 2175 -390
rect 899 -525 1251 -494
rect 1696 -463 1728 -456
rect 1696 -483 1703 -463
rect 1724 -483 1728 -463
rect 1696 -548 1728 -483
rect 2066 -548 2106 -547
rect 1696 -550 2108 -548
rect 1696 -576 2076 -550
rect 2102 -576 2108 -550
rect 1696 -584 2108 -576
rect 1130 -599 1162 -598
rect 1127 -604 1162 -599
rect 1127 -624 1134 -604
rect 1154 -624 1162 -604
rect 1127 -632 1162 -624
rect 683 -697 715 -690
rect 683 -717 690 -697
rect 711 -717 715 -697
rect 683 -782 715 -717
rect 1053 -782 1093 -781
rect 683 -784 1095 -782
rect 683 -810 1063 -784
rect 1089 -810 1095 -784
rect 683 -818 1095 -810
rect 683 -846 715 -818
rect 683 -866 688 -846
rect 709 -866 715 -846
rect 683 -873 715 -866
rect 883 -846 933 -837
rect 1128 -838 1162 -632
rect 1696 -612 1728 -584
rect 1696 -632 1701 -612
rect 1722 -632 1728 -612
rect 1696 -639 1728 -632
rect 1903 -611 1945 -603
rect 2141 -604 2175 -398
rect 1903 -631 1912 -611
rect 1936 -631 1945 -611
rect 1903 -643 1945 -631
rect 2119 -609 2175 -604
rect 2119 -629 2126 -609
rect 2146 -629 2175 -609
rect 2119 -636 2175 -629
rect 2119 -637 2154 -636
rect 1905 -672 1940 -643
rect 1905 -673 2215 -672
rect 1790 -679 1826 -675
rect 1790 -698 1798 -679
rect 1818 -698 1826 -679
rect 1790 -701 1826 -698
rect 1791 -729 1825 -701
rect 1905 -707 2232 -673
rect 883 -867 895 -846
rect 917 -867 933 -846
rect 883 -875 933 -867
rect 1106 -843 1162 -838
rect 1106 -863 1113 -843
rect 1133 -863 1162 -843
rect 1106 -870 1162 -863
rect 1263 -757 1826 -729
rect 1106 -871 1141 -870
rect 888 -908 929 -875
rect 1263 -908 1303 -757
rect 888 -937 1303 -908
rect 2192 -931 2232 -707
rect 888 -938 1297 -937
rect 2192 -951 2202 -931
rect 2222 -951 2232 -931
rect 2192 -961 2232 -951
rect 1751 -1024 1783 -1017
rect 1751 -1044 1758 -1024
rect 1779 -1044 1783 -1024
rect 1751 -1109 1783 -1044
rect 2121 -1109 2161 -1108
rect 1751 -1111 2163 -1109
rect 1751 -1137 2131 -1111
rect 2157 -1137 2163 -1111
rect 1751 -1145 2163 -1137
rect 1136 -1165 1168 -1164
rect 1133 -1170 1168 -1165
rect 1133 -1190 1140 -1170
rect 1160 -1190 1168 -1170
rect 1133 -1198 1168 -1190
rect 689 -1263 721 -1256
rect 689 -1283 696 -1263
rect 717 -1283 721 -1263
rect 689 -1348 721 -1283
rect 1059 -1348 1099 -1347
rect 689 -1350 1101 -1348
rect 689 -1376 1069 -1350
rect 1095 -1376 1101 -1350
rect 689 -1384 1101 -1376
rect 689 -1412 721 -1384
rect 1134 -1404 1168 -1198
rect 1751 -1173 1783 -1145
rect 1751 -1193 1756 -1173
rect 1777 -1193 1783 -1173
rect 1751 -1200 1783 -1193
rect 1962 -1174 2000 -1162
rect 2196 -1165 2230 -961
rect 1962 -1191 1971 -1174
rect 1995 -1191 2000 -1174
rect 1962 -1234 2000 -1191
rect 2174 -1170 2230 -1165
rect 2174 -1190 2181 -1170
rect 2201 -1190 2230 -1170
rect 2174 -1197 2230 -1190
rect 2174 -1198 2209 -1197
rect 2308 -1234 2392 -1229
rect 1962 -1263 2392 -1234
rect 689 -1432 694 -1412
rect 715 -1432 721 -1412
rect 689 -1439 721 -1432
rect 898 -1410 938 -1405
rect 898 -1431 910 -1410
rect 932 -1431 938 -1410
rect 898 -1443 938 -1431
rect 1112 -1409 1168 -1404
rect 1112 -1429 1119 -1409
rect 1139 -1429 1168 -1409
rect 1112 -1436 1168 -1429
rect 1225 -1335 2182 -1316
rect 1112 -1437 1147 -1436
rect 904 -1475 932 -1443
rect 1225 -1475 1256 -1335
rect 2145 -1351 2180 -1335
rect 2145 -1371 2152 -1351
rect 2172 -1371 2180 -1351
rect 2145 -1379 2180 -1371
rect 904 -1506 1256 -1475
rect 1701 -1444 1733 -1437
rect 1701 -1464 1708 -1444
rect 1729 -1464 1733 -1444
rect 1701 -1529 1733 -1464
rect 2071 -1529 2111 -1528
rect 1701 -1531 2113 -1529
rect 1701 -1557 2081 -1531
rect 2107 -1557 2113 -1531
rect 1701 -1565 2113 -1557
rect 1135 -1580 1167 -1579
rect 1132 -1585 1167 -1580
rect 1132 -1605 1139 -1585
rect 1159 -1605 1167 -1585
rect 1132 -1613 1167 -1605
rect 688 -1678 720 -1671
rect 688 -1698 695 -1678
rect 716 -1698 720 -1678
rect 688 -1763 720 -1698
rect 1058 -1763 1098 -1762
rect 688 -1765 1100 -1763
rect 688 -1791 1068 -1765
rect 1094 -1791 1100 -1765
rect 688 -1799 1100 -1791
rect 688 -1827 720 -1799
rect 688 -1847 693 -1827
rect 714 -1847 720 -1827
rect 688 -1854 720 -1847
rect 888 -1827 938 -1818
rect 1133 -1819 1167 -1613
rect 1701 -1593 1733 -1565
rect 1701 -1613 1706 -1593
rect 1727 -1613 1733 -1593
rect 1906 -1591 1948 -1582
rect 2146 -1585 2180 -1379
rect 1906 -1605 1916 -1591
rect 1701 -1620 1733 -1613
rect 1905 -1611 1916 -1605
rect 1940 -1611 1948 -1591
rect 1905 -1622 1948 -1611
rect 2124 -1590 2180 -1585
rect 2124 -1610 2131 -1590
rect 2151 -1610 2180 -1590
rect 2124 -1617 2180 -1610
rect 2124 -1618 2159 -1617
rect 1905 -1652 1945 -1622
rect 1795 -1660 1831 -1656
rect 1795 -1679 1803 -1660
rect 1823 -1679 1831 -1660
rect 1795 -1682 1831 -1679
rect 1905 -1657 2252 -1652
rect 1796 -1710 1830 -1682
rect 1905 -1683 2224 -1657
rect 2243 -1683 2252 -1657
rect 1905 -1687 2252 -1683
rect 888 -1848 900 -1827
rect 922 -1848 938 -1827
rect 888 -1856 938 -1848
rect 1111 -1824 1167 -1819
rect 1111 -1844 1118 -1824
rect 1138 -1844 1167 -1824
rect 1111 -1851 1167 -1844
rect 1268 -1738 1831 -1710
rect 1111 -1852 1146 -1851
rect 893 -1889 934 -1856
rect 1268 -1889 1308 -1738
rect 2357 -1857 2392 -1263
rect 2357 -1863 2395 -1857
rect 2357 -1883 2367 -1863
rect 2387 -1883 2395 -1863
rect 2357 -1885 2395 -1883
rect 893 -1918 1308 -1889
rect 2360 -1891 2395 -1885
rect 893 -1919 1302 -1918
rect 1916 -1956 1948 -1949
rect 1916 -1976 1923 -1956
rect 1944 -1976 1948 -1956
rect 1916 -2041 1948 -1976
rect 2286 -2041 2326 -2040
rect 1916 -2043 2328 -2041
rect 1916 -2069 2296 -2043
rect 2322 -2069 2328 -2043
rect 1916 -2077 2328 -2069
rect 1916 -2105 1948 -2077
rect 2361 -2097 2395 -1891
rect 1916 -2125 1921 -2105
rect 1942 -2125 1948 -2105
rect 1916 -2132 1948 -2125
rect 2125 -2104 2164 -2098
rect 2125 -2123 2136 -2104
rect 2159 -2123 2164 -2104
rect 2125 -2136 2164 -2123
rect 2339 -2102 2395 -2097
rect 2339 -2122 2346 -2102
rect 2366 -2122 2395 -2102
rect 2339 -2129 2395 -2122
rect 2339 -2130 2374 -2129
rect 1143 -2144 1175 -2143
rect 1140 -2149 1175 -2144
rect 1140 -2169 1147 -2149
rect 1167 -2169 1175 -2149
rect 1140 -2177 1175 -2169
rect 696 -2242 728 -2235
rect 696 -2262 703 -2242
rect 724 -2262 728 -2242
rect 696 -2327 728 -2262
rect 1066 -2327 1106 -2326
rect 696 -2329 1108 -2327
rect 696 -2355 1076 -2329
rect 1102 -2355 1108 -2329
rect 696 -2363 1108 -2355
rect 696 -2391 728 -2363
rect 1141 -2383 1175 -2177
rect 2132 -2167 2162 -2136
rect 2442 -2167 2479 -2161
rect 2132 -2172 2479 -2167
rect 2132 -2191 2448 -2172
rect 2471 -2191 2479 -2172
rect 2132 -2197 2479 -2191
rect 2442 -2202 2479 -2197
rect 696 -2411 701 -2391
rect 722 -2411 728 -2391
rect 696 -2418 728 -2411
rect 905 -2389 945 -2384
rect 905 -2410 917 -2389
rect 939 -2410 945 -2389
rect 905 -2422 945 -2410
rect 1119 -2388 1175 -2383
rect 1119 -2408 1126 -2388
rect 1146 -2408 1175 -2388
rect 1119 -2415 1175 -2408
rect 1232 -2314 2189 -2295
rect 1119 -2416 1154 -2415
rect 911 -2454 939 -2422
rect 1232 -2454 1263 -2314
rect 2152 -2330 2187 -2314
rect 2152 -2350 2159 -2330
rect 2179 -2350 2187 -2330
rect 2152 -2358 2187 -2350
rect 911 -2485 1263 -2454
rect 1708 -2423 1740 -2416
rect 1708 -2443 1715 -2423
rect 1736 -2443 1740 -2423
rect 1708 -2508 1740 -2443
rect 2078 -2508 2118 -2507
rect 1708 -2510 2120 -2508
rect 1708 -2536 2088 -2510
rect 2114 -2536 2120 -2510
rect 1708 -2544 2120 -2536
rect 1142 -2559 1174 -2558
rect 1139 -2564 1174 -2559
rect 1139 -2584 1146 -2564
rect 1166 -2584 1174 -2564
rect 1139 -2592 1174 -2584
rect 695 -2657 727 -2650
rect 695 -2677 702 -2657
rect 723 -2677 727 -2657
rect 695 -2742 727 -2677
rect 1065 -2742 1105 -2741
rect 695 -2744 1107 -2742
rect 695 -2770 1075 -2744
rect 1101 -2770 1107 -2744
rect 695 -2778 1107 -2770
rect 695 -2806 727 -2778
rect 695 -2826 700 -2806
rect 721 -2826 727 -2806
rect 695 -2833 727 -2826
rect 895 -2806 945 -2797
rect 1140 -2798 1174 -2592
rect 1708 -2572 1740 -2544
rect 1708 -2592 1713 -2572
rect 1734 -2592 1740 -2572
rect 1708 -2599 1740 -2592
rect 1915 -2571 1957 -2563
rect 2153 -2564 2187 -2358
rect 1915 -2591 1924 -2571
rect 1948 -2591 1957 -2571
rect 1915 -2603 1957 -2591
rect 2131 -2569 2187 -2564
rect 2131 -2589 2138 -2569
rect 2158 -2589 2187 -2569
rect 2131 -2596 2187 -2589
rect 2131 -2597 2166 -2596
rect 1917 -2632 1952 -2603
rect 1917 -2633 2227 -2632
rect 1802 -2639 1838 -2635
rect 1802 -2658 1810 -2639
rect 1830 -2658 1838 -2639
rect 1802 -2661 1838 -2658
rect 1803 -2689 1837 -2661
rect 1917 -2667 2244 -2633
rect 895 -2827 907 -2806
rect 929 -2827 945 -2806
rect 895 -2835 945 -2827
rect 1118 -2803 1174 -2798
rect 1118 -2823 1125 -2803
rect 1145 -2823 1174 -2803
rect 1118 -2830 1174 -2823
rect 1275 -2717 1838 -2689
rect 1118 -2831 1153 -2830
rect 900 -2868 941 -2835
rect 1275 -2868 1315 -2717
rect 900 -2897 1315 -2868
rect 2204 -2891 2244 -2667
rect 900 -2898 1309 -2897
rect 2204 -2911 2214 -2891
rect 2234 -2911 2244 -2891
rect 2204 -2921 2244 -2911
rect 1763 -2984 1795 -2977
rect 1763 -3004 1770 -2984
rect 1791 -3004 1795 -2984
rect 1763 -3069 1795 -3004
rect 2133 -3069 2173 -3068
rect 1763 -3071 2175 -3069
rect 1763 -3097 2143 -3071
rect 2169 -3097 2175 -3071
rect 1763 -3105 2175 -3097
rect 1148 -3125 1180 -3124
rect 1145 -3130 1180 -3125
rect 1145 -3150 1152 -3130
rect 1172 -3150 1180 -3130
rect 1145 -3158 1180 -3150
rect 701 -3223 733 -3216
rect 701 -3243 708 -3223
rect 729 -3243 733 -3223
rect 701 -3308 733 -3243
rect 1071 -3308 1111 -3307
rect 701 -3310 1113 -3308
rect 701 -3336 1081 -3310
rect 1107 -3336 1113 -3310
rect 701 -3344 1113 -3336
rect 701 -3372 733 -3344
rect 1146 -3364 1180 -3158
rect 1763 -3133 1795 -3105
rect 2208 -3125 2242 -2921
rect 1763 -3153 1768 -3133
rect 1789 -3153 1795 -3133
rect 1763 -3160 1795 -3153
rect 1974 -3133 2011 -3127
rect 1974 -3152 1980 -3133
rect 2003 -3152 2011 -3133
rect 1974 -3157 2011 -3152
rect 2186 -3130 2242 -3125
rect 2186 -3150 2193 -3130
rect 2213 -3150 2242 -3130
rect 2186 -3157 2242 -3150
rect 1982 -3194 2006 -3157
rect 2186 -3158 2221 -3157
rect 1982 -3196 2350 -3194
rect 1982 -3201 2355 -3196
rect 1982 -3219 2328 -3201
rect 2348 -3219 2355 -3201
rect 1982 -3224 2355 -3219
rect 2326 -3226 2355 -3224
rect 701 -3392 706 -3372
rect 727 -3392 733 -3372
rect 701 -3399 733 -3392
rect 910 -3370 950 -3365
rect 910 -3391 922 -3370
rect 944 -3391 950 -3370
rect 910 -3403 950 -3391
rect 1124 -3369 1180 -3364
rect 1124 -3389 1131 -3369
rect 1151 -3389 1180 -3369
rect 1124 -3396 1180 -3389
rect 1237 -3295 2194 -3276
rect 1124 -3397 1159 -3396
rect 916 -3435 944 -3403
rect 1237 -3435 1268 -3295
rect 2157 -3311 2192 -3295
rect 2157 -3331 2164 -3311
rect 2184 -3331 2192 -3311
rect 2157 -3339 2192 -3331
rect 916 -3466 1268 -3435
rect 1713 -3404 1745 -3397
rect 1713 -3424 1720 -3404
rect 1741 -3424 1745 -3404
rect 1713 -3489 1745 -3424
rect 2083 -3489 2123 -3488
rect 1713 -3491 2125 -3489
rect 1713 -3517 2093 -3491
rect 2119 -3517 2125 -3491
rect 1713 -3525 2125 -3517
rect 1147 -3540 1179 -3539
rect 1144 -3545 1179 -3540
rect 1144 -3565 1151 -3545
rect 1171 -3565 1179 -3545
rect 1144 -3573 1179 -3565
rect 700 -3638 732 -3631
rect 700 -3658 707 -3638
rect 728 -3658 732 -3638
rect 700 -3723 732 -3658
rect 1070 -3723 1110 -3722
rect 700 -3725 1112 -3723
rect 700 -3751 1080 -3725
rect 1106 -3751 1112 -3725
rect 700 -3759 1112 -3751
rect 700 -3787 732 -3759
rect 700 -3807 705 -3787
rect 726 -3807 732 -3787
rect 700 -3814 732 -3807
rect 900 -3787 950 -3778
rect 1145 -3779 1179 -3573
rect 1713 -3553 1745 -3525
rect 1713 -3573 1718 -3553
rect 1739 -3573 1745 -3553
rect 1918 -3551 1960 -3542
rect 2158 -3545 2192 -3339
rect 1918 -3565 1928 -3551
rect 1713 -3580 1745 -3573
rect 1917 -3571 1928 -3565
rect 1952 -3571 1960 -3551
rect 1917 -3582 1960 -3571
rect 2136 -3550 2192 -3545
rect 2136 -3570 2143 -3550
rect 2163 -3570 2192 -3550
rect 2136 -3577 2192 -3570
rect 2136 -3578 2171 -3577
rect 1917 -3612 1957 -3582
rect 1807 -3620 1843 -3616
rect 1807 -3639 1815 -3620
rect 1835 -3639 1843 -3620
rect 1807 -3642 1843 -3639
rect 1917 -3617 2264 -3612
rect 1808 -3670 1842 -3642
rect 1917 -3643 2236 -3617
rect 2255 -3643 2264 -3617
rect 1917 -3647 2264 -3643
rect 900 -3808 912 -3787
rect 934 -3808 950 -3787
rect 900 -3816 950 -3808
rect 1123 -3784 1179 -3779
rect 1123 -3804 1130 -3784
rect 1150 -3804 1179 -3784
rect 1123 -3811 1179 -3804
rect 1280 -3698 1843 -3670
rect 1123 -3812 1158 -3811
rect 905 -3849 946 -3816
rect 1280 -3849 1320 -3698
rect 905 -3878 1320 -3849
rect 905 -3879 1314 -3878
<< labels >>
rlabel locali 304 3712 333 3718 1 vdd
rlabel locali 517 3709 546 3715 1 vdd
rlabel locali 250 3524 272 3539 1 d0
rlabel nwell 671 3679 694 3682 1 vdd
rlabel locali 301 3413 330 3419 1 gnd
rlabel locali 514 3413 543 3419 1 gnd
rlabel space 611 3408 640 3417 1 gnd
rlabel locali 303 3297 332 3303 1 vdd
rlabel locali 516 3294 545 3300 1 vdd
rlabel locali 249 3109 271 3124 1 d0
rlabel nwell 670 3264 693 3267 1 vdd
rlabel locali 300 2998 329 3004 1 gnd
rlabel locali 513 2998 542 3004 1 gnd
rlabel space 610 2993 639 3002 1 gnd
rlabel locali 1316 3531 1345 3537 1 vdd
rlabel locali 1529 3528 1558 3534 1 vdd
rlabel nwell 1683 3498 1706 3501 1 vdd
rlabel locali 1313 3232 1342 3238 1 gnd
rlabel locali 1526 3232 1555 3238 1 gnd
rlabel space 1623 3227 1652 3236 1 gnd
rlabel locali 1254 3342 1301 3363 1 d1
rlabel locali 116 3904 141 3913 1 vref
rlabel locali 309 2731 338 2737 1 vdd
rlabel locali 522 2728 551 2734 1 vdd
rlabel locali 255 2543 277 2558 1 d0
rlabel nwell 676 2698 699 2701 1 vdd
rlabel locali 306 2432 335 2438 1 gnd
rlabel locali 519 2432 548 2438 1 gnd
rlabel space 616 2427 645 2436 1 gnd
rlabel locali 308 2316 337 2322 1 vdd
rlabel locali 521 2313 550 2319 1 vdd
rlabel locali 254 2128 276 2143 1 d0
rlabel nwell 675 2283 698 2286 1 vdd
rlabel locali 305 2017 334 2023 1 gnd
rlabel locali 518 2017 547 2023 1 gnd
rlabel locali 1321 2550 1350 2556 1 vdd
rlabel locali 1534 2547 1563 2553 1 vdd
rlabel nwell 1688 2517 1711 2520 1 vdd
rlabel locali 1318 2251 1347 2257 1 gnd
rlabel locali 1531 2251 1560 2257 1 gnd
rlabel space 1628 2246 1657 2255 1 gnd
rlabel locali 1259 2361 1306 2382 1 d1
rlabel locali 1371 2970 1400 2976 1 vdd
rlabel locali 1584 2967 1613 2973 1 vdd
rlabel nwell 1738 2937 1761 2940 1 vdd
rlabel locali 1368 2671 1397 2677 1 gnd
rlabel locali 1581 2671 1610 2677 1 gnd
rlabel space 1678 2666 1707 2675 1 gnd
rlabel locali 1314 2782 1337 2797 1 d2
rlabel space 615 2012 644 2021 1 gnd
rlabel locali 1326 822 1349 837 1 d2
rlabel space 1690 706 1719 715 1 gnd
rlabel locali 1593 711 1622 717 1 gnd
rlabel locali 1380 711 1409 717 1 gnd
rlabel nwell 1750 977 1773 980 1 vdd
rlabel locali 1596 1007 1625 1013 1 vdd
rlabel locali 1383 1010 1412 1016 1 vdd
rlabel locali 1271 401 1318 422 1 d1
rlabel space 1640 286 1669 295 1 gnd
rlabel locali 1543 291 1572 297 1 gnd
rlabel locali 1330 291 1359 297 1 gnd
rlabel nwell 1700 557 1723 560 1 vdd
rlabel locali 1546 587 1575 593 1 vdd
rlabel locali 1333 590 1362 596 1 vdd
rlabel space 627 52 656 61 1 gnd
rlabel locali 530 57 559 63 1 gnd
rlabel locali 317 57 346 63 1 gnd
rlabel nwell 687 323 710 326 1 vdd
rlabel locali 266 168 288 183 1 d0
rlabel locali 533 353 562 359 1 vdd
rlabel locali 320 356 349 362 1 vdd
rlabel space 628 467 657 476 1 gnd
rlabel locali 531 472 560 478 1 gnd
rlabel locali 318 472 347 478 1 gnd
rlabel nwell 688 738 711 741 1 vdd
rlabel locali 267 583 289 598 1 d0
rlabel locali 534 768 563 774 1 vdd
rlabel locali 321 771 350 777 1 vdd
rlabel locali 1266 1382 1313 1403 1 d1
rlabel space 1635 1267 1664 1276 1 gnd
rlabel locali 1538 1272 1567 1278 1 gnd
rlabel locali 1325 1272 1354 1278 1 gnd
rlabel nwell 1695 1538 1718 1541 1 vdd
rlabel locali 1541 1568 1570 1574 1 vdd
rlabel locali 1328 1571 1357 1577 1 vdd
rlabel space 622 1033 651 1042 1 gnd
rlabel locali 525 1038 554 1044 1 gnd
rlabel locali 312 1038 341 1044 1 gnd
rlabel nwell 682 1304 705 1307 1 vdd
rlabel locali 261 1149 283 1164 1 d0
rlabel locali 528 1334 557 1340 1 vdd
rlabel locali 315 1337 344 1343 1 vdd
rlabel space 623 1448 652 1457 1 gnd
rlabel locali 526 1453 555 1459 1 gnd
rlabel locali 313 1453 342 1459 1 gnd
rlabel nwell 683 1719 706 1722 1 vdd
rlabel locali 262 1564 284 1579 1 d0
rlabel locali 529 1749 558 1755 1 vdd
rlabel locali 316 1752 345 1758 1 vdd
rlabel locali 1536 2038 1565 2044 1 vdd
rlabel locali 1749 2035 1778 2041 1 vdd
rlabel nwell 1903 2005 1926 2008 1 vdd
rlabel locali 1533 1739 1562 1745 1 gnd
rlabel locali 1746 1739 1775 1745 1 gnd
rlabel space 1843 1734 1872 1743 1 gnd
rlabel locali 1474 1848 1506 1867 1 d3
rlabel locali 1494 -2069 1526 -2050 1 d3
rlabel space 1863 -2183 1892 -2174 1 gnd
rlabel locali 1766 -2178 1795 -2172 1 gnd
rlabel locali 1553 -2178 1582 -2172 1 gnd
rlabel nwell 1923 -1912 1946 -1909 1 vdd
rlabel locali 1769 -1882 1798 -1876 1 vdd
rlabel locali 1556 -1879 1585 -1873 1 vdd
rlabel locali 336 -2165 365 -2159 1 vdd
rlabel locali 549 -2168 578 -2162 1 vdd
rlabel locali 282 -2353 304 -2338 1 d0
rlabel nwell 703 -2198 726 -2195 1 vdd
rlabel locali 333 -2464 362 -2458 1 gnd
rlabel locali 546 -2464 575 -2458 1 gnd
rlabel space 643 -2469 672 -2460 1 gnd
rlabel locali 335 -2580 364 -2574 1 vdd
rlabel locali 548 -2583 577 -2577 1 vdd
rlabel locali 281 -2768 303 -2753 1 d0
rlabel nwell 702 -2613 725 -2610 1 vdd
rlabel locali 332 -2879 361 -2873 1 gnd
rlabel locali 545 -2879 574 -2873 1 gnd
rlabel space 642 -2884 671 -2875 1 gnd
rlabel locali 1348 -2346 1377 -2340 1 vdd
rlabel locali 1561 -2349 1590 -2343 1 vdd
rlabel nwell 1715 -2379 1738 -2376 1 vdd
rlabel locali 1345 -2645 1374 -2639 1 gnd
rlabel locali 1558 -2645 1587 -2639 1 gnd
rlabel space 1655 -2650 1684 -2641 1 gnd
rlabel locali 1286 -2535 1333 -2514 1 d1
rlabel locali 341 -3146 370 -3140 1 vdd
rlabel locali 554 -3149 583 -3143 1 vdd
rlabel locali 287 -3334 309 -3319 1 d0
rlabel nwell 708 -3179 731 -3176 1 vdd
rlabel locali 338 -3445 367 -3439 1 gnd
rlabel locali 551 -3445 580 -3439 1 gnd
rlabel space 648 -3450 677 -3441 1 gnd
rlabel locali 340 -3561 369 -3555 1 vdd
rlabel locali 553 -3564 582 -3558 1 vdd
rlabel locali 286 -3749 308 -3734 1 d0
rlabel nwell 707 -3594 730 -3591 1 vdd
rlabel locali 337 -3860 366 -3854 1 gnd
rlabel locali 550 -3860 579 -3854 1 gnd
rlabel space 647 -3865 676 -3856 1 gnd
rlabel locali 1353 -3327 1382 -3321 1 vdd
rlabel locali 1566 -3330 1595 -3324 1 vdd
rlabel nwell 1720 -3360 1743 -3357 1 vdd
rlabel locali 1350 -3626 1379 -3620 1 gnd
rlabel locali 1563 -3626 1592 -3620 1 gnd
rlabel space 1660 -3631 1689 -3622 1 gnd
rlabel locali 1291 -3516 1338 -3495 1 d1
rlabel locali 158 -3909 185 -3896 1 gnd
rlabel locali 1403 -2907 1432 -2901 1 vdd
rlabel locali 1616 -2910 1645 -2904 1 vdd
rlabel nwell 1770 -2940 1793 -2937 1 vdd
rlabel locali 1400 -3206 1429 -3200 1 gnd
rlabel locali 1613 -3206 1642 -3200 1 gnd
rlabel space 1710 -3211 1739 -3202 1 gnd
rlabel locali 1346 -3095 1369 -3080 1 d2
rlabel space 635 -1905 664 -1896 1 gnd
rlabel locali 1334 -1135 1357 -1120 1 d2
rlabel space 1698 -1251 1727 -1242 1 gnd
rlabel locali 1601 -1246 1630 -1240 1 gnd
rlabel locali 1388 -1246 1417 -1240 1 gnd
rlabel nwell 1758 -980 1781 -977 1 vdd
rlabel locali 1604 -950 1633 -944 1 vdd
rlabel locali 1391 -947 1420 -941 1 vdd
rlabel locali 1279 -1556 1326 -1535 1 d1
rlabel space 1648 -1671 1677 -1662 1 gnd
rlabel locali 1551 -1666 1580 -1660 1 gnd
rlabel locali 1338 -1666 1367 -1660 1 gnd
rlabel nwell 1708 -1400 1731 -1397 1 vdd
rlabel locali 1554 -1370 1583 -1364 1 vdd
rlabel locali 1341 -1367 1370 -1361 1 vdd
rlabel locali 538 -1900 567 -1894 1 gnd
rlabel locali 325 -1900 354 -1894 1 gnd
rlabel nwell 695 -1634 718 -1631 1 vdd
rlabel locali 274 -1789 296 -1774 1 d0
rlabel locali 541 -1604 570 -1598 1 vdd
rlabel locali 328 -1601 357 -1595 1 vdd
rlabel space 636 -1490 665 -1481 1 gnd
rlabel locali 539 -1485 568 -1479 1 gnd
rlabel locali 326 -1485 355 -1479 1 gnd
rlabel nwell 696 -1219 719 -1216 1 vdd
rlabel locali 275 -1374 297 -1359 1 d0
rlabel locali 542 -1189 571 -1183 1 vdd
rlabel locali 329 -1186 358 -1180 1 vdd
rlabel locali 1274 -575 1321 -554 1 d1
rlabel space 1643 -690 1672 -681 1 gnd
rlabel locali 1546 -685 1575 -679 1 gnd
rlabel locali 1333 -685 1362 -679 1 gnd
rlabel nwell 1703 -419 1726 -416 1 vdd
rlabel locali 1549 -389 1578 -383 1 vdd
rlabel locali 1336 -386 1365 -380 1 vdd
rlabel space 630 -924 659 -915 1 gnd
rlabel locali 533 -919 562 -913 1 gnd
rlabel locali 320 -919 349 -913 1 gnd
rlabel nwell 690 -653 713 -650 1 vdd
rlabel locali 269 -808 291 -793 1 d0
rlabel locali 536 -623 565 -617 1 vdd
rlabel locali 323 -620 352 -614 1 vdd
rlabel space 631 -509 660 -500 1 gnd
rlabel locali 534 -504 563 -498 1 gnd
rlabel locali 321 -504 350 -498 1 gnd
rlabel nwell 691 -238 714 -235 1 vdd
rlabel locali 270 -393 292 -378 1 d0
rlabel locali 537 -208 566 -202 1 vdd
rlabel locali 324 -205 353 -199 1 vdd
rlabel locali 1631 46 1660 52 1 vdd
rlabel locali 1844 43 1873 49 1 vdd
rlabel nwell 1998 13 2021 16 1 vdd
rlabel locali 1628 -253 1657 -247 1 gnd
rlabel locali 1841 -253 1870 -247 1 gnd
rlabel space 1938 -258 1967 -249 1 gnd
rlabel locali 2207 -107 2229 -92 1 vout
rlabel locali 1573 -148 1595 -124 1 d4
<< end >>
