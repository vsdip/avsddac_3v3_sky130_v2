magic
tech sky130A
timestamp 1616157560
<< nwell >>
rect 278 611 1089 761
rect 1290 430 2101 580
rect 277 196 1088 346
rect 1345 -131 2156 19
rect 283 -370 1094 -220
rect 1295 -551 2106 -401
rect 282 -785 1093 -635
<< nmos >>
rect 342 510 392 552
rect 555 510 605 552
rect 763 510 813 552
rect 971 510 1021 552
rect 1354 329 1404 371
rect 1567 329 1617 371
rect 1775 329 1825 371
rect 1983 329 2033 371
rect 341 95 391 137
rect 554 95 604 137
rect 762 95 812 137
rect 970 95 1020 137
rect 1409 -232 1459 -190
rect 1622 -232 1672 -190
rect 1830 -232 1880 -190
rect 2038 -232 2088 -190
rect 347 -471 397 -429
rect 560 -471 610 -429
rect 768 -471 818 -429
rect 976 -471 1026 -429
rect 1359 -652 1409 -610
rect 1572 -652 1622 -610
rect 1780 -652 1830 -610
rect 1988 -652 2038 -610
rect 346 -886 396 -844
rect 559 -886 609 -844
rect 767 -886 817 -844
rect 975 -886 1025 -844
<< pmos >>
rect 342 629 392 729
rect 555 629 605 729
rect 763 629 813 729
rect 971 629 1021 729
rect 1354 448 1404 548
rect 1567 448 1617 548
rect 1775 448 1825 548
rect 1983 448 2033 548
rect 341 214 391 314
rect 554 214 604 314
rect 762 214 812 314
rect 970 214 1020 314
rect 1409 -113 1459 -13
rect 1622 -113 1672 -13
rect 1830 -113 1880 -13
rect 2038 -113 2088 -13
rect 347 -352 397 -252
rect 560 -352 610 -252
rect 768 -352 818 -252
rect 976 -352 1026 -252
rect 1359 -533 1409 -433
rect 1572 -533 1622 -433
rect 1780 -533 1830 -433
rect 1988 -533 2038 -433
rect 346 -767 396 -667
rect 559 -767 609 -667
rect 767 -767 817 -667
rect 975 -767 1025 -667
<< ndiff >>
rect 293 542 342 552
rect 293 522 304 542
rect 324 522 342 542
rect 293 510 342 522
rect 392 546 436 552
rect 392 526 407 546
rect 427 526 436 546
rect 392 510 436 526
rect 506 542 555 552
rect 506 522 517 542
rect 537 522 555 542
rect 506 510 555 522
rect 605 546 649 552
rect 605 526 620 546
rect 640 526 649 546
rect 605 510 649 526
rect 714 542 763 552
rect 714 522 725 542
rect 745 522 763 542
rect 714 510 763 522
rect 813 546 857 552
rect 813 526 828 546
rect 848 526 857 546
rect 813 510 857 526
rect 927 546 971 552
rect 927 526 936 546
rect 956 526 971 546
rect 927 510 971 526
rect 1021 542 1070 552
rect 1021 522 1039 542
rect 1059 522 1070 542
rect 1021 510 1070 522
rect 1305 361 1354 371
rect 1305 341 1316 361
rect 1336 341 1354 361
rect 1305 329 1354 341
rect 1404 365 1448 371
rect 1404 345 1419 365
rect 1439 345 1448 365
rect 1404 329 1448 345
rect 1518 361 1567 371
rect 1518 341 1529 361
rect 1549 341 1567 361
rect 1518 329 1567 341
rect 1617 365 1661 371
rect 1617 345 1632 365
rect 1652 345 1661 365
rect 1617 329 1661 345
rect 1726 361 1775 371
rect 1726 341 1737 361
rect 1757 341 1775 361
rect 1726 329 1775 341
rect 1825 365 1869 371
rect 1825 345 1840 365
rect 1860 345 1869 365
rect 1825 329 1869 345
rect 1939 365 1983 371
rect 1939 345 1948 365
rect 1968 345 1983 365
rect 1939 329 1983 345
rect 2033 361 2082 371
rect 2033 341 2051 361
rect 2071 341 2082 361
rect 2033 329 2082 341
rect 292 127 341 137
rect 292 107 303 127
rect 323 107 341 127
rect 292 95 341 107
rect 391 131 435 137
rect 391 111 406 131
rect 426 111 435 131
rect 391 95 435 111
rect 505 127 554 137
rect 505 107 516 127
rect 536 107 554 127
rect 505 95 554 107
rect 604 131 648 137
rect 604 111 619 131
rect 639 111 648 131
rect 604 95 648 111
rect 713 127 762 137
rect 713 107 724 127
rect 744 107 762 127
rect 713 95 762 107
rect 812 131 856 137
rect 812 111 827 131
rect 847 111 856 131
rect 812 95 856 111
rect 926 131 970 137
rect 926 111 935 131
rect 955 111 970 131
rect 926 95 970 111
rect 1020 127 1069 137
rect 1020 107 1038 127
rect 1058 107 1069 127
rect 1020 95 1069 107
rect 1360 -200 1409 -190
rect 1360 -220 1371 -200
rect 1391 -220 1409 -200
rect 1360 -232 1409 -220
rect 1459 -196 1503 -190
rect 1459 -216 1474 -196
rect 1494 -216 1503 -196
rect 1459 -232 1503 -216
rect 1573 -200 1622 -190
rect 1573 -220 1584 -200
rect 1604 -220 1622 -200
rect 1573 -232 1622 -220
rect 1672 -196 1716 -190
rect 1672 -216 1687 -196
rect 1707 -216 1716 -196
rect 1672 -232 1716 -216
rect 1781 -200 1830 -190
rect 1781 -220 1792 -200
rect 1812 -220 1830 -200
rect 1781 -232 1830 -220
rect 1880 -196 1924 -190
rect 1880 -216 1895 -196
rect 1915 -216 1924 -196
rect 1880 -232 1924 -216
rect 1994 -196 2038 -190
rect 1994 -216 2003 -196
rect 2023 -216 2038 -196
rect 1994 -232 2038 -216
rect 2088 -200 2137 -190
rect 2088 -220 2106 -200
rect 2126 -220 2137 -200
rect 2088 -232 2137 -220
rect 298 -439 347 -429
rect 298 -459 309 -439
rect 329 -459 347 -439
rect 298 -471 347 -459
rect 397 -435 441 -429
rect 397 -455 412 -435
rect 432 -455 441 -435
rect 397 -471 441 -455
rect 511 -439 560 -429
rect 511 -459 522 -439
rect 542 -459 560 -439
rect 511 -471 560 -459
rect 610 -435 654 -429
rect 610 -455 625 -435
rect 645 -455 654 -435
rect 610 -471 654 -455
rect 719 -439 768 -429
rect 719 -459 730 -439
rect 750 -459 768 -439
rect 719 -471 768 -459
rect 818 -435 862 -429
rect 818 -455 833 -435
rect 853 -455 862 -435
rect 818 -471 862 -455
rect 932 -435 976 -429
rect 932 -455 941 -435
rect 961 -455 976 -435
rect 932 -471 976 -455
rect 1026 -439 1075 -429
rect 1026 -459 1044 -439
rect 1064 -459 1075 -439
rect 1026 -471 1075 -459
rect 1310 -620 1359 -610
rect 1310 -640 1321 -620
rect 1341 -640 1359 -620
rect 1310 -652 1359 -640
rect 1409 -616 1453 -610
rect 1409 -636 1424 -616
rect 1444 -636 1453 -616
rect 1409 -652 1453 -636
rect 1523 -620 1572 -610
rect 1523 -640 1534 -620
rect 1554 -640 1572 -620
rect 1523 -652 1572 -640
rect 1622 -616 1666 -610
rect 1622 -636 1637 -616
rect 1657 -636 1666 -616
rect 1622 -652 1666 -636
rect 1731 -620 1780 -610
rect 1731 -640 1742 -620
rect 1762 -640 1780 -620
rect 1731 -652 1780 -640
rect 1830 -616 1874 -610
rect 1830 -636 1845 -616
rect 1865 -636 1874 -616
rect 1830 -652 1874 -636
rect 1944 -616 1988 -610
rect 1944 -636 1953 -616
rect 1973 -636 1988 -616
rect 1944 -652 1988 -636
rect 2038 -620 2087 -610
rect 2038 -640 2056 -620
rect 2076 -640 2087 -620
rect 2038 -652 2087 -640
rect 297 -854 346 -844
rect 297 -874 308 -854
rect 328 -874 346 -854
rect 297 -886 346 -874
rect 396 -850 440 -844
rect 396 -870 411 -850
rect 431 -870 440 -850
rect 396 -886 440 -870
rect 510 -854 559 -844
rect 510 -874 521 -854
rect 541 -874 559 -854
rect 510 -886 559 -874
rect 609 -850 653 -844
rect 609 -870 624 -850
rect 644 -870 653 -850
rect 609 -886 653 -870
rect 718 -854 767 -844
rect 718 -874 729 -854
rect 749 -874 767 -854
rect 718 -886 767 -874
rect 817 -850 861 -844
rect 817 -870 832 -850
rect 852 -870 861 -850
rect 817 -886 861 -870
rect 931 -850 975 -844
rect 931 -870 940 -850
rect 960 -870 975 -850
rect 931 -886 975 -870
rect 1025 -854 1074 -844
rect 1025 -874 1043 -854
rect 1063 -874 1074 -854
rect 1025 -886 1074 -874
<< pdiff >>
rect 298 691 342 729
rect 298 671 310 691
rect 330 671 342 691
rect 298 629 342 671
rect 392 691 434 729
rect 392 671 406 691
rect 426 671 434 691
rect 392 629 434 671
rect 511 691 555 729
rect 511 671 523 691
rect 543 671 555 691
rect 511 629 555 671
rect 605 691 647 729
rect 605 671 619 691
rect 639 671 647 691
rect 605 629 647 671
rect 719 691 763 729
rect 719 671 731 691
rect 751 671 763 691
rect 719 629 763 671
rect 813 691 855 729
rect 813 671 827 691
rect 847 671 855 691
rect 813 629 855 671
rect 929 691 971 729
rect 929 671 937 691
rect 957 671 971 691
rect 929 629 971 671
rect 1021 698 1066 729
rect 1021 691 1065 698
rect 1021 671 1033 691
rect 1053 671 1065 691
rect 1021 629 1065 671
rect 1310 510 1354 548
rect 1310 490 1322 510
rect 1342 490 1354 510
rect 1310 448 1354 490
rect 1404 510 1446 548
rect 1404 490 1418 510
rect 1438 490 1446 510
rect 1404 448 1446 490
rect 1523 510 1567 548
rect 1523 490 1535 510
rect 1555 490 1567 510
rect 1523 448 1567 490
rect 1617 510 1659 548
rect 1617 490 1631 510
rect 1651 490 1659 510
rect 1617 448 1659 490
rect 1731 510 1775 548
rect 1731 490 1743 510
rect 1763 490 1775 510
rect 1731 448 1775 490
rect 1825 510 1867 548
rect 1825 490 1839 510
rect 1859 490 1867 510
rect 1825 448 1867 490
rect 1941 510 1983 548
rect 1941 490 1949 510
rect 1969 490 1983 510
rect 1941 448 1983 490
rect 2033 517 2078 548
rect 2033 510 2077 517
rect 2033 490 2045 510
rect 2065 490 2077 510
rect 2033 448 2077 490
rect 297 276 341 314
rect 297 256 309 276
rect 329 256 341 276
rect 297 214 341 256
rect 391 276 433 314
rect 391 256 405 276
rect 425 256 433 276
rect 391 214 433 256
rect 510 276 554 314
rect 510 256 522 276
rect 542 256 554 276
rect 510 214 554 256
rect 604 276 646 314
rect 604 256 618 276
rect 638 256 646 276
rect 604 214 646 256
rect 718 276 762 314
rect 718 256 730 276
rect 750 256 762 276
rect 718 214 762 256
rect 812 276 854 314
rect 812 256 826 276
rect 846 256 854 276
rect 812 214 854 256
rect 928 276 970 314
rect 928 256 936 276
rect 956 256 970 276
rect 928 214 970 256
rect 1020 283 1065 314
rect 1020 276 1064 283
rect 1020 256 1032 276
rect 1052 256 1064 276
rect 1020 214 1064 256
rect 1365 -51 1409 -13
rect 1365 -71 1377 -51
rect 1397 -71 1409 -51
rect 1365 -113 1409 -71
rect 1459 -51 1501 -13
rect 1459 -71 1473 -51
rect 1493 -71 1501 -51
rect 1459 -113 1501 -71
rect 1578 -51 1622 -13
rect 1578 -71 1590 -51
rect 1610 -71 1622 -51
rect 1578 -113 1622 -71
rect 1672 -51 1714 -13
rect 1672 -71 1686 -51
rect 1706 -71 1714 -51
rect 1672 -113 1714 -71
rect 1786 -51 1830 -13
rect 1786 -71 1798 -51
rect 1818 -71 1830 -51
rect 1786 -113 1830 -71
rect 1880 -51 1922 -13
rect 1880 -71 1894 -51
rect 1914 -71 1922 -51
rect 1880 -113 1922 -71
rect 1996 -51 2038 -13
rect 1996 -71 2004 -51
rect 2024 -71 2038 -51
rect 1996 -113 2038 -71
rect 2088 -44 2133 -13
rect 2088 -51 2132 -44
rect 2088 -71 2100 -51
rect 2120 -71 2132 -51
rect 2088 -113 2132 -71
rect 303 -290 347 -252
rect 303 -310 315 -290
rect 335 -310 347 -290
rect 303 -352 347 -310
rect 397 -290 439 -252
rect 397 -310 411 -290
rect 431 -310 439 -290
rect 397 -352 439 -310
rect 516 -290 560 -252
rect 516 -310 528 -290
rect 548 -310 560 -290
rect 516 -352 560 -310
rect 610 -290 652 -252
rect 610 -310 624 -290
rect 644 -310 652 -290
rect 610 -352 652 -310
rect 724 -290 768 -252
rect 724 -310 736 -290
rect 756 -310 768 -290
rect 724 -352 768 -310
rect 818 -290 860 -252
rect 818 -310 832 -290
rect 852 -310 860 -290
rect 818 -352 860 -310
rect 934 -290 976 -252
rect 934 -310 942 -290
rect 962 -310 976 -290
rect 934 -352 976 -310
rect 1026 -283 1071 -252
rect 1026 -290 1070 -283
rect 1026 -310 1038 -290
rect 1058 -310 1070 -290
rect 1026 -352 1070 -310
rect 1315 -471 1359 -433
rect 1315 -491 1327 -471
rect 1347 -491 1359 -471
rect 1315 -533 1359 -491
rect 1409 -471 1451 -433
rect 1409 -491 1423 -471
rect 1443 -491 1451 -471
rect 1409 -533 1451 -491
rect 1528 -471 1572 -433
rect 1528 -491 1540 -471
rect 1560 -491 1572 -471
rect 1528 -533 1572 -491
rect 1622 -471 1664 -433
rect 1622 -491 1636 -471
rect 1656 -491 1664 -471
rect 1622 -533 1664 -491
rect 1736 -471 1780 -433
rect 1736 -491 1748 -471
rect 1768 -491 1780 -471
rect 1736 -533 1780 -491
rect 1830 -471 1872 -433
rect 1830 -491 1844 -471
rect 1864 -491 1872 -471
rect 1830 -533 1872 -491
rect 1946 -471 1988 -433
rect 1946 -491 1954 -471
rect 1974 -491 1988 -471
rect 1946 -533 1988 -491
rect 2038 -464 2083 -433
rect 2038 -471 2082 -464
rect 2038 -491 2050 -471
rect 2070 -491 2082 -471
rect 2038 -533 2082 -491
rect 302 -705 346 -667
rect 302 -725 314 -705
rect 334 -725 346 -705
rect 302 -767 346 -725
rect 396 -705 438 -667
rect 396 -725 410 -705
rect 430 -725 438 -705
rect 396 -767 438 -725
rect 515 -705 559 -667
rect 515 -725 527 -705
rect 547 -725 559 -705
rect 515 -767 559 -725
rect 609 -705 651 -667
rect 609 -725 623 -705
rect 643 -725 651 -705
rect 609 -767 651 -725
rect 723 -705 767 -667
rect 723 -725 735 -705
rect 755 -725 767 -705
rect 723 -767 767 -725
rect 817 -705 859 -667
rect 817 -725 831 -705
rect 851 -725 859 -705
rect 817 -767 859 -725
rect 933 -705 975 -667
rect 933 -725 941 -705
rect 961 -725 975 -705
rect 933 -767 975 -725
rect 1025 -698 1070 -667
rect 1025 -705 1069 -698
rect 1025 -725 1037 -705
rect 1057 -725 1069 -705
rect 1025 -767 1069 -725
<< ndiffc >>
rect 118 906 136 924
rect 120 807 138 825
rect 116 692 134 710
rect 118 593 136 611
rect 304 522 324 542
rect 407 526 427 546
rect 517 522 537 542
rect 620 526 640 546
rect 725 522 745 542
rect 828 526 848 546
rect 936 526 956 546
rect 1039 522 1059 542
rect 116 410 134 428
rect 1316 341 1336 361
rect 1419 345 1439 365
rect 1529 341 1549 361
rect 1632 345 1652 365
rect 1737 341 1757 361
rect 1840 345 1860 365
rect 1948 345 1968 365
rect 2051 341 2071 361
rect 118 311 136 329
rect 123 209 141 227
rect 125 110 143 128
rect 303 107 323 127
rect 406 111 426 131
rect 516 107 536 127
rect 619 111 639 131
rect 724 107 744 127
rect 827 111 847 131
rect 935 111 955 131
rect 1038 107 1058 127
rect 123 -75 141 -57
rect 125 -174 143 -156
rect 1371 -220 1391 -200
rect 1474 -216 1494 -196
rect 1584 -220 1604 -200
rect 1687 -216 1707 -196
rect 1792 -220 1812 -200
rect 1895 -216 1915 -196
rect 2003 -216 2023 -196
rect 2106 -220 2126 -200
rect 121 -289 139 -271
rect 123 -388 141 -370
rect 309 -459 329 -439
rect 412 -455 432 -435
rect 522 -459 542 -439
rect 625 -455 645 -435
rect 730 -459 750 -439
rect 833 -455 853 -435
rect 941 -455 961 -435
rect 1044 -459 1064 -439
rect 121 -571 139 -553
rect 1321 -640 1341 -620
rect 1424 -636 1444 -616
rect 1534 -640 1554 -620
rect 1637 -636 1657 -616
rect 1742 -640 1762 -620
rect 1845 -636 1865 -616
rect 1953 -636 1973 -616
rect 2056 -640 2076 -620
rect 123 -670 141 -652
rect 128 -772 146 -754
rect 130 -871 148 -853
rect 308 -874 328 -854
rect 411 -870 431 -850
rect 521 -874 541 -854
rect 624 -870 644 -850
rect 729 -874 749 -854
rect 832 -870 852 -850
rect 940 -870 960 -850
rect 1043 -874 1063 -854
<< pdiffc >>
rect 310 671 330 691
rect 406 671 426 691
rect 523 671 543 691
rect 619 671 639 691
rect 731 671 751 691
rect 827 671 847 691
rect 937 671 957 691
rect 1033 671 1053 691
rect 1322 490 1342 510
rect 1418 490 1438 510
rect 1535 490 1555 510
rect 1631 490 1651 510
rect 1743 490 1763 510
rect 1839 490 1859 510
rect 1949 490 1969 510
rect 2045 490 2065 510
rect 309 256 329 276
rect 405 256 425 276
rect 522 256 542 276
rect 618 256 638 276
rect 730 256 750 276
rect 826 256 846 276
rect 936 256 956 276
rect 1032 256 1052 276
rect 1377 -71 1397 -51
rect 1473 -71 1493 -51
rect 1590 -71 1610 -51
rect 1686 -71 1706 -51
rect 1798 -71 1818 -51
rect 1894 -71 1914 -51
rect 2004 -71 2024 -51
rect 2100 -71 2120 -51
rect 315 -310 335 -290
rect 411 -310 431 -290
rect 528 -310 548 -290
rect 624 -310 644 -290
rect 736 -310 756 -290
rect 832 -310 852 -290
rect 942 -310 962 -290
rect 1038 -310 1058 -290
rect 1327 -491 1347 -471
rect 1423 -491 1443 -471
rect 1540 -491 1560 -471
rect 1636 -491 1656 -471
rect 1748 -491 1768 -471
rect 1844 -491 1864 -471
rect 1954 -491 1974 -471
rect 2050 -491 2070 -471
rect 314 -725 334 -705
rect 410 -725 430 -705
rect 527 -725 547 -705
rect 623 -725 643 -705
rect 735 -725 755 -705
rect 831 -725 851 -705
rect 941 -725 961 -705
rect 1037 -725 1057 -705
<< poly >>
rect 342 729 392 742
rect 555 729 605 742
rect 763 729 813 742
rect 971 729 1021 742
rect 342 601 392 629
rect 342 581 355 601
rect 375 581 392 601
rect 342 552 392 581
rect 555 600 605 629
rect 555 576 566 600
rect 590 576 605 600
rect 555 552 605 576
rect 763 605 813 629
rect 763 581 775 605
rect 799 581 813 605
rect 763 552 813 581
rect 971 603 1021 629
rect 971 577 989 603
rect 1015 577 1021 603
rect 971 552 1021 577
rect 1354 548 1404 561
rect 1567 548 1617 561
rect 1775 548 1825 561
rect 1983 548 2033 561
rect 342 494 392 510
rect 555 494 605 510
rect 763 494 813 510
rect 971 494 1021 510
rect 1354 420 1404 448
rect 1354 400 1367 420
rect 1387 400 1404 420
rect 1354 371 1404 400
rect 1567 419 1617 448
rect 1567 395 1578 419
rect 1602 395 1617 419
rect 1567 371 1617 395
rect 1775 424 1825 448
rect 1775 400 1787 424
rect 1811 400 1825 424
rect 1775 371 1825 400
rect 1983 422 2033 448
rect 1983 396 2001 422
rect 2027 396 2033 422
rect 1983 371 2033 396
rect 341 314 391 327
rect 554 314 604 327
rect 762 314 812 327
rect 970 314 1020 327
rect 1354 313 1404 329
rect 1567 313 1617 329
rect 1775 313 1825 329
rect 1983 313 2033 329
rect 341 186 391 214
rect 341 166 354 186
rect 374 166 391 186
rect 341 137 391 166
rect 554 185 604 214
rect 554 161 565 185
rect 589 161 604 185
rect 554 137 604 161
rect 762 190 812 214
rect 762 166 774 190
rect 798 166 812 190
rect 762 137 812 166
rect 970 188 1020 214
rect 970 162 988 188
rect 1014 162 1020 188
rect 970 137 1020 162
rect 341 79 391 95
rect 554 79 604 95
rect 762 79 812 95
rect 970 79 1020 95
rect 1409 -13 1459 0
rect 1622 -13 1672 0
rect 1830 -13 1880 0
rect 2038 -13 2088 0
rect 1409 -141 1459 -113
rect 1409 -161 1422 -141
rect 1442 -161 1459 -141
rect 1409 -190 1459 -161
rect 1622 -142 1672 -113
rect 1622 -166 1633 -142
rect 1657 -166 1672 -142
rect 1622 -190 1672 -166
rect 1830 -137 1880 -113
rect 1830 -161 1842 -137
rect 1866 -161 1880 -137
rect 1830 -190 1880 -161
rect 2038 -139 2088 -113
rect 2038 -165 2056 -139
rect 2082 -165 2088 -139
rect 2038 -190 2088 -165
rect 347 -252 397 -239
rect 560 -252 610 -239
rect 768 -252 818 -239
rect 976 -252 1026 -239
rect 1409 -248 1459 -232
rect 1622 -248 1672 -232
rect 1830 -248 1880 -232
rect 2038 -248 2088 -232
rect 347 -380 397 -352
rect 347 -400 360 -380
rect 380 -400 397 -380
rect 347 -429 397 -400
rect 560 -381 610 -352
rect 560 -405 571 -381
rect 595 -405 610 -381
rect 560 -429 610 -405
rect 768 -376 818 -352
rect 768 -400 780 -376
rect 804 -400 818 -376
rect 768 -429 818 -400
rect 976 -378 1026 -352
rect 976 -404 994 -378
rect 1020 -404 1026 -378
rect 976 -429 1026 -404
rect 1359 -433 1409 -420
rect 1572 -433 1622 -420
rect 1780 -433 1830 -420
rect 1988 -433 2038 -420
rect 347 -487 397 -471
rect 560 -487 610 -471
rect 768 -487 818 -471
rect 976 -487 1026 -471
rect 1359 -561 1409 -533
rect 1359 -581 1372 -561
rect 1392 -581 1409 -561
rect 1359 -610 1409 -581
rect 1572 -562 1622 -533
rect 1572 -586 1583 -562
rect 1607 -586 1622 -562
rect 1572 -610 1622 -586
rect 1780 -557 1830 -533
rect 1780 -581 1792 -557
rect 1816 -581 1830 -557
rect 1780 -610 1830 -581
rect 1988 -559 2038 -533
rect 1988 -585 2006 -559
rect 2032 -585 2038 -559
rect 1988 -610 2038 -585
rect 346 -667 396 -654
rect 559 -667 609 -654
rect 767 -667 817 -654
rect 975 -667 1025 -654
rect 1359 -668 1409 -652
rect 1572 -668 1622 -652
rect 1780 -668 1830 -652
rect 1988 -668 2038 -652
rect 346 -795 396 -767
rect 346 -815 359 -795
rect 379 -815 396 -795
rect 346 -844 396 -815
rect 559 -796 609 -767
rect 559 -820 570 -796
rect 594 -820 609 -796
rect 559 -844 609 -820
rect 767 -791 817 -767
rect 767 -815 779 -791
rect 803 -815 817 -791
rect 767 -844 817 -815
rect 975 -793 1025 -767
rect 975 -819 993 -793
rect 1019 -819 1025 -793
rect 975 -844 1025 -819
rect 346 -902 396 -886
rect 559 -902 609 -886
rect 767 -902 817 -886
rect 975 -902 1025 -886
<< polycont >>
rect 355 581 375 601
rect 566 576 590 600
rect 775 581 799 605
rect 989 577 1015 603
rect 1367 400 1387 420
rect 1578 395 1602 419
rect 1787 400 1811 424
rect 2001 396 2027 422
rect 354 166 374 186
rect 565 161 589 185
rect 774 166 798 190
rect 988 162 1014 188
rect 1422 -161 1442 -141
rect 1633 -166 1657 -142
rect 1842 -161 1866 -137
rect 2056 -165 2082 -139
rect 360 -400 380 -380
rect 571 -405 595 -381
rect 780 -400 804 -376
rect 994 -404 1020 -378
rect 1372 -581 1392 -561
rect 1583 -586 1607 -562
rect 1792 -581 1816 -557
rect 2006 -585 2032 -559
rect 359 -815 379 -795
rect 570 -820 594 -796
rect 779 -815 803 -791
rect 993 -819 1019 -793
<< ndiffres >>
rect 97 924 154 943
rect 97 921 118 924
rect 3 906 118 921
rect 136 906 154 924
rect 3 883 154 906
rect 3 847 45 883
rect 2 846 102 847
rect 2 825 158 846
rect 2 807 120 825
rect 138 807 158 825
rect 2 803 158 807
rect 97 787 158 803
rect 95 710 152 729
rect 95 707 116 710
rect 1 692 116 707
rect 134 692 152 710
rect 1 669 152 692
rect 1 633 43 669
rect 0 632 100 633
rect 0 611 156 632
rect 0 593 118 611
rect 136 593 156 611
rect 0 589 156 593
rect 95 573 156 589
rect 95 428 152 447
rect 95 425 116 428
rect 1 410 116 425
rect 134 410 152 428
rect 1 387 152 410
rect 1 351 43 387
rect 0 350 100 351
rect 0 329 156 350
rect 0 311 118 329
rect 136 311 156 329
rect 0 307 156 311
rect 95 291 156 307
rect 102 227 159 246
rect 102 224 123 227
rect 8 209 123 224
rect 141 209 159 227
rect 8 186 159 209
rect 8 150 50 186
rect 7 149 107 150
rect 7 128 163 149
rect 7 110 125 128
rect 143 110 163 128
rect 7 106 163 110
rect 102 90 163 106
rect 102 -57 159 -38
rect 102 -60 123 -57
rect 8 -75 123 -60
rect 141 -75 159 -57
rect 8 -98 159 -75
rect 8 -134 50 -98
rect 7 -135 107 -134
rect 7 -156 163 -135
rect 7 -174 125 -156
rect 143 -174 163 -156
rect 7 -178 163 -174
rect 102 -194 163 -178
rect 100 -271 157 -252
rect 100 -274 121 -271
rect 6 -289 121 -274
rect 139 -289 157 -271
rect 6 -312 157 -289
rect 6 -348 48 -312
rect 5 -349 105 -348
rect 5 -370 161 -349
rect 5 -388 123 -370
rect 141 -388 161 -370
rect 5 -392 161 -388
rect 100 -408 161 -392
rect 100 -553 157 -534
rect 100 -556 121 -553
rect 6 -571 121 -556
rect 139 -571 157 -553
rect 6 -594 157 -571
rect 6 -630 48 -594
rect 5 -631 105 -630
rect 5 -652 161 -631
rect 5 -670 123 -652
rect 141 -670 161 -652
rect 5 -674 161 -670
rect 100 -690 161 -674
rect 107 -754 164 -735
rect 107 -757 128 -754
rect 13 -772 128 -757
rect 146 -772 164 -754
rect 13 -795 164 -772
rect 13 -831 55 -795
rect 12 -832 112 -831
rect 12 -853 168 -832
rect 12 -871 130 -853
rect 148 -871 168 -853
rect 12 -875 168 -871
rect 107 -891 168 -875
<< locali >>
rect 110 933 145 981
rect 108 924 145 933
rect 108 906 118 924
rect 136 906 145 924
rect 108 896 145 906
rect 111 832 148 834
rect 111 831 759 832
rect 110 825 759 831
rect 110 807 120 825
rect 138 811 759 825
rect 138 807 148 811
rect 589 810 759 811
rect 110 797 148 807
rect 110 719 145 797
rect 722 787 759 810
rect 106 710 145 719
rect 106 692 116 710
rect 134 692 145 710
rect 106 686 145 692
rect 301 762 551 786
rect 301 691 338 762
rect 453 701 484 702
rect 106 682 143 686
rect 301 671 310 691
rect 330 671 338 691
rect 301 661 338 671
rect 397 691 484 701
rect 397 671 406 691
rect 426 671 484 691
rect 397 662 484 671
rect 397 661 434 662
rect 109 611 146 620
rect 107 593 118 611
rect 136 593 146 611
rect 453 609 484 662
rect 514 691 551 762
rect 722 767 1115 787
rect 1135 767 1138 787
rect 722 762 1138 767
rect 722 761 1063 762
rect 666 701 697 702
rect 514 671 523 691
rect 543 671 551 691
rect 514 661 551 671
rect 610 694 697 701
rect 610 691 671 694
rect 610 671 619 691
rect 639 674 671 691
rect 692 674 697 694
rect 639 671 697 674
rect 610 664 697 671
rect 722 691 759 761
rect 1025 760 1062 761
rect 874 701 910 702
rect 722 671 731 691
rect 751 671 759 691
rect 610 662 666 664
rect 610 661 647 662
rect 722 661 759 671
rect 818 691 966 701
rect 1066 698 1162 700
rect 818 671 827 691
rect 847 671 937 691
rect 957 671 966 691
rect 818 662 966 671
rect 1024 691 1162 698
rect 1024 671 1033 691
rect 1053 671 1162 691
rect 1024 662 1162 671
rect 818 661 855 662
rect 874 610 910 662
rect 929 661 966 662
rect 1025 661 1062 662
rect 345 608 386 609
rect 107 444 146 593
rect 237 601 386 608
rect 237 581 355 601
rect 375 581 386 601
rect 237 573 386 581
rect 453 605 812 609
rect 453 600 775 605
rect 453 576 566 600
rect 590 581 775 600
rect 799 581 812 605
rect 590 576 812 581
rect 453 573 812 576
rect 874 573 909 610
rect 977 607 1077 610
rect 977 603 1044 607
rect 977 577 989 603
rect 1015 581 1044 603
rect 1070 581 1077 607
rect 1015 577 1077 581
rect 977 573 1077 577
rect 453 552 484 573
rect 874 552 910 573
rect 296 551 333 552
rect 295 542 333 551
rect 295 522 304 542
rect 324 522 333 542
rect 295 514 333 522
rect 399 546 484 552
rect 509 551 546 552
rect 399 526 407 546
rect 427 526 484 546
rect 399 518 484 526
rect 508 542 546 551
rect 508 522 517 542
rect 537 522 546 542
rect 399 517 435 518
rect 508 514 546 522
rect 612 546 697 552
rect 717 551 754 552
rect 612 526 620 546
rect 640 545 697 546
rect 640 526 669 545
rect 612 525 669 526
rect 690 525 697 545
rect 612 518 697 525
rect 716 542 754 551
rect 716 522 725 542
rect 745 522 754 542
rect 612 517 648 518
rect 716 514 754 522
rect 820 547 964 552
rect 820 546 885 547
rect 820 526 828 546
rect 848 526 885 546
rect 907 546 964 547
rect 907 526 936 546
rect 956 526 964 546
rect 820 518 964 526
rect 820 517 856 518
rect 928 517 964 518
rect 1030 551 1067 552
rect 1030 550 1068 551
rect 1030 542 1094 550
rect 1030 522 1039 542
rect 1059 528 1094 542
rect 1114 528 1117 548
rect 1059 523 1117 528
rect 1059 522 1094 523
rect 296 485 333 514
rect 297 483 333 485
rect 509 483 546 514
rect 297 461 546 483
rect 717 482 754 514
rect 1030 510 1094 522
rect 1134 484 1161 662
rect 993 482 1161 484
rect 717 456 1161 482
rect 1313 581 1563 605
rect 1313 510 1350 581
rect 1465 520 1496 521
rect 1313 490 1322 510
rect 1342 490 1350 510
rect 1313 480 1350 490
rect 1409 510 1496 520
rect 1409 490 1418 510
rect 1438 490 1496 510
rect 1409 481 1496 490
rect 1409 480 1446 481
rect 717 446 739 456
rect 993 455 1161 456
rect 677 444 739 446
rect 107 437 739 444
rect 106 428 739 437
rect 1465 428 1496 481
rect 1526 510 1563 581
rect 1734 586 2127 606
rect 2147 586 2150 606
rect 1734 581 2150 586
rect 1734 580 2075 581
rect 1678 520 1709 521
rect 1526 490 1535 510
rect 1555 490 1563 510
rect 1526 480 1563 490
rect 1622 513 1709 520
rect 1622 510 1683 513
rect 1622 490 1631 510
rect 1651 493 1683 510
rect 1704 493 1709 513
rect 1651 490 1709 493
rect 1622 483 1709 490
rect 1734 510 1771 580
rect 2037 579 2074 580
rect 1886 520 1922 521
rect 1734 490 1743 510
rect 1763 490 1771 510
rect 1622 481 1678 483
rect 1622 480 1659 481
rect 1734 480 1771 490
rect 1830 510 1978 520
rect 2078 517 2174 519
rect 1830 490 1839 510
rect 1859 490 1949 510
rect 1969 490 1978 510
rect 1830 481 1978 490
rect 2036 510 2174 517
rect 2036 490 2045 510
rect 2065 490 2174 510
rect 2036 481 2174 490
rect 1830 480 1867 481
rect 1886 429 1922 481
rect 1941 480 1978 481
rect 2037 480 2074 481
rect 106 410 116 428
rect 134 427 739 428
rect 1357 427 1398 428
rect 134 422 155 427
rect 134 410 146 422
rect 1249 420 1398 427
rect 106 402 146 410
rect 189 409 215 410
rect 106 400 143 402
rect 189 391 743 409
rect 1249 400 1367 420
rect 1387 400 1398 420
rect 1249 392 1398 400
rect 1465 424 1824 428
rect 1465 419 1787 424
rect 1465 395 1578 419
rect 1602 400 1787 419
rect 1811 400 1824 424
rect 1602 395 1824 400
rect 1465 392 1824 395
rect 1886 392 1921 429
rect 1989 426 2089 429
rect 1989 422 2056 426
rect 1989 396 2001 422
rect 2027 400 2056 422
rect 2082 400 2089 426
rect 2027 396 2089 400
rect 1989 392 2089 396
rect 109 332 146 338
rect 189 332 215 391
rect 722 372 743 391
rect 109 329 215 332
rect 109 311 118 329
rect 136 315 215 329
rect 300 347 550 371
rect 136 313 212 315
rect 136 311 146 313
rect 109 301 146 311
rect 114 236 145 301
rect 300 276 337 347
rect 452 286 483 287
rect 300 256 309 276
rect 329 256 337 276
rect 300 246 337 256
rect 396 276 483 286
rect 396 256 405 276
rect 425 256 483 276
rect 396 247 483 256
rect 396 246 433 247
rect 113 227 150 236
rect 113 209 123 227
rect 141 209 150 227
rect 113 199 150 209
rect 452 194 483 247
rect 513 276 550 347
rect 721 352 1114 372
rect 1134 352 1137 372
rect 1465 371 1496 392
rect 1886 371 1922 392
rect 1308 370 1345 371
rect 721 347 1137 352
rect 1307 361 1345 370
rect 721 346 1062 347
rect 665 286 696 287
rect 513 256 522 276
rect 542 256 550 276
rect 513 246 550 256
rect 609 279 696 286
rect 609 276 670 279
rect 609 256 618 276
rect 638 259 670 276
rect 691 259 696 279
rect 638 256 696 259
rect 609 249 696 256
rect 721 276 758 346
rect 1024 345 1061 346
rect 1307 341 1316 361
rect 1336 341 1345 361
rect 1307 333 1345 341
rect 1411 365 1496 371
rect 1521 370 1558 371
rect 1411 345 1419 365
rect 1439 345 1496 365
rect 1411 337 1496 345
rect 1520 361 1558 370
rect 1520 341 1529 361
rect 1549 341 1558 361
rect 1411 336 1447 337
rect 1520 333 1558 341
rect 1624 365 1709 371
rect 1729 370 1766 371
rect 1624 345 1632 365
rect 1652 364 1709 365
rect 1652 345 1681 364
rect 1624 344 1681 345
rect 1702 344 1709 364
rect 1624 337 1709 344
rect 1728 361 1766 370
rect 1728 341 1737 361
rect 1757 341 1766 361
rect 1624 336 1660 337
rect 1728 333 1766 341
rect 1832 365 1976 371
rect 1832 345 1840 365
rect 1860 345 1892 365
rect 1916 345 1948 365
rect 1968 345 1976 365
rect 1832 337 1976 345
rect 1832 336 1868 337
rect 1940 336 1976 337
rect 2042 370 2079 371
rect 2042 369 2080 370
rect 2042 361 2106 369
rect 2042 341 2051 361
rect 2071 347 2106 361
rect 2126 347 2129 367
rect 2071 342 2129 347
rect 2071 341 2106 342
rect 1308 304 1345 333
rect 1309 302 1345 304
rect 1521 302 1558 333
rect 873 286 909 287
rect 721 256 730 276
rect 750 256 758 276
rect 609 247 665 249
rect 609 246 646 247
rect 721 246 758 256
rect 817 276 965 286
rect 1065 283 1161 285
rect 817 256 826 276
rect 846 256 936 276
rect 956 256 965 276
rect 817 247 965 256
rect 1023 276 1161 283
rect 1309 280 1558 302
rect 1729 301 1766 333
rect 2042 329 2106 341
rect 2146 303 2173 481
rect 2005 301 2173 303
rect 1729 297 2173 301
rect 1023 256 1032 276
rect 1052 256 1161 276
rect 1729 278 1778 297
rect 1798 278 2173 297
rect 1729 275 2173 278
rect 2005 274 2173 275
rect 1023 247 1161 256
rect 817 246 854 247
rect 873 195 909 247
rect 928 246 965 247
rect 1024 246 1061 247
rect 344 193 385 194
rect 236 186 385 193
rect 236 166 354 186
rect 374 166 385 186
rect 236 158 385 166
rect 452 190 811 194
rect 452 185 774 190
rect 452 161 565 185
rect 589 166 774 185
rect 798 166 811 190
rect 589 161 811 166
rect 452 158 811 161
rect 873 158 908 195
rect 976 192 1076 195
rect 976 188 1043 192
rect 976 162 988 188
rect 1014 166 1043 188
rect 1069 166 1076 192
rect 1014 162 1076 166
rect 976 158 1076 162
rect 452 137 483 158
rect 873 137 909 158
rect 116 128 153 137
rect 295 136 332 137
rect 116 110 125 128
rect 143 110 153 128
rect 116 100 153 110
rect 117 65 153 100
rect 294 127 332 136
rect 294 107 303 127
rect 323 107 332 127
rect 294 99 332 107
rect 398 131 483 137
rect 508 136 545 137
rect 398 111 406 131
rect 426 111 483 131
rect 398 103 483 111
rect 507 127 545 136
rect 507 107 516 127
rect 536 107 545 127
rect 398 102 434 103
rect 507 99 545 107
rect 611 131 696 137
rect 716 136 753 137
rect 611 111 619 131
rect 639 130 696 131
rect 639 111 668 130
rect 611 110 668 111
rect 689 110 696 130
rect 611 103 696 110
rect 715 127 753 136
rect 715 107 724 127
rect 744 107 753 127
rect 611 102 647 103
rect 715 99 753 107
rect 819 131 963 137
rect 819 111 827 131
rect 847 130 935 131
rect 847 111 875 130
rect 819 109 875 111
rect 897 111 935 130
rect 955 111 963 131
rect 897 109 963 111
rect 819 103 963 109
rect 819 102 855 103
rect 927 102 963 103
rect 1029 136 1066 137
rect 1029 135 1067 136
rect 1029 127 1093 135
rect 1029 107 1038 127
rect 1058 113 1093 127
rect 1113 113 1116 133
rect 1058 108 1116 113
rect 1058 107 1093 108
rect 295 70 332 99
rect 115 24 153 65
rect 296 68 332 70
rect 508 68 545 99
rect 296 46 545 68
rect 716 67 753 99
rect 1029 95 1093 107
rect 1133 69 1160 247
rect 992 67 1160 69
rect 716 41 1160 67
rect 717 24 741 41
rect 992 40 1160 41
rect 115 6 742 24
rect 1368 20 1618 44
rect 115 0 153 6
rect 115 -24 152 0
rect 115 -48 150 -24
rect 113 -57 150 -48
rect 113 -75 123 -57
rect 141 -75 150 -57
rect 113 -85 150 -75
rect 1368 -51 1405 20
rect 1520 -41 1551 -40
rect 1368 -71 1377 -51
rect 1397 -71 1405 -51
rect 1368 -81 1405 -71
rect 1464 -51 1551 -41
rect 1464 -71 1473 -51
rect 1493 -71 1551 -51
rect 1464 -80 1551 -71
rect 1464 -81 1501 -80
rect 1520 -133 1551 -80
rect 1581 -51 1618 20
rect 1789 25 2182 45
rect 2202 25 2205 45
rect 1789 20 2205 25
rect 1789 19 2130 20
rect 1733 -41 1764 -40
rect 1581 -71 1590 -51
rect 1610 -71 1618 -51
rect 1581 -81 1618 -71
rect 1677 -48 1764 -41
rect 1677 -51 1738 -48
rect 1677 -71 1686 -51
rect 1706 -68 1738 -51
rect 1759 -68 1764 -48
rect 1706 -71 1764 -68
rect 1677 -78 1764 -71
rect 1789 -51 1826 19
rect 2092 18 2129 19
rect 1941 -41 1977 -40
rect 1789 -71 1798 -51
rect 1818 -71 1826 -51
rect 1677 -80 1733 -78
rect 1677 -81 1714 -80
rect 1789 -81 1826 -71
rect 1885 -51 2033 -41
rect 2133 -44 2229 -42
rect 1885 -71 1894 -51
rect 1914 -71 2004 -51
rect 2024 -71 2033 -51
rect 1885 -80 2033 -71
rect 2091 -51 2229 -44
rect 2091 -71 2100 -51
rect 2120 -71 2229 -51
rect 2091 -80 2229 -71
rect 1885 -81 1922 -80
rect 1941 -132 1977 -80
rect 1996 -81 2033 -80
rect 2092 -81 2129 -80
rect 1412 -134 1453 -133
rect 1304 -141 1453 -134
rect 116 -149 153 -147
rect 116 -150 764 -149
rect 115 -156 764 -150
rect 115 -174 125 -156
rect 143 -170 764 -156
rect 1304 -161 1422 -141
rect 1442 -161 1453 -141
rect 1304 -169 1453 -161
rect 1520 -137 1879 -133
rect 1520 -142 1842 -137
rect 1520 -166 1633 -142
rect 1657 -161 1842 -142
rect 1866 -161 1879 -137
rect 1657 -166 1879 -161
rect 1520 -169 1879 -166
rect 1941 -169 1976 -132
rect 2044 -135 2144 -132
rect 2044 -139 2111 -135
rect 2044 -165 2056 -139
rect 2082 -161 2111 -139
rect 2137 -161 2144 -135
rect 2082 -165 2144 -161
rect 2044 -169 2144 -165
rect 143 -174 153 -170
rect 594 -171 764 -170
rect 115 -184 153 -174
rect 115 -262 150 -184
rect 727 -194 764 -171
rect 1520 -190 1551 -169
rect 1941 -190 1977 -169
rect 1363 -191 1400 -190
rect 111 -271 150 -262
rect 111 -289 121 -271
rect 139 -289 150 -271
rect 111 -295 150 -289
rect 306 -219 556 -195
rect 306 -290 343 -219
rect 458 -280 489 -279
rect 111 -299 148 -295
rect 306 -310 315 -290
rect 335 -310 343 -290
rect 306 -320 343 -310
rect 402 -290 489 -280
rect 402 -310 411 -290
rect 431 -310 489 -290
rect 402 -319 489 -310
rect 402 -320 439 -319
rect 114 -370 151 -361
rect 112 -388 123 -370
rect 141 -388 151 -370
rect 458 -372 489 -319
rect 519 -290 556 -219
rect 727 -214 1120 -194
rect 1140 -214 1143 -194
rect 727 -219 1143 -214
rect 1362 -200 1400 -191
rect 727 -220 1068 -219
rect 1362 -220 1371 -200
rect 1391 -220 1400 -200
rect 671 -280 702 -279
rect 519 -310 528 -290
rect 548 -310 556 -290
rect 519 -320 556 -310
rect 615 -287 702 -280
rect 615 -290 676 -287
rect 615 -310 624 -290
rect 644 -307 676 -290
rect 697 -307 702 -287
rect 644 -310 702 -307
rect 615 -317 702 -310
rect 727 -290 764 -220
rect 1030 -221 1067 -220
rect 1362 -228 1400 -220
rect 1466 -196 1551 -190
rect 1576 -191 1613 -190
rect 1466 -216 1474 -196
rect 1494 -216 1551 -196
rect 1466 -224 1551 -216
rect 1575 -200 1613 -191
rect 1575 -220 1584 -200
rect 1604 -220 1613 -200
rect 1466 -225 1502 -224
rect 1575 -228 1613 -220
rect 1679 -196 1764 -190
rect 1784 -191 1821 -190
rect 1679 -216 1687 -196
rect 1707 -197 1764 -196
rect 1707 -216 1736 -197
rect 1679 -217 1736 -216
rect 1757 -217 1764 -197
rect 1679 -224 1764 -217
rect 1783 -200 1821 -191
rect 1783 -220 1792 -200
rect 1812 -220 1821 -200
rect 1679 -225 1715 -224
rect 1783 -228 1821 -220
rect 1887 -196 2031 -190
rect 1887 -216 1895 -196
rect 1915 -216 2003 -196
rect 2023 -216 2031 -196
rect 1887 -224 2031 -216
rect 1887 -225 1923 -224
rect 1995 -225 2031 -224
rect 2097 -191 2134 -190
rect 2097 -192 2135 -191
rect 2097 -200 2161 -192
rect 2097 -220 2106 -200
rect 2126 -214 2161 -200
rect 2181 -214 2184 -194
rect 2126 -219 2184 -214
rect 2126 -220 2161 -219
rect 1363 -257 1400 -228
rect 1364 -259 1400 -257
rect 1576 -259 1613 -228
rect 879 -280 915 -279
rect 727 -310 736 -290
rect 756 -310 764 -290
rect 615 -319 671 -317
rect 615 -320 652 -319
rect 727 -320 764 -310
rect 823 -290 971 -280
rect 1364 -281 1613 -259
rect 1784 -260 1821 -228
rect 2097 -232 2161 -220
rect 2201 -258 2228 -80
rect 2060 -260 2228 -258
rect 1784 -271 2228 -260
rect 1071 -283 1167 -281
rect 823 -310 832 -290
rect 852 -310 942 -290
rect 962 -310 971 -290
rect 823 -319 971 -310
rect 1029 -290 1167 -283
rect 1784 -286 2230 -271
rect 2060 -287 2230 -286
rect 1029 -310 1038 -290
rect 1058 -310 1167 -290
rect 1029 -319 1167 -310
rect 823 -320 860 -319
rect 879 -371 915 -319
rect 934 -320 971 -319
rect 1030 -320 1067 -319
rect 350 -373 391 -372
rect 112 -537 151 -388
rect 242 -380 391 -373
rect 242 -400 360 -380
rect 380 -400 391 -380
rect 242 -408 391 -400
rect 458 -376 817 -372
rect 458 -381 780 -376
rect 458 -405 571 -381
rect 595 -400 780 -381
rect 804 -400 817 -376
rect 595 -405 817 -400
rect 458 -408 817 -405
rect 879 -408 914 -371
rect 982 -374 1082 -371
rect 982 -378 1049 -374
rect 982 -404 994 -378
rect 1020 -400 1049 -378
rect 1075 -400 1082 -374
rect 1020 -404 1082 -400
rect 982 -408 1082 -404
rect 458 -429 489 -408
rect 879 -429 915 -408
rect 301 -430 338 -429
rect 300 -439 338 -430
rect 300 -459 309 -439
rect 329 -459 338 -439
rect 300 -467 338 -459
rect 404 -435 489 -429
rect 514 -430 551 -429
rect 404 -455 412 -435
rect 432 -455 489 -435
rect 404 -463 489 -455
rect 513 -439 551 -430
rect 513 -459 522 -439
rect 542 -459 551 -439
rect 404 -464 440 -463
rect 513 -467 551 -459
rect 617 -435 702 -429
rect 722 -430 759 -429
rect 617 -455 625 -435
rect 645 -436 702 -435
rect 645 -455 674 -436
rect 617 -456 674 -455
rect 695 -456 702 -436
rect 617 -463 702 -456
rect 721 -439 759 -430
rect 721 -459 730 -439
rect 750 -459 759 -439
rect 617 -464 653 -463
rect 721 -467 759 -459
rect 825 -434 969 -429
rect 825 -435 890 -434
rect 825 -455 833 -435
rect 853 -455 890 -435
rect 912 -435 969 -434
rect 912 -455 941 -435
rect 961 -455 969 -435
rect 825 -463 969 -455
rect 825 -464 861 -463
rect 933 -464 969 -463
rect 1035 -430 1072 -429
rect 1035 -431 1073 -430
rect 1035 -439 1099 -431
rect 1035 -459 1044 -439
rect 1064 -453 1099 -439
rect 1119 -453 1122 -433
rect 1064 -458 1122 -453
rect 1064 -459 1099 -458
rect 301 -496 338 -467
rect 302 -498 338 -496
rect 514 -498 551 -467
rect 302 -520 551 -498
rect 722 -499 759 -467
rect 1035 -471 1099 -459
rect 1139 -497 1166 -319
rect 998 -499 1166 -497
rect 722 -525 1166 -499
rect 1318 -400 1568 -376
rect 1318 -471 1355 -400
rect 1470 -461 1501 -460
rect 1318 -491 1327 -471
rect 1347 -491 1355 -471
rect 1318 -501 1355 -491
rect 1414 -471 1501 -461
rect 1414 -491 1423 -471
rect 1443 -491 1501 -471
rect 1414 -500 1501 -491
rect 1414 -501 1451 -500
rect 722 -535 744 -525
rect 998 -526 1166 -525
rect 682 -537 744 -535
rect 112 -544 744 -537
rect 111 -553 744 -544
rect 1470 -553 1501 -500
rect 1531 -471 1568 -400
rect 1739 -395 2132 -375
rect 2152 -395 2155 -375
rect 1739 -400 2155 -395
rect 1739 -401 2080 -400
rect 1683 -461 1714 -460
rect 1531 -491 1540 -471
rect 1560 -491 1568 -471
rect 1531 -501 1568 -491
rect 1627 -468 1714 -461
rect 1627 -471 1688 -468
rect 1627 -491 1636 -471
rect 1656 -488 1688 -471
rect 1709 -488 1714 -468
rect 1656 -491 1714 -488
rect 1627 -498 1714 -491
rect 1739 -471 1776 -401
rect 2042 -402 2079 -401
rect 1891 -461 1927 -460
rect 1739 -491 1748 -471
rect 1768 -491 1776 -471
rect 1627 -500 1683 -498
rect 1627 -501 1664 -500
rect 1739 -501 1776 -491
rect 1835 -471 1983 -461
rect 2083 -464 2179 -462
rect 1835 -491 1844 -471
rect 1864 -491 1954 -471
rect 1974 -491 1983 -471
rect 1835 -500 1983 -491
rect 2041 -471 2179 -464
rect 2041 -491 2050 -471
rect 2070 -491 2179 -471
rect 2041 -500 2179 -491
rect 1835 -501 1872 -500
rect 1891 -552 1927 -500
rect 1946 -501 1983 -500
rect 2042 -501 2079 -500
rect 111 -571 121 -553
rect 139 -554 744 -553
rect 1362 -554 1403 -553
rect 139 -559 160 -554
rect 139 -571 151 -559
rect 1254 -561 1403 -554
rect 111 -579 151 -571
rect 194 -572 220 -571
rect 111 -581 148 -579
rect 194 -590 748 -572
rect 1254 -581 1372 -561
rect 1392 -581 1403 -561
rect 1254 -589 1403 -581
rect 1470 -557 1829 -553
rect 1470 -562 1792 -557
rect 1470 -586 1583 -562
rect 1607 -581 1792 -562
rect 1816 -581 1829 -557
rect 1607 -586 1829 -581
rect 1470 -589 1829 -586
rect 1891 -589 1926 -552
rect 1994 -555 2094 -552
rect 1994 -559 2061 -555
rect 1994 -585 2006 -559
rect 2032 -581 2061 -559
rect 2087 -581 2094 -555
rect 2032 -585 2094 -581
rect 1994 -589 2094 -585
rect 114 -649 151 -643
rect 194 -649 220 -590
rect 727 -609 748 -590
rect 114 -652 220 -649
rect 114 -670 123 -652
rect 141 -666 220 -652
rect 305 -634 555 -610
rect 141 -668 217 -666
rect 141 -670 151 -668
rect 114 -680 151 -670
rect 119 -745 150 -680
rect 305 -705 342 -634
rect 457 -695 488 -694
rect 305 -725 314 -705
rect 334 -725 342 -705
rect 305 -735 342 -725
rect 401 -705 488 -695
rect 401 -725 410 -705
rect 430 -725 488 -705
rect 401 -734 488 -725
rect 401 -735 438 -734
rect 118 -754 155 -745
rect 118 -772 128 -754
rect 146 -772 155 -754
rect 118 -782 155 -772
rect 457 -787 488 -734
rect 518 -705 555 -634
rect 726 -629 1119 -609
rect 1139 -629 1142 -609
rect 1470 -610 1501 -589
rect 1891 -610 1927 -589
rect 1313 -611 1350 -610
rect 726 -634 1142 -629
rect 1312 -620 1350 -611
rect 726 -635 1067 -634
rect 670 -695 701 -694
rect 518 -725 527 -705
rect 547 -725 555 -705
rect 518 -735 555 -725
rect 614 -702 701 -695
rect 614 -705 675 -702
rect 614 -725 623 -705
rect 643 -722 675 -705
rect 696 -722 701 -702
rect 643 -725 701 -722
rect 614 -732 701 -725
rect 726 -705 763 -635
rect 1029 -636 1066 -635
rect 1312 -640 1321 -620
rect 1341 -640 1350 -620
rect 1312 -648 1350 -640
rect 1416 -616 1501 -610
rect 1526 -611 1563 -610
rect 1416 -636 1424 -616
rect 1444 -636 1501 -616
rect 1416 -644 1501 -636
rect 1525 -620 1563 -611
rect 1525 -640 1534 -620
rect 1554 -640 1563 -620
rect 1416 -645 1452 -644
rect 1525 -648 1563 -640
rect 1629 -616 1714 -610
rect 1734 -611 1771 -610
rect 1629 -636 1637 -616
rect 1657 -617 1714 -616
rect 1657 -636 1686 -617
rect 1629 -637 1686 -636
rect 1707 -637 1714 -617
rect 1629 -644 1714 -637
rect 1733 -620 1771 -611
rect 1733 -640 1742 -620
rect 1762 -640 1771 -620
rect 1629 -645 1665 -644
rect 1733 -648 1771 -640
rect 1837 -615 1981 -610
rect 1837 -616 1896 -615
rect 1837 -636 1845 -616
rect 1865 -635 1896 -616
rect 1920 -616 1981 -615
rect 1920 -635 1953 -616
rect 1865 -636 1953 -635
rect 1973 -636 1981 -616
rect 1837 -644 1981 -636
rect 1837 -645 1873 -644
rect 1945 -645 1981 -644
rect 2047 -611 2084 -610
rect 2047 -612 2085 -611
rect 2047 -620 2111 -612
rect 2047 -640 2056 -620
rect 2076 -634 2111 -620
rect 2131 -634 2134 -614
rect 2076 -639 2134 -634
rect 2076 -640 2111 -639
rect 1313 -677 1350 -648
rect 1314 -679 1350 -677
rect 1526 -679 1563 -648
rect 878 -695 914 -694
rect 726 -725 735 -705
rect 755 -725 763 -705
rect 614 -734 670 -732
rect 614 -735 651 -734
rect 726 -735 763 -725
rect 822 -705 970 -695
rect 1070 -698 1166 -696
rect 822 -725 831 -705
rect 851 -725 941 -705
rect 961 -725 970 -705
rect 822 -734 970 -725
rect 1028 -705 1166 -698
rect 1314 -701 1563 -679
rect 1734 -680 1771 -648
rect 2047 -652 2111 -640
rect 2151 -678 2178 -500
rect 2010 -680 2178 -678
rect 1734 -684 2178 -680
rect 1028 -725 1037 -705
rect 1057 -725 1166 -705
rect 1734 -703 1783 -684
rect 1803 -703 2178 -684
rect 1734 -706 2178 -703
rect 2010 -707 2178 -706
rect 2199 -681 2230 -287
rect 2199 -707 2204 -681
rect 2223 -707 2230 -681
rect 2199 -710 2230 -707
rect 1028 -734 1166 -725
rect 822 -735 859 -734
rect 878 -786 914 -734
rect 933 -735 970 -734
rect 1029 -735 1066 -734
rect 349 -788 390 -787
rect 241 -795 390 -788
rect 241 -815 359 -795
rect 379 -815 390 -795
rect 241 -823 390 -815
rect 457 -791 816 -787
rect 457 -796 779 -791
rect 457 -820 570 -796
rect 594 -815 779 -796
rect 803 -815 816 -791
rect 594 -820 816 -815
rect 457 -823 816 -820
rect 878 -823 913 -786
rect 981 -789 1081 -786
rect 981 -793 1048 -789
rect 981 -819 993 -793
rect 1019 -815 1048 -793
rect 1074 -815 1081 -789
rect 1019 -819 1081 -815
rect 981 -823 1081 -819
rect 457 -844 488 -823
rect 878 -844 914 -823
rect 121 -853 158 -844
rect 300 -845 337 -844
rect 121 -871 130 -853
rect 148 -871 158 -853
rect 121 -881 158 -871
rect 122 -916 158 -881
rect 299 -854 337 -845
rect 299 -874 308 -854
rect 328 -874 337 -854
rect 299 -882 337 -874
rect 403 -850 488 -844
rect 513 -845 550 -844
rect 403 -870 411 -850
rect 431 -870 488 -850
rect 403 -878 488 -870
rect 512 -854 550 -845
rect 512 -874 521 -854
rect 541 -874 550 -854
rect 403 -879 439 -878
rect 512 -882 550 -874
rect 616 -850 701 -844
rect 721 -845 758 -844
rect 616 -870 624 -850
rect 644 -851 701 -850
rect 644 -870 673 -851
rect 616 -871 673 -870
rect 694 -871 701 -851
rect 616 -878 701 -871
rect 720 -854 758 -845
rect 720 -874 729 -854
rect 749 -874 758 -854
rect 616 -879 652 -878
rect 720 -882 758 -874
rect 824 -850 968 -844
rect 824 -870 832 -850
rect 852 -851 940 -850
rect 852 -870 880 -851
rect 824 -872 880 -870
rect 902 -870 940 -851
rect 960 -870 968 -850
rect 902 -872 968 -870
rect 824 -878 968 -872
rect 824 -879 860 -878
rect 932 -879 968 -878
rect 1034 -845 1071 -844
rect 1034 -846 1072 -845
rect 1034 -854 1098 -846
rect 1034 -874 1043 -854
rect 1063 -868 1098 -854
rect 1118 -868 1121 -848
rect 1063 -873 1121 -868
rect 1063 -874 1098 -873
rect 300 -911 337 -882
rect 120 -957 158 -916
rect 301 -913 337 -911
rect 513 -913 550 -882
rect 301 -935 550 -913
rect 721 -914 758 -882
rect 1034 -886 1098 -874
rect 1138 -912 1165 -734
rect 997 -914 1165 -912
rect 721 -940 1165 -914
rect 722 -957 746 -940
rect 997 -941 1165 -940
rect 120 -975 747 -957
rect 120 -981 158 -975
<< viali >>
rect 1115 767 1135 787
rect 671 674 692 694
rect 1044 581 1070 607
rect 669 525 690 545
rect 885 526 907 547
rect 1094 528 1114 548
rect 2127 586 2147 606
rect 1683 493 1704 513
rect 2056 400 2082 426
rect 1114 352 1134 372
rect 670 259 691 279
rect 1681 344 1702 364
rect 1892 345 1916 365
rect 2106 347 2126 367
rect 1778 278 1798 297
rect 1043 166 1069 192
rect 668 110 689 130
rect 875 109 897 130
rect 1093 113 1113 133
rect 2182 25 2202 45
rect 1738 -68 1759 -48
rect 2111 -161 2137 -135
rect 1120 -214 1140 -194
rect 676 -307 697 -287
rect 1736 -217 1757 -197
rect 2161 -214 2181 -194
rect 1049 -400 1075 -374
rect 674 -456 695 -436
rect 890 -455 912 -434
rect 1099 -453 1119 -433
rect 2132 -395 2152 -375
rect 1688 -488 1709 -468
rect 2061 -581 2087 -555
rect 1119 -629 1139 -609
rect 675 -722 696 -702
rect 1686 -637 1707 -617
rect 1896 -635 1920 -615
rect 2111 -634 2131 -614
rect 1783 -703 1803 -684
rect 2204 -707 2223 -681
rect 1048 -815 1074 -789
rect 673 -871 694 -851
rect 880 -872 902 -851
rect 1098 -868 1118 -848
<< metal1 >>
rect 1111 792 1143 793
rect 1108 787 1143 792
rect 1108 767 1115 787
rect 1135 767 1143 787
rect 1108 759 1143 767
rect 664 694 696 701
rect 664 674 671 694
rect 692 674 696 694
rect 664 609 696 674
rect 1034 609 1074 610
rect 664 607 1076 609
rect 664 581 1044 607
rect 1070 581 1076 607
rect 664 573 1076 581
rect 664 545 696 573
rect 1109 553 1143 759
rect 664 525 669 545
rect 690 525 696 545
rect 664 518 696 525
rect 873 547 913 552
rect 873 526 885 547
rect 907 526 913 547
rect 873 514 913 526
rect 1087 548 1143 553
rect 1087 528 1094 548
rect 1114 528 1143 548
rect 1087 521 1143 528
rect 1200 622 2157 641
rect 1087 520 1122 521
rect 879 482 907 514
rect 1200 482 1231 622
rect 2120 606 2155 622
rect 2120 586 2127 606
rect 2147 586 2155 606
rect 2120 578 2155 586
rect 879 451 1231 482
rect 1676 513 1708 520
rect 1676 493 1683 513
rect 1704 493 1708 513
rect 1676 428 1708 493
rect 2046 428 2086 429
rect 1676 426 2088 428
rect 1676 400 2056 426
rect 2082 400 2088 426
rect 1676 392 2088 400
rect 1110 377 1142 378
rect 1107 372 1142 377
rect 1107 352 1114 372
rect 1134 352 1142 372
rect 1107 344 1142 352
rect 663 279 695 286
rect 663 259 670 279
rect 691 259 695 279
rect 663 194 695 259
rect 1033 194 1073 195
rect 663 192 1075 194
rect 663 166 1043 192
rect 1069 166 1075 192
rect 663 158 1075 166
rect 663 130 695 158
rect 663 110 668 130
rect 689 110 695 130
rect 663 103 695 110
rect 863 130 913 139
rect 1108 138 1142 344
rect 1676 364 1708 392
rect 1676 344 1681 364
rect 1702 344 1708 364
rect 1676 337 1708 344
rect 1883 365 1925 373
rect 2121 372 2155 578
rect 1883 345 1892 365
rect 1916 345 1925 365
rect 1883 333 1925 345
rect 2099 367 2155 372
rect 2099 347 2106 367
rect 2126 347 2155 367
rect 2099 340 2155 347
rect 2099 339 2134 340
rect 1885 304 1920 333
rect 1885 303 2195 304
rect 1770 297 1806 301
rect 1770 278 1778 297
rect 1798 278 1806 297
rect 1770 275 1806 278
rect 1771 247 1805 275
rect 1885 269 2212 303
rect 863 109 875 130
rect 897 109 913 130
rect 863 101 913 109
rect 1086 133 1142 138
rect 1086 113 1093 133
rect 1113 113 1142 133
rect 1086 106 1142 113
rect 1243 219 1806 247
rect 1086 105 1121 106
rect 868 68 909 101
rect 1243 68 1283 219
rect 868 39 1283 68
rect 2172 45 2212 269
rect 868 38 1277 39
rect 2172 25 2182 45
rect 2202 25 2212 45
rect 2172 15 2212 25
rect 1731 -48 1763 -41
rect 1731 -68 1738 -48
rect 1759 -68 1763 -48
rect 1731 -133 1763 -68
rect 2101 -133 2141 -132
rect 1731 -135 2143 -133
rect 1731 -161 2111 -135
rect 2137 -161 2143 -135
rect 1731 -169 2143 -161
rect 1116 -189 1148 -188
rect 1113 -194 1148 -189
rect 1113 -214 1120 -194
rect 1140 -214 1148 -194
rect 1113 -222 1148 -214
rect 669 -287 701 -280
rect 669 -307 676 -287
rect 697 -307 701 -287
rect 669 -372 701 -307
rect 1039 -372 1079 -371
rect 669 -374 1081 -372
rect 669 -400 1049 -374
rect 1075 -400 1081 -374
rect 669 -408 1081 -400
rect 669 -436 701 -408
rect 1114 -428 1148 -222
rect 1731 -197 1763 -169
rect 2176 -189 2210 15
rect 1731 -217 1736 -197
rect 1757 -217 1763 -197
rect 1731 -224 1763 -217
rect 2154 -194 2210 -189
rect 2154 -214 2161 -194
rect 2181 -214 2210 -194
rect 2154 -221 2210 -214
rect 2154 -222 2189 -221
rect 669 -456 674 -436
rect 695 -456 701 -436
rect 669 -463 701 -456
rect 878 -434 918 -429
rect 878 -455 890 -434
rect 912 -455 918 -434
rect 878 -467 918 -455
rect 1092 -433 1148 -428
rect 1092 -453 1099 -433
rect 1119 -453 1148 -433
rect 1092 -460 1148 -453
rect 1205 -359 2162 -340
rect 1092 -461 1127 -460
rect 884 -499 912 -467
rect 1205 -499 1236 -359
rect 2125 -375 2160 -359
rect 2125 -395 2132 -375
rect 2152 -395 2160 -375
rect 2125 -403 2160 -395
rect 884 -530 1236 -499
rect 1681 -468 1713 -461
rect 1681 -488 1688 -468
rect 1709 -488 1713 -468
rect 1681 -553 1713 -488
rect 2051 -553 2091 -552
rect 1681 -555 2093 -553
rect 1681 -581 2061 -555
rect 2087 -581 2093 -555
rect 1681 -589 2093 -581
rect 1115 -604 1147 -603
rect 1112 -609 1147 -604
rect 1112 -629 1119 -609
rect 1139 -629 1147 -609
rect 1112 -637 1147 -629
rect 668 -702 700 -695
rect 668 -722 675 -702
rect 696 -722 700 -702
rect 668 -787 700 -722
rect 1038 -787 1078 -786
rect 668 -789 1080 -787
rect 668 -815 1048 -789
rect 1074 -815 1080 -789
rect 668 -823 1080 -815
rect 668 -851 700 -823
rect 668 -871 673 -851
rect 694 -871 700 -851
rect 668 -878 700 -871
rect 868 -851 918 -842
rect 1113 -843 1147 -637
rect 1681 -617 1713 -589
rect 1681 -637 1686 -617
rect 1707 -637 1713 -617
rect 1886 -615 1928 -606
rect 2126 -609 2160 -403
rect 1886 -629 1896 -615
rect 1681 -644 1713 -637
rect 1885 -635 1896 -629
rect 1920 -635 1928 -615
rect 1885 -646 1928 -635
rect 2104 -614 2160 -609
rect 2104 -634 2111 -614
rect 2131 -634 2160 -614
rect 2104 -641 2160 -634
rect 2104 -642 2139 -641
rect 1885 -676 1925 -646
rect 1775 -684 1811 -680
rect 1775 -703 1783 -684
rect 1803 -703 1811 -684
rect 1775 -706 1811 -703
rect 1885 -681 2232 -676
rect 1776 -734 1810 -706
rect 1885 -707 2204 -681
rect 2223 -707 2232 -681
rect 1885 -711 2232 -707
rect 868 -872 880 -851
rect 902 -872 918 -851
rect 868 -880 918 -872
rect 1091 -848 1147 -843
rect 1091 -868 1098 -848
rect 1118 -868 1147 -848
rect 1091 -875 1147 -868
rect 1248 -762 1811 -734
rect 1091 -876 1126 -875
rect 873 -913 914 -880
rect 1248 -913 1288 -762
rect 873 -942 1288 -913
rect 873 -943 1282 -942
<< labels >>
rlabel locali 304 771 333 777 1 vdd
rlabel locali 517 768 546 774 1 vdd
rlabel locali 250 583 272 598 1 d0
rlabel nwell 671 738 694 741 1 vdd
rlabel locali 301 472 330 478 1 gnd
rlabel locali 514 472 543 478 1 gnd
rlabel space 611 467 640 476 1 gnd
rlabel locali 303 356 332 362 1 vdd
rlabel locali 516 353 545 359 1 vdd
rlabel locali 249 168 271 183 1 d0
rlabel nwell 670 323 693 326 1 vdd
rlabel locali 300 57 329 63 1 gnd
rlabel locali 513 57 542 63 1 gnd
rlabel space 610 52 639 61 1 gnd
rlabel locali 1316 590 1345 596 1 vdd
rlabel locali 1529 587 1558 593 1 vdd
rlabel nwell 1683 557 1706 560 1 vdd
rlabel locali 1313 291 1342 297 1 gnd
rlabel locali 1526 291 1555 297 1 gnd
rlabel space 1623 286 1652 295 1 gnd
rlabel locali 1254 401 1301 422 1 d1
rlabel locali 116 963 141 972 1 vref
rlabel locali 309 -210 338 -204 1 vdd
rlabel locali 522 -213 551 -207 1 vdd
rlabel locali 255 -398 277 -383 1 d0
rlabel nwell 676 -243 699 -240 1 vdd
rlabel locali 306 -509 335 -503 1 gnd
rlabel locali 519 -509 548 -503 1 gnd
rlabel space 616 -514 645 -505 1 gnd
rlabel locali 308 -625 337 -619 1 vdd
rlabel locali 521 -628 550 -622 1 vdd
rlabel locali 254 -813 276 -798 1 d0
rlabel nwell 675 -658 698 -655 1 vdd
rlabel locali 305 -924 334 -918 1 gnd
rlabel locali 518 -924 547 -918 1 gnd
rlabel space 615 -929 644 -920 1 gnd
rlabel locali 1321 -391 1350 -385 1 vdd
rlabel locali 1534 -394 1563 -388 1 vdd
rlabel nwell 1688 -424 1711 -421 1 vdd
rlabel locali 1318 -690 1347 -684 1 gnd
rlabel locali 1531 -690 1560 -684 1 gnd
rlabel space 1628 -695 1657 -686 1 gnd
rlabel locali 1259 -580 1306 -559 1 d1
rlabel locali 126 -973 153 -960 1 gnd
rlabel locali 1371 29 1400 35 1 vdd
rlabel locali 1584 26 1613 32 1 vdd
rlabel locali 1947 -124 1969 -109 1 vout
rlabel nwell 1738 -4 1761 -1 1 vdd
rlabel locali 1368 -270 1397 -264 1 gnd
rlabel locali 1581 -270 1610 -264 1 gnd
rlabel space 1678 -275 1707 -266 1 gnd
rlabel locali 1314 -159 1337 -144 1 d2
<< end >>
