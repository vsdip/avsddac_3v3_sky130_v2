* SPICE3 file created from 7bit_DAC.ext - technology: sky130A

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_2745_8212# a_2998_8199# a_2776_7096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 a_3822_2038# a_3828_1312# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2 a_5490_2942# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3 a_5705_1290# a_5492_1290# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4 a_7799_4018# a_7989_3236# a_7944_3249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5 a_120_1130# a_649_1249# a_857_1249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6 a_119_3752# a_119_3565# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7 a_5704_736# a_5491_736# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_7830_2902# a_7849_1622# a_7800_1812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9 a_1586_2108# a_1373_2108# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X10 a_1808_4963# a_1481_7044# a_1803_7044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X11 a_6849_5458# a_6428_5458# a_5910_5148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 a_8878_4839# a_9135_4649# a_7943_4352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X13 gnd a_3001_1581# a_2793_1581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X14 a_2888_2105# a_3141_2092# a_2748_1594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_7937_8941# a_8924_8507# a_8875_8697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_5909_6251# a_6640_6561# a_6848_6561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X17 a_2774_5061# a_3031_4871# a_2004_136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X18 a_5700_8457# a_5487_8457# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X19 a_6864_5004# a_6750_4885# a_6958_4885# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 a_8882_1902# a_9135_1889# a_7940_2323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X21 a_5702_4045# a_5489_4045# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X22 a_7939_4529# a_8926_4095# a_8877_4285# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X23 a_7830_2902# a_7849_1622# a_7804_1635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X24 a_5172_9121# a_5172_8892# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X25 a_3821_7004# a_4078_6814# a_2886_6517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X26 vdd a_3001_1581# a_2793_1581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X27 a_7941_8764# a_8194_8751# a_7801_8253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X28 a_854_5107# a_1585_5417# a_1793_5417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X29 a_6640_7664# a_6427_7664# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X30 a_1371_6520# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X31 a_6641_4355# a_6428_4355# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X32 a_5175_3606# a_5704_3496# a_5912_3496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_856_2352# a_1586_2108# a_1794_2108# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X34 a_6861_2673# a_6752_2673# a_6859_4885# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X35 a_8879_3736# a_8882_3005# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X36 a_5173_6915# a_5173_6686# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X37 a_5492_1290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X38 a_856_695# a_1587_1005# a_1795_1005# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X39 a_1726_3722# a_1513_3722# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X40 a_6642_3252# a_6429_3252# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X41 a_3823_935# a_122_801# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X42 a_1373_2108# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X43 a_7937_8941# a_8194_8751# a_7801_8253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X44 a_852_8416# a_431_8416# a_116_8621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X45 a_6864_5004# a_6537_7085# a_6864_7204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X46 a_5913_1290# a_5492_1290# a_5176_1171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X47 a_8877_5388# a_9134_5198# a_7939_5632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X48 a_6849_5458# a_6781_5969# a_6859_7085# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X49 a_647_1798# a_434_1798# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X50 a_8883_2456# a_9136_2443# a_7944_2146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_6864_7204# a_6567_8175# a_6847_8767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X52 a_7939_4529# a_8196_4339# a_7803_3841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X53 a_854_4004# a_433_4004# a_118_4209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X54 a_5175_3147# a_5703_2942# a_5911_2942# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X55 a_5174_5999# a_5701_6251# a_5909_6251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X56 gnd d0 a_4080_745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X57 a_5908_8457# a_6639_8767# a_6847_8767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X58 a_8877_7045# a_9134_6855# a_7942_6558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X59 a_2887_4311# a_3140_4298# a_2747_3800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 gnd a_3000_3787# a_2792_3787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X61 a_8882_5765# a_8878_5942# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X62 a_117_7748# a_117_7518# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X63 a_2746_6006# a_2931_6504# a_2882_6694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X64 a_1895_136# a_1682_136# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X65 vout a_4632_116# a_2103_136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X66 a_8879_2633# a_9136_2443# a_7944_2146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X67 a_5910_4045# a_6641_4355# a_6849_4355# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X68 a_3820_7553# a_3825_6827# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X69 a_2004_136# a_2823_4871# a_2778_4884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X70 a_7943_4352# a_8927_4649# a_8882_4662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X71 a_5174_4250# a_5175_3793# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X72 a_3827_3518# a_4080_3505# a_2888_3208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 a_6782_3763# a_6569_3763# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X74 vdd d0 a_4080_745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X75 vdd d0 a_4079_1848# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X76 a_2748_1594# a_2933_2092# a_2884_2282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 a_1513_3722# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 a_6958_4885# a_6537_4885# a_6859_4885# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_7940_2323# a_8927_1889# a_8878_2079# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X80 a_119_2649# a_119_2462# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X81 a_3827_758# a_3823_935# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X82 a_5175_2044# a_5176_1587# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X83 a_2886_7620# a_3870_7917# a_3821_8107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X84 a_7942_6558# a_8195_6545# a_7802_6047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X85 a_6641_5458# a_6428_5458# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X86 a_434_1798# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X87 a_6642_2149# a_6429_2149# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X88 a_1725_5928# a_1512_5928# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X89 a_647_5661# a_434_5661# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_3823_2592# a_3826_1861# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X91 a_5488_9011# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_7801_8253# a_7986_8751# a_7937_8941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 a_117_6415# a_645_6210# a_853_6210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 a_5912_3496# a_5491_3496# a_5175_3377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X95 a_8876_7594# a_9133_7404# a_7938_7838# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X96 a_7830_5102# a_8087_4912# a_7060_177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X97 a_6643_1046# a_6430_1046# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X98 a_7944_2146# a_8197_2133# a_7804_1635# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X99 a_8882_4662# a_9135_4649# a_7943_4352# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X100 a_1727_1516# a_1514_1516# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_7938_6735# a_8195_6545# a_7802_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X102 a_853_6210# a_432_6210# a_117_6415# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X103 a_8883_799# a_9136_786# a_7941_1220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X104 gnd d0 a_9136_786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X105 a_5173_8205# a_5700_8457# a_5908_8457# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X106 gnd d4 a_8087_4912# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X107 a_5702_6805# a_5489_6805# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X108 a_8878_3182# a_9135_2992# a_7940_3426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X109 a_7801_8253# a_7986_8751# a_7941_8764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X110 a_6958_4885# a_6951_177# a_4954_116# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_8879_2633# a_8882_1902# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X112 a_2776_7096# a_2790_8199# a_2745_8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X113 a_117_6645# a_646_6764# a_854_6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X114 a_6859_7085# a_6568_5969# a_6848_6561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X115 a_7939_5632# a_8926_5198# a_8881_5211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X116 a_5175_3793# a_5702_4045# a_5910_4045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X117 a_7940_2323# a_8197_2133# a_7804_1635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X118 a_3822_3141# a_4079_2951# a_2884_3385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X119 a_6750_4885# a_6537_4885# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X120 a_5704_2393# a_5491_2393# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X121 a_7944_2146# a_8928_2443# a_8879_2633# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X122 a_5909_6251# a_5488_6251# a_5173_6456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X123 a_7803_3841# a_7988_4339# a_7943_4352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X124 a_8879_976# a_9136_786# a_7941_1220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X125 vdd d0 a_9136_786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X126 a_6781_5969# a_6568_5969# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X127 a_119_2233# a_648_2352# a_856_2352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X128 a_7942_6558# a_8926_6855# a_8881_6868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X129 a_2747_3800# a_2932_4298# a_2883_4488# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_6848_6561# a_6427_6561# a_5909_6251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X131 a_1512_5928# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X132 a_434_5661# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X133 a_1694_4844# a_1481_4844# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X134 a_2103_136# a_1682_136# a_2004_136# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 a_5911_1839# a_6642_2149# a_6850_2149# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X136 a_6783_1557# a_6570_1557# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 a_6430_1046# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X138 a_3828_1312# a_4081_1299# a_2889_1002# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_7944_2146# a_8928_2443# a_8883_2456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X140 a_8882_4662# a_8878_4839# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X141 a_1514_1516# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X142 a_2888_3208# a_3872_3505# a_3823_3695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X143 a_116_8621# a_644_8416# a_852_8416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 a_646_7867# a_433_7867# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X145 a_117_6645# a_117_6415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X146 gnd d0 a_4078_7917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X147 a_7943_4352# a_8196_4339# a_7803_3841# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X148 a_2883_5591# a_3140_5401# a_2742_6183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X149 a_117_7061# a_645_7313# a_853_7313# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X150 a_7802_6047# a_7987_6545# a_7938_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X151 a_3820_6450# a_3826_5724# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X152 a_118_4209# a_646_4004# a_854_4004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 a_648_3455# a_435_3455# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 a_2741_8389# a_2931_7607# a_2886_7620# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X155 a_5491_2393# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X156 gnd a_3139_6504# a_2931_6504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X157 gnd d2 a_2999_5993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X158 a_6951_177# a_6738_177# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X159 a_5176_1400# a_5176_1171# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X160 a_5173_7559# a_5173_7102# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X161 a_2885_1179# a_3142_989# a_2744_1771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X162 a_7938_7838# a_8925_7404# a_8880_7417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X163 a_8880_1530# a_8883_799# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X164 vdd d0 a_9135_1889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X165 a_7804_1635# a_7989_2133# a_7940_2323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_119_2649# a_647_2901# a_855_2901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X167 a_1481_4844# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X168 a_7060_177# a_7879_4912# a_7834_4925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X169 a_118_5958# a_118_5771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X170 vdd a_3031_4871# a_2823_4871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X171 a_7943_4352# a_8927_4649# a_8878_4839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X172 a_6849_4355# a_6782_3763# a_6866_2792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 gnd a_3141_2092# a_2933_2092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X174 a_7802_6047# a_7987_6545# a_7942_6558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X175 a_5703_4599# a_5490_4599# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X176 a_5176_941# a_5178_842# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X177 a_6570_1557# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X178 a_5908_8457# a_5487_8457# a_5172_8662# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X179 a_2772_7273# a_2791_5993# a_2746_6006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X180 a_2743_3977# a_3000_3787# a_2778_2684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X181 a_7940_3426# a_8927_2992# a_8882_3005# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X182 a_118_4439# a_647_4558# a_855_4558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X183 a_6847_8767# a_6426_8767# a_5908_8457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X184 gnd d0 a_9134_7958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X185 a_3822_5901# a_3825_5170# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X186 gnd a_4078_7917# a_3870_7917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X187 a_433_7867# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_120_1130# a_120_900# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X189 a_7804_1635# a_7989_2133# a_7944_2146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X190 a_1803_7044# a_1694_7044# a_1808_4963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X191 gnd d2 a_8054_8240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X192 a_6848_7664# a_6427_7664# a_5910_7908# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X193 a_4845_116# a_4632_116# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X194 a_6849_4355# a_6428_4355# a_5910_4045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X195 a_435_3455# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X196 vdd a_9135_1889# a_8927_1889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X197 vdd d2 a_8054_8240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X198 a_5173_6686# a_5702_6805# a_5910_6805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X199 a_2889_1002# a_3873_1299# a_3824_1489# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X200 a_645_8970# a_432_8970# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X201 a_5490_4599# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X202 a_6640_6561# a_6427_6561# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X203 a_854_4004# a_1585_4314# a_1793_4314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X204 a_2774_2861# a_2793_1581# a_2744_1771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X205 a_5175_2503# a_5704_2393# a_5912_2393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 a_5489_7908# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X207 a_118_4855# a_646_5107# a_854_5107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X208 a_6859_4885# a_6750_4885# a_6958_4885# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X209 a_649_1249# a_436_1249# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X210 a_2884_3385# a_3141_3195# a_2743_3977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X211 gnd a_9134_7958# a_8926_7958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X212 a_7803_3841# a_7988_4339# a_7939_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X213 a_6848_6561# a_6781_5969# a_6859_7085# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 a_2742_6183# a_2932_5401# a_2887_5414# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X215 gnd a_3140_4298# a_2932_4298# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X216 a_8875_8697# a_9132_8507# a_7937_8941# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X217 gnd a_8054_8240# a_7846_8240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X218 a_1792_7623# a_1371_7623# a_853_7313# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X219 a_8877_5388# a_8882_4662# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X220 a_2778_2684# a_3031_2671# a_2774_5061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X221 a_2744_1771# a_2934_989# a_2889_1002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X222 a_6850_2149# a_6783_1557# a_6861_2673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X223 a_2774_2861# a_2793_1581# a_2748_1594# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X224 a_5488_7354# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X225 gnd a_4080_3505# a_3872_3505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X226 a_5175_3606# a_5175_3377# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X227 a_1794_3211# a_1373_3211# a_855_2901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X228 a_5173_6456# a_5174_5999# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X229 vdd a_8054_8240# a_7846_8240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X230 a_432_8970# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X231 a_2774_2861# a_3031_2671# a_2774_5061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X232 a_118_4855# a_118_4668# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X233 vdd d1 a_8195_7648# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X234 gnd d2 a_8055_6034# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X235 a_5704_736# a_5491_736# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X236 vdd a_3139_7607# a_2931_7607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X237 a_1808_4963# a_1481_7044# a_1808_7163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X238 a_6849_5458# a_6428_5458# a_5911_5702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X239 a_436_1249# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_5703_1839# a_5490_1839# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X241 a_3822_4798# a_3825_4067# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X242 a_119_2003# a_647_1798# a_855_1798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X243 a_3827_2415# a_4080_2402# a_2888_2105# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X244 a_853_6210# a_1584_6520# a_1792_6520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X245 a_2778_2684# a_2792_3787# a_2743_3977# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 gnd d0 a_4077_9020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 a_645_8970# a_432_8970# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 vdd d2 a_8055_6034# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X249 a_5174_4480# a_5703_4599# a_5911_4599# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X250 a_5172_8892# a_5172_8662# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X251 a_6537_7085# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X252 a_2886_6517# a_3870_6814# a_3821_7004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X253 a_855_1798# a_1586_2108# a_1794_2108# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X254 a_6850_3252# a_6429_3252# a_5911_2942# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X255 a_8879_8520# a_8875_8697# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X256 a_2741_8389# a_2998_8199# a_2776_7096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X257 a_6641_4355# a_6428_4355# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X258 a_5912_2393# a_5491_2393# a_5175_2274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X259 a_8876_6491# a_9133_6301# a_7938_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X260 a_6958_4885# a_6537_4885# a_6864_5004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X261 a_2743_3977# a_2933_3195# a_2888_3208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X262 vdd d0 a_4077_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X263 a_1726_3722# a_1513_3722# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X264 a_7937_8941# a_8924_8507# a_8879_8520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X265 a_5910_7908# a_5489_7908# a_5173_8018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X266 vdd a_8195_7648# a_7987_7648# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X267 gnd a_8055_6034# a_7847_6034# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X268 a_6859_7085# a_6568_5969# a_6849_5458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X269 a_1793_5417# a_1372_5417# a_854_5107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X270 a_5490_1839# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X271 gnd d1 a_8196_5442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_2774_5061# a_2823_2671# a_2774_2861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X273 gnd a_4081_1299# a_3873_1299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 a_5489_5148# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 a_1795_1005# a_1374_1005# a_856_695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X276 gnd d0 a_9133_9061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X277 a_3822_2038# a_4079_1848# a_2884_2282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X278 gnd a_4077_9020# a_3869_9020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X279 a_432_8970# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 a_8881_6868# a_8877_7045# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X281 vdd a_8055_6034# a_7847_6034# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X282 a_8877_4285# a_8883_3559# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X283 gnd d1 a_8198_1030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X284 gnd d2 a_8056_3828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 vdd d1 a_8196_5442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X286 a_2774_5061# a_2823_2671# a_2778_2684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X287 vdd a_3140_5401# a_2932_5401# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X288 gnd d4 a_3031_4871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X289 a_6782_3763# a_6569_3763# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X290 a_5175_2503# a_5175_2274# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X291 a_7834_2725# a_8087_2712# a_7830_5102# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X292 vdd d0 a_9133_9061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X293 a_3819_8656# a_3825_7930# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X294 vdd a_4077_9020# a_3869_9020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X295 a_1791_8726# a_1724_8134# a_1808_7163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_2883_5591# a_3870_5157# a_3825_5170# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X297 a_1513_3722# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X298 vdd d1 a_8198_1030# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X299 a_2888_2105# a_3872_2402# a_3823_2592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X300 a_646_6764# a_433_6764# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X301 gnd d0 a_4078_6814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X302 a_5911_4599# a_5490_4599# a_5174_4480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X303 gnd d3 a_8085_7124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X304 gnd a_8196_5442# a_7988_5442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X305 a_6851_1046# a_6430_1046# a_5912_736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X306 a_6642_2149# a_6429_2149# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X307 a_7830_2902# a_8087_2712# a_7830_5102# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X308 a_119_3106# a_647_2901# a_855_2901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X309 a_5488_9011# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X310 a_2742_6183# a_2999_5993# a_2772_7273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X311 a_647_5661# a_434_5661# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X312 a_2883_4488# a_3140_4298# a_2747_3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X313 vdd a_3000_3787# a_2792_3787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X314 a_648_2352# a_435_2352# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X315 gnd a_9133_9061# a_8925_9061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X316 gnd a_8198_1030# a_7990_1030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X317 a_3821_8107# a_3824_7376# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X318 gnd d1 a_8195_7648# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X319 a_8877_4285# a_9134_4095# a_7939_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X320 a_8884_1353# a_8880_1530# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X321 a_1727_1516# a_1514_1516# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X322 vdd a_8196_5442# a_7988_5442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X323 a_8881_4108# a_8877_4285# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X324 gnd a_8056_3828# a_7848_3828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 a_119_3336# a_119_3106# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X326 vdd d3 a_8085_7124# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X327 a_7938_6735# a_8925_6301# a_8880_6314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X328 a_5175_2044# a_5703_1839# a_5911_1839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X329 a_6567_8175# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X330 a_7060_177# a_6951_177# a_4954_116# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X331 gnd d1 a_8197_3236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X332 vdd a_9133_9061# a_8925_9061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X333 a_3823_8479# a_3819_8656# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X334 vdd a_8198_1030# a_7990_1030# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X335 gnd d0 a_9134_6855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_433_6764# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 a_856_695# a_435_695# a_120_900# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X338 a_2884_3385# a_3871_2951# a_3822_3141# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X339 a_645_7313# a_432_7313# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 gnd a_4078_6814# a_3870_6814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X341 a_1810_2751# a_1696_2632# a_1803_4844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X342 a_5910_5148# a_5489_5148# a_5174_4896# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X343 a_5173_7102# a_5173_6915# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X344 a_2103_136# a_1682_136# a_1902_4844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X345 vdd d1 a_8197_3236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X346 a_2745_8212# a_2930_8710# a_2881_8900# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X347 a_6848_6561# a_6427_6561# a_5910_6805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X348 a_434_5661# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X349 a_435_2352# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X350 vdd a_3141_3195# a_2933_3195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X351 a_2887_4311# a_3871_4608# a_3822_4798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X352 vdd d0 a_4078_5157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X353 a_6783_1557# a_6570_1557# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X354 gnd a_8195_7648# a_7987_7648# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_1514_1516# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X356 a_7830_5102# a_7879_2712# a_7830_2902# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X357 a_646_7867# a_433_7867# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X358 a_5489_7908# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X359 a_117_8164# a_644_8416# a_852_8416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X360 a_1808_7163# a_1511_8134# a_1792_7623# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X361 a_647_4558# a_434_4558# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X362 gnd a_3031_2671# a_2823_2671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X363 a_2745_8212# a_2930_8710# a_2885_8723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X364 gnd a_8197_3236# a_7989_3236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_648_3455# a_435_3455# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X366 a_122_801# a_648_695# a_856_695# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X367 a_2884_2282# a_3141_2092# a_2748_1594# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X368 a_119_3752# a_646_4004# a_854_4004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X369 gnd a_9134_6855# a_8926_6855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X370 a_2747_3800# a_2932_4298# a_2887_4311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X371 a_7830_5102# a_7879_2712# a_7834_2725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X372 vref a_116_9080# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X373 a_432_7313# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X374 a_5911_5702# a_5490_5702# a_5174_5583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 vdd a_3031_2671# a_2823_2671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X376 a_2886_7620# a_3870_7917# a_3825_7930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X377 a_7939_4529# a_8926_4095# a_8881_4108# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X378 vdd a_8197_3236# a_7989_3236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X379 gnd d0 a_4077_7363# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X380 a_1792_6520# a_1371_6520# a_853_6210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X381 a_6850_3252# a_6782_3763# a_6866_2792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X382 a_435_695# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X383 a_3824_1489# a_4081_1299# a_2889_1002# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X384 a_2883_5591# a_3870_5157# a_3821_5347# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X385 vdd a_4078_5157# a_3870_5157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X386 a_6570_1557# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X387 a_2885_1179# a_3872_745# a_3823_935# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 gnd a_4080_2402# a_3872_2402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 a_3821_7004# a_3824_6273# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X390 a_5488_6251# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X391 a_6847_8767# a_6426_8767# a_5909_9011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X392 a_433_7867# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X393 a_434_4558# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X394 a_1682_136# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X395 a_2103_136# a_4845_116# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X396 a_119_2233# a_119_2003# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X397 vdd d0 a_4077_7363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X398 a_646_5107# a_433_5107# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X399 a_648_695# a_435_695# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X400 gnd d1 a_3138_8710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_8880_7417# a_8876_7594# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X402 a_4845_116# a_4632_116# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X403 a_6849_4355# a_6428_4355# a_5911_4599# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X404 a_435_3455# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X405 a_1803_4844# a_1483_2632# a_1805_2632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X406 a_2885_1179# a_3872_745# a_3827_758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X407 gnd a_8087_4912# a_7879_4912# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X408 a_5175_3147# a_5175_2690# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X409 gnd d0 a_9133_7404# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 vdd d1 a_3138_8710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X411 gnd a_4077_7363# a_3869_7363# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X412 a_118_5958# a_645_6210# a_853_6210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X413 a_2887_5414# a_3871_5711# a_3822_5901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X414 a_120_1546# a_120_1359# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X415 a_2746_6006# a_2931_6504# a_2886_6517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X416 a_5910_7908# a_5489_7908# a_5173_7789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 gnd d0 a_9135_2992# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X418 a_649_1249# a_436_1249# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X419 gnd a_4079_2951# a_3871_2951# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X420 a_1791_8726# a_1370_8726# a_852_8416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X421 a_3824_1489# a_3827_758# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X422 a_3823_3695# a_4080_3505# a_2888_3208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X423 a_2748_1594# a_2933_2092# a_2888_2105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X424 gnd d1 a_8194_8751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X425 vdd d0 a_4078_7917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X426 vdd a_4077_7363# a_3869_7363# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X427 a_433_5107# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_6859_4885# a_6539_2673# a_6861_2673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X429 gnd a_3138_8710# a_2930_8710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X430 a_2776_7096# a_3029_7083# a_2778_4884# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 a_2887_5414# a_3871_5711# a_3826_5724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X432 a_5487_8457# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_1792_7623# a_1371_7623# a_854_7867# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X434 gnd a_4079_4608# a_3871_4608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X435 a_1793_4314# a_1372_4314# a_854_4004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X436 gnd d0 a_4078_5157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X437 a_6738_177# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X438 a_6851_1046# a_6783_1557# a_6861_2673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X439 a_2889_1002# a_3873_1299# a_3828_1312# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X440 a_2886_7620# a_3139_7607# a_2741_8389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 a_5488_7354# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X442 a_5489_4045# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X443 a_1794_3211# a_1373_3211# a_856_3455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X444 vdd d1 a_8194_8751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X445 gnd a_9133_7404# a_8925_7404# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X446 vdd a_3138_8710# a_2930_8710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X447 a_2772_7273# a_3029_7083# a_2778_4884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X448 a_6427_7664# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X449 vdd d1 a_8196_4339# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X450 gnd a_9135_2992# a_8927_2992# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X451 vdd a_3140_4298# a_2932_4298# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X452 a_436_1249# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X453 a_116_8621# a_117_8164# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X454 vdd d0 a_9134_7958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X455 gnd d1 a_3140_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X456 a_5703_1839# a_5490_1839# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X457 a_6429_3252# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X458 gnd a_8194_8751# a_7986_8751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X459 vdd a_4078_7917# a_3870_7917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X460 gnd a_8876_9251# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X461 gnd d0 a_9134_5198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X462 a_8883_3559# a_8879_3736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X463 a_8880_6314# a_8876_6491# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X464 gnd a_4078_5157# a_3870_5157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X465 a_1694_7044# a_1481_7044# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X466 gnd d0 a_4080_3505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X467 a_6850_3252# a_6429_3252# a_5912_3496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X468 vdd a_8194_8751# a_7986_8751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X469 a_3821_5347# a_3826_4621# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X470 gnd d1 a_8195_6545# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X471 a_855_1798# a_434_1798# a_119_2003# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X472 a_1793_5417# a_1372_5417# a_855_5661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X473 vdd a_8196_4339# a_7988_4339# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X474 a_2888_3208# a_3872_3505# a_3827_3518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X475 a_1794_2108# a_1373_2108# a_855_1798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 vdd a_9134_7958# a_8926_7958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X477 a_5490_1839# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X478 gnd d3 a_3029_7083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 vdd d4 a_8087_4912# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X480 a_2778_2684# a_2792_3787# a_2747_3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X481 gnd d1 a_8197_2133# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X482 vdd d1 a_8195_6545# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X483 gnd d0 a_9135_5752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X484 a_5489_5148# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X485 gnd a_9134_5198# a_8926_5198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X486 a_1795_1005# a_1374_1005# a_857_1249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X487 a_5176_1171# a_5176_941# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X488 a_7800_1812# a_7990_1030# a_7941_1220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X489 a_6750_7085# a_6537_7085# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X490 vdd d2 a_2999_5993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X491 gnd a_4079_5711# a_3871_5711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X492 vdd a_3139_6504# a_2931_6504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X493 a_645_6210# a_432_6210# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_6428_5458# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X495 a_5705_1290# a_5492_1290# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 gnd d1 a_3139_7607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X497 a_1481_7044# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X498 a_5174_4480# a_5174_4250# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X499 a_5910_4045# a_5489_4045# a_5175_3793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X500 gnd d0 a_9137_1340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 vdd d3 a_3029_7083# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X502 vdd d1 a_8197_2133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X503 vdd a_3141_2092# a_2933_2092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X504 vdd d0 a_9135_5752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X505 a_7800_1812# a_7990_1030# a_7945_1043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X506 a_5911_2942# a_5490_2942# a_5175_3147# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X507 gnd d1 a_3141_3195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X508 gnd a_8195_6545# a_7987_6545# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X509 vdd a_4079_5711# a_3871_5711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X510 a_3825_5170# a_3821_5347# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X511 a_1792_7623# a_1724_8134# a_1808_7163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X512 a_6850_2149# a_6429_2149# a_5911_1839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X513 a_5489_6805# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X514 a_855_5661# a_434_5661# a_118_5542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X515 a_3827_2415# a_3823_2592# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X516 a_646_6764# a_433_6764# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X517 vdd d0 a_9137_1340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X518 vdd a_4081_1299# a_3873_1299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X519 gnd a_8197_2133# a_7989_2133# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X520 a_6851_1046# a_6430_1046# a_5913_1290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X521 gnd d0 a_4081_1299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X522 vdd a_8195_6545# a_7987_6545# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X523 gnd a_9135_5752# a_8927_5752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X524 a_648_2352# a_435_2352# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X525 gnd d2 a_3001_1581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X526 a_432_6210# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_5492_1290# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_8883_2456# a_8879_2633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X529 gnd d1 a_8196_4339# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X530 a_116_9080# a_116_8851# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X531 a_3824_9033# a_3820_9210# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X532 a_1808_4963# a_1694_4844# a_1902_4844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X533 gnd a_9137_1340# a_8929_1340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X534 vdd a_8197_2133# a_7989_2133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X535 a_5176_1587# a_5703_1839# a_5911_1839# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X536 a_6567_8175# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X537 gnd d0 a_4077_6260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 vdd a_9135_5752# a_8927_5752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X539 a_2883_4488# a_3870_4054# a_3821_4244# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X540 a_5704_3496# a_5491_3496# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X541 a_644_8416# a_431_8416# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 a_3825_6827# a_3821_7004# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X543 vdd d2 a_3001_1581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X544 gnd d0 a_9136_3546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X545 a_5912_736# a_5491_736# a_5178_842# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X546 a_5491_736# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X547 a_433_6764# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X548 a_5174_5353# a_5174_4896# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X549 vdd a_9137_1340# a_8929_1340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X550 a_645_7313# a_432_7313# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X551 a_646_4004# a_433_4004# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 a_1805_2632# a_1696_2632# a_1803_4844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X553 vdd d0 a_4077_6260# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X554 a_5910_5148# a_5489_5148# a_5174_5353# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X555 a_2883_4488# a_3870_4054# a_3825_4067# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X556 gnd a_4080_745# a_3872_745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_435_2352# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X558 a_854_7867# a_433_7867# a_117_7748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 vdd d0 a_9136_3546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X560 gnd d1 a_3142_989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_647_2901# a_434_2901# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X562 a_853_8970# a_1583_8726# a_1791_8726# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_1793_5417# a_1725_5928# a_1803_7044# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X564 gnd a_8196_4339# a_7988_4339# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X565 vdd a_4080_3505# a_3872_3505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X566 a_3823_3695# a_3826_2964# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X567 gnd d0 a_9133_6301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X568 vdd d2 a_8056_3828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X569 a_1808_7163# a_1511_8134# a_1791_8726# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X570 a_647_4558# a_434_4558# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X571 a_856_3455# a_435_3455# a_119_3336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X572 gnd a_4077_6260# a_3869_6260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X573 gnd d2 a_3000_3787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X574 vdd a_4080_745# a_3872_745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X575 a_5173_7789# a_5173_7559# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X576 a_5491_3496# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X577 a_431_8416# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X578 a_6864_7204# a_6750_7085# a_6864_5004# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_5910_6805# a_5489_6805# a_5173_6686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X580 a_3825_4067# a_3821_4244# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X581 gnd a_9136_3546# a_8928_3546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X582 a_5175_3377# a_5704_3496# a_5912_3496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X583 gnd d0 a_4076_8466# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X584 a_432_7313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X585 vdd a_4077_6260# a_3869_6260# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X586 a_5911_5702# a_5490_5702# a_5174_5812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X587 a_433_4004# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X588 a_3823_2592# a_4080_2402# a_2888_2105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X589 a_3826_5724# a_3822_5901# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X590 a_2887_4311# a_3871_4608# a_3826_4621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X591 a_5175_2690# a_5175_2503# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X592 a_6568_5969# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X593 gnd d0 a_4078_4054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X594 a_1902_4844# a_1481_4844# a_1803_4844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X595 vdd a_9136_3546# a_8928_3546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X596 gnd a_3142_989# a_2934_989# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X597 a_434_2901# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X598 a_2884_2282# a_3871_1848# a_3822_2038# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X599 vdd d0 a_4076_8466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X600 a_8881_7971# a_8877_8148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X601 a_2886_6517# a_3139_6504# a_2746_6006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X602 a_5488_6251# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X603 gnd a_8085_7124# a_7877_7124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X604 gnd a_9133_6301# a_8925_6301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X605 vdd a_8056_3828# a_7848_3828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X606 a_5701_9011# a_5488_9011# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X607 a_434_4558# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X608 a_1682_136# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X609 a_6427_6561# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X610 a_646_5107# a_433_5107# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X611 a_4954_116# a_4845_116# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X612 vdd d0 a_4078_4054# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X613 gnd d2 a_8057_1622# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X614 a_1803_4844# a_1483_2632# a_1810_2751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X615 a_3824_9033# a_5172_9121# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X616 gnd d0 a_9132_8507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X617 a_853_8970# a_432_8970# a_116_9080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X618 gnd a_4076_8466# a_3868_8466# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X619 vdd a_8085_7124# a_7877_7124# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X620 a_6639_8767# a_6426_8767# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X621 a_3825_7930# a_4078_7917# a_2886_7620# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X622 gnd d0 a_9134_4095# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X623 a_857_1249# a_436_1249# a_120_1130# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X624 vdd d2 a_8057_1622# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X625 a_1803_7044# a_1512_5928# a_1792_6520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X626 gnd a_4078_4054# a_3870_4054# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_6539_2673# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X628 gnd d0 a_4080_2402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X629 vdd a_4076_8466# a_3868_8466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X630 a_2886_6517# a_3870_6814# a_3825_6827# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X631 a_118_5312# a_118_4855# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X632 a_1791_8726# a_1370_8726# a_853_8970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X633 gnd a_9136_786# a_8928_786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_5176_1171# a_5705_1290# a_5913_1290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X635 a_8878_2079# a_9135_1889# a_7940_2323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X636 a_119_2462# a_119_2233# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X637 a_6864_5004# a_6537_7085# a_6859_7085# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X638 a_433_5107# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X639 vdd a_4078_4054# a_3870_4054# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X640 a_5912_3496# a_5491_3496# a_5175_3606# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X641 gnd a_8057_1622# a_7849_1622# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X642 a_6859_4885# a_6539_2673# a_6866_2792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X643 a_2888_2105# a_3872_2402# a_3827_2415# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X644 a_8882_3005# a_8878_3182# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X645 a_5487_8457# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X646 a_5173_6686# a_5173_6456# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X647 a_1793_4314# a_1372_4314# a_855_4558# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X648 a_647_1798# a_434_1798# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X649 gnd a_9132_8507# a_8924_8507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X650 a_6738_177# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X651 a_8881_7971# a_9134_7958# a_7942_7661# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X652 a_6426_8767# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_3827_758# a_4080_745# a_2885_1179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X654 vdd a_9136_786# a_8928_786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X655 a_5489_4045# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X656 a_7801_8253# a_8054_8240# a_7832_7137# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X657 a_3824_7376# a_3820_7553# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X658 gnd a_9134_4095# a_8926_4095# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X659 a_1902_4844# a_1895_136# a_2103_136# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X660 vdd a_8057_1622# a_7849_1622# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X661 a_1584_7623# a_1371_7623# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 a_6427_7664# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X663 gnd d1 a_3139_6504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_3826_4621# a_3822_4798# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X665 a_6428_4355# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X666 a_5911_2942# a_5490_2942# a_5175_2690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X667 gnd d0 a_4079_2951# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X668 a_5174_5999# a_5174_5812# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X669 a_3823_935# a_4080_745# a_2885_1179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X670 a_6429_3252# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X671 a_1586_3211# a_1373_3211# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_853_8970# a_432_8970# a_116_8851# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X673 vdd d0 a_9135_4649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X674 gnd d1 a_3141_2092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_7797_8430# a_8054_8240# a_7832_7137# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X676 vdd d4 a_3031_4871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X677 a_1793_4314# a_1726_3722# a_1810_2751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X678 gnd d0 a_4079_4608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 vdd a_4079_4608# a_3871_4608# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X680 gnd d0 a_9135_1889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X681 a_434_1798# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X682 a_2882_7797# a_3139_7607# a_2741_8389# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X683 a_1694_7044# a_1481_7044# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X684 gnd a_4079_1848# a_3871_1848# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X685 gnd d3 a_8087_2712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X686 vdd d0 a_4078_6814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X687 a_5172_9121# a_5701_9011# a_5909_9011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X688 a_1792_6520# a_1371_6520# a_854_6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X689 a_1371_7623# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 a_117_8164# a_117_7977# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X691 a_5913_1290# a_5492_1290# a_5176_1400# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X692 a_7940_2323# a_8927_1889# a_8882_1902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X693 vdd d3 a_8087_2712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X694 a_6569_3763# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X695 a_1794_2108# a_1373_2108# a_856_2352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X696 a_1373_3211# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X697 vdd a_9135_4649# a_8927_4649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X698 a_118_4209# a_119_3752# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X699 vdd d0 a_9134_5198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X700 a_5704_2393# a_5491_2393# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_7942_7661# a_8926_7958# a_8877_8148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X702 a_4954_116# a_6738_177# a_7060_177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 gnd a_9135_1889# a_8927_1889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X704 gnd d0 a_9136_2443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X705 a_5702_7908# a_5489_7908# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X706 a_7802_6047# a_8055_6034# a_7828_7314# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X707 a_4632_116# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 a_119_2003# a_120_1546# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X709 a_647_2901# a_434_2901# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X710 a_1481_7044# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X711 a_118_5771# a_118_5542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X712 a_1585_5417# a_1372_5417# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X713 a_6428_5458# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X714 a_8882_1902# a_8878_2079# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X715 a_6429_2149# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X716 a_7832_7137# a_7846_8240# a_7797_8430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X717 vdd d0 a_9134_6855# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X718 gnd d1 a_3140_4298# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X719 a_5910_4045# a_5489_4045# a_5174_4250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X720 a_2884_3385# a_3871_2951# a_3826_2964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X721 vdd a_4078_6814# a_3870_6814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X722 a_1792_6520# a_1725_5928# a_1803_7044# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X723 a_854_6764# a_433_6764# a_117_6645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X724 a_1587_1005# a_1374_1005# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 vdd d0 a_9136_2443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X726 a_3824_6273# a_3820_6450# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X727 a_7798_6224# a_8055_6034# a_7828_7314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X728 a_8879_976# a_5178_842# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X729 a_1794_2108# a_1727_1516# a_1805_2632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 vdd a_4080_2402# a_3872_2402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X731 a_3824_9033# a_4077_9020# a_2885_8723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X732 a_6850_2149# a_6429_2149# a_5912_2393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X733 a_7832_7137# a_7846_8240# a_7801_8253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X734 a_5701_7354# a_5488_7354# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X735 a_5489_6805# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X736 a_855_5661# a_434_5661# a_118_5771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X737 a_1810_2751# a_1513_3722# a_1794_3211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 a_5176_1587# a_5176_1400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X739 a_856_2352# a_435_2352# a_119_2233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 vdd a_9134_5198# a_8926_5198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X741 a_5174_4896# a_5174_4709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X742 a_5491_2393# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X743 a_3820_9210# a_4077_9020# a_2885_8723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X744 gnd d0 a_4079_5711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X745 gnd a_9136_2443# a_8928_2443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X746 vdd d1 a_3139_7607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X747 a_6568_5969# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X748 a_5175_2274# a_5704_2393# a_5912_2393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X749 a_434_2901# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X750 a_5909_9011# a_5488_9011# a_5172_8892# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_1372_5417# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X752 vdd a_9134_6855# a_8926_6855# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X753 a_5703_4599# a_5490_4599# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X754 vdd d0 a_9133_7404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X755 a_1803_4844# a_1694_4844# a_1902_4844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X756 gnd d0 a_9135_4649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X757 a_1374_1005# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X758 gnd a_9133_9061# a_7941_8764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X759 a_853_7313# a_432_7313# a_117_7061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X760 vdd d0 a_4079_5711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X761 vdd a_9136_2443# a_8928_2443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X762 a_644_8416# a_431_8416# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X763 vdd d0 a_9135_2992# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X764 a_6866_2792# a_6569_3763# a_6850_3252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X765 a_5491_736# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X766 a_5912_736# a_5491_736# a_5176_941# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X767 a_8883_799# a_8879_976# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X768 a_7803_3841# a_8056_3828# a_7834_2725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X769 vdd d0 a_4081_1299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X770 a_2778_4884# a_3031_4871# a_2004_136# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X771 a_646_4004# a_433_4004# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X772 a_7828_7314# a_7847_6034# a_7798_6224# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 a_8876_9251# a_9133_9061# a_7941_8764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X774 a_5910_7908# a_6640_7664# a_6848_7664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 gnd a_2999_5993# a_2791_5993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_854_7867# a_433_7867# a_117_7977# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X777 a_8878_5942# a_8881_5211# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X778 a_852_8416# a_1583_8726# a_1791_8726# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X779 a_1803_7044# a_1512_5928# a_1793_5417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X780 a_855_4558# a_434_4558# a_118_4439# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X781 a_117_7518# a_117_7061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X782 a_8876_9251# a_8879_8520# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X783 a_3825_6827# a_4078_6814# a_2886_6517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X784 a_5490_4599# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X785 a_5912_3496# a_6642_3252# a_6850_3252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 vdd a_9133_7404# a_8925_7404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X787 a_7828_7314# a_7847_6034# a_7802_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X788 a_5702_5148# a_5489_5148# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 vdd a_8087_4912# a_7879_4912# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X790 a_118_4668# a_118_4439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X791 a_856_3455# a_435_3455# a_119_3565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X792 a_2885_8723# a_3869_9020# a_3820_9210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X793 gnd d2 a_2998_8199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X794 gnd a_9135_4649# a_8927_4649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 a_1805_2632# a_1514_1516# a_1795_1005# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X796 a_120_1546# a_647_1798# a_855_1798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X797 a_8881_5211# a_8877_5388# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X798 a_431_8416# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X799 a_6537_7085# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X800 a_5910_6805# a_5489_6805# a_5173_6915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X801 vdd a_9135_2992# a_8927_2992# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X802 a_5173_7789# a_5702_7908# a_5910_7908# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X803 vdd d1 a_3140_5401# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X804 vdd a_4079_2951# a_3871_2951# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X805 a_2885_8723# a_3869_9020# a_3824_9033# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X806 a_1724_8134# a_1511_8134# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 a_433_4004# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X808 a_5912_2393# a_5491_2393# a_5175_2503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X809 vdd d1 a_3142_989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X810 a_8878_3182# a_8883_2456# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X811 a_854_5107# a_433_5107# a_118_4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X812 a_1902_4844# a_1481_4844# a_1808_4963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X813 vdd d0 a_4080_3505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X814 a_8881_6868# a_9134_6855# a_7942_6558# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X815 a_645_6210# a_432_6210# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X816 a_5173_7559# a_5701_7354# a_5909_7354# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_5176_941# a_5704_736# a_5912_736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X818 a_6861_2673# a_6570_1557# a_6851_1046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X819 a_7941_8764# a_8925_9061# a_8876_9251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X820 a_5703_5702# a_5490_5702# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X821 vdd d2 a_3000_3787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X822 a_5701_9011# a_5488_9011# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X823 gnd a_2998_8199# a_2790_8199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X824 a_118_5771# a_647_5661# a_855_5661# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X825 a_1584_6520# a_1371_6520# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X826 a_6427_6561# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X827 a_6537_4885# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X828 a_7834_2725# a_7848_3828# a_7799_4018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X829 a_5175_3377# a_5175_3147# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X830 a_5911_5702# a_6641_5458# a_6849_5458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X831 a_3821_5347# a_4078_5157# a_2883_5591# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X832 a_2004_136# a_2823_4871# a_2774_5061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 a_7941_8764# a_8925_9061# gnd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X834 a_6639_8767# a_6426_8767# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X835 a_6780_8175# a_6567_8175# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X836 a_5174_4709# a_5703_4599# a_5911_4599# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 a_1511_8134# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X838 a_5913_1290# a_6643_1046# a_6851_1046# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 vdd a_3142_989# a_2934_989# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X840 a_3828_1312# a_3824_1489# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X841 a_857_1249# a_436_1249# a_120_1359# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X842 a_1696_2632# a_1483_2632# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X843 a_6539_2673# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X844 a_432_6210# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X845 a_8878_4839# a_8881_4108# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X846 a_117_6415# a_118_5958# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X847 a_7834_4925# a_8087_4912# a_7060_177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X848 a_5911_4599# a_5490_4599# a_5174_4709# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X849 a_5490_5702# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X850 vdd d1 a_3141_3195# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X851 a_3824_7376# a_4077_7363# a_2882_7797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X852 a_1371_6520# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 vdd d0 a_9132_8507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X854 a_117_7977# a_117_7748# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X855 a_3825_7930# a_3821_8107# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X856 a_5702_7908# a_5489_7908# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 gnd d3 a_3031_2671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_3826_2964# a_4079_2951# a_2884_3385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X859 a_1583_8726# a_1370_8726# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 a_6426_8767# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X861 a_117_7977# a_646_7867# a_854_7867# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X862 a_5174_5353# a_5702_5148# a_5910_5148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 a_3820_7553# a_4077_7363# a_2882_7797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X864 a_7942_6558# a_8926_6855# a_8877_7045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X865 a_6752_2673# a_6539_2673# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X866 a_2885_8723# a_3138_8710# a_2745_8212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_5909_7354# a_5488_7354# a_5173_7102# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X868 a_2004_136# a_1895_136# a_2103_136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X869 a_116_8851# a_116_8621# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X870 a_1584_7623# a_1371_7623# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X871 a_3826_4621# a_4079_4608# a_2887_4311# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X872 a_1585_4314# a_1372_4314# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 a_6428_4355# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X874 a_119_3565# a_648_3455# a_856_3455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X875 a_1483_2632# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X876 a_8878_2079# a_8884_1353# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X877 a_2884_2282# a_3871_1848# a_3826_1861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X878 vdd d3 a_3031_2671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X879 a_1586_3211# a_1373_3211# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X880 a_8880_7417# a_9133_7404# a_7938_7838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X881 a_2881_8900# a_3138_8710# a_2745_8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X882 a_1794_3211# a_1726_3722# a_1810_2751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X883 vdd a_9132_8507# a_8924_8507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X884 a_5701_6251# a_5488_6251# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X885 a_5175_2274# a_5175_2044# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X886 a_8882_3005# a_9135_2992# a_7940_3426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 a_854_7867# a_1584_7623# a_1792_7623# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X888 a_1370_8726# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X889 a_5172_8892# a_5701_9011# a_5909_9011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X890 a_5174_5812# a_5703_5702# a_5911_5702# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 a_3821_8107# a_4078_7917# a_2886_7620# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X892 a_3826_2964# a_3822_3141# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X893 a_856_3455# a_1586_3211# a_1794_3211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_1371_7623# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X895 a_7060_177# a_7879_4912# a_7830_5102# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X896 a_1372_4314# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X897 a_3825_5170# a_4078_5157# a_2883_5591# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X898 gnd a_3031_4871# a_2823_4871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 vdd d0 a_9133_6301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X900 a_6847_8767# a_6780_8175# a_6864_7204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X901 a_2882_7797# a_3869_7363# a_3820_7553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X902 a_6569_3763# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X903 a_1373_3211# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X904 a_853_6210# a_432_6210# a_118_5958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X905 vdd d0 a_4079_4608# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X906 a_856_695# a_435_695# a_122_801# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X907 a_116_8851# a_645_8970# a_853_8970# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X908 a_8877_8148# a_8880_7417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X909 a_5911_1839# a_5490_1839# a_5176_1587# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 a_435_695# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X911 a_4632_116# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X912 a_4954_116# a_6738_177# a_6958_4885# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X913 gnd d0 a_4079_1848# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X914 a_2882_7797# a_3869_7363# a_3824_7376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X915 a_117_6874# a_117_6645# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X916 a_1585_5417# a_1372_5417# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X917 a_120_1359# a_649_1249# a_857_1249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X918 a_6429_2149# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X919 a_1586_2108# a_1373_2108# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X920 a_8877_8148# a_9134_7958# a_7942_7661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X921 a_2887_5414# a_3140_5401# a_2742_6183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 a_5910_6805# a_6640_6561# a_6848_6561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 a_5700_8457# a_5487_8457# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X924 a_5173_8205# a_5173_8018# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X925 a_854_6764# a_433_6764# a_117_6874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X926 a_8881_5211# a_9134_5198# a_7939_5632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X927 a_1587_1005# a_1374_1005# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X928 a_3826_5724# a_4079_5711# a_2887_5414# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X929 a_2882_6694# a_3139_6504# a_2746_6006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X930 a_1795_1005# a_1727_1516# a_1805_2632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X931 a_5173_8018# a_5702_7908# a_5910_7908# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X932 a_5701_7354# a_5488_7354# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X933 a_7938_7838# a_8925_7404# a_8876_7594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X934 a_8876_7594# a_8881_6868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X935 vdd a_9133_6301# a_8925_6301# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X936 a_5702_4045# a_5489_4045# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X937 a_1810_2751# a_1513_3722# a_1793_4314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X938 a_120_900# a_648_695# a_856_695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X939 a_856_2352# a_435_2352# a_119_2462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X940 a_6640_7664# a_6427_7664# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X941 a_2772_7273# a_2791_5993# a_2742_6183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 a_855_5661# a_1585_5417# a_1793_5417# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X943 a_6866_2792# a_6752_2673# a_6859_4885# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X944 a_7940_3426# a_8927_2992# a_8878_3182# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_5703_2942# a_5490_2942# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X946 a_3822_5901# a_4079_5711# a_2887_5414# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X947 a_5174_5812# a_5174_5583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X948 a_5172_8662# a_5173_8205# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X949 a_5909_9011# a_5488_9011# a_5172_9121# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X950 vdd d1 a_3140_4298# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X951 a_857_1249# a_1587_1005# a_1795_1005# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_6642_3252# a_6429_3252# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X953 a_1372_5417# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X954 a_120_1359# a_120_1130# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X955 vdd a_4079_1848# a_3871_1848# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X956 a_1373_2108# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X957 a_852_8416# a_431_8416# a_117_8164# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X958 a_117_7061# a_117_6874# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X959 vdd d0 a_9134_4095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X960 a_7941_1220# a_8928_786# a_8879_976# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_5174_5583# a_5174_5353# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X962 a_8882_5765# a_9135_5752# a_7943_5455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X963 a_1374_1005# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X964 a_116_9080# a_645_8970# a_853_8970# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_6864_7204# a_6567_8175# a_6848_7664# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X966 a_7938_7838# a_8195_7648# a_7797_8430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X967 a_853_7313# a_432_7313# a_117_7518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X968 a_854_4004# a_433_4004# a_119_3752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X969 vdd d0 a_4080_2402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X970 a_5173_6456# a_5701_6251# a_5909_6251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X971 a_6866_2792# a_6569_3763# a_6849_4355# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X972 a_648_695# a_435_695# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 a_3826_1861# a_3822_2038# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X974 gnd a_8087_2712# a_7879_2712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_5909_9011# a_6639_8767# a_6847_8767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X976 a_8884_1353# a_9137_1340# a_7945_1043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X977 a_7941_1220# a_8928_786# a_8883_799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X978 a_855_2901# a_434_2901# a_119_3106# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X979 a_3827_3518# a_3823_3695# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X980 a_8878_5942# a_9135_5752# a_7943_5455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X981 a_1895_136# a_1682_136# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_5490_2942# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X983 a_2888_3208# a_3141_3195# a_2743_3977# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X984 a_5909_7354# a_6640_7664# a_6848_7664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X985 a_5911_4599# a_6641_4355# a_6849_4355# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X986 vout a_4632_116# a_4954_116# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X987 a_7942_7661# a_8926_7958# a_8881_7971# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X988 a_8877_7045# a_8880_6314# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X989 a_2742_6183# a_2932_5401# a_2883_5591# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X990 a_855_4558# a_434_4558# a_118_4668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X991 vdd a_8087_2712# a_7879_2712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X992 a_8880_1530# a_9137_1340# a_7945_1043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X993 a_2776_7096# a_2790_8199# a_2741_8389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 a_7939_5632# a_8926_5198# a_8877_5388# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_5911_2942# a_6642_3252# a_6850_3252# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X996 a_5702_5148# a_5489_5148# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X997 vdd a_9134_4095# a_8926_4095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X998 a_120_900# a_122_801# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X999 a_1805_2632# a_1514_1516# a_1794_2108# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1000 a_6537_4885# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1001 vdd d1 a_3139_6504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1002 a_6641_5458# a_6428_5458# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1003 a_2748_1594# a_3001_1581# a_2774_2861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1004 a_7943_5455# a_8196_5442# a_7798_6224# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 vdd d1 a_3141_2092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1006 a_8876_6491# a_8882_5765# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1007 a_6643_1046# a_6430_1046# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1008 a_1724_8134# a_1511_8134# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1009 a_3824_6273# a_4077_6260# a_2882_6694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 a_5172_8662# a_5700_8457# a_5908_8457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1011 a_7945_1043# a_8198_1030# a_7800_1812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1012 a_2744_1771# a_3001_1581# a_2774_2861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1013 a_5702_6805# a_5489_6805# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1014 a_8883_3559# a_9136_3546# a_7944_3249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 a_2778_4884# a_2821_7083# a_2772_7273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 a_117_6874# a_646_6764# a_854_6764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1017 a_854_5107# a_433_5107# a_118_5312# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1018 a_5174_4709# a_5174_4480# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1019 a_5173_7102# a_5701_7354# a_5909_7354# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1020 a_7939_5632# a_8196_5442# a_7798_6224# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1021 a_119_3106# a_119_2649# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1022 vdd d2 a_2998_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1023 a_7943_5455# a_8927_5752# a_8878_5942# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1024 a_5703_5702# a_5490_5702# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1025 a_5174_4250# a_5702_4045# a_5910_4045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1026 a_5178_842# a_5704_736# a_5912_736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1027 a_6861_2673# a_6570_1557# a_6850_2149# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1028 a_7797_8430# a_7987_7648# a_7942_7661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1029 a_3820_6450# a_4077_6260# a_2882_6694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1030 a_5909_6251# a_5488_6251# a_5174_5999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1031 a_118_5542# a_647_5661# a_855_5661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1032 a_119_2462# a_648_2352# a_856_2352# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_2741_8389# a_2931_7607# a_2882_7797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1034 a_7941_1220# a_8198_1030# a_7800_1812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1035 a_5175_2690# a_5703_2942# a_5911_2942# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1036 a_6750_7085# a_6537_7085# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1037 a_1694_4844# a_1481_4844# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1038 a_8879_3736# a_9136_3546# a_7944_3249# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1039 a_2889_1002# a_3142_989# a_2744_1771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_7945_1043# a_8929_1340# a_8880_1530# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1041 a_2778_4884# a_2821_7083# a_2776_7096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1042 a_5910_5148# a_6641_5458# a_6849_5458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1043 a_5912_2393# a_6642_2149# a_6850_2149# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1044 a_6780_8175# a_6567_8175# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1045 a_7832_7137# a_8085_7124# a_7834_4925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1046 a_8880_6314# a_9133_6301# a_7938_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1047 a_7943_5455# a_8927_5752# a_8882_5765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1048 a_7799_4018# a_8056_3828# a_7834_2725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1049 vdd d0 a_4079_2951# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1050 a_2743_3977# a_2933_3195# a_2884_3385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1051 a_6430_1046# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1052 a_1511_8134# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1053 a_2747_3800# a_3000_3787# a_2778_2684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1054 a_5912_736# a_6643_1046# a_6851_1046# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1055 a_118_5542# a_118_5312# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1056 a_7945_1043# a_8929_1340# a_8884_1353# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1057 a_7942_7661# a_8195_7648# a_7797_8430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1058 a_1696_2632# a_1483_2632# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1059 a_854_6764# a_1584_6520# a_1792_6520# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1060 a_3823_8479# a_4076_8466# a_2881_8900# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 a_117_7518# a_645_7313# a_853_7313# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1062 a_7828_7314# a_8085_7124# a_7834_4925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1063 a_5175_3793# a_5175_3606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1064 vdd a_2998_8199# a_2790_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1065 a_5490_5702# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1066 a_6951_177# a_6738_177# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1067 a_855_1798# a_434_1798# a_120_1546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1068 a_7944_3249# a_8197_3236# a_7799_4018# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1069 a_1725_5928# a_1512_5928# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1070 a_7798_6224# a_7988_5442# a_7939_5632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1071 a_6750_4885# a_6537_4885# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1072 a_3825_4067# a_4078_4054# a_2883_4488# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1073 a_3822_3141# a_3827_2415# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1074 a_1481_4844# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1075 a_2882_6694# a_3869_6260# a_3820_6450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1076 gnd a_3140_5401# a_2932_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1077 a_3819_8656# a_4076_8466# a_2881_8900# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1078 a_5908_8457# a_5487_8457# a_5173_8205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 a_1583_8726# a_1370_8726# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1080 a_117_7748# a_646_7867# a_854_7867# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1081 a_118_4668# a_647_4558# a_855_4558# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1082 a_7940_3426# a_8197_3236# a_7799_4018# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1083 a_8875_8697# a_8881_7971# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1084 a_5174_4896# a_5702_5148# a_5910_5148# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1085 a_7944_3249# a_8928_3546# a_8879_3736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1086 a_7798_6224# a_7988_5442# a_7943_5455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1087 a_3821_4244# a_4078_4054# a_2883_4488# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1088 a_5704_3496# a_5491_3496# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1089 a_7804_1635# a_8057_1622# a_7830_2902# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1090 a_6752_2673# a_6539_2673# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1091 a_5909_7354# a_5488_7354# a_5173_7559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1092 a_1483_2632# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1093 a_1808_7163# a_1694_7044# a_1808_4963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1094 a_2882_6694# a_3869_6260# a_3824_6273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1095 a_1585_4314# a_1372_4314# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1096 a_119_3336# a_648_3455# a_856_3455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1097 a_8879_8520# a_9132_8507# a_7937_8941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_6848_7664# a_6427_7664# a_5909_7354# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1099 a_2746_6006# a_2999_5993# a_2772_7273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1100 a_7944_3249# a_8928_3546# a_8883_3559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1101 a_2744_1771# a_2934_989# a_2885_1179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1102 a_5173_8018# a_5173_7789# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1103 a_6781_5969# a_6568_5969# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1104 a_8881_4108# a_9134_4095# a_7939_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_7800_1812# a_8057_1622# a_7830_2902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1106 a_1512_5928# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1107 a_7834_4925# a_7877_7124# a_7828_7314# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1108 a_7938_6735# a_8925_6301# a_8876_6491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_7834_2725# a_7848_3828# a_7803_3841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1110 a_5703_2942# a_5490_2942# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1111 a_5173_6915# a_5702_6805# a_5910_6805# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1112 a_5701_6251# a_5488_6251# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1113 a_119_3565# a_119_3336# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1114 gnd a_3029_7083# a_2821_7083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1115 a_853_7313# a_1584_7623# a_1792_7623# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1116 a_6640_6561# a_6427_6561# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1117 a_855_4558# a_1585_4314# a_1793_4314# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1118 a_1370_8726# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1119 a_5174_5583# a_5703_5702# a_5911_5702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1120 a_7797_8430# a_7987_7648# a_7938_7838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1121 vdd a_2999_5993# a_2791_5993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1122 a_118_5312# a_646_5107# a_854_5107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1123 a_3820_9210# a_3823_8479# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1124 gnd a_3139_7607# a_2931_7607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_3822_4798# a_4079_4608# a_2887_4311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1126 a_5491_3496# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1127 a_2881_8900# a_3868_8466# a_3819_8656# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 a_7834_4925# a_7877_7124# a_7832_7137# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1129 a_5176_1400# a_5705_1290# a_5913_1290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1130 a_855_2901# a_1586_3211# a_1794_3211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1131 a_6859_7085# a_6750_7085# a_6864_5004# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1132 vdd a_3029_7083# a_2821_7083# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1133 a_118_4439# a_118_4209# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1134 a_1372_4314# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1135 a_3826_1861# a_4079_1848# a_2884_2282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1136 a_7799_4018# a_7989_3236# a_7940_3426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1137 a_6848_7664# a_6780_8175# a_6864_7204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1138 gnd a_3141_3195# a_2933_3195# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1139 a_3821_4244# a_3827_3518# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1140 a_855_2901# a_434_2901# a_119_2649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1141 a_2881_8900# a_3868_8466# a_3823_8479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1142 a_1584_6520# a_1371_6520# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1143 a_5911_1839# a_5490_1839# a_5175_2044# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
C0 d0 vdd 2.11fF
C1 a_1902_4844# a_2004_136# 8.08fF
C2 a_7060_177# a_6958_4885# 8.08fF
C3 a_4954_116# gnd 3.40fF
C4 a_2103_136# gnd 4.59fF
C5 a_8879_976# gnd 2.22fF
C6 a_5178_842# gnd 6.43fF
C7 d0 gnd 23.88fF
C8 a_3823_935# gnd 2.22fF
C9 a_122_801# gnd 6.43fF
C10 a_8883_799# gnd 2.38fF
C11 a_5176_941# gnd 2.23fF
C12 a_3827_758# gnd 2.38fF
C13 a_7941_1220# gnd 2.38fF
C14 d1 gnd 11.78fF
C15 a_5912_736# gnd 2.52fF
C16 a_120_900# gnd 2.23fF
C17 a_2885_1179# gnd 2.38fF
C18 a_856_695# gnd 2.52fF
C19 a_5176_1171# gnd 2.38fF
C20 a_5913_1290# gnd 2.18fF
C21 a_5176_1400# gnd 2.28fF
C22 a_120_1130# gnd 2.38fF
C23 a_857_1249# gnd 2.18fF
C24 a_120_1359# gnd 2.28fF
C25 a_7945_1043# gnd 2.52fF
C26 a_8880_1530# gnd 2.23fF
C27 a_2889_1002# gnd 2.52fF
C28 a_3824_1489# gnd 2.23fF
C29 a_8884_1353# gnd 2.49fF
C30 d2 gnd 6.13fF
C31 a_3828_1312# gnd 2.49fF
C32 a_8878_2079# gnd 2.28fF
C33 a_5176_1587# gnd 2.49fF
C34 a_3822_2038# gnd 2.28fF
C35 a_120_1546# gnd 2.49fF
C36 a_8882_1902# gnd 2.38fF
C37 a_5175_2044# gnd 2.23fF
C38 a_3826_1861# gnd 2.38fF
C39 a_7940_2323# gnd 2.18fF
C40 a_5911_1839# gnd 2.52fF
C41 a_119_2003# gnd 2.23fF
C42 a_2884_2282# gnd 2.18fF
C43 a_855_1798# gnd 2.52fF
C44 a_5175_2274# gnd 2.38fF
C45 a_5912_2393# gnd 2.45fF
C46 a_5175_2503# gnd 2.28fF
C47 a_119_2233# gnd 2.38fF
C48 a_856_2352# gnd 2.45fF
C49 a_119_2462# gnd 2.28fF
C50 a_7944_2146# gnd 2.52fF
C51 a_8879_2633# gnd 2.23fF
C52 a_2888_2105# gnd 2.52fF
C53 a_3823_2592# gnd 2.23fF
C54 a_6861_2673# gnd 2.28fF
C55 a_1805_2632# gnd 2.28fF
C56 a_8883_2456# gnd 2.49fF
C57 d3 gnd 3.32fF
C58 a_3827_2415# gnd 2.49fF
C59 a_7830_2902# gnd 2.04fF
C60 a_2774_2861# gnd 2.04fF
C61 a_8878_3182# gnd 2.28fF
C62 a_5175_2690# gnd 2.49fF
C63 a_3822_3141# gnd 2.28fF
C64 a_119_2649# gnd 2.49fF
C65 a_8882_3005# gnd 2.38fF
C66 a_5175_3147# gnd 2.23fF
C67 a_3826_2964# gnd 2.38fF
C68 a_7940_3426# gnd 2.45fF
C69 a_5911_2942# gnd 2.52fF
C70 a_119_3106# gnd 2.23fF
C71 a_2884_3385# gnd 2.45fF
C72 a_855_2901# gnd 2.52fF
C73 a_5175_3377# gnd 2.38fF
C74 a_5912_3496# gnd 2.18fF
C75 a_5175_3606# gnd 2.28fF
C76 a_119_3336# gnd 2.38fF
C77 a_856_3455# gnd 2.18fF
C78 a_119_3565# gnd 2.28fF
C79 a_7944_3249# gnd 2.52fF
C80 a_8879_3736# gnd 2.23fF
C81 a_2888_3208# gnd 2.52fF
C82 a_3823_3695# gnd 2.23fF
C83 a_8883_3559# gnd 2.49fF
C84 a_6866_2792# gnd 2.45fF
C85 a_3827_3518# gnd 2.49fF
C86 a_1810_2751# gnd 2.45fF
C87 a_7834_2725# gnd 2.34fF
C88 a_2778_2684# gnd 2.34fF
C89 a_8877_4285# gnd 2.28fF
C90 a_5175_3793# gnd 2.49fF
C91 a_3821_4244# gnd 2.28fF
C92 a_119_3752# gnd 2.49fF
C93 a_8881_4108# gnd 2.38fF
C94 a_5174_4250# gnd 2.23fF
C95 a_3825_4067# gnd 2.38fF
C96 a_7939_4529# gnd 2.18fF
C97 a_5910_4045# gnd 2.52fF
C98 a_118_4209# gnd 2.23fF
C99 a_2883_4488# gnd 2.18fF
C100 a_854_4004# gnd 2.52fF
C101 a_5174_4480# gnd 2.38fF
C102 a_5911_4599# gnd 2.45fF
C103 a_5174_4709# gnd 2.28fF
C104 a_118_4439# gnd 2.38fF
C105 a_855_4558# gnd 2.45fF
C106 a_118_4668# gnd 2.28fF
C107 a_7943_4352# gnd 2.52fF
C108 a_8878_4839# gnd 2.23fF
C109 a_2887_4311# gnd 2.52fF
C110 a_3822_4798# gnd 2.23fF
C111 a_8882_4662# gnd 2.50fF
C112 a_7060_177# gnd 6.48fF
C113 a_6859_4885# gnd 3.68fF
C114 a_6958_4885# gnd 5.48fF
C115 a_3826_4621# gnd 2.50fF
C116 a_7830_5102# gnd 3.32fF
C117 a_2004_136# gnd 6.48fF
C118 a_1803_4844# gnd 3.68fF
C119 a_1902_4844# gnd 5.48fF
C120 a_2774_5061# gnd 3.32fF
C121 a_8877_5388# gnd 2.28fF
C122 a_5174_4896# gnd 2.50fF
C123 a_3821_5347# gnd 2.28fF
C124 a_118_4855# gnd 2.50fF
C125 a_8881_5211# gnd 2.38fF
C126 a_5174_5353# gnd 2.23fF
C127 a_3825_5170# gnd 2.38fF
C128 a_7939_5632# gnd 2.45fF
C129 a_5910_5148# gnd 2.52fF
C130 a_118_5312# gnd 2.23fF
C131 a_2883_5591# gnd 2.45fF
C132 a_854_5107# gnd 2.52fF
C133 a_5174_5583# gnd 2.38fF
C134 a_5911_5702# gnd 2.18fF
C135 a_5174_5812# gnd 2.28fF
C136 a_118_5542# gnd 2.38fF
C137 a_855_5661# gnd 2.18fF
C138 a_118_5771# gnd 2.28fF
C139 a_7943_5455# gnd 2.52fF
C140 a_8878_5942# gnd 2.23fF
C141 a_2887_5414# gnd 2.52fF
C142 a_3822_5901# gnd 2.23fF
C143 a_8882_5765# gnd 2.49fF
C144 a_3826_5724# gnd 2.49fF
C145 a_8876_6491# gnd 2.28fF
C146 a_5174_5999# gnd 2.49fF
C147 a_3820_6450# gnd 2.28fF
C148 a_118_5958# gnd 2.49fF
C149 a_8880_6314# gnd 2.38fF
C150 a_5173_6456# gnd 2.23fF
C151 a_3824_6273# gnd 2.38fF
C152 a_7938_6735# gnd 2.18fF
C153 a_5909_6251# gnd 2.52fF
C154 a_117_6415# gnd 2.23fF
C155 a_2882_6694# gnd 2.18fF
C156 a_853_6210# gnd 2.52fF
C157 a_5173_6686# gnd 2.38fF
C158 a_5910_6805# gnd 2.45fF
C159 a_5173_6915# gnd 2.28fF
C160 a_117_6645# gnd 2.38fF
C161 a_854_6764# gnd 2.45fF
C162 a_117_6874# gnd 2.28fF
C163 a_7942_6558# gnd 2.52fF
C164 a_8877_7045# gnd 2.23fF
C165 a_2886_6517# gnd 2.52fF
C166 a_3821_7004# gnd 2.23fF
C167 a_6859_7085# gnd 2.34fF
C168 a_6864_5004# gnd 3.32fF
C169 a_1803_7044# gnd 2.34fF
C170 a_1808_4963# gnd 3.32fF
C171 a_8881_6868# gnd 2.49fF
C172 a_7834_4925# gnd 3.68fF
C173 a_3825_6827# gnd 2.49fF
C174 a_7828_7314# gnd 2.45fF
C175 a_2778_4884# gnd 3.68fF
C176 a_2772_7273# gnd 2.45fF
C177 a_8876_7594# gnd 2.28fF
C178 a_5173_7102# gnd 2.49fF
C179 a_3820_7553# gnd 2.28fF
C180 a_117_7061# gnd 2.49fF
C181 a_8880_7417# gnd 2.38fF
C182 a_5173_7559# gnd 2.23fF
C183 a_3824_7376# gnd 2.38fF
C184 a_7938_7838# gnd 2.45fF
C185 a_5909_7354# gnd 2.52fF
C186 a_117_7518# gnd 2.23fF
C187 a_2882_7797# gnd 2.45fF
C188 a_853_7313# gnd 2.52fF
C189 a_5173_7789# gnd 2.38fF
C190 a_5910_7908# gnd 2.18fF
C191 a_5173_8018# gnd 2.28fF
C192 a_117_7748# gnd 2.38fF
C193 a_854_7867# gnd 2.18fF
C194 a_117_7977# gnd 2.28fF
C195 a_7942_7661# gnd 2.52fF
C196 a_8877_8148# gnd 2.23fF
C197 a_2886_7620# gnd 2.52fF
C198 a_3821_8107# gnd 2.23fF
C199 a_8881_7971# gnd 2.49fF
C200 a_6864_7204# gnd 2.04fF
C201 a_3825_7930# gnd 2.49fF
C202 a_1808_7163# gnd 2.04fF
C203 a_7832_7137# gnd 2.28fF
C204 a_2776_7096# gnd 2.28fF
C205 a_8875_8697# gnd 2.28fF
C206 a_5173_8205# gnd 2.49fF
C207 a_3819_8656# gnd 2.28fF
C208 a_117_8164# gnd 2.49fF
C209 a_8879_8520# gnd 2.38fF
C210 a_5172_8662# gnd 2.23fF
C211 a_3823_8479# gnd 2.38fF
C212 a_7937_8941# gnd 2.18fF
C213 a_5908_8457# gnd 2.52fF
C214 a_116_8621# gnd 2.23fF
C215 a_2881_8900# gnd 2.18fF
C216 a_852_8416# gnd 2.52fF
C217 a_5172_8892# gnd 2.38fF
C218 a_5909_9011# gnd 2.38fF
C219 a_5172_9121# gnd 2.22fF
C220 a_116_8851# gnd 2.38fF
C221 a_853_8970# gnd 2.38fF
C222 a_116_9080# gnd 2.22fF
C223 a_7941_8764# gnd 2.79fF
C224 a_8876_9251# gnd 2.75fF
C225 a_2885_8723# gnd 2.52fF
C226 a_3820_9210# gnd 2.23fF
C227 a_3824_9033# gnd 2.98fF
C228 vdd gnd 224.08fF

Vdd vdd 0 dc 3.3
Vin1 vref 0 3.3
Vd0 d0 0 pulse(0 1.8 0 0 0 5us 10us)
Vd1 d1 0 pulse(0 1.8 0 0 0 10us 20us)
Vd2 d2 0 pulse(0 1.8 0 0 0 20us 40us)
Vd3 d3 0 pulse(0 1.8 0 0 0 40us 80us)
Vd4 d4 0 pulse(0 1.8 0 0 0 80us 160us)
Vd5 d5 0 pulse(0 1.8 0 0 0 160us 320us)
Vd6 d6 0 pulse(0 1.8 0 0 0 320us 640us)

.tran 0.1us 640us
.control
run
plot V(vout) V(d0) V(d1) V(d2) V(d3) V(d4) V(d5) V(d6)
.endc
.end
