* SPICE3 file created from 10bit_DAC.ext - technology: sky130A

.option scale=10000u

X0 a_83962_n11746# a_85059_n11940# a_85010_n11750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 gnd a_8707_n14895# a_8499_n14895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 vdd a_85270_n8899# a_85062_n8899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3 a_18898_3272# a_19155_3082# a_17451_3952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4 a_54739_n12639# a_54739_n13034# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5 vdd d1 a_51581_9096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6 a_73258_n10470# a_74351_n9808# a_74306_n9795# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7 a_49838_11234# a_49925_12743# a_49876_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_12227_n11877# a_12014_n11877# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9 a_66325_n14161# a_66112_n14161# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X10 a_52630_n14709# a_53698_n15020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X11 a_33019_8565# a_33643_9145# a_33851_9145# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X12 a_58107_n5872# a_57686_n5872# a_58013_n5753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X13 a_65851_6110# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X14 gnd a_82514_12735# a_82306_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 vdd d1 a_41089_n4481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X16 a_20205_n11748# a_20210_n12766# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X17 a_76412_n14738# a_75371_n15022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X18 a_44031_n14730# a_42947_n15028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X19 a_14511_n4427# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X20 vdd a_51579_3088# a_51371_3088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X21 a_9238_4721# a_9242_3776# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X22 a_30122_n11740# a_31219_n11934# a_31174_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X23 a_34108_n9753# a_33687_n9753# a_33279_n10069# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_8454_n14882# a_9547_n14220# a_9498_n14030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X25 vdd a_63337_9086# a_63129_9086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X26 a_83965_n8705# a_85062_n8899# a_85013_n8709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_76154_9903# a_76154_9508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X28 a_30129_n7429# a_30382_n7442# a_28682_n8196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_66535_n8153# a_67375_n8157# a_67583_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_41619_5392# a_41876_5202# a_40575_4540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X31 a_60546_11228# a_60633_12737# a_60584_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X32 a_33019_7659# a_33640_7551# a_33848_7551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_33280_n14738# a_33901_n14846# a_34109_n14846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X34 a_1521_n5863# a_1308_n5863# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X35 a_641_9911# a_1262_9832# a_1470_9832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X36 vdd a_84221_n5928# a_84013_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X37 gnd a_19415_n14901# a_19207_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_16257_n5742# a_16651_n9803# a_16606_n9790# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X39 a_55147_n13397# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X40 a_65706_n8074# a_65706_n8469# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X41 a_57753_12230# a_57383_13556# a_56357_14236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X42 a_82262_9781# a_83754_10535# a_83709_10548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X43 a_33903_n6712# a_33690_n6712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X44 gnd d0 a_20465_n6771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X45 a_54478_6469# a_55099_6785# a_55307_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X46 vdd a_30119_7500# a_29911_7500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X47 a_17412_5220# a_17499_6729# a_17450_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_67160_n12718# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X49 a_24027_n9751# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X50 a_30914_7509# a_31167_7496# a_29862_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_33851_10592# a_34691_11267# a_34899_11267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X52 a_1730_n8830# a_2570_n8155# a_2778_n8155# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X53 a_71810_n8019# a_72067_n8209# a_71767_n6574# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X54 a_28637_n12759# a_28890_n12772# a_27567_n9609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X55 a_56615_n11202# a_56194_n11202# a_55567_n11877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X56 vdd d0 a_85269_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X57 a_37454_9136# a_37033_9136# a_36388_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X58 a_41878_n10303# a_42135_n10493# a_40830_n10299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X59 a_44602_9832# a_44181_9832# a_43773_9516# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 a_6746_6748# a_8238_7502# a_8193_7515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X61 gnd a_73251_6053# a_73043_6053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X62 gnd a_52626_7498# a_52418_7498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X63 a_41880_n3616# a_42137_n3806# a_40836_n4468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X64 gnd d0 a_20463_n12779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 vdd a_84219_n11936# a_84011_n11936# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X66 a_65852_4590# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X67 a_27091_5271# a_26670_5271# a_26746_9142# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X68 vdd a_74302_10537# a_74094_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X69 a_65703_n11510# a_65703_n11765# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X70 a_55568_n12718# a_55147_n12718# a_54739_n13034# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X71 a_66534_n4418# a_66113_n4418# a_65705_n4851# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 gnd a_28932_n11250# a_28724_n11250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 a_67583_n6710# a_67162_n6710# a_66535_n7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X74 a_16027_5267# a_16391_8180# a_16346_8193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X75 a_1467_6791# a_1046_6791# a_638_6870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X76 a_56358_11269# a_55937_11269# a_55310_10594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 a_65854_10598# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 a_44861_n4416# a_44440_n4416# a_44032_n4308# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X79 a_641_9911# a_641_9516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X80 a_12436_n14844# a_13276_n14169# a_13484_n14169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X81 vdd d0 a_9495_4531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X82 a_76775_9145# a_76562_9145# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X83 a_51324_10733# a_52421_10539# a_52376_10552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X84 a_71550_9964# a_71807_9774# a_71507_11409# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X85 a_81151_8191# a_82264_11213# a_82219_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X86 a_83966_n11923# a_85059_n11261# a_85014_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X87 vdd d6 a_53885_n1645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X88 a_36554_n5755# a_36440_n5874# a_36648_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X89 gnd a_38187_n5934# a_37979_n5934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_11347_3247# a_11968_3139# a_12176_3139# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X91 a_76413_n4316# a_77034_n4424# a_77242_n4424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_54740_n5506# a_55361_n5190# a_55569_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X93 a_66114_n7385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X94 a_1728_n13391# a_1307_n13391# a_899_n13283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X95 a_2354_n9749# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X96 a_25470_6107# a_25257_6107# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X97 a_76772_7551# a_76559_7551# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X98 a_23400_n11194# a_22979_n11194# a_22571_n11510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X99 a_13485_n5194# a_13064_n5194# a_12437_n5869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X100 a_44391_6791# a_44178_6791# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X101 a_51588_n8874# a_52681_n8212# a_52632_n8022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 a_51581_n11738# a_52678_n11932# a_52629_n11742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X103 a_56618_n6714# a_56197_n6714# a_55570_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X104 a_51328_9109# a_51581_9096# a_49877_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X105 a_35157_n14171# a_36396_n13404# a_36547_n11882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X106 a_83969_n8882# a_85062_n8220# a_85017_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X107 a_1469_13567# a_1048_13567# a_640_13675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X108 a_62032_9280# a_62289_9090# a_60585_9960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X109 a_7003_n14025# a_8499_n14895# a_8450_n14705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 gnd a_41875_6043# a_41667_6043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_22721_12118# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X112 vdd d0 a_52887_n13452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X113 a_2355_n14163# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X114 a_71808_n14027# a_72065_n14217# a_71765_n12582# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X115 gnd a_41087_n11936# a_40879_n11936# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X116 a_47298_n11874# a_46934_n13396# a_45908_n14163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 a_76775_10592# a_76562_10592# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 a_66112_n14161# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X119 a_1468_5271# a_2308_5267# a_2516_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X120 a_1262_10600# a_1049_10600# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X121 a_5894_n9607# a_7009_n12770# a_6964_n12757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X122 a_52632_n6575# a_52889_n6765# a_51588_n7427# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X123 a_1730_n6704# a_1309_n6704# a_901_n7020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X124 a_12177_14240# a_11756_14240# a_11348_14319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X125 vdd a_70611_n5928# a_70403_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X126 a_51321_7692# a_52418_7498# a_52373_7511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X127 a_65704_n14082# a_65704_n14477# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X128 a_68971_n11876# a_68862_n11876# a_69070_n11876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X129 a_36398_n7396# a_36185_n7396# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_55569_n3743# a_55148_n3743# a_54740_n3664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X131 gnd a_1520_n14838# a_1728_n14838# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X132 a_25732_n5868# a_25519_n5868# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X133 a_13277_n3747# a_13064_n3747# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X134 a_36136_4579# a_35923_4579# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 gnd a_6999_6735# a_6791_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_67581_n14165# a_67160_n14165# a_66533_n14840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 gnd d0 a_63335_5204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X138 a_22934_14244# a_22721_14244# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X139 a_56356_3814# a_57595_4581# a_57746_6103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X140 a_18898_4719# a_19995_4525# a_19946_4715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X141 vdd d0 a_74299_6728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X142 vdd a_82774_n5248# a_82566_n5248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X143 gnd d1 a_83960_4527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 a_49838_11234# a_49925_12743# a_49880_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X145 a_22314_11356# a_22314_10961# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X146 a_12017_n7389# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X147 a_33642_12112# a_33429_12112# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X148 a_40574_7507# a_40827_7494# a_39127_6740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X149 vdd a_82514_12735# a_82306_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X150 gnd a_85268_n14907# a_85060_n14907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X151 a_68348_13560# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X152 a_83703_3270# a_84800_3076# a_84751_3266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 gnd d0 a_85008_3755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 a_10566_n15020# a_12228_n14844# a_12436_n14844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X155 a_66066_12797# a_65853_12797# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 a_76982_12112# a_76561_12112# a_76154_11606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X157 a_67321_3818# a_66900_3818# a_66273_3143# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X158 a_23767_6785# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X159 a_43773_3154# a_44392_3145# a_44600_3145# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X160 a_66113_n3739# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X161 a_44602_10600# a_44181_10600# a_43773_10708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X162 a_76561_12791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X163 gnd a_7259_n11248# a_7051_n11248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X164 a_34897_5259# a_34476_5259# a_33849_5263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X165 a_19950_4538# a_20203_4525# a_18898_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_76153_13922# a_76153_13667# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X167 vdd d0 a_31428_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X168 a_55148_n5869# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X169 a_65443_8315# a_66064_8236# a_66272_8236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X170 a_11347_4694# a_11347_4153# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X171 a_3755_4587# a_3542_4587# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X172 a_9241_6064# a_9237_6241# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X173 a_41622_6735# a_41875_6722# a_40574_6060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X174 gnd a_39598_n12778# a_39390_n12778# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X175 a_20208_n7260# a_20212_n8205# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X176 a_16257_n5742# a_16514_n5932# a_10496_n1455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X177 a_13017_12789# a_12804_12789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X178 a_33687_n11200# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X179 a_2777_n5188# a_2356_n5188# a_1729_n5863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X180 a_66326_n5865# a_66113_n5865# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X181 vdd a_73251_6053# a_73043_6053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X182 a_34475_8226# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X183 vdd a_73514_n8889# a_73306_n8889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X184 a_74045_9959# a_74302_9769# a_73001_9107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X185 a_1727_n11192# a_1306_n11192# a_898_n11508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X186 gnd a_17967_n11254# a_17759_n11254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X187 gnd d0 a_74559_n9808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_76819_n11879# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X189 a_67323_9826# a_68562_10593# a_68713_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X190 a_13223_6781# a_14462_7548# a_14619_6222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X191 a_4168_n5866# a_3804_n7388# a_2778_n8155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X192 a_84750_7680# a_84754_6735# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X193 vdd a_27824_n9799# a_27616_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X194 a_44181_11279# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X195 a_63340_n8028# a_63344_n8884# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X196 a_2095_5267# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X197 gnd a_28890_n12772# a_28682_n12772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X198 a_70699_n9609# a_71814_n12772# a_71765_n12582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_11348_12477# a_11969_12793# a_12177_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X200 a_83703_4717# a_83960_4527# a_82260_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X201 a_23193_n12714# a_22980_n12714# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X202 a_46889_10595# a_46676_10595# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X203 a_23140_6110# a_23980_6785# a_24188_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X204 a_78083_n8163# a_77870_n8163# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X205 a_55567_n10430# a_55146_n10430# a_54738_n10322# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X206 a_16606_n9790# a_16859_n9803# a_16257_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X207 a_78030_12787# a_77609_12787# a_76982_12791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X208 a_22313_13673# a_22313_13132# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X209 a_41878_n11750# a_41883_n12768# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X210 vdd a_85268_n14228# a_85060_n14228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X211 a_33641_5263# a_33428_5263# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X212 a_77868_n14171# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X213 a_76414_n8730# a_76411_n9418# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X214 gnd a_9495_4531# a_9287_4531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_67580_n11198# a_68819_n10431# a_68976_n11757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X216 a_51323_13700# a_52420_13506# a_52371_13696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X217 a_76154_11350# a_76775_11271# a_76983_11271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X218 a_11608_n5111# a_11608_n5506# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X219 a_77032_n9753# a_76819_n9753# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X220 vdd a_8449_9096# a_8241_9096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X221 a_73254_n10293# a_74351_n10487# a_74306_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X222 vdd a_31427_n9808# a_31219_n9808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X223 a_41623_3089# a_41619_3266# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X224 vdd a_41875_6043# a_41667_6043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X225 a_65706_n8074# a_66327_n8153# a_66535_n8153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X226 a_49030_n9784# a_50143_n6762# a_50098_n6749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X227 a_22573_n5757# a_23194_n5865# a_23402_n5865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X228 a_34478_11267# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X229 a_77241_n14846# a_76820_n14846# a_76412_n14738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X230 gnd d3 a_50089_5213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X231 a_22571_n10318# a_22571_n10859# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X232 gnd d0 a_63596_n5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X233 a_44440_n4416# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X234 a_17711_n14031# a_17968_n14221# a_17668_n12586# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X235 a_55102_11273# a_54889_11273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X236 a_9502_n12760# a_9755_n12773# a_8454_n13435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X237 a_901_n7275# a_901_n7816# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X238 a_63079_12922# a_63083_12066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X239 gnd a_42138_n8899# a_41930_n8899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_45229_11275# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X241 a_44031_n12377# a_44651_n11871# a_44859_n11871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X242 vdd d0 a_42135_n9814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X243 a_901_n8467# a_1522_n8151# a_1730_n8151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X244 a_11757_9147# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X245 gnd d2 a_39381_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_55307_7553# a_54886_7553# a_54478_7120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 a_76981_3816# a_76560_3816# a_76152_3500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 a_44862_n8830# a_44441_n8830# a_44030_n9410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X249 a_22314_9259# a_22935_9151# a_23143_9151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X250 vdd a_6999_6735# a_6791_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X251 vdd a_7262_n8207# a_7054_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X252 a_52635_n4464# a_52888_n4477# a_51583_n4283# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X253 a_23142_13565# a_22721_13565# a_22313_13132# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X254 a_84756_12743# a_84752_12920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X255 a_84754_7503# a_85007_7490# a_83702_7684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X256 a_68819_n10431# a_68606_n10431# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X257 a_5418_5273# a_4997_5273# a_5073_9144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X258 a_18898_4719# a_19995_4525# a_19950_4538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X259 a_30914_8188# a_30910_8365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X260 a_66899_8232# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X261 a_11754_7553# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X262 a_53727_n1632# a_64921_n1634# a_43231_n1412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X263 a_51321_7692# a_51578_7502# a_49878_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X264 vdd d0 a_31168_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X265 a_66535_n6706# a_66114_n6706# a_65706_n7022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X266 vdd d3 a_7219_n6762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X267 a_29869_10554# a_30122_10541# a_28422_9787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X268 a_3053_n1225# a_2944_n1225# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X269 a_56356_3814# a_55935_3814# a_55308_3139# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X270 a_52375_12072# a_52628_12059# a_51323_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X271 a_58705_9138# a_58492_9138# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X272 a_21608_973# a_21395_973# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X273 a_1729_n3737# a_2569_n3741# a_2777_n3741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 gnd d1 a_30380_n14897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 gnd a_63596_n4483# a_63388_n4483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X276 a_83703_3270# a_84800_3076# a_84755_3089# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X277 a_44862_n6704# a_44441_n6704# a_44033_n6625# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X278 vdd d0 a_85008_3755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X279 a_1469_12799# a_2309_12795# a_2517_12795# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 a_50139_n14202# a_51631_n13448# a_51582_n13258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X281 a_74308_n5234# a_74304_n5057# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X282 a_71553_12754# a_73045_13508# a_73000_13521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X283 a_57847_12111# a_57426_12111# a_57748_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X284 a_25839_n11876# a_25475_n13398# a_24449_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X285 a_48342_5273# a_48129_5273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X286 a_3797_6109# a_3584_6109# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X287 vdd a_52629_9092# a_52421_9092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X288 a_83706_7507# a_84799_8169# a_84750_8359# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X289 a_76414_n6633# a_77035_n6712# a_77243_n6712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 a_29867_3099# a_30120_3086# a_28416_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X291 a_79527_n10437# a_79314_n10437# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X292 a_1306_n9745# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X293 a_19160_n7256# a_20257_n7450# a_20208_n7260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X294 a_30126_n11917# a_30379_n11930# a_28675_n11060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X295 vdd d0 a_63596_n5930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X296 a_19946_4715# a_20203_4525# a_18898_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X297 a_76822_n8159# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X298 a_76980_6104# a_76559_6104# a_76151_6212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X299 a_78028_6779# a_79267_7546# a_79424_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X300 gnd d0 a_74559_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X301 a_52373_8190# a_52626_8177# a_51325_7515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X302 a_41618_6912# a_41875_6722# a_40574_6060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X303 a_77242_n4424# a_78082_n3749# a_78290_n3749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X304 a_43150_941# a_64527_973# a_64849_973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X305 a_25429_13560# a_25216_13560# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X306 a_24190_12793# a_23769_12793# a_23142_12118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X307 a_64527_973# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X308 a_78031_11267# a_79270_10587# a_79421_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X309 a_63082_3091# a_63335_3078# a_62030_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 vdd d0 a_20464_n4483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X311 a_55359_n11877# a_55146_n11877# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X312 vdd a_63594_n9812# a_63386_n9812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X313 a_44601_12120# a_45441_12795# a_45649_12795# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X314 vdd a_42138_n8220# a_41930_n8220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X315 gnd d0 a_31170_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X316 a_44861_n5184# a_45701_n5188# a_45909_n5188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X317 a_35156_n11204# a_34735_n11204# a_34108_n11879# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 a_76412_n13036# a_76412_n13291# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X319 a_57597_10589# a_57384_10589# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X320 a_48044_n8839# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X321 a_67323_11273# a_66902_11273# a_66275_11277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X322 a_68713_12115# a_68604_12115# a_68812_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X323 a_12229_n3743# a_12016_n3743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X324 a_41621_11400# a_41625_10544# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X325 a_46931_12117# a_46718_12117# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X326 a_55309_14240# a_54888_14240# a_54480_13924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X327 a_8453_n10468# a_9546_n9806# a_9497_n9616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X328 vdd d2 a_50132_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X329 a_72999_4546# a_74092_5208# a_74047_5221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X330 vdd a_9495_4531# a_9287_4531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X331 a_2097_11275# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X332 a_76562_9145# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X333 gnd d1 a_73254_9094# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X334 vdd d3 a_50089_5213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X335 a_66065_5269# a_65852_5269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_1047_3824# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 a_22933_5269# a_22720_5269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X338 gnd a_52629_11218# a_52421_11218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X339 a_82518_n8025# a_84014_n8895# a_83969_n8882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X340 vdd a_62287_4529# a_62079_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X341 a_44180_12120# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X342 a_30122_n11740# a_31219_n11934# a_31170_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X343 vdd d0 a_74559_n11255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X344 a_17451_3952# a_18947_3082# a_18898_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X345 a_76983_10592# a_76562_10592# a_76154_10700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X346 a_19945_6235# a_19950_5217# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X347 a_71509_5224# a_71596_6733# a_71547_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X348 a_46976_n11874# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X349 a_68973_n5868# a_68864_n5868# a_69072_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X350 a_7004_n5050# a_8500_n5920# a_8455_n5907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X351 vdd d2 a_39381_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X352 gnd a_84221_n5928# a_84013_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X353 a_14723_n13402# a_14510_n13402# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X354 a_1467_6791# a_2307_6787# a_2515_6787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_76412_n13036# a_77033_n12720# a_77241_n12720# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X356 a_65445_13928# a_66066_14244# a_66274_14244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X357 a_22311_7920# a_22311_7665# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X358 a_1261_13567# a_1048_13567# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X359 vdd a_61101_n5246# a_60893_n5246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X360 a_79314_n10437# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X361 a_1729_n5184# a_1308_n5184# a_900_n5500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X362 a_11348_14319# a_11348_13924# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X363 a_63337_n11748# a_63594_n11938# a_62289_n11744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X364 a_85016_n5919# a_85269_n5932# a_83964_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_76154_11606# a_76774_12112# a_76982_12112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X366 a_11756_12793# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X367 a_44393_14246# a_44180_14246# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X368 a_29865_10731# a_30122_10541# a_28422_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X369 a_44599_7559# a_44178_7559# a_43770_7667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X370 a_44860_n14838# a_45700_n14163# a_45908_n14163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X371 gnd a_63335_5204# a_63127_5204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 gnd d0 a_63337_11212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X373 a_43041_941# a_42828_941# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X374 gnd a_83959_7494# a_83751_7494# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 a_55101_12114# a_54888_12114# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X376 a_1046_6112# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X377 gnd a_84219_n11936# a_84011_n11936# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X378 a_33019_8565# a_33019_8309# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X379 a_6743_3958# a_7000_3768# a_6700_5403# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X380 a_76562_11271# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X381 gnd a_20464_n3804# a_20256_n3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X382 a_29863_3276# a_30120_3086# a_28416_3956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X383 a_54479_3897# a_55100_3818# a_55308_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X384 gnd d0 a_85267_n10493# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X385 a_66274_12797# a_65853_12797# a_65445_12876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X386 a_22573_n5502# a_22573_n5757# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X387 a_22981_n5865# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 gnd a_85008_3755# a_84800_3755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 gnd a_73253_12061# a_73045_12061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X390 gnd d2 a_7002_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X391 gnd a_19417_n8893# a_19209_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_8190_4725# a_9287_4531# a_9238_4721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X393 a_60800_n12586# a_60892_n14221# a_60843_n14031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X394 gnd d6 a_53885_n1645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X395 a_65443_6473# a_65443_6218# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X396 a_34111_n8159# a_34951_n8163# a_35159_n8163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 a_76981_4584# a_77821_5259# a_78029_5259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X398 a_45647_6787# a_45226_6787# a_44599_6791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X399 a_33850_14238# a_34690_14234# a_34898_14234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X400 a_55309_12793# a_56149_12789# a_56357_12789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_12227_n11198# a_12014_n11198# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X402 a_74303_n12585# a_74307_n13441# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X403 a_31177_n8880# a_31430_n8893# a_30125_n8699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X404 gnd a_60799_11215# a_60591_11215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X405 a_54740_n5761# a_54741_n6375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X406 a_40834_n10476# a_41927_n9814# a_41882_n9801# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X407 a_65706_n8724# a_65703_n9412# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X408 a_34896_6779# a_34475_6779# a_33848_6783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X409 a_49876_12933# a_51372_12063# a_51323_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 gnd d0 a_52886_n9806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X411 a_44441_n6704# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X412 a_9240_9282# a_9241_8190# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X413 a_30126_n11917# a_31219_n11255# a_31174_n11242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X414 a_39126_9958# a_39383_9768# a_39083_11403# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X415 a_78290_n3749# a_79529_n4429# a_79686_n5755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X416 a_1468_3824# a_1047_3824# a_639_3508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_83969_n8882# a_85062_n8220# a_85013_n8030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X418 gnd a_41090_n8895# a_40882_n8895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X419 a_73256_n4285# a_74353_n4479# a_74308_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X420 vdd d0 a_52889_n8891# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X421 a_33280_n14088# a_33901_n14167# a_34109_n14167# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X422 a_1521_n5184# a_1308_n5184# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X423 a_641_9261# a_1262_9153# a_1470_9153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 a_8450_n13258# a_8707_n13448# a_7007_n14202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X425 a_53698_n15020# a_55360_n14844# a_55568_n14844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X426 a_3053_n1225# a_43280_n1602# a_21631_n1621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X427 a_76822_n7391# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_60540_5397# a_60797_5207# a_59474_8370# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X429 a_71812_n14204# a_72065_n14217# a_71765_n12582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X430 a_11349_11352# a_11970_11273# a_12178_11273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 a_66534_n5865# a_67374_n5190# a_67582_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X432 a_41884_n5240# a_41880_n5063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X433 a_65705_n4851# a_66326_n4418# a_66534_n4418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X434 a_3541_7554# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X435 a_71551_6746# a_73043_7500# a_72994_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X436 a_54479_5600# a_55099_6106# a_55307_6106# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X437 a_30912_13694# a_30916_12749# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X438 a_5894_n9607# a_7009_n12770# a_6960_n12580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X439 a_52636_n6752# a_52889_n6765# a_51588_n7427# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X440 a_48257_n8839# a_48044_n8839# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X441 gnd a_70611_n5928# a_70403_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X442 a_78031_11267# a_77610_11267# a_76983_10592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X443 a_35159_n6716# a_34738_n6716# a_34111_n7391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X444 a_44179_5271# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X445 a_54738_n9672# a_54738_n10067# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X446 a_33021_12220# a_33022_11606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X447 a_25430_10593# a_25217_10593# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X448 vdd d0 a_85269_n5253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X449 a_67322_12793# a_68561_13560# a_68718_12234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X450 a_74303_n14711# a_74560_n14901# a_73255_n14707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X451 a_44392_3824# a_44179_3824# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X452 a_56408_n14169# a_56195_n14169# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X453 a_55359_n9751# a_55146_n9751# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X454 a_24243_n8157# a_24030_n8157# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X455 a_44602_9153# a_44181_9153# a_43770_8573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X456 gnd d0 a_20204_13500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X457 a_22572_n12635# a_22572_n13030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X458 a_19158_n13264# a_19415_n13454# a_17715_n14208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X459 gnd a_63597_n6771# a_63389_n6771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X460 a_11968_5265# a_11755_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X461 a_67113_5265# a_66900_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X462 a_74049_9103# a_74302_9090# a_72997_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X463 a_85011_n13270# a_85015_n14215# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X464 a_45229_9828# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X465 a_5648_n5913# a_5598_n5926# a_5333_n8839# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X466 a_24190_14240# a_23769_14240# a_23142_14244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X467 gnd a_82774_n5248# a_82566_n5248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_1467_6112# a_1046_6112# a_638_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X469 a_33640_6783# a_33427_6783# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X470 a_79268_4579# a_79055_4579# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X471 a_54741_n6375# a_55361_n5869# a_55569_n5869# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X472 a_55099_8232# a_54886_8232# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X473 a_67582_n3743# a_67161_n3743# a_66534_n3739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X474 a_898_n10316# a_1519_n10424# a_1727_n10424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X475 a_77869_n3749# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X476 a_2516_3820# a_3755_4587# a_3906_6109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X477 a_79528_n13404# a_79315_n13404# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X478 a_17712_n5056# a_17969_n5246# a_17674_n6755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X479 a_82473_n12588# a_82730_n12778# a_81407_n9615# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X480 a_36184_n4429# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X481 a_17451_3952# a_18947_3082# a_18902_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X482 a_37700_5265# a_37591_5265# a_32753_984# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X483 vdd a_30121_13508# a_29913_13508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X484 a_639_4159# a_639_3903# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X485 a_71509_5224# a_71596_6733# a_71551_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X486 a_57641_n10435# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X487 a_31173_n8024# a_31430_n8214# a_30129_n8876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X488 a_30125_n7252# a_30382_n7442# a_28682_n8196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X489 gnd a_31428_n14901# a_31220_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X490 a_44031_n12633# a_44031_n13028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X491 a_76412_n12641# a_76412_n13036# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X492 a_29865_10731# a_30962_10537# a_30913_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X493 a_65851_7557# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X494 a_45488_n5188# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X495 a_49875_3958# a_51371_3088# a_51322_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 a_44391_6112# a_44178_6112# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X497 a_47043_6228# a_46673_7554# a_45647_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X498 a_52631_n5734# a_52888_n5924# a_51583_n5730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X499 a_41625_10544# a_41621_10721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X500 a_51585_n11915# a_52678_n11253# a_52629_n11063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 a_9497_n11742# a_9502_n12760# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X502 a_66112_n14840# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X503 vdd d0 a_20465_n6771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X504 a_65704_n14732# a_64406_n15026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X505 gnd a_19156_12057# a_18948_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X506 a_33279_n11771# a_33280_n12385# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X507 a_33020_4947# a_33641_5263# a_33849_5263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X508 a_69457_9142# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X509 a_28633_n12582# a_28890_n12772# a_27567_n9609# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X510 a_76821_n3745# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X511 vdd a_28892_n6764# a_28684_n6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X512 a_35157_n14171# a_34736_n14171# a_34109_n14846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X513 a_9504_n8878# a_9757_n8891# a_8452_n8697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X514 vdd d0 a_63337_11212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X515 a_14975_n5872# a_15833_n8845# a_16041_n8845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X516 a_63339_n4293# a_63343_n5238# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X517 a_52375_14198# a_52371_14375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X518 a_29862_7690# a_30959_7496# a_30910_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 gnd a_73514_n8889# a_73306_n8889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X520 a_69070_n11876# a_69930_n8841# a_70138_n8841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X521 a_13225_14236# a_14464_13556# a_14621_12230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X522 vdd a_31168_4529# a_30960_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X523 a_66112_n12714# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X524 vdd a_50394_n8207# a_50186_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X525 a_29863_4723# a_30960_4529# a_30911_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X526 a_29868_13521# a_30121_13508# a_28421_12754# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_899_n14475# a_1520_n14159# a_1728_n14159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X528 a_17414_11228# a_17667_11215# a_16346_8193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X529 a_58492_9138# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X530 vdd a_64921_n1634# a_64713_n1634# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X531 a_21395_973# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X532 a_63337_n11748# a_63342_n12766# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X533 a_68810_6107# a_69670_9142# a_69878_9142# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X534 a_54738_n11769# a_54739_n12383# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X535 vdd a_85008_3755# a_84800_3755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X536 vdd d2 a_7002_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X537 gnd d1 a_84222_n8895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 a_77034_n5871# a_76821_n5871# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X539 vdd a_73253_12061# a_73045_12061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X540 a_40830_n10299# a_41087_n10489# a_39387_n11243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X541 a_8190_4725# a_9287_4531# a_9242_4544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X542 a_26883_5271# a_26670_5271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X543 a_67581_n12718# a_67160_n12718# a_66533_n12714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X544 vdd d0 a_74299_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X545 a_22979_n11873# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X546 a_11606_n9416# a_12230_n8836# a_12438_n8836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X547 a_3584_6109# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X548 vdd a_63336_13500# a_63128_13500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X549 vdd a_60799_11215# a_60591_11215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X550 gnd a_85268_n14228# a_85060_n14228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_49876_12933# a_51372_12063# a_51327_12076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X552 vdd d0 a_41875_7490# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X553 a_33019_6862# a_33019_6467# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X554 a_68651_n5868# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X555 a_44602_11279# a_45442_11275# a_45650_11275# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X556 a_56195_n14169# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_73260_n5909# a_73513_n5922# a_71809_n5052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X558 a_22311_7665# a_22932_7557# a_23140_7557# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 vdd d0 a_42135_n10493# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X560 gnd d0 a_85008_3076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_11607_n14481# a_12228_n14165# a_12436_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X562 a_9238_5400# a_9242_4544# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X563 a_9241_6743# a_9237_6920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X564 a_59050_5267# a_58837_5267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X565 a_65853_14244# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X566 a_11348_13924# a_11348_13669# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X567 a_51581_n11738# a_52678_n11932# a_52633_n11919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X568 a_40831_n14713# a_41928_n14907# a_41879_n14717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X569 a_73254_n10293# a_74351_n10487# a_74302_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 gnd d4 a_5891_8186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X571 a_71507_11409# a_71764_11219# a_70443_8197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X572 a_76773_5263# a_76560_5263# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X573 a_54889_9826# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X574 a_17711_n14031# a_19207_n14901# a_19162_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X575 a_76561_12112# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X576 a_55570_n6710# a_56410_n6714# a_56618_n6714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X577 gnd d0 a_52629_10539# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X578 a_23141_3822# a_23981_3818# a_24189_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_30916_13517# a_31169_13504# a_29864_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X580 a_65446_9909# a_66067_9830# a_66275_9830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X581 a_33687_n11879# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X582 a_57748_12111# a_57384_10589# a_56358_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X583 a_85011_n13270# a_85268_n13460# a_83963_n13266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X584 a_11349_9255# a_11346_8567# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X585 gnd d0 a_42135_n9814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X586 a_41622_6056# a_41875_6043# a_40570_6237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_14505_6103# a_14292_6103# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X588 a_38015_8368# a_38272_8178# a_37700_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X589 a_63338_n14715# a_63595_n14905# a_62290_n14711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X590 a_23401_n14840# a_22980_n14840# a_22572_n14732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X591 a_19162_n13441# a_20255_n12779# a_20210_n12766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X592 a_63080_9955# a_63084_9099# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X593 a_31175_n12762# a_31171_n12585# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X594 a_34478_9820# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X595 a_41882_n11248# a_42135_n11261# a_40834_n11923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X596 a_77240_n10432# a_76819_n10432# a_76411_n10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X597 a_66326_n5186# a_66113_n5186# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X598 a_6966_n6749# a_7219_n6762# a_5898_n9784# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X599 a_37506_n8847# a_37293_n8847# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X600 a_76819_n11200# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X601 vdd a_74560_n12775# a_74352_n12775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X602 a_23403_n7385# a_22982_n7385# a_22574_n7818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X603 a_18898_4719# a_19155_4529# a_17455_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X604 a_72998_6066# a_74091_6728# a_74046_6741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X605 a_41624_14190# a_41620_14367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X606 vdd a_50132_3768# a_49924_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X607 a_2776_n14163# a_2355_n14163# a_1728_n14159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X608 vdd d2 a_72065_n14217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X609 a_34477_14234# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X610 a_12435_n11877# a_12014_n11877# a_11607_n12383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X611 a_11349_11608# a_11969_12114# a_12177_12114# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X612 a_66533_n14161# a_66112_n14161# a_65704_n14477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X613 a_82213_5395# a_82470_5205# a_81147_8368# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X614 vdd d1 a_41089_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X615 gnd a_73254_9094# a_73046_9094# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X616 a_21631_n1621# a_43488_n1602# a_3053_n1225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X617 a_41623_3768# a_41619_3945# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X618 a_66064_6789# a_65851_6789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X619 gnd d0 a_63594_n10491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X620 vdd a_53885_n1645# a_53677_n1645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X621 a_13065_n6714# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X622 a_1470_9832# a_1049_9832# a_641_9911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X623 a_78083_n6716# a_77870_n6716# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X624 a_22720_5269# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X625 gnd d0 a_63596_n5930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 a_49836_5226# a_49923_6735# a_49874_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_55147_n14844# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X628 gnd a_28935_n8209# a_28727_n8209# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X629 gnd a_17665_5207# a_17457_5207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X630 a_11757_11273# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X631 vdd d2 a_60839_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X632 a_76982_13559# a_76561_13559# a_76153_13667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X633 a_79099_12109# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X634 a_40835_n14890# a_41928_n14228# a_41883_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X635 vdd d1 a_51841_n8887# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X636 a_25687_n10431# a_25474_n10431# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X637 a_78288_n9757# a_77867_n9757# a_77240_n9753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X638 a_62292_n8703# a_62549_n8893# a_60845_n8023# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X639 a_22573_n5107# a_23194_n5186# a_23402_n5186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X640 a_73261_n7429# a_74354_n6767# a_74309_n6754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X641 a_75301_n1457# a_75558_n1647# a_64664_n1444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X642 a_77241_n14167# a_76820_n14167# a_76412_n14088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X643 a_65705_n5757# a_65706_n6371# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X644 a_65706_n7022# a_66327_n6706# a_66535_n6706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X645 a_77034_n4424# a_76821_n4424# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X646 a_41878_n11750# a_42135_n11940# a_40830_n11746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X647 a_62292_n8703# a_63389_n8897# a_63344_n8884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X648 gnd a_42138_n8220# a_41930_n8220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X649 a_34737_n5196# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X650 gnd a_74561_n3800# a_74353_n3800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X651 a_82217_5218# a_82304_6727# a_82255_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X652 gnd a_52627_5210# a_52419_5210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_33640_8230# a_33427_8230# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X654 a_44030_n11508# a_44651_n11192# a_44859_n11192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X655 vdd a_31429_n4479# a_31221_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X656 a_33901_n13399# a_33688_n13399# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X657 a_63078_4715# a_63082_3770# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X658 a_66275_11277# a_65854_11277# a_65446_10961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X659 a_22979_n10426# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X660 a_33281_n4061# a_33281_n4316# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X661 a_76981_3137# a_76560_3137# a_76154_3146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 a_17410_11405# a_17667_11215# a_16346_8193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X663 a_78029_5259# a_79268_4579# a_79419_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_71511_11232# a_71598_12741# a_71549_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X665 a_14249_7548# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X666 gnd d0 a_20202_7492# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X667 gnd d0 a_63336_14179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X668 vdd a_28890_n12772# a_28682_n12772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X669 a_44861_n5863# a_44440_n5863# a_44032_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X670 a_23140_6110# a_22719_6110# a_22312_5604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 a_66533_n12714# a_67373_n12718# a_67581_n12718# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_74308_n5913# a_74304_n5736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X673 a_70699_n9609# a_71814_n12772# a_71769_n12759# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X674 a_57855_n13402# a_57642_n13402# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_28633_n12582# a_28725_n14217# a_28680_n14204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X676 a_36294_12228# a_35924_13554# a_34898_12787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X677 a_77240_n9753# a_76819_n9753# a_76411_n10069# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X678 a_45702_n8155# a_45489_n8155# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 a_23402_n3739# a_22981_n3739# a_22573_n4055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X680 a_5333_n8839# a_4912_n8839# a_4267_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X681 vdd d0 a_9754_n9806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X682 gnd a_41878_10531# a_41670_10531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X683 a_79310_6101# a_79097_6101# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X684 a_66114_n8832# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X685 vdd d0 a_85008_3076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X686 gnd a_7002_9776# a_6794_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X687 a_50096_n12757# a_50183_n11248# a_50138_n11235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X688 a_899_n13283# a_1520_n13391# a_1728_n13391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 a_12437_n5869# a_12016_n5869# a_11609_n6375# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 a_24242_n3743# a_24029_n3743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X691 a_76980_6104# a_77820_6779# a_78028_6779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X692 a_44032_n4849# a_44653_n4416# a_44861_n4416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X693 a_16342_8370# a_17457_5207# a_17412_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X694 vdd d4 a_5891_8186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X695 a_55570_n7389# a_55149_n7389# a_54741_n7822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X696 a_41878_n11071# a_41882_n11927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X697 a_76414_n6633# a_76414_n7028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X698 a_67322_14240# a_66901_14240# a_66274_13565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X699 a_57642_n13402# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X700 a_24028_n14165# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_57426_12111# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X702 vdd d0 a_63596_n5251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X703 a_52376_9784# a_52629_9771# a_51328_9109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X704 gnd d0 a_74559_n11255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X705 a_9498_n12583# a_9755_n12773# a_8454_n13435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X706 a_9239_13696# a_9496_13506# a_8191_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X707 a_41618_6233# a_41875_6043# a_40570_6237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X708 a_7004_n5050# a_8500_n5920# a_8451_n5730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X709 a_33851_11271# a_33430_11271# a_33022_11350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X710 a_23141_4590# a_22720_4590# a_22312_4157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X711 a_68560_4585# a_68347_4585# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X712 a_1308_n4416# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X713 a_39081_5395# a_39173_3760# a_39124_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 a_78081_n14171# a_77868_n14171# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X715 a_2357_n6708# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X716 a_63079_12243# a_63084_11225# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X717 a_62032_10727# a_62289_10537# a_60589_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X718 gnd a_61101_n5246# a_60893_n5246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X719 a_2096_14242# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X720 a_55359_n11198# a_55146_n11198# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X721 a_44178_6791# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X722 a_14767_n5872# a_14554_n5872# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X723 a_63341_n11925# a_63594_n11938# a_62289_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X724 a_55361_n4422# a_55148_n4422# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 a_26798_n8841# a_26585_n8841# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X726 a_640_13930# a_640_13675# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X727 a_55308_5265# a_54887_5265# a_54479_5344# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X728 a_25474_n10431# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X729 a_12017_n8836# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X730 a_33020_4692# a_33020_4151# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X731 a_37930_n5744# a_38324_n9805# a_38275_n9615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X732 vdd a_63596_n4483# a_63388_n4483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X733 a_58013_n5753# a_57643_n4427# a_56617_n3747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X734 a_11755_5265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X735 a_9242_4544# a_9238_4721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X736 a_83703_4717# a_84800_4523# a_84751_4713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X737 gnd d0 a_9755_n14899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 gnd a_74302_10537# a_74094_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X739 a_65703_n10318# a_65703_n10859# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X740 a_79055_4579# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X741 a_20209_n9799# a_20462_n9812# a_19161_n10474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X742 a_43771_4159# a_44392_4592# a_44600_4592# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X743 a_25259_12115# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X744 a_49836_5226# a_49923_6735# a_49878_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X745 a_19950_3091# a_19946_3268# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X746 a_51324_10733# a_52421_10539# a_52372_10729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X747 a_30911_5398# a_31168_5208# a_29867_4546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X748 a_36182_n10437# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X749 a_20205_n9622# a_20209_n10478# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X750 a_22934_12797# a_22721_12797# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_85014_n10480# a_85010_n10303# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X752 a_79530_n7396# a_79317_n7396# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X753 a_51582_n14705# a_52679_n14899# a_52634_n14886# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X754 a_55308_5265# a_56148_5261# a_56356_5261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X755 a_76151_7659# a_76772_7551# a_76980_7551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X756 a_40834_n10476# a_41927_n9814# a_41878_n9624# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X757 a_1047_3145# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X758 vdd a_20462_n10491# a_20254_n10491# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X759 a_76154_11350# a_76154_10955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X760 a_33427_6783# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X761 a_4171_n11755# a_3801_n10429# a_2775_n11196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X762 vdd d0 a_31170_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X763 a_30126_n11917# a_31219_n11255# a_31170_n11065# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X764 a_66324_n10426# a_66111_n10426# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X765 a_40833_n8705# a_41930_n8899# a_41885_n8886# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X766 vdd a_41088_n14903# a_40880_n14903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X767 vdd a_52627_5210# a_52419_5210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X768 vdd a_73251_7500# a_73043_7500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X769 a_60806_n6755# a_60893_n5246# a_60848_n5233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X770 a_73256_n4285# a_74353_n4479# a_74304_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X771 a_74046_7509# a_74299_7496# a_72994_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X772 a_8454_n13435# a_8707_n13448# a_7007_n14202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 gnd d0 a_85010_10531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X774 a_71511_11232# a_71598_12741# a_71553_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X775 vdd d1 a_40827_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X776 a_68978_n5749# a_68608_n4423# a_67582_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X777 a_85016_n5240# a_85269_n5253# a_83968_n5915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X778 a_63337_n11069# a_63594_n11259# a_62293_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X779 a_59734_n9613# a_60849_n12776# a_60804_n12763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X780 a_11756_12114# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X781 a_19951_12745# a_20204_12732# a_18903_12070# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 vdd a_20465_n7450# a_20257_n7450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X783 vdd a_41878_10531# a_41670_10531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X784 a_66067_9151# a_65854_9151# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X785 a_43770_8317# a_44391_8238# a_44599_8238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 a_34109_n13399# a_33688_n13399# a_33280_n13832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X787 a_56194_n9755# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X788 a_48770_8199# a_49883_11221# a_49834_11411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 vdd a_7002_9776# a_6794_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X790 a_19162_n13441# a_19415_n13454# a_17715_n14208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X791 a_65444_5348# a_65444_4953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X792 a_26670_5271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X793 a_58965_n8845# a_58752_n8845# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X794 gnd a_82472_11213# a_82264_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 gnd a_74299_8175# a_74091_8175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X796 a_5898_n9784# a_6151_n9797# a_5549_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X797 vdd d0 a_9755_n14220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X798 a_5648_n5913# a_5598_n5926# a_5549_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X799 a_3799_12117# a_3586_12117# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X800 gnd d0 a_74299_6728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X801 a_54479_3247# a_55100_3139# a_55308_3139# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X802 a_73254_n11740# a_74351_n11934# a_74306_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X803 a_67159_n11198# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X804 a_66274_12118# a_65853_12118# a_65445_12226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X805 vdd a_41875_7490# a_41667_7490# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X806 vdd d0 a_31430_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X807 a_54479_3502# a_54479_3247# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X808 a_67372_n9751# a_67159_n9751# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X809 a_50137_n8017# a_51633_n8887# a_51588_n8874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X810 a_68602_6107# a_68389_6107# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X811 a_22981_n5186# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X812 gnd a_85008_3076# a_84800_3076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 a_59478_8193# a_60591_11215# a_60542_11405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X814 a_52372_9961# a_52629_9771# a_51328_9109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X815 a_82477_n12765# a_82730_n12778# a_81407_n9615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X816 a_17716_n5233# a_17969_n5246# a_17674_n6755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_76982_12112# a_77822_12787# a_78030_12787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X818 a_76151_8309# a_76151_7914# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X819 a_39388_n14210# a_39641_n14223# a_39341_n12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X820 a_45910_n6708# a_47149_n7388# a_47300_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X821 a_80638_n8847# a_80425_n8847# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X822 a_40577_10548# a_41670_11210# a_41621_11400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X823 a_31177_n8201# a_31430_n8214# a_30129_n8876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X824 a_83962_n10299# a_84219_n10489# a_82519_n11243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X825 a_54738_n10067# a_54738_n10322# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X826 a_76560_5263# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X827 a_41884_n5919# a_41880_n5742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X828 a_34111_n7391# a_34951_n6716# a_35159_n6716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X829 a_39081_5395# a_39173_3760# a_39128_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X830 a_56149_12789# a_55936_12789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X831 a_31177_n7433# a_31173_n7256# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X832 gnd d0 a_20464_n5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 a_52635_n5911# a_52888_n5924# a_51583_n5730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X834 a_76153_13667# a_76153_13126# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X835 a_1468_3145# a_1047_3145# a_641_3154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X836 a_12175_8232# a_13015_8228# a_13223_8228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 a_85012_n5742# a_85269_n5932# a_83964_n5738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X838 a_14292_6103# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 vdd d0 a_52889_n8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X840 vdd a_30381_n4475# a_30173_n4475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X841 a_41879_n14717# a_42136_n14907# a_40831_n14713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X842 a_9239_13696# a_9243_12751# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X843 a_54739_n14481# a_55360_n14165# a_55568_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X844 vdd a_31430_n6767# a_31222_n6767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X845 a_59738_n9790# a_59991_n9803# a_59389_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X846 vdd a_30380_n13450# a_30172_n13450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X847 gnd a_28892_n6764# a_28684_n6764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X848 a_38015_8368# a_39130_5205# a_39085_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X849 a_62035_13517# a_62288_13504# a_60588_12750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X850 a_11348_12222# a_11349_11608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X851 a_40575_4540# a_41668_5202# a_41619_5392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X852 a_47305_n5747# a_46935_n4421# a_45909_n5188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 a_83703_4717# a_84800_4523# a_84755_4536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X854 a_41882_n9801# a_41878_n9624# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X855 a_50135_n14025# a_51631_n14895# a_51582_n14705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X856 a_44392_3145# a_44179_3145# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 a_74049_9782# a_74302_9769# a_73001_9107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_47038_6109# a_46674_4587# a_45648_3820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X859 a_29866_7513# a_30119_7500# a_28419_6746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 gnd a_64921_n1634# a_64713_n1634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X861 a_77610_11267# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X862 a_83706_7507# a_83959_7494# a_82259_6740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 a_29867_4546# a_30120_4533# a_28420_3779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X864 a_40834_n10476# a_41087_n10489# a_39387_n11243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X865 a_19160_n8703# a_20257_n8897# a_20208_n8707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X866 a_79684_n11763# a_79314_n10437# a_78288_n11204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_83707_4540# a_83960_4527# a_82260_3773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X868 a_60800_n12586# a_60892_n14221# a_60847_n14208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X869 gnd d2 a_61102_n8213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X870 gnd a_42135_n10493# a_41927_n10493# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 vdd a_20204_14179# a_19996_14179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X872 a_66899_6785# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 a_44178_8238# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X874 a_67162_n8157# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X875 a_79681_n5874# a_79572_n5874# a_79780_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X876 a_24189_5265# a_23768_5265# a_23141_5269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X877 vdd d2 a_17709_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X878 a_66900_3818# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X879 a_78029_5259# a_77608_5259# a_76981_5263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X880 a_52372_9961# a_52376_9105# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X881 a_63082_4538# a_63335_4525# a_62030_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X882 vdd d0 a_20464_n5930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X883 a_56617_n5194# a_56196_n5194# a_55569_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X884 a_54740_n3664# a_54740_n4059# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X885 a_65706_n6627# a_65706_n7022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X886 a_55567_n11877# a_55146_n11877# a_54739_n12383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 vdd d0 a_85010_10531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X888 gnd a_31428_n14222# a_31220_n14222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X889 a_14462_7548# a_14249_7548# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X890 a_44600_4592# a_45440_5267# a_45648_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X891 a_64849_973# a_75563_984# a_75885_984# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X892 a_84754_7503# a_84750_7680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X893 a_1309_n6704# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_12178_10594# a_13018_11269# a_13226_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X895 a_52631_n5055# a_52888_n5245# a_51587_n5907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X896 gnd a_52626_6730# a_52418_6730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X897 a_85015_n13447# a_85268_n13460# a_83963_n13266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X898 a_75563_984# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 a_65444_4157# a_66065_4590# a_66273_4590# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X900 a_77607_8226# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X901 a_12436_n13397# a_12015_n13397# a_11607_n13289# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X902 a_19947_12922# a_20204_12732# a_18903_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X903 a_19162_n13441# a_20255_n12779# a_20206_n12589# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X904 a_52635_n4464# a_52631_n4287# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X905 gnd a_20202_7492# a_19994_7492# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X906 a_9504_n8199# a_9757_n8212# a_8456_n8874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X907 a_31171_n13264# a_31428_n13454# a_30123_n13260# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X908 a_48770_8199# a_49883_11221# a_49838_11234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X909 a_71814_n8196# a_73306_n7442# a_73257_n7252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 a_76413_n3410# a_85012_n3616# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X911 vdd a_62548_n4479# a_62340_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X912 a_56409_n3747# a_56196_n3747# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X913 a_639_5350# a_1260_5271# a_1468_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X914 vdd a_82472_11213# a_82264_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X915 vdd a_74299_8175# a_74091_8175# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X916 vdd a_63597_n6771# a_63389_n6771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X917 a_13063_n14169# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X918 a_66272_6110# a_67112_6785# a_67320_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X919 gnd d0 a_31168_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X920 gnd a_74560_n12775# a_74352_n12775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X921 a_12177_13561# a_11756_13561# a_11348_13128# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 gnd a_41877_13498# a_41669_13498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 gnd d2 a_72065_n14217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X924 a_47399_n5866# a_46978_n5866# a_47300_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X925 a_47139_12117# a_46718_12117# a_47045_12236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X926 vdd a_85008_3076# a_84800_3076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X927 a_59478_8193# a_60591_11215# a_60546_11228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X928 a_77034_n5192# a_76821_n5192# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X929 a_76154_10955# a_76154_10700# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X930 a_19164_n8880# a_20257_n8218# a_20212_n8205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X931 gnd d1 a_41089_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X932 vdd d1 a_73513_n4475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X933 a_19952_11225# a_19948_11402# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X934 a_65443_7124# a_65443_6868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X935 a_1470_9153# a_2310_9828# a_2518_9828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X936 a_46935_n4421# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X937 a_36552_n11763# a_36438_n11882# a_36646_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X938 a_22979_n11194# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X939 a_11609_n8473# a_12230_n8157# a_12438_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X940 a_40577_10548# a_41670_11210# a_41625_11223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X941 a_75885_984# a_80510_5265# a_80832_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 a_44600_5271# a_44179_5271# a_43771_4955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X943 vdd d0 a_74560_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X944 gnd a_53885_n1645# a_53677_n1645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_36183_n13404# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X946 a_3906_6109# a_3542_4587# a_2516_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X947 a_56148_5261# a_55935_5261# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X948 a_83705_10725# a_84802_10531# a_84753_10721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X949 a_11349_9905# a_11349_9510# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X950 vdd d1 a_19415_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X951 a_4166_n11874# a_3802_n13396# a_2776_n14163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_51585_n11915# a_52678_n11253# a_52633_n11240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X953 a_39386_n8025# a_40882_n8895# a_40837_n8882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X954 a_66325_n13393# a_66112_n13393# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X955 a_40835_n14890# a_41928_n14228# a_41879_n14038# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X956 gnd a_52886_n9806# a_52678_n9806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X957 a_74048_14196# a_74301_14183# a_73000_13521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X958 gnd d1 a_51841_n8887# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X959 a_35159_n6716# a_36398_n7396# a_36549_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X960 a_73261_n7429# a_74354_n6767# a_74305_n6577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_70453_n5915# a_75558_n1647# a_64664_n1444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X962 a_66273_3822# a_65852_3822# a_65444_3506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X963 a_54889_9147# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X964 a_46886_7554# a_46673_7554# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X965 a_12437_n3743# a_13277_n3747# a_13485_n3747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X966 a_9497_n11063# a_9501_n11919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X967 a_47137_6109# a_46716_6109# a_47043_6228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X968 a_52371_13696# a_52628_13506# a_51323_13700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X969 a_65704_n12635# a_65704_n13030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X970 a_30912_14373# a_30916_13517# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X971 a_65446_9259# a_66067_9151# a_66275_9151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X972 a_44859_n10424# a_44438_n10424# a_44030_n10857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 a_22313_13132# a_22934_13565# a_23142_13565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X974 a_1307_n14838# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X975 a_41882_n11927# a_42135_n11940# a_40830_n11746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X976 a_65444_4953# a_65444_4698# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X977 a_84757_9097# a_84753_9274# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X978 a_74306_n9795# a_74559_n9808# a_73258_n10470# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X979 gnd a_31429_n4479# a_31221_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X980 a_23770_11273# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X981 a_54886_7553# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_23401_n14161# a_22980_n14161# a_22572_n14082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X983 a_83968_n4468# a_84221_n4481# a_82521_n5235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X984 a_22571_n11765# a_22572_n12379# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X985 vdd d0 a_74561_n3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X986 a_74305_n8703# a_74562_n8893# a_73257_n8699# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X987 gnd d1 a_8446_6055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X988 a_4997_5273# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X989 a_29863_4723# a_30120_4533# a_28420_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X990 a_52634_n13439# a_52887_n13452# a_51582_n13258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X991 a_55146_n9751# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X992 a_28633_n12582# a_28725_n14217# a_28676_n14027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X993 a_65445_12876# a_66066_12797# a_66274_12797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 gnd d0 a_20205_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_76151_7914# a_76151_7659# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X996 a_66533_n14840# a_66112_n14840# a_64406_n15026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X997 a_47191_n5866# a_46978_n5866# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X998 a_81407_n9615# a_81664_n9805# a_81062_n5744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X999 a_77609_12787# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1000 a_72994_6243# a_74091_6049# a_74046_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1001 a_33282_n8730# a_33903_n8838# a_34111_n8838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1002 a_39347_n6757# a_39434_n5248# a_39389_n5235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1003 a_23192_n9747# a_22979_n9747# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1004 a_72999_3099# a_73252_3086# a_71548_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 a_12435_n11198# a_12014_n11198# a_11606_n11514# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1006 gnd d2 a_50132_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1007 a_44393_12799# a_44180_12799# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1008 a_52629_n11742# a_52634_n12760# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1009 a_24451_n6710# a_24030_n6710# a_23403_n6706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1010 a_49880_12756# a_51372_13510# a_51323_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1011 a_50096_n12757# a_50183_n11248# a_50134_n11058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1012 a_73256_n5732# a_73513_n5922# a_71809_n5052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1013 a_30910_6918# a_31167_6728# a_29866_6066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1014 a_63078_4715# a_63335_4525# a_62030_4719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1015 a_44030_n11763# a_44031_n12377# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1016 a_76411_n11771# a_76412_n12385# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1017 a_24448_n11198# a_24027_n11198# a_23400_n11194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1018 a_20211_n4470# a_20207_n4293# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1019 a_12435_n11198# a_13275_n11202# a_13483_n11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1020 a_1260_3824# a_1047_3824# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1021 a_55307_6785# a_56147_6781# a_56355_6781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1022 a_66533_n12714# a_66112_n12714# a_65704_n12635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1023 a_73256_n5732# a_74353_n5926# a_74308_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1024 a_1470_9153# a_1049_9153# a_641_9261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1025 a_23400_n10426# a_24240_n9751# a_24448_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1026 a_33282_n7028# a_33903_n6712# a_34111_n6712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1027 gnd d5 a_16514_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1028 a_22312_4953# a_22933_5269# a_23141_5269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1029 gnd d0 a_52887_n14899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 a_60542_11405# a_60634_9770# a_60585_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1031 gnd a_28673_3766# a_28465_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1032 vdd a_52626_6730# a_52418_6730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1033 a_55147_n14165# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1034 a_65706_n6371# a_66326_n5865# a_66534_n5865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1035 a_25730_n11876# a_25517_n11876# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1036 a_44654_n7383# a_44441_n7383# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1037 gnd a_62287_4529# a_62079_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1038 a_33282_n8080# a_33282_n8475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1039 a_23192_n11873# a_22979_n11873# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 gnd d0 a_85009_13498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1041 a_36438_n11882# a_36225_n11882# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1042 a_30128_n4462# a_31221_n3800# a_22573_n3404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1043 a_8196_9109# a_8449_9096# a_6745_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1044 a_638_7922# a_638_7667# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1045 vdd a_40827_6047# a_40619_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1046 a_22311_7665# a_22311_7124# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1047 a_11606_n11119# a_11606_n11514# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1048 a_56616_n14169# a_56195_n14169# a_55568_n14844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1049 a_41878_n11071# a_42135_n11261# a_40834_n11923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1050 a_13278_n8161# a_13065_n8161# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1051 a_33643_9824# a_33430_9824# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1052 vdd a_63594_n10491# a_63386_n10491# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1053 a_34950_n3749# a_34737_n3749# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1054 a_63080_9276# a_63081_8184# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1055 a_6962_n6572# a_7219_n6762# a_5898_n9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1056 a_64740_973# a_64527_973# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1057 a_2567_n11196# a_2354_n11196# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1058 a_76983_11271# a_77823_11267# a_78031_11267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1059 vdd a_84220_n14903# a_84012_n14903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1060 vdd d0 a_9494_8177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1061 a_44861_n5184# a_44440_n5184# a_44032_n5105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1062 a_34111_n8838# a_33690_n8838# a_33282_n8730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1063 vdd d0 a_85268_n13460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1064 a_1259_7559# a_1046_7559# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1065 a_17455_3775# a_18947_4529# a_18902_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1066 a_17414_11228# a_17501_12737# a_17456_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1067 a_41624_12064# a_41620_12241# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1068 a_2777_n3741# a_4016_n4421# a_4173_n5747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1069 a_6747_3781# a_7000_3768# a_6700_5403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1070 vdd a_52886_n10485# a_52678_n10485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1071 a_45702_n6708# a_45489_n6708# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1072 a_7004_n5050# a_7261_n5240# a_6966_n6749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1073 a_66114_n8153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1074 a_30917_11229# a_30913_11406# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1075 a_58011_n11761# a_57641_n10435# a_56615_n11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1076 a_83705_10725# a_84802_10531# a_84757_10544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1077 gnd d0 a_42135_n11261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1078 a_12437_n5190# a_12016_n5190# a_11608_n5506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 a_36648_n5874# a_36227_n5874# a_36549_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1080 a_22573_n4310# a_22573_n4851# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1081 a_49879_3781# a_51371_4535# a_51322_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1082 a_77242_n4424# a_76821_n4424# a_76413_n4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 a_16346_8193# a_16599_8180# a_16027_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1084 a_74044_14373# a_74301_14183# a_73000_13521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1085 a_78291_n6716# a_77870_n6716# a_77243_n7391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1086 a_12805_11269# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1087 a_45907_n9749# a_45486_n9749# a_44859_n9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1088 a_36386_6101# a_35965_6101# a_36287_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1089 a_74307_n12762# a_74303_n12585# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1090 vdd d1 a_62549_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1091 a_51326_3101# a_52419_3763# a_52370_3953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1092 a_65706_n8469# a_65706_n8724# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1093 vdd d0 a_9756_n4477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1094 vdd d0 a_52887_n14220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1095 a_82518_n8025# a_82775_n8215# a_82475_n6580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1096 a_48681_n5736# a_48938_n5926# a_48780_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1097 a_52376_9105# a_52629_9092# a_51324_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_44653_n3737# a_44440_n3737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1099 a_82255_6917# a_83751_6047# a_83706_6060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1100 vdd d7 a_21789_n1634# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1101 a_67161_n3743# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1102 a_24028_n12718# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1103 a_60806_n6755# a_60893_n5246# a_60844_n5056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 a_39130_9781# a_39383_9768# a_39083_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 vdd d1 a_8446_6055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1106 a_33429_12791# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1107 a_18901_7509# a_19994_8171# a_19945_8361# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1108 a_63341_n11246# a_63594_n11259# a_62293_n11921# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_59734_n9613# a_60849_n12776# a_60800_n12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1110 vdd d0 a_20205_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1111 a_2356_n3741# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1112 a_43771_3508# a_43771_3253# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1113 a_40830_n11746# a_41087_n11936# a_39383_n11066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1114 vdd a_73253_13508# a_73045_13508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1115 a_19945_7682# a_19949_6737# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1116 a_12228_n12718# a_12015_n12718# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1117 a_33428_3816# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1118 a_77240_n11879# a_78080_n11204# a_78288_n11204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1119 a_85017_n8207# a_85013_n8030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1120 a_12017_n8157# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1121 gnd a_20465_n7450# a_20257_n7450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1122 a_65705_n3404# a_74304_n3610# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1123 a_72995_3276# a_73252_3086# a_71548_3956# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1124 a_1519_n11871# a_1306_n11871# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_19950_3770# a_19946_3947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1126 a_22932_6110# a_22719_6110# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1127 a_25584_6226# a_25214_7552# a_24188_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 a_8455_n4460# a_9548_n3798# a_900_n3402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1129 vdd a_21789_n1634# a_21581_n1634# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1130 a_74048_14196# a_74044_14373# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1131 a_49880_12756# a_51372_13510# a_51327_13523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1132 a_9244_9105# a_9240_9282# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1133 a_23140_7557# a_22719_7557# a_22311_7665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1134 a_48550_5273# a_54103_986# a_54311_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1135 vdd a_81319_n5934# a_81111_n5934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1136 vdd d0 a_42135_n11940# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1137 gnd a_17708_3762# a_17500_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1138 gnd d0 a_85008_4523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1139 gnd d0 a_9755_n14220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1140 a_66066_13565# a_65853_13565# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1141 a_62289_n10297# a_63386_n10491# a_63341_n10478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1142 a_23192_n10426# a_22979_n10426# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1143 a_24190_14240# a_25429_13560# a_25586_12234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1144 a_36440_n5874# a_36227_n5874# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1145 a_73254_n11740# a_74351_n11934# a_74302_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1146 gnd d0 a_31430_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1147 a_52369_7688# a_52373_6743# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1148 a_50137_n8017# a_51633_n8887# a_51584_n8697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1149 a_60542_11405# a_60634_9770# a_60589_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1150 a_19949_8184# a_20202_8171# a_18901_7509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1151 vdd a_28673_3766# a_28465_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1152 a_78028_6779# a_77607_6779# a_76980_6783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1153 vdd d0 a_31169_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1154 a_43772_13930# a_43772_13675# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1155 a_83966_n10476# a_84219_n10489# a_82519_n11243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1156 a_56358_11269# a_57597_10589# a_57748_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1157 a_37033_9136# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1158 a_47139_12117# a_47997_9144# a_48205_9144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1159 a_11608_n3664# a_12229_n3743# a_12437_n3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1160 a_33427_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1161 a_63078_5394# a_63082_4538# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1162 gnd a_30381_n4475# a_30173_n4475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1163 a_22933_4590# a_22720_4590# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1164 a_7002_n11058# a_7259_n11248# a_6964_n12757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1165 a_33903_n7391# a_33690_n7391# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1166 gnd a_31430_n6767# a_31222_n6767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1167 a_54481_10702# a_54481_10161# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1168 a_65853_12797# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1169 gnd a_30380_n13450# a_30172_n13450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1170 gnd a_9754_n9806# a_9546_n9806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1171 a_33282_n6377# a_33282_n6633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1172 a_24241_n14165# a_24028_n14165# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1173 a_23403_n8832# a_22982_n8832# a_22571_n9412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1174 a_51327_12076# a_52420_12738# a_52375_12751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1175 a_638_6870# a_1259_6791# a_1467_6791# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1176 a_66067_9830# a_65854_9830# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1177 a_55307_7553# a_56147_8228# a_56355_8228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1178 a_901_n7275# a_1522_n7383# a_1730_n7383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1179 a_1728_n14159# a_2568_n14163# a_2776_n14163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 a_37591_5265# a_37378_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1181 a_20207_n3614# a_20211_n4470# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1182 a_55100_4586# a_54887_4586# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1183 gnd a_31168_4529# a_30960_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1184 a_19951_12066# a_20204_12053# a_18899_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1185 a_44860_n12712# a_44439_n12712# a_44031_n13028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1186 a_76152_5598# a_76152_5342# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1187 a_36180_12109# a_35967_12109# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1188 a_55568_n13397# a_55147_n13397# a_54739_n13289# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1189 vdd a_84222_n8895# a_84014_n8895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1190 a_49879_3781# a_51371_4535# a_51326_4548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1191 a_26992_5271# a_26883_5271# a_27091_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1192 a_74049_9782# a_74045_9959# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1193 a_16342_8370# a_16599_8180# a_16027_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1194 a_67581_n14165# a_68820_n13398# a_68971_n11876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1195 a_14252_10589# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 gnd d0 a_74299_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1197 vdd a_19156_13504# a_18948_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1198 a_73258_n11917# a_74351_n11255# a_74306_n11242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1199 a_51326_3101# a_52419_3763# a_52374_3776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1200 gnd d0 a_31429_n3800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1201 a_76774_12791# a_76561_12791# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1202 a_1048_12120# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1203 a_56147_6781# a_55934_6781# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1204 a_77243_n8838# a_78083_n8163# a_78291_n8163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1205 a_83704_13692# a_84801_13498# a_84752_13688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1206 a_3844_n11874# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1207 a_4057_n11874# a_3844_n11874# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1208 a_25844_n11757# a_25474_n10431# a_24448_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1209 a_67582_n3743# a_68821_n4423# a_68978_n5749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1210 a_85011_n14717# a_84756_14190# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1211 gnd d0 a_20464_n5930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1212 vdd d0 a_52888_n3798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1213 a_25678_6107# a_25257_6107# a_25584_6226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1214 vdd a_31429_n5926# a_31221_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1215 a_76152_4947# a_76773_5263# a_76981_5263# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1216 a_71511_11232# a_71764_11219# a_70443_8197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1217 a_46673_7554# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1218 a_44599_6791# a_44178_6791# a_43770_6870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1219 a_33901_n14846# a_33688_n14846# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1220 a_77870_n8163# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1221 gnd d1 a_8708_n4473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1222 gnd a_51581_9096# a_51373_9096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1223 a_1519_n10424# a_1306_n10424# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1224 a_52635_n5232# a_52888_n5245# a_51587_n5907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1225 a_18901_7509# a_19994_8171# a_19949_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1226 a_12178_9826# a_13018_9822# a_13226_9822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1227 a_78289_n12724# a_77868_n12724# a_77241_n12720# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1228 vdd d4 a_59991_n9803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1229 a_62034_4542# a_63127_5204# a_63082_5217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1230 a_85012_n5063# a_85269_n5253# a_83968_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1231 gnd d1 a_83961_12055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1232 a_33902_n3745# a_33689_n3745# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1233 a_12175_7553# a_11754_7553# a_11346_7661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1234 a_51585_n10468# a_51838_n10481# a_50138_n11235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1235 a_36552_n11763# a_36182_n10437# a_35156_n9757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1236 a_8195_12076# a_8448_12063# a_6744_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1237 a_1730_n7383# a_1309_n7383# a_901_n7275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1238 a_63344_n8884# a_63340_n8707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1239 a_38019_8191# a_38272_8178# a_37700_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1240 gnd a_8446_6055# a_8238_6055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1241 a_31175_n13441# a_31428_n13454# a_30123_n13260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1242 a_64527_973# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1243 a_62029_6239# a_62286_6049# a_60582_6919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1244 a_3803_n4421# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1245 vdd d2 a_39640_n11256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1246 a_46933_n10429# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1247 a_900_n3658# a_1521_n3737# a_1729_n3737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 gnd a_63596_n5251# a_63388_n5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 gnd a_62548_n4479# a_62340_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1250 a_83962_n10299# a_85059_n10493# a_85010_n10303# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1251 vdd a_17708_3762# a_17500_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1252 vdd d0 a_85008_4523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1253 gnd a_72066_n5242# a_71858_n5242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1254 a_70015_5271# a_69802_5271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1255 a_12227_n10430# a_12014_n10430# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1256 a_44601_12799# a_44180_12799# a_43772_12878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1257 a_898_n11113# a_898_n11508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1258 a_44033_n6369# a_44653_n5863# a_44861_n5863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1259 a_3913_12236# a_3543_13562# a_2517_12795# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1260 a_55570_n8836# a_55149_n8836# a_54738_n9416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1261 a_63343_n4470# a_63596_n4483# a_62291_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1262 a_72998_6066# a_74091_6728# a_74042_6918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_65444_3251# a_65446_3152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1264 a_18902_4542# a_19155_4529# a_17455_3775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1265 a_19945_8361# a_20202_8171# a_18901_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1266 gnd a_50132_3768# a_49924_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1267 vdd d0 a_63595_n13458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1268 a_19164_n8880# a_20257_n8218# a_20208_n8028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1269 a_13223_6781# a_12802_6781# a_12175_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1270 gnd d1 a_73513_n4475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1271 a_12177_14240# a_13017_14236# a_13225_14236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1272 a_39384_n14033# a_39641_n14223# a_39341_n12588# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1273 a_41619_3945# a_41623_3089# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1274 a_77243_n6712# a_76822_n6712# a_76414_n7028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 a_41618_7680# a_41875_7490# a_40570_7684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1276 a_79316_n4429# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1277 a_33429_14238# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1278 a_76151_6212# a_76152_5598# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1279 gnd a_20205_11212# a_19997_11212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_55570_n6710# a_55149_n6710# a_54741_n6631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1281 vdd d0 a_9757_n6765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1282 a_65446_11356# a_65446_10961# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1283 a_47397_n11874# a_48257_n8839# a_48465_n8839# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1284 a_66273_3822# a_67113_3818# a_67321_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1285 a_22313_12226# a_22934_12118# a_23142_12118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1286 gnd d1 a_19415_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1287 vdd d0 a_20464_n5251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1288 a_54480_13128# a_55101_13561# a_55309_13561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1289 gnd d2 a_60839_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1290 a_55567_n11198# a_55146_n11198# a_54738_n11514# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1291 a_52632_n8022# a_52636_n8878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1292 a_11606_n10322# a_12227_n10430# a_12435_n10430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1293 a_57637_6103# a_57424_6103# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1294 a_54738_n10067# a_55359_n9751# a_55567_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1295 a_63337_n9622# a_63594_n9812# a_62293_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1296 a_33022_10955# a_33643_11271# a_33851_11271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1297 a_13483_n9755# a_13062_n9755# a_12435_n10430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1298 a_45649_12795# a_45228_12795# a_44601_12799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1299 gnd a_52626_6051# a_52418_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1300 a_33430_9824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1301 a_25841_n5868# a_25477_n7390# a_24451_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1302 a_641_11358# a_641_10963# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1303 vdd a_63596_n5930# a_63388_n5930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1304 a_19947_12243# a_20204_12053# a_18899_12247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1305 a_68862_n11876# a_68649_n11876# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1306 a_28418_9964# a_29914_9094# a_29865_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1307 vdd a_9494_8177# a_9286_8177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1308 a_1306_n10424# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1309 a_85013_n7262# a_85017_n8207# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1310 a_46887_4587# a_46674_4587# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1311 a_29864_12251# a_30961_12057# a_30916_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1312 a_14881_n5753# a_14511_n4427# a_13485_n3747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1313 vdd d0 a_42136_n14907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1314 a_74309_n8201# a_74305_n8024# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1315 a_39347_n6757# a_39434_n5248# a_39385_n5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 a_3846_n5866# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1317 a_23193_n13393# a_22980_n13393# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1318 a_2516_3820# a_2095_3820# a_1468_3824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1319 vdd a_20462_n11938# a_20254_n11938# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1320 a_44031_n12633# a_44652_n12712# a_44860_n12712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1321 a_11080_986# a_15705_5267# a_16027_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 a_12016_n3743# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1323 a_69930_n8841# a_69717_n8841# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1324 a_33849_5263# a_33428_5263# a_33020_4947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1325 a_73256_n5732# a_74353_n5926# a_74304_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1326 a_638_7922# a_1259_8238# a_1467_8238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1327 vdd a_31428_n14222# a_31220_n14222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1328 gnd d1 a_30119_7500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1329 a_8454_n14882# a_8707_n14895# a_7003_n14025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1330 vdd d2 a_72067_n8209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1331 a_45227_5267# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1332 a_84757_9776# a_84753_9953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1333 a_45440_3820# a_45227_3820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1334 vdd d1 a_83961_12055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1335 a_11347_4153# a_11347_3897# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1336 a_9239_14375# a_9243_13519# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1337 a_66273_3143# a_65852_3143# a_65446_3152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1338 a_8191_12253# a_8448_12063# a_6744_12933# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1339 vdd d0 a_42137_n3806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1340 a_41881_n8709# a_42138_n8899# a_40833_n8705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1341 vdd a_8446_6055# a_8238_6055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1342 a_76413_n5113# a_76413_n5508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1343 a_68391_12115# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1344 gnd d0 a_63334_7492# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1345 a_1307_n14159# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1346 a_62036_10550# a_62289_10537# a_60589_9783# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1347 a_62033_6062# a_63126_6724# a_63077_6914# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1348 a_71814_n8196# a_73306_n7442# a_73261_n7429# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1349 a_34109_n14846# a_33688_n14846# a_32239_n15022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1350 a_19162_n14888# a_19415_n14901# a_17711_n14031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1351 a_76774_14238# a_76561_14238# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1352 a_640_13675# a_640_13134# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1353 a_56147_8228# a_55934_8228# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1354 a_34898_12787# a_36137_13554# a_36294_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1355 a_24451_n8157# a_24030_n8157# a_23403_n8832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1356 a_27567_n9609# a_28682_n12772# a_28633_n12582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1357 a_45649_14242# a_46888_13562# a_47045_12236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_66535_n7385# a_66114_n7385# a_65706_n7277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1359 a_66272_6789# a_65851_6789# a_65443_6868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1360 a_56407_n11202# a_56194_n11202# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1361 a_2775_n9749# a_2354_n9749# a_1727_n10424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1362 a_20208_n8028# a_20212_n8884# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1363 a_33020_3500# a_33020_3245# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1364 a_14464_13556# a_14251_13556# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1365 gnd d0 a_85268_n13460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1366 gnd a_85008_4523# a_84800_4523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1367 a_68608_n4423# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1368 a_11347_3502# a_11968_3818# a_12176_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1369 a_33282_n8080# a_33903_n8159# a_34111_n8159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 gnd a_52886_n10485# a_52678_n10485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1371 a_7008_n5227# a_7261_n5240# a_6966_n6749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1372 a_65445_14323# a_65445_13928# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1373 vdd a_20205_11212# a_19997_11212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1374 a_83962_n11746# a_84219_n11936# a_82515_n11066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1375 a_33282_n6377# a_33902_n5871# a_34110_n5871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1376 a_78082_n5196# a_77869_n5196# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1377 vdd d0 a_31428_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1378 a_55148_n4422# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1379 a_33282_n8730# a_33279_n9418# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1380 a_30910_6239# a_31167_6049# a_29862_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1381 gnd d0 a_31169_12736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1382 a_76414_n7824# a_77035_n7391# a_77243_n7391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1383 a_1260_3145# a_1047_3145# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1384 a_25680_12115# a_26538_9142# a_26746_9142# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1385 a_13484_n14169# a_13063_n14169# a_12436_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1386 gnd a_30120_3086# a_29912_3086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 a_81147_8368# a_82262_5205# a_82213_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 vdd a_9754_n10485# a_9546_n10485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1389 gnd d1 a_62549_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 a_73260_n5909# a_74353_n5247# a_74308_n5234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1391 a_23194_n4418# a_22981_n4418# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1392 a_82257_12925# a_83753_12055# a_83704_12245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1393 gnd d0 a_9756_n4477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1394 gnd d0 a_52887_n14220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1395 a_82522_n8202# a_82775_n8215# a_82475_n6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1396 a_48465_n8839# a_48938_n5926# a_48780_n5913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1397 a_31170_n10297# a_31174_n11242# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1398 a_65705_n5502# a_66326_n5186# a_66534_n5186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1399 vdd a_52626_6051# a_52418_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1400 gnd d7 a_21789_n1634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1401 a_6743_3958# a_8239_3088# a_8190_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1402 a_11969_12793# a_11756_12793# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1403 a_23192_n11194# a_22979_n11194# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1404 a_22720_4590# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1405 a_44651_n11871# a_44438_n11871# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1406 a_55147_n12718# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1407 a_76819_n10432# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1408 a_36646_n11882# a_37506_n8847# a_37714_n8847# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1409 a_51587_n4460# a_51840_n4473# a_50140_n5227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1410 a_57897_n11880# a_57684_n11880# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1411 a_46929_6109# a_46716_6109# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1412 a_83964_n4291# a_84221_n4481# a_82521_n5235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1413 a_36547_n11882# a_36183_n13404# a_35157_n12724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1414 gnd a_70956_n9799# a_70748_n9799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1415 gnd d0 a_63594_n9812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1416 gnd d1 a_40827_6047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1417 a_33643_9145# a_33430_9145# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1418 a_52630_n13262# a_52887_n13452# a_51582_n13258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1419 a_40834_n11923# a_41087_n11936# a_39383_n11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1420 a_54887_5265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1421 a_41624_12743# a_41620_12920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1422 a_46934_n13396# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1423 a_83964_n4291# a_85061_n4485# a_85016_n4472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1424 a_71550_9964# a_73046_9094# a_73001_9107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1425 a_13278_n6714# a_13065_n6714# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1426 a_12804_14236# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1427 a_85010_n10303# a_85014_n11248# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1428 a_63079_13690# a_63083_12745# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1429 a_33640_7551# a_33427_7551# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1430 a_63344_n6758# a_63597_n6771# a_62296_n7433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1431 gnd a_21789_n1634# a_21581_n1634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1432 a_76154_11606# a_76154_11350# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1433 a_34111_n8159# a_33690_n8159# a_33282_n8080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1434 a_66534_n3739# a_66113_n3739# a_65705_n3660# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1435 gnd a_81319_n5934# a_81111_n5934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1436 a_1728_n14838# a_1307_n14838# a_899_n14730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1437 a_76982_12791# a_76561_12791# a_76153_12870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1438 gnd d0 a_42135_n11940# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1439 a_4059_n5866# a_3846_n5866# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1440 a_9244_11231# a_9240_11408# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1441 a_67373_n14165# a_67160_n14165# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1442 vdd a_74562_n6767# a_74354_n6767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1443 a_66275_9151# a_67115_9826# a_67323_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1444 a_52629_n11063# a_52633_n11919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1445 a_54888_13561# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1446 a_68716_6226# a_68346_7552# a_67320_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1447 a_29866_6066# a_30959_6728# a_30914_6741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1448 vdd d5 a_16514_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1449 a_24030_n8157# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1450 a_76413_n4061# a_77034_n3745# a_77242_n3745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1451 a_21816_973# a_43041_941# a_3058_n1106# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1452 a_641_10963# a_641_10708# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1453 a_85015_n14894# a_85268_n14907# a_83963_n14713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1454 a_65703_n11765# a_65704_n12379# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1455 a_51322_3278# a_52419_3084# a_52370_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1456 a_74049_11229# a_74302_11216# a_73001_10554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1457 a_12436_n14844# a_12015_n14844# a_11607_n14736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1458 a_2517_12795# a_3756_13562# a_3913_12236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1459 a_11607_n13289# a_12228_n13397# a_12436_n13397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1460 a_62033_6062# a_63126_6724# a_63081_6737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1461 a_12435_n9751# a_12014_n9751# a_11606_n10067# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1462 a_65444_5604# a_65444_5348# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1463 a_44602_11279# a_44181_11279# a_43773_10963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1464 a_22314_10165# a_22935_10598# a_23143_10598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1465 a_76153_12475# a_76153_12220# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1466 a_7006_n11235# a_7259_n11248# a_6964_n12757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 vdd a_62548_n5926# a_62340_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1468 a_40833_n7258# a_41090_n7448# a_39390_n8202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1469 vdd a_50349_n12770# a_50141_n12770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1470 a_57899_n5872# a_57686_n5872# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1471 a_40570_6237# a_40827_6047# a_39123_6917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1472 a_56196_n5194# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1473 a_22719_8236# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1474 a_8193_7515# a_9286_8177# a_9241_8190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1475 gnd d0 a_41876_3755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1476 a_74042_7686# a_74046_6741# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1477 vdd a_85008_4523# a_84800_4523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1478 a_50137_n8017# a_50394_n8207# a_50094_n6572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1479 a_69802_5271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1480 a_33428_3137# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1481 vdd a_62546_n10487# a_62338_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1482 a_1307_n13391# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1483 a_44859_n9745# a_45699_n9749# a_45907_n9749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1484 a_1519_n11192# a_1306_n11192# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1485 vdd a_42136_n13460# a_41928_n13460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1486 a_20207_n3614# a_20464_n3804# a_19163_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1487 gnd d1 a_8449_9096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1488 a_34899_11267# a_34478_11267# a_33851_11271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1489 a_74305_n7256# a_74309_n8201# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1490 vdd d0 a_31169_12736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1491 vdd d0 a_42135_n11261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1492 vdd a_7000_3768# a_6792_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1493 a_71767_n6574# a_71859_n8209# a_71814_n8196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1494 a_45910_n6708# a_45489_n6708# a_44862_n7383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1495 vdd a_20463_n14905# a_20255_n14905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1496 vdd a_30120_3086# a_29912_3086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1497 vdd a_82772_n11256# a_82564_n11256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1498 a_73258_n11917# a_74351_n11255# a_74302_n11065# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1499 a_82257_12925# a_83753_12055# a_83708_12068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1500 gnd a_20204_14179# a_19996_14179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1501 a_79269_13554# a_79056_13554# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1502 a_40836_n4468# a_41929_n3806# a_33281_n3410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1503 a_55359_n10430# a_55146_n10430# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1504 a_6704_5226# a_6791_6735# a_6742_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1505 gnd d2 a_17709_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1506 a_85011_n14038# a_85268_n14228# a_83967_n14890# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1507 a_30913_9959# a_31170_9769# a_29869_9107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1508 a_44441_n7383# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1509 a_12175_6106# a_11754_6106# a_11347_5600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1510 gnd a_31429_n5926# a_31221_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1511 a_57424_6103# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1512 a_77033_n12720# a_76820_n12720# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1513 a_34690_12787# a_34477_12787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1514 gnd d1 a_30122_10541# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1515 vdd d2 a_28932_n11250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1516 gnd a_38532_n9805# a_38324_n9805# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1517 a_77241_n13399# a_76820_n13399# a_76412_n13832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1518 a_46675_13562# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1519 a_8454_n13435# a_9547_n12773# a_9498_n12583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1520 a_51323_12253# a_52420_12059# a_52375_12072# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1521 a_45700_n14163# a_45487_n14163# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1522 a_23403_n8153# a_22982_n8153# a_22574_n8469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1523 a_55310_9147# a_56150_9822# a_56358_9822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1524 a_31177_n8880# a_31173_n8703# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1525 gnd d2 a_39640_n11256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1526 a_54738_n10322# a_55359_n10430# a_55567_n10430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1527 a_2515_8234# a_2094_8234# a_1467_7559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1528 a_72999_4546# a_73252_4533# a_71552_3779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1529 a_1727_n9745# a_1306_n9745# a_898_n10061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1530 gnd a_85270_n7452# a_85062_n7452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1531 a_33689_n5871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1532 a_24241_n12718# a_24028_n12718# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1533 a_14725_n7394# a_14512_n7394# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1534 a_46674_4587# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1535 a_29868_12074# a_30961_12736# a_30912_12926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1536 a_1728_n13391# a_2568_n12716# a_2776_n12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1537 a_66064_7557# a_65851_7557# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1538 a_43772_14325# a_44393_14246# a_44601_14246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1539 a_1470_11279# a_1049_11279# a_641_11358# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1540 a_22932_7557# a_22719_7557# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1541 a_76411_n11516# a_77032_n11200# a_77240_n11200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1542 gnd d0 a_63595_n13458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1543 a_12176_4586# a_11755_4586# a_11347_4153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1544 a_11969_14240# a_11756_14240# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1545 vdd d2 a_82512_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1546 a_44654_n8830# a_44441_n8830# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1547 a_33848_6783# a_33427_6783# a_33019_6467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1548 a_54480_12222# a_55101_12114# a_55309_12114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1549 a_51322_3278# a_52419_3084# a_52374_3097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1550 a_74045_11406# a_74302_11216# a_73001_10554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1551 a_34111_n7391# a_33690_n7391# a_33282_n7824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1552 a_23768_5265# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1553 a_26538_9142# a_26325_9142# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 a_34110_n5871# a_34950_n5196# a_35158_n5196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1555 a_1261_12120# a_1048_12120# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1556 a_57594_7548# a_57381_7548# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1557 a_23195_n6706# a_22982_n6706# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1558 a_23981_3818# a_23768_3818# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1559 gnd d0 a_9757_n6765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1560 a_25688_n13398# a_25475_n13398# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1561 a_44440_n3737# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1562 vdd a_31429_n5247# a_31221_n5247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1563 vdd a_63594_n11938# a_63386_n11938# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1564 a_51326_3101# a_51579_3088# a_49875_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1565 a_33901_n14167# a_33688_n14167# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1566 vdd d1 a_51839_n14895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1567 a_44599_6112# a_44178_6112# a_43770_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1568 a_14507_12111# a_14294_12111# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1569 a_8452_n8697# a_8709_n8887# a_7005_n8017# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1570 a_13224_3814# a_12803_3814# a_12176_3139# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 a_14509_n10435# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1572 gnd a_63334_7492# a_63126_7492# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1573 a_34688_8226# a_34475_8226# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1574 vdd d0 a_41876_3755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1575 a_45648_3820# a_46887_4587# a_47038_6109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1576 a_77870_n6716# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1577 a_2310_9828# a_2097_9828# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1578 gnd a_63596_n5930# a_63388_n5930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1579 a_2518_11275# a_2097_11275# a_1470_11279# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1580 a_34897_3812# a_36136_4579# a_36287_6101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1581 a_11346_8311# a_11967_8232# a_12175_8232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1582 a_80586_9136# a_80165_9136# a_79518_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1583 a_35158_n3749# a_34737_n3749# a_34110_n3745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1584 a_82258_9958# a_82515_9768# a_82215_11403# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1585 a_34735_n11204# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 gnd a_85269_n3806# a_85061_n3806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 a_22722_11277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1588 a_85010_n9624# a_85267_n9814# a_83966_n10476# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1589 vdd a_42137_n4485# a_41929_n4485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1590 a_38019_8191# a_39132_11213# a_39083_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1591 a_70223_5271# a_69802_5271# a_70124_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1592 a_44601_12120# a_44180_12120# a_43772_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1593 a_44032_n5500# a_44653_n5184# a_44861_n5184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1594 a_55570_n8157# a_55149_n8157# a_54741_n8473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_33688_n12720# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1596 a_70439_8374# a_71554_5211# a_71505_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1597 a_72994_6243# a_74091_6049# a_74042_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1598 a_52369_8367# a_52373_7511# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1599 a_25680_12115# a_25259_12115# a_25586_12234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1600 gnd a_20462_n11938# a_20254_n11938# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1601 vdd d0 a_9756_n5924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1602 a_6704_5226# a_6791_6735# a_6746_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1603 a_56410_n8161# a_56197_n8161# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1604 vdd d0 a_52889_n7444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1605 a_30914_6741# a_31167_6728# a_29866_6066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_34110_n3745# a_33689_n3745# a_33281_n4061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1607 a_27567_n9609# a_27824_n9799# a_27222_n5738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1608 a_4017_n7388# a_3804_n7388# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1609 a_1048_13567# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1610 a_54212_986# a_58837_5267# a_58913_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1611 vdd d1 a_30122_10541# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1612 vdd d1 a_8446_7502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1613 vdd d2 a_17967_n11254# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1614 vdd d1 a_8708_n4473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1615 a_65443_8571# a_65443_8315# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1616 a_33643_11271# a_33430_11271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1617 a_65852_3822# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1618 a_74303_n13264# a_74560_n13454# a_73255_n13260# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1619 a_640_13930# a_1261_14246# a_1469_14246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1620 a_51581_n10291# a_51838_n10481# a_50138_n11235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1621 a_46716_6109# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1622 a_55362_n6710# a_55149_n6710# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1623 a_79270_10587# a_79057_10587# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1624 a_638_7667# a_638_7126# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1625 gnd a_40827_6047# a_40619_6047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1626 a_76983_11271# a_76562_11271# a_76154_10955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1627 a_45486_n9749# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1628 a_33430_9145# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1629 gnd a_20465_n8897# a_20257_n8897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1630 a_72995_4723# a_73252_4533# a_71552_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1631 a_24449_n12718# a_24028_n12718# a_23401_n13393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1632 a_11967_7553# a_11754_7553# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1633 a_22311_6473# a_22311_6218# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1634 a_25475_n13398# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1635 vdd a_63596_n5251# a_63388_n5251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1636 a_63344_n6758# a_63340_n6581# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1637 vdd a_72066_n5242# a_71858_n5242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1638 a_20207_n4293# a_20211_n5238# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1639 a_4005_6109# a_4865_9144# a_5073_9144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1640 gnd d4 a_49023_8186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1641 a_29868_12074# a_30961_12736# a_30916_12749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1642 a_76559_8230# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1643 a_54740_n4855# a_55361_n4422# a_55569_n4422# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1644 a_62289_n11744# a_63386_n11938# a_63341_n11925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1645 a_23400_n10426# a_22979_n10426# a_22571_n10859# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1646 a_63339_n4293# a_63596_n4483# a_62291_n4289# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1647 gnd d0 a_9494_8177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1648 gnd d0 a_31430_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_6749_9789# a_8241_10543# a_8192_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1650 a_44394_10600# a_44181_10600# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1651 a_74042_6918# a_74299_6728# a_72998_6066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1652 a_1469_12799# a_1048_12799# a_640_12878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1653 a_17455_3775# a_18947_4529# a_18898_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1654 a_17414_11228# a_17501_12737# a_17452_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1655 a_22934_13565# a_22721_13565# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1656 a_11346_8311# a_11346_7916# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1657 a_83966_n11923# a_84219_n11936# a_82515_n11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1658 vdd a_82470_5205# a_82262_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1659 a_13015_6781# a_12802_6781# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1660 gnd d0 a_31428_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1661 vdd a_20462_n11259# a_20254_n11259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1662 a_41619_3266# a_33022_3146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1663 a_74047_5221# a_74300_5208# a_72999_4546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1664 a_43773_11358# a_43773_10963# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1665 a_84751_5392# a_85008_5202# a_83707_4540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1666 a_33019_7118# a_33640_7551# a_33848_7551# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1667 a_641_9516# a_1262_9832# a_1470_9832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1668 gnd a_9754_n10485# a_9546_n10485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1669 a_73260_n5909# a_74353_n5247# a_74304_n5057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1670 vdd a_52888_n3798# a_52680_n3798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1671 gnd d1 a_19154_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1672 gnd a_30381_n5922# a_30173_n5922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1673 vdd a_83959_6047# a_83751_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1674 a_25844_n11757# a_25730_n11876# a_25938_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1675 a_34949_n14171# a_34736_n14171# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1676 gnd a_30380_n14897# a_30172_n14897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1677 a_78291_n8163# a_79530_n7396# a_79681_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1678 gnd a_73514_n7442# a_73306_n7442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1679 a_82255_6917# a_83751_6047# a_83702_6237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1680 a_55569_n4422# a_56409_n3747# a_56617_n3747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1681 gnd d2 a_28672_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1682 a_29868_12074# a_30121_12061# a_28417_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1683 a_13485_n3747# a_14724_n4427# a_14881_n5753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1684 gnd a_41877_12730# a_41669_12730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1685 a_30910_6918# a_30914_6062# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1686 a_44602_9832# a_44181_9832# a_43773_9911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1687 vdd a_20465_n8218# a_20257_n8218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1688 a_62029_6239# a_63126_6045# a_63077_6235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1689 a_33848_8230# a_33427_8230# a_33019_8309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1690 a_34109_n14167# a_33688_n14167# a_33280_n14483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1691 gnd a_41876_3755# a_41668_3755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1692 a_55568_n14844# a_55147_n14844# a_54739_n14736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1693 a_54739_n13289# a_55360_n13397# a_55568_n13397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1694 a_83964_n4291# a_85061_n4485# a_85012_n4295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1695 a_17716_n5233# a_19208_n4479# a_19163_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1696 a_38019_8191# a_39132_11213# a_39087_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1697 a_43771_3253# a_43773_3154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1698 a_36554_n5755# a_36184_n4429# a_35158_n5196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1699 a_23982_12793# a_23769_12793# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1700 a_56358_11269# a_55937_11269# a_55310_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1701 a_70439_8374# a_71554_5211# a_71509_5224# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1702 a_54888_12114# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1703 a_22311_6218# a_22932_6110# a_23140_6110# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1704 vdd d0 a_31430_n8214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1705 a_73255_n14707# a_74352_n14901# a_74307_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1706 a_66272_6110# a_65851_6110# a_65443_6218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1707 a_66324_n9747# a_66111_n9747# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1708 a_24450_n5190# a_24029_n5190# a_23402_n5186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1709 a_23402_n4418# a_22981_n4418# a_22573_n4310# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1710 a_45909_n5188# a_45488_n5188# a_44861_n5863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_11349_3148# a_11968_3139# a_12176_3139# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1712 a_81147_8368# a_81404_8178# a_80832_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1713 a_11609_n7822# a_11609_n8078# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1714 a_54478_6214# a_54479_5600# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1715 a_78031_9820# a_77610_9820# a_76983_9145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1716 a_34691_11267# a_34478_11267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1717 a_17715_n14208# a_19207_n13454# a_19162_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1718 gnd a_74562_n6767# a_74354_n6767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 a_79518_6101# a_79097_6101# a_79419_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1720 a_76772_7551# a_76559_7551# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1721 a_36185_n7396# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1722 a_33281_n5508# a_33902_n5192# a_34110_n5192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1723 a_33687_n10432# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1724 a_44032_n4053# a_44032_n4308# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1725 a_15918_5267# a_15705_5267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1726 gnd a_61100_n14221# a_60892_n14221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1727 a_76822_n8838# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1728 a_13064_n3747# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1729 gnd d0 a_31169_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1730 vdd a_39600_n6770# a_39392_n6770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1731 a_35965_6101# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_84756_13511# a_85009_13498# a_83704_13692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 a_19949_7505# a_19945_7682# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1734 a_1727_n10424# a_1306_n10424# a_898_n10857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1735 a_43772_13675# a_43772_13134# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1736 gnd d1 a_51581_10543# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1737 a_77241_n12720# a_78081_n12724# a_78289_n12724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1738 a_54481_10161# a_55102_10594# a_55310_10594# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1739 a_81407_n9615# a_82522_n12778# a_82477_n12765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1740 a_49836_5226# a_50089_5213# a_48766_8376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1741 a_25217_10593# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1742 vdd a_63595_n14905# a_63387_n14905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1743 a_1468_4592# a_2308_5267# a_2516_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1744 a_8195_13523# a_8448_13510# a_6748_12756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1745 a_1730_n8830# a_1309_n8830# a_901_n8722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1746 gnd d1 a_30121_13508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1747 a_35156_n9757# a_36395_n10437# a_36552_n11763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1748 a_56618_n6714# a_57857_n7394# a_58008_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1749 a_22573_n5757# a_22574_n6371# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1750 a_31175_n14888# a_31428_n14901# a_30123_n14707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1751 a_76822_n6712# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1752 a_30917_9103# a_31170_9090# a_29865_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1753 a_44651_n11192# a_44438_n11192# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1754 a_68711_6107# a_68347_4585# a_67321_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1755 a_22312_4698# a_22933_4590# a_23141_4590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1756 gnd a_62548_n5926# a_62340_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1757 vdd d4 a_49023_8186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1758 a_40837_n7435# a_41090_n7448# a_39390_n8202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1759 gnd a_50349_n12770# a_50141_n12770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1760 vdd a_39642_n5248# a_39434_n5248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1761 a_36136_4579# a_35923_4579# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1762 a_47148_n4421# a_46935_n4421# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1763 a_52373_7511# a_52369_7688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1764 a_51327_12076# a_52420_12738# a_52371_12928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_55936_12789# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1766 a_27567_n9609# a_28682_n12772# a_28637_n12759# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1767 a_6749_9789# a_8241_10543# a_8196_10556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1768 gnd a_51581_10543# a_51373_10543# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_34736_n14171# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1770 a_34735_n9757# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1771 gnd d1 a_73513_n5922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1772 gnd a_62546_n10487# a_62338_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1773 a_45701_n5188# a_45488_n5188# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1774 a_54479_3897# a_54479_3502# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1775 a_33850_14238# a_33429_14238# a_33021_13922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1776 a_13062_n11202# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1777 a_24029_n3743# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1778 gnd a_42136_n13460# a_41928_n13460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1779 a_23980_8232# a_23767_8232# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1780 vdd a_82512_6727# a_82304_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1781 a_63081_8184# a_63334_8171# a_62033_7509# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1782 a_1728_n14159# a_1307_n14159# a_899_n14080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1783 a_76982_12112# a_76561_12112# a_76153_12220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1784 a_67321_3818# a_66900_3818# a_66273_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1785 gnd d1 a_19415_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1786 gnd d0 a_85009_12730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1787 a_57753_12230# a_57639_12111# a_57847_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1788 gnd a_82772_n11256# a_82564_n11256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1789 a_62292_n7256# a_62549_n7446# a_60849_n8200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1790 a_65445_12226# a_65446_11612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1791 a_26325_9142# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1792 a_57381_7548# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1793 a_67373_n12718# a_67160_n12718# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1794 a_63083_13513# a_63336_13500# a_62031_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1795 a_33282_n6633# a_33282_n7028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1796 a_29862_6243# a_30959_6049# a_30914_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1797 a_65443_7920# a_66064_8236# a_66272_8236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1798 a_12438_n8157# a_13278_n8161# a_13486_n8161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1799 a_11609_n7281# a_12230_n7389# a_12438_n7389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1800 a_84754_6735# a_85007_6722# a_83706_6060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1801 a_66532_n11194# a_67372_n11198# a_67580_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1802 a_54311_986# a_53890_986# a_54212_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1803 vdd d2 a_28672_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1804 a_85015_n14215# a_85268_n14228# a_83967_n14890# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1805 a_29864_12251# a_30121_12061# a_28417_12931# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1806 a_12436_n14165# a_12015_n14165# a_11607_n14086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1807 a_51583_n4283# a_51840_n4473# a_50140_n5227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1808 gnd a_50091_11221# a_49883_11221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1809 vdd a_41877_12730# a_41669_12730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1810 a_8192_10733# a_9289_10539# a_9244_10552# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1811 a_19947_13690# a_20204_13500# a_18899_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1812 a_19952_9099# a_19948_9276# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1813 a_62029_6239# a_63126_6045# a_63081_6058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1814 a_34475_8226# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1815 gnd d2 a_28932_n11250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1816 a_44438_n9745# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 vdd a_41876_3755# a_41668_3755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1818 a_85010_n9624# a_85014_n10480# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1819 a_34898_14234# a_34477_14234# a_33850_13559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1820 a_51583_n4283# a_52680_n4477# a_52635_n4464# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1821 a_14552_n11880# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1822 gnd d0 a_31167_8175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1823 gnd d5 a_59646_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1824 a_34899_9820# a_36138_10587# a_36289_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1825 a_44181_11279# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1826 vdd d0 a_74299_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1827 a_2310_11275# a_2097_11275# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1828 a_11346_7916# a_11346_7661# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1829 a_48550_5273# a_48129_5273# a_48451_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1830 a_12437_n4422# a_12016_n4422# a_11608_n4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_62290_n14711# a_63387_n14905# a_63342_n14892# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1832 a_23193_n14840# a_22980_n14840# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1833 gnd d0 a_41876_3076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1834 a_33020_4151# a_33020_3895# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1835 a_62033_6062# a_62286_6049# a_60582_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1836 a_63340_n6581# a_63597_n6771# a_62296_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1837 a_13486_n6714# a_13065_n6714# a_12438_n7389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1838 a_23401_n13393# a_22980_n13393# a_22572_n13826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1839 a_43773_10963# a_43773_10708# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1840 a_14465_10589# a_14252_10589# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1841 a_68562_10593# a_68349_10593# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1842 a_82213_5395# a_82305_3760# a_82256_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1843 a_33641_5263# a_33428_5263# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1844 a_30912_12247# a_31169_12057# a_29864_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1845 a_74302_n10297# a_74306_n11242# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1846 a_76154_10955# a_76775_11271# a_76983_11271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1847 a_55568_n13397# a_56408_n12722# a_56616_n12722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1848 vdd d6 a_75558_n1647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1849 a_68973_n5868# a_68609_n7390# a_67583_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1850 a_2568_n14163# a_2355_n14163# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1851 a_3058_n1106# a_42828_941# a_43150_941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1852 vdd d1 a_51581_10543# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1853 a_77867_n11204# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 vdd d1 a_83961_13502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1855 a_12227_n11877# a_12014_n11877# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1856 a_66325_n14161# a_66112_n14161# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1857 a_49832_5403# a_50089_5213# a_48766_8376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1858 a_58107_n5872# a_57686_n5872# a_58008_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1859 a_55102_11273# a_54889_11273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1860 a_8191_13700# a_8448_13510# a_6748_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1861 a_14511_n4427# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1862 vdd a_8446_7502# a_8238_7502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1863 a_9241_7511# a_9494_7498# a_8189_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1864 a_63341_n10478# a_63594_n10491# a_62289_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1865 a_73000_13521# a_74093_14183# a_74044_14373# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1866 a_45229_11275# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1867 a_23982_14240# a_23769_14240# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1868 a_39384_n14033# a_40880_n14903# a_40835_n14890# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1869 a_1521_n5863# a_1308_n5863# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1870 gnd a_31429_n5247# a_31221_n5247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1871 gnd a_63594_n11938# a_63386_n11938# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1872 a_34951_n8163# a_34738_n8163# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1873 a_55307_7553# a_54886_7553# a_54478_7661# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1874 a_76981_3816# a_76560_3816# a_76152_3895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1875 a_22311_8571# a_22935_9151# a_23143_9151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1876 a_8456_n8874# a_8709_n8887# a_7005_n8017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1877 a_23142_13565# a_22721_13565# a_22313_13673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1878 vdd a_9756_n3798# a_9548_n3798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1879 vdd d1 a_19157_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1880 a_52375_14198# a_54480_14319# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1881 a_11754_7553# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1882 vdd a_51581_10543# a_51373_10543# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1883 a_66535_n8832# a_66114_n8832# a_65706_n8724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1884 a_1730_n8151# a_2570_n8155# a_2778_n8155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1885 a_65445_13673# a_66066_13565# a_66274_13565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1886 a_33022_10700# a_33022_10159# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1887 gnd d0 a_85268_n14907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1888 a_39081_5395# a_39338_5205# a_38015_8368# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1889 gnd a_49023_8186# a_48815_8186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1890 a_83969_n7435# a_85062_n6773# a_85013_n6583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1891 a_56356_3814# a_55935_3814# a_55308_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1892 a_63079_14369# a_63083_13513# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1893 gnd a_9494_8177# a_9286_8177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1894 a_21532_n1444# a_32218_n1647# a_27321_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1895 a_18899_13694# a_19996_13500# a_19947_13690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1896 gnd a_52886_n11932# a_52678_n11932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1897 a_63077_8361# a_63334_8171# a_62033_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1898 a_76412_n12385# a_77032_n11879# a_77240_n11879# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1899 a_44032_n3658# a_44032_n4053# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1900 gnd d1 a_40830_9088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 a_44393_13567# a_44180_13567# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1902 a_33689_n5192# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1903 gnd a_42137_n4485# a_41929_n4485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1904 a_85014_n9801# a_85267_n9814# a_83966_n10476# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1905 a_57847_12111# a_57426_12111# a_57753_12230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1906 a_23403_n6706# a_22982_n6706# a_22574_n6627# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1907 vdd d0 a_85009_12730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1908 a_22573_n3404# a_31429_n3800# a_30128_n4462# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1909 a_29864_12251# a_30961_12057# a_30912_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 vdd d2 a_17707_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1911 a_1260_4592# a_1047_4592# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1912 vdd d0 a_85269_n3806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1913 gnd a_30120_4533# a_29912_4533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1914 a_34689_5259# a_34476_5259# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1915 a_85013_n8709# a_85270_n8899# a_83965_n8705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1916 a_12436_n14165# a_13276_n14169# a_13484_n14169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1917 a_12802_6781# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1918 gnd d1 a_62549_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1919 a_24243_n6710# a_24030_n6710# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1920 gnd d0 a_9756_n5924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1921 a_54889_10594# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1922 a_22571_n10063# a_23192_n9747# a_23400_n9747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1923 vdd a_41088_n13456# a_40880_n13456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1924 a_1729_n4416# a_1308_n4416# a_900_n4849# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1925 a_84750_6912# a_85007_6722# a_83706_6060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1926 a_2778_n6708# a_2357_n6708# a_1730_n7383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1927 a_641_11614# a_641_11358# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1928 vdd a_52626_7498# a_52418_7498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1929 a_44654_n8151# a_44441_n8151# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1930 gnd d0 a_52889_n7444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1931 a_2517_14242# a_2096_14242# a_1469_13567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1932 gnd d4 a_16859_n9803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1933 a_24448_n9751# a_24027_n9751# a_23400_n9747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1934 a_66114_n7385# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1935 a_6747_3781# a_8239_4535# a_8190_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1936 vdd a_50091_11221# a_49883_11221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1937 gnd a_19154_7496# a_18946_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1938 a_1728_n13391# a_1307_n13391# a_899_n13824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1939 a_2518_9828# a_3757_10595# a_3908_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1940 gnd d2 a_17967_n11254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1941 a_83964_n5738# a_84221_n5928# a_82517_n5058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1942 a_68718_12234# a_68348_13560# a_67322_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1943 a_29869_9107# a_30962_9769# a_30917_9782# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1944 a_84753_9953# a_84757_9097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1945 a_76153_13126# a_76153_12870# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1946 a_49832_5403# a_49924_3768# a_49879_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1947 a_11967_6106# a_11754_6106# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 a_22721_14244# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1949 vdd d0 a_31167_8175# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1950 a_74307_n13441# a_74560_n13454# a_73255_n13260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1951 a_1309_n7383# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1952 vdd a_63594_n11259# a_63386_n11259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1953 a_8191_13700# a_9288_13506# a_9239_13696# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1954 a_8454_n13435# a_9547_n12773# a_9502_n12760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1955 a_2355_n14163# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1956 a_52371_12928# a_52375_12072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1957 gnd a_51840_n4473# a_51632_n4473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1958 vdd d0 a_41876_3076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1959 a_74042_8365# a_74046_7509# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1960 gnd d0 a_20462_n9812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1961 a_59474_8370# a_60589_5207# a_60540_5397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1962 vdd d0 a_85268_n14228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1963 vdd a_85270_n7452# a_85062_n7452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1964 a_68976_n11757# a_68862_n11876# a_69070_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1965 a_55569_n3743# a_55148_n3743# a_54740_n4059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1966 a_899_n14730# a_1520_n14838# a_1728_n14838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 a_25732_n5868# a_25519_n5868# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1968 a_82213_5395# a_82305_3760# a_82260_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1969 a_640_12483# a_640_12228# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1970 a_62289_n11744# a_63386_n11938# a_63337_n11748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1971 a_83708_12068# a_84801_12730# a_84752_12920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_56150_11269# a_55937_11269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1973 a_15833_n8845# a_15620_n8845# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1974 a_12017_n7389# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1975 a_33019_6212# a_33640_6104# a_33848_6104# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1976 a_66065_5269# a_65852_5269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1977 a_10758_986# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1978 a_1047_3824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1979 a_899_n13028# a_1520_n12712# a_1728_n12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1980 a_9498_n14030# a_9502_n14886# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1981 a_51322_4725# a_52419_4531# a_52370_4721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1982 a_11968_4586# a_11755_4586# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1983 a_15705_5267# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1984 vdd d0 a_9756_n5245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1985 gnd d1 a_73251_7500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1986 a_11607_n14736# a_12228_n14844# a_12436_n14844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1987 gnd a_20462_n11259# a_20254_n11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1988 a_73000_13521# a_74093_14183# a_74048_14196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1989 a_43771_5350# a_44392_5271# a_44600_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1990 a_30914_6062# a_31167_6049# a_29862_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1991 a_66113_n3739# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1992 a_56410_n6714# a_56197_n6714# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1993 gnd a_72022_n12772# a_71814_n12772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 a_1261_13567# a_1048_13567# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1995 a_55937_11269# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1996 a_84751_4713# a_84755_3768# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1997 a_40570_7684# a_41667_7490# a_41618_7680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1998 gnd a_85268_n12781# a_85060_n12781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1999 gnd d0 a_74300_3761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 a_22312_5348# a_22312_4953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2001 a_55148_n5869# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2002 a_25428_4585# a_25215_4585# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2003 gnd d0 a_20204_12732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2004 gnd d2 a_82773_n14223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2005 a_65852_3143# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2006 a_20205_n10301# a_20462_n10491# a_19157_n10297# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2007 a_56615_n9755# a_56194_n9755# a_55567_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2008 a_51588_n7427# a_52681_n6765# a_52636_n6752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2009 a_1308_n3737# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2010 vdd a_49023_8186# a_48815_8186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2011 a_53628_n1455# a_53885_n1645# a_53727_n1632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2012 a_13016_3814# a_12803_3814# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2013 a_82475_n6580# a_82732_n6770# a_81411_n9792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2014 gnd d4 a_6151_n9797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2015 a_70354_n5738# a_70611_n5928# a_70453_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2016 vdd a_62546_n11934# a_62338_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2017 a_40831_n14713# a_41088_n14903# a_39384_n14033# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2018 a_55361_n3743# a_55148_n3743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2019 a_28682_n8196# a_28935_n8209# a_28635_n6574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2020 a_66326_n5865# a_66113_n5865# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2021 a_9503_n4464# a_9499_n4287# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2022 gnd a_20465_n8218# a_20257_n8218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2023 a_33020_4692# a_33641_4584# a_33849_4584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2024 a_40577_10548# a_40830_10535# a_39130_9781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2025 a_17716_n5233# a_19208_n4479# a_19159_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2026 a_11347_5600# a_11347_5344# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2027 a_76562_11271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2028 a_67320_8232# a_66899_8232# a_66272_7557# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2029 a_54479_3502# a_55100_3818# a_55308_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2030 a_54480_12872# a_54480_12477# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2031 a_62293_n11921# a_63386_n11259# a_63341_n11246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2032 vdd a_30120_4533# a_29912_4533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2033 a_12176_5265# a_13016_5261# a_13224_5261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2034 gnd d0 a_9497_9771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2035 a_76772_6104# a_76559_6104# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2036 a_79424_6220# a_79054_7546# a_78028_6779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2037 gnd d0 a_52628_13506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2038 a_65851_6789# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2039 a_82261_12748# a_83753_13502# a_83708_13515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2040 gnd d0 a_31430_n8214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2041 a_25689_n4423# a_25476_n4423# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2042 a_74042_6239# a_74299_6049# a_72994_6243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2043 a_33850_13559# a_34690_14234# a_34898_14234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2044 a_1469_12120# a_1048_12120# a_640_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2045 a_6747_3781# a_8239_4535# a_8194_4548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2046 a_17715_n14208# a_19207_n13454# a_19158_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2047 a_84752_13688# a_84756_12743# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2048 a_44441_n8830# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2049 a_44862_n6704# a_45702_n6708# a_45910_n6708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2050 a_33849_3816# a_34689_3812# a_34897_3812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2051 a_77868_n14171# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2052 a_67580_n9751# a_68819_n10431# a_68976_n11757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2053 a_54741_n8473# a_54741_n8728# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2054 a_52632_n6575# a_52636_n7431# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2055 a_77032_n9753# a_76819_n9753# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2056 a_1468_3824# a_1047_3824# a_639_3903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2057 vdd d0 a_20203_5204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2058 vdd d1 a_40827_7494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2059 a_29866_6066# a_30959_6728# a_30910_6918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2060 a_50135_n14025# a_50392_n14215# a_50092_n12580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2061 gnd a_39600_n6770# a_39392_n6770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2062 a_30915_5221# a_30911_5398# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2063 a_638_8573# a_1262_9153# a_1470_9153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2064 a_81407_n9615# a_82522_n12778# a_82473_n12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2065 a_39341_n12588# a_39433_n14223# a_39384_n14033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2066 a_77241_n14846# a_76820_n14846# a_75371_n15022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2067 a_11349_10957# a_11970_11273# a_12178_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2068 a_41625_10544# a_41878_10531# a_40573_10725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2069 a_21717_973# a_21608_973# a_21816_973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2070 a_56357_14236# a_55936_14236# a_55309_13561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2071 a_65853_13565# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2072 a_19951_14192# a_22313_14323# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2073 a_3541_7554# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2074 a_41884_n4472# a_41880_n4295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2075 a_63083_13513# a_63079_13690# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2076 a_47298_n11874# a_47189_n11874# a_47397_n11874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2077 gnd a_31169_14183# a_30961_14183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2078 a_43771_3903# a_43771_3508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2079 a_78031_11267# a_77610_11267# a_76983_11271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2080 a_44179_5271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2081 a_44030_n11763# a_44651_n11871# a_44859_n11871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2082 a_76773_4584# a_76560_4584# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2083 a_901_n8072# a_1522_n8151# a_1730_n8151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2084 gnd a_31167_8175# a_30959_8175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2085 a_41622_8182# a_41618_8359# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2086 a_44392_3824# a_44179_3824# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2087 gnd d2 a_28674_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2088 a_11970_9826# a_11757_9826# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2089 a_9240_9282# a_9497_9092# a_8192_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2090 gnd a_39642_n5248# a_39434_n5248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2091 gnd a_41877_12051# a_41669_12051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2092 a_40574_6060# a_40827_6047# a_39123_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2093 a_83708_12068# a_84801_12730# a_84756_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2094 a_44602_9153# a_44181_9153# a_43773_9261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2095 a_68713_12115# a_68349_10593# a_67323_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2096 a_9240_9961# a_9244_9105# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2097 vdd a_73512_n14897# a_73304_n14897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2098 a_65703_n9412# a_65703_n9668# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2099 gnd a_41876_3076# a_41668_3076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2100 a_14463_4581# a_14250_4581# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2101 a_55568_n14165# a_55147_n14165# a_54739_n14086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2102 a_8193_7515# a_9286_8177# a_9237_8367# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2103 a_67583_n8157# a_67162_n8157# a_66535_n8153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2104 gnd d0 a_63595_n14905# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2105 gnd a_41089_n4481# a_40881_n4481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2106 a_22979_n9747# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2107 gnd a_42138_n6773# a_41930_n6773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2108 gnd a_40829_13502# a_40621_13502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2109 vdd d0 a_74560_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2110 a_3058_n1106# a_2944_n1225# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2111 a_55099_8232# a_54886_8232# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2112 a_44033_n8072# a_44033_n8467# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2113 a_70443_8197# a_70696_8184# a_70124_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2114 a_51322_4725# a_52419_4531# a_52374_4544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2115 a_16257_n5742# a_16651_n9803# a_16602_n9613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2116 a_34109_n13399# a_34949_n12724# a_35157_n12724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2117 a_77821_3812# a_77608_3812# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2118 a_30916_12749# a_31169_12736# a_29868_12074# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2119 a_79312_12109# a_79099_12109# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2120 vdd d0 a_9497_10539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2121 a_25839_n11876# a_25475_n13398# a_24449_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2122 gnd a_7000_3768# a_6792_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2123 a_62296_n7433# a_62549_n7446# a_60849_n8200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2124 a_79527_n10437# a_79314_n10437# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2125 a_62031_12247# a_62288_12057# a_60584_12927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2126 a_43770_8573# a_43770_8317# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2127 vdd a_30381_n5922# a_30173_n5922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2128 a_76980_8230# a_76559_8230# a_76151_7914# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2129 a_51326_4548# a_51579_4535# a_49879_3781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2130 vdd d0 a_74300_3761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2131 a_1049_10600# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2132 a_57856_n4427# a_57643_n4427# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2133 vdd d0 a_20204_12732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2134 a_41882_n10480# a_42135_n10493# a_40830_n10299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2135 a_76822_n8159# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2136 a_14876_n5872# a_14767_n5872# a_14975_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2137 vdd a_73514_n7442# a_73306_n7442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2138 a_25938_n11876# a_26798_n8841# a_27006_n8841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2139 a_76821_n5871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2140 a_77242_n3745# a_78082_n3749# a_78290_n3749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2141 a_69457_9142# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2142 a_30917_9782# a_31170_9769# a_29869_9107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2143 a_74305_n7256# a_74562_n7446# a_73257_n7252# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2144 a_83702_6237# a_83959_6047# a_82255_6917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2145 gnd d1 a_8706_n10481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2146 a_63080_10723# a_63084_9778# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2147 a_1730_n8151# a_1309_n8151# a_901_n8072# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2148 a_55359_n11877# a_55146_n11877# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2149 vdd a_19157_9090# a_18949_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2150 a_22311_7124# a_22311_6868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2151 a_31175_n14209# a_31428_n14222# a_30127_n14884# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2152 a_40573_10725# a_40830_10535# a_39130_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2153 vdd d0 a_85007_8169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2154 a_51583_n4283# a_52680_n4477# a_52631_n4287# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2155 vdd d0 a_63596_n3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2156 a_13225_12789# a_14464_13556# a_14621_12230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2157 vdd a_39640_n11256# a_39432_n11256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2158 a_30910_6239# a_30915_5221# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2159 a_13277_n5194# a_13064_n5194# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2160 a_65444_5348# a_66065_5269# a_66273_5269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2161 vdd d0 a_9497_9771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2162 a_41623_3768# a_41876_3755# a_40575_3093# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2163 a_12228_n13397# a_12015_n13397# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2164 a_63343_n5238# a_63596_n5251# a_62295_n5913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2165 a_51323_12253# a_52420_12059# a_52371_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2166 a_33430_10592# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2167 vdd d0 a_63595_n14226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2168 gnd a_8708_n4473# a_8500_n4473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2169 a_33280_n13832# a_33280_n14088# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2170 a_28375_11409# a_28632_11219# a_27311_8197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2171 a_34688_6779# a_34475_6779# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2172 a_23400_n11873# a_24240_n11198# a_24448_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2173 vdd d3 a_17927_n6768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2174 a_22573_n4310# a_23194_n4418# a_23402_n4418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2175 a_34476_5259# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2176 vdd d2 a_39643_n8215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2177 gnd d0 a_74301_14183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2178 a_44602_10600# a_45442_11275# a_45650_11275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2179 a_22311_7124# a_22932_7557# a_23140_7557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2180 a_20210_n13445# a_20206_n13268# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2181 gnd d6 a_75558_n1647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2182 a_22312_4953# a_22312_4698# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2183 vdd a_61100_n14221# a_60892_n14221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2184 a_54103_986# a_53890_986# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2185 gnd d2 a_82512_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2186 a_44030_n10857# a_44651_n10424# a_44859_n10424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2187 vdd d1 a_8708_n5920# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2188 gnd d0 a_85009_12051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2189 a_22574_n6371# a_22574_n6627# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2190 a_41621_10721# a_41878_10531# a_40573_10725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2191 a_55307_6106# a_54886_6106# a_54479_5600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2192 a_19952_9778# a_19948_9955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2193 a_23141_3143# a_23981_3818# a_24189_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2194 a_44180_14246# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2195 a_51581_n11738# a_51838_n11928# a_50134_n11058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2196 a_73258_n10470# a_73511_n10483# a_71811_n11237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2197 a_78290_n3749# a_77869_n3749# a_77242_n3745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2198 a_23142_12118# a_22721_12118# a_22314_11612# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 gnd d0 a_20202_6724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2200 a_54739_n13830# a_54739_n14086# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2201 a_62295_n4466# a_63388_n3804# a_63339_n3614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2202 a_56150_9822# a_55937_9822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2203 a_31173_n8703# a_31174_n9795# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2204 gnd d1 a_84221_n4481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2205 vdd a_31169_14183# a_30961_14183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2206 a_28375_11409# a_28467_9774# a_28418_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2207 a_5549_n5736# a_5943_n9797# a_5894_n9607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2208 vdd d2 a_17969_n5246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2209 a_84754_6056# a_85007_6043# a_83702_6237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2210 vdd d0 a_74562_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2211 a_11607_n12383# a_11607_n12639# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2212 a_11754_6106# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2213 a_14505_6103# a_14292_6103# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2214 vdd a_31167_8175# a_30959_8175# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2215 a_68978_n5749# a_68864_n5868# a_69072_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2216 vdd d2 a_28674_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2217 gnd a_74301_13504# a_74093_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2218 a_12438_n7389# a_13278_n6714# a_13486_n6714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2219 vdd a_84220_n13456# a_84012_n13456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2220 vdd a_41877_12051# a_41669_12051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2221 vdd a_41876_3076# a_41668_3076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2222 a_9497_n9616# a_9754_n9806# a_8453_n10468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2223 a_58105_n11880# a_58965_n8845# a_59173_n8845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2224 a_18904_9103# a_19997_9765# a_19948_9955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2225 a_33851_10592# a_33430_10592# a_33022_10159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2226 a_29865_9284# a_30962_9090# a_30913_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2227 a_63339_n5740# a_63596_n5930# a_62291_n5736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2228 a_4168_n5866# a_4059_n5866# a_4267_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2229 a_1259_6112# a_1046_6112# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2230 a_52376_9784# a_52372_9961# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2231 a_898_n11508# a_898_n11763# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2232 vdd d1 a_73513_n5922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2233 a_70439_8374# a_70696_8184# a_70124_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2234 a_44860_n14159# a_45700_n14163# a_45908_n14163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2235 a_34477_14234# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2236 a_67374_n5190# a_67161_n5190# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2237 a_55101_14240# a_54888_14240# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2238 a_21532_n1444# a_32218_n1647# a_32169_n1457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2239 a_32753_984# a_37378_5265# a_37700_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2240 a_640_12878# a_1261_12799# a_1469_12799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2241 a_23193_n14161# a_22980_n14161# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2242 a_30912_12926# a_31169_12736# a_29868_12074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2243 a_57684_n11880# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2244 vdd d0 a_41877_14177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2245 a_45489_n6708# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_82262_9781# a_82515_9768# a_82215_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2247 a_44860_n13391# a_44439_n13391# a_44031_n13283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2248 a_55308_4586# a_54887_4586# a_54479_4153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2249 gnd d0 a_31428_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2250 a_45228_14242# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2251 a_31175_n14209# a_31171_n14032# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2252 a_39124_3950# a_40620_3080# a_40571_3270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2253 a_51582_n13258# a_52679_n13452# a_52630_n13262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2254 vdd a_61102_n8213# a_60894_n8213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2255 a_30126_n10470# a_31219_n9808# a_31170_n9618# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2256 a_19160_n8703# a_19417_n8893# a_17713_n8023# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2257 a_23141_3822# a_22720_3822# a_22312_3506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2258 a_66325_n14840# a_66112_n14840# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2259 a_2569_n5188# a_2356_n5188# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2260 a_51322_4725# a_51579_4535# a_49879_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2261 a_11755_4586# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2262 a_19952_9778# a_20205_9765# a_18904_9103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2263 gnd a_9754_n11932# a_9546_n11932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2264 a_22572_n12379# a_23192_n11873# a_23400_n11873# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2265 a_40833_n7258# a_41930_n7452# a_41881_n7262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_11757_11273# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2267 a_43770_6870# a_44391_6791# a_44599_6791# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2268 gnd a_41088_n13456# a_40880_n13456# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 a_30125_n8699# a_31222_n8893# a_31177_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2270 a_78289_n12724# a_79528_n13404# a_79679_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2271 a_50098_n6749# a_50185_n5240# a_50140_n5227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2272 a_85012_n3616# a_85016_n4472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2273 gnd d0 a_9496_13506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2274 a_12227_n11198# a_12014_n11198# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2275 a_22314_9514# a_22935_9830# a_23143_9830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2276 a_28379_11232# a_28466_12741# a_28417_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2277 a_85015_n14215# a_85011_n14038# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2278 a_13483_n11202# a_13062_n11202# a_12435_n11877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2279 a_66325_n12714# a_66112_n12714# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2280 a_83968_n5915# a_84221_n5928# a_82517_n5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2281 a_25215_4585# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2282 a_6962_n6572# a_7054_n8207# a_7005_n8017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2283 a_43770_6870# a_43770_6475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2284 a_52634_n14886# a_52887_n14899# a_51582_n14705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2285 a_60844_n5056# a_61101_n5246# a_60806_n6755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2286 a_66275_11277# a_65854_11277# a_65446_11356# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2287 vdd d1 a_30122_9094# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2288 a_12803_3814# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2289 gnd a_63594_n11259# a_63386_n11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2290 a_899_n14080# a_899_n14475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2291 a_1521_n5184# a_1308_n5184# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2292 a_54739_n14736# a_55360_n14844# a_55568_n14844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2293 a_83964_n5738# a_85061_n5932# a_85012_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2294 a_17712_n5056# a_19208_n5926# a_19163_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2295 a_76981_3137# a_76560_3137# a_76152_3245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2296 a_78029_3812# a_79268_4579# a_79419_6101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2297 a_52631_n5734# a_52636_n6752# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2298 a_54481_10161# a_54481_9905# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2299 a_54478_8311# a_55099_8232# a_55307_8232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2300 vdd d5 a_59646_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2301 a_11349_10702# a_11349_10161# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2302 a_41619_3945# a_41876_3755# a_40575_3093# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2303 a_72994_7690# a_74091_7496# a_74046_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2304 a_48257_n8839# a_48044_n8839# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2305 a_638_6475# a_638_6220# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2306 vdd d2 a_7261_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2307 a_36294_12228# a_35924_13554# a_34898_14234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2308 a_66535_n8153# a_66114_n8153# a_65706_n8074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2309 gnd d0 a_85268_n14228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2310 a_23402_n5865# a_22981_n5865# a_22573_n5757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2311 a_2308_3820# a_2095_3820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2312 a_56408_n14169# a_56195_n14169# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2313 a_12175_6785# a_13015_6781# a_13223_6781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2314 a_55359_n9751# a_55146_n9751# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2315 a_24243_n8157# a_24030_n8157# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2316 a_11347_4153# a_11968_4586# a_12176_4586# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2317 a_900_n4849# a_1521_n4416# a_1729_n4416# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2318 gnd a_9497_9771# a_9289_9771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2319 a_1730_n7383# a_2570_n6708# a_2778_n6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2320 a_79310_6101# a_79097_6101# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2321 vdd d0 a_74301_14183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2322 a_78030_14234# a_79269_13554# a_79426_12228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2323 gnd a_52886_n11253# a_52678_n11253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2324 a_82522_n8202# a_84014_n7448# a_83969_n7435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2325 a_30916_14196# a_30912_14373# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2326 vdd d0 a_85009_12051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2327 a_14973_n11880# a_14552_n11880# a_14879_n11761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2328 a_68820_n13398# a_68607_n13398# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2329 a_14554_n5872# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2330 a_74046_6741# a_74299_6728# a_72998_6066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2331 a_57596_13556# a_57383_13556# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2332 a_26585_n8841# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2333 a_54740_n5761# a_55361_n5869# a_55569_n5869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2334 a_63343_n5238# a_63339_n5061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2335 a_67582_n3743# a_67161_n3743# a_66534_n4418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2336 a_77869_n3749# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2337 vdd d0 a_20202_6724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2338 gnd d0 a_9756_n5245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2339 a_54740_n3408# a_54740_n3664# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2340 a_28375_11409# a_28467_9774# a_28422_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2341 a_77243_n7391# a_76822_n7391# a_76414_n7283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2342 a_18900_10727# a_19157_10537# a_17457_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2343 vdd a_20203_5204# a_19995_5204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2344 a_84750_6233# a_85007_6043# a_83702_6237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2345 a_36294_12228# a_36180_12109# a_36388_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2346 vdd a_40827_7494# a_40619_7494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2347 a_63084_10546# a_63337_10533# a_62032_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2348 vdd d2 a_50391_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2349 a_57641_n10435# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2350 a_49030_n9784# a_49283_n9797# a_48681_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2351 a_11969_13561# a_11756_13561# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2352 a_2777_n3741# a_2356_n3741# a_1729_n3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2353 a_41624_13511# a_41877_13498# a_40572_13692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2354 a_40837_n8882# a_41090_n8895# a_39386_n8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2355 gnd d2 a_17710_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2356 a_76413_n5508# a_76413_n5763# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2357 a_55310_9826# a_54889_9826# a_54481_9510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2358 a_2096_14242# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2359 a_67162_n6710# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2360 a_18904_9103# a_19997_9765# a_19952_9778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2361 gnd a_83959_6047# a_83751_6047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2362 a_76560_4584# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2363 a_52630_n14030# a_52887_n14220# a_51586_n14882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2364 a_84757_9776# a_85010_9763# a_83709_9101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2365 a_26992_5271# a_27356_8184# a_27307_8374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2366 a_51588_n7427# a_52681_n6765# a_52632_n6575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2367 a_8452_n8697# a_9549_n8891# a_9504_n8878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2368 a_48780_n5913# a_53885_n1645# a_53727_n1632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2369 a_78080_n11204# a_77867_n11204# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2370 a_82479_n6757# a_82732_n6770# a_81411_n9792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2371 a_17713_n8023# a_17970_n8213# a_17670_n6578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2372 a_70138_n8841# a_70611_n5928# a_70453_n5915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2373 a_12229_n5190# a_12016_n5190# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2374 a_67114_12793# a_66901_12793# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2375 gnd a_62546_n11934# a_62338_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2376 a_83969_n7435# a_85062_n6773# a_85017_n6760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2377 a_59173_n8845# a_59646_n5932# a_53628_n1455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2378 a_9237_7688# a_9241_6743# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2379 a_49875_3958# a_51371_3088# a_51326_3101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2380 a_20212_n8884# a_20208_n8707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2381 a_16606_n9790# a_17719_n6768# a_17674_n6755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2382 a_22981_n4418# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2383 a_71505_5401# a_71597_3766# a_71548_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2384 a_33020_3895# a_33020_3500# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2385 a_14250_4581# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2386 a_2355_n12716# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2387 a_69072_n5868# a_69930_n8841# a_70138_n8841# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2388 a_900_n4053# a_900_n4308# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2389 vdd a_52886_n11932# a_52678_n11932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2390 a_52633_n9793# a_52886_n9806# a_51585_n10468# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2391 gnd a_42136_n14907# a_41928_n14907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2392 a_76820_n12720# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2393 a_39124_3950# a_40620_3080# a_40575_3093# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2394 a_43773_11614# a_43773_11358# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2395 a_1262_9832# a_1049_9832# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2396 a_899_n14080# a_1520_n14159# a_1728_n14159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 a_62293_n11921# a_63386_n11259# a_63337_n11069# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2398 a_83704_12245# a_84801_12051# a_84752_12241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2399 a_25259_12115# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2400 a_19948_9955# a_20205_9765# a_18904_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2401 a_41883_n13447# a_41879_n13270# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2402 a_22574_n6627# a_23195_n6706# a_23403_n6706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2403 a_78288_n11204# a_77867_n11204# a_77240_n11200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2404 a_33021_14317# a_33642_14238# a_33850_14238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2405 gnd a_63594_n9812# a_63386_n9812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2406 a_82259_6740# a_83751_7494# a_83706_7507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2407 a_11609_n8728# a_12230_n8836# a_12438_n8836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2408 a_14619_6222# a_14505_6103# a_14713_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2409 a_17674_n6755# a_17761_n5246# a_17716_n5233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2410 a_81151_8191# a_81404_8178# a_80832_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2411 a_34738_n6716# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2412 a_55308_4586# a_56148_5261# a_56356_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2413 a_29864_13698# a_30121_13508# a_28421_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2414 a_76151_7118# a_76772_7551# a_76980_7551# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2415 a_44031_n13824# a_44652_n13391# a_44860_n13391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2416 a_1047_3145# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2417 a_14621_12230# a_14507_12111# a_14715_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2418 a_68651_n5868# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2419 a_28379_11232# a_28466_12741# a_28421_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2420 a_51583_n5730# a_51840_n5920# a_50136_n5050# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2421 a_77242_n3745# a_76821_n3745# a_76413_n3666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2422 a_79570_n11882# a_79357_n11882# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2423 a_11607_n14086# a_12228_n14165# a_12436_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2424 a_71547_6923# a_73043_6053# a_72994_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2425 a_51582_n14705# a_51839_n14895# a_50135_n14025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2426 a_50139_n14202# a_50392_n14215# a_50092_n12580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2427 a_62029_7686# a_63126_7492# a_63081_7505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2428 a_73001_10554# a_74094_11216# a_74045_11406# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2429 a_44178_7559# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2430 a_58752_n8845# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2431 a_51583_n5730# a_52680_n5924# a_52635_n5911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2432 a_11609_n7026# a_12230_n6710# a_12438_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2433 a_43772_12483# a_43772_12228# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2434 a_9500_n8022# a_9504_n8878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2435 a_84753_9274# a_84754_8182# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2436 gnd d0 a_74300_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2437 a_33687_n11879# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2438 a_55148_n5190# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2439 a_45648_3820# a_45227_3820# a_44600_3824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2440 gnd d0 a_20204_12053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2441 vdd a_9497_11218# a_9289_11218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2442 a_23143_10598# a_22722_10598# a_22314_10706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2443 a_28419_6746# a_28672_6733# a_28377_5224# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2444 vdd a_51840_n4473# a_51632_n4473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2445 vdd a_85007_8169# a_84799_8169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2446 gnd d0 a_41876_4523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2447 a_52371_12249# a_52376_11231# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2448 a_40576_13515# a_41669_14177# a_41624_14190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2449 a_65443_6868# a_66064_6789# a_66272_6789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2450 a_40835_n13443# a_41928_n12781# a_41879_n12591# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2451 a_80425_n8847# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2452 vdd a_9497_9771# a_9289_9771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2453 a_43770_7922# a_44391_8238# a_44599_8238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2454 a_14616_12111# a_14252_10589# a_13226_9822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2455 a_66326_n5186# a_66113_n5186# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2456 a_899_n12377# a_899_n12633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2457 vdd a_42136_n14228# a_41928_n14228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2458 a_18900_10727# a_19997_10533# a_19948_10723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 a_3913_12236# a_3799_12117# a_4007_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2460 a_24448_n11198# a_25687_n10431# a_25844_n11757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2461 a_37506_n8847# a_37293_n8847# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2462 vdd d0 a_31169_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2463 gnd d0 a_74560_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2464 a_54481_3148# a_55100_3139# a_55308_3139# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2465 a_3542_4587# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2466 a_34475_6779# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2467 a_2776_n14163# a_2355_n14163# a_1728_n14838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2468 gnd d0 a_9497_9092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2469 a_23402_n5186# a_24242_n5190# a_24450_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2470 a_11348_14319# a_11969_14240# a_12177_14240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2471 a_65851_6110# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2472 a_31171_n13264# a_31175_n14209# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2473 a_23140_8236# a_23980_8232# a_24188_8232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2474 a_63080_10723# a_63337_10533# a_62032_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2475 a_44652_n12712# a_44439_n12712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2476 a_28678_n8019# a_30174_n8889# a_30129_n8876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2477 a_9242_5223# a_9495_5210# a_8194_4548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2478 gnd a_82512_6727# a_82304_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2479 a_43771_4700# a_43771_4159# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2480 a_45650_11275# a_45229_11275# a_44602_10600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2481 a_78030_14234# a_77609_14234# a_76982_13559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2482 a_24451_n6710# a_25690_n7390# a_25841_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2483 a_41881_n8030# a_41885_n8886# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2484 a_44441_n8151# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2485 a_67583_n8157# a_68822_n7390# a_68973_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2486 vdd d2 a_17710_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2487 a_33903_n8838# a_33690_n8838# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2488 gnd a_20202_6724# a_19994_6724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2489 a_18903_13517# a_19156_13504# a_17456_12750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2490 vdd a_72022_n12772# a_71814_n12772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2491 a_56616_n12722# a_57855_n13402# a_58006_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2492 vdd a_28933_n14217# a_28725_n14217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2493 a_44861_n4416# a_45701_n3741# a_45909_n3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2494 a_1468_3145# a_1047_3145# a_639_3253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2495 gnd d1 a_8448_12063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2496 a_29862_6243# a_30959_6049# a_30910_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2497 vdd a_85268_n12781# a_85060_n12781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2498 a_72999_3099# a_74092_3761# a_74043_3951# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2499 a_12175_7553# a_13015_8228# a_13223_8228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2500 a_14292_6103# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2501 a_84753_9953# a_85010_9763# a_83709_9101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2502 a_54478_7661# a_54478_7120# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2503 vdd d2 a_82773_n14223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2504 a_26992_5271# a_27356_8184# a_27311_8197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2505 a_25687_n10431# a_25474_n10431# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2506 a_78288_n9757# a_77867_n9757# a_77240_n10432# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2507 a_77241_n14167# a_76820_n14167# a_76412_n14483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2508 a_901_n8722# a_1522_n8830# a_1730_n8830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2509 a_74309_n7433# a_74562_n7446# a_73257_n7252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2510 a_22312_3251# a_22314_3152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2511 a_8192_10733# a_9289_10539# a_9240_10729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2512 a_71505_5401# a_71597_3766# a_71552_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2513 a_35159_n8163# a_34738_n8163# a_34111_n8159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2514 a_77034_n4424# a_76821_n4424# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2515 gnd d4 a_16599_8180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2516 a_44030_n11113# a_44651_n11192# a_44859_n11192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2517 a_33281_n5113# a_33281_n5508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2518 a_43773_10708# a_44394_10600# a_44602_10600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2519 vdd a_17665_5207# a_17457_5207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2520 gnd a_39640_n11256# a_39432_n11256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2521 a_22979_n10426# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2522 a_44392_3145# a_44179_3145# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2523 a_11970_10594# a_11757_10594# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2524 gnd a_42137_n5932# a_41929_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2525 a_11970_9147# a_11757_9147# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2526 a_640_13134# a_640_12878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2527 a_44033_n8722# a_44030_n9410# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2528 a_52630_n14030# a_52634_n14886# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2529 a_5898_n9784# a_7011_n6762# a_6962_n6572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2530 a_83704_12245# a_84801_12051# a_84756_12064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2531 a_901_n7020# a_1522_n6704# a_1730_n6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2532 gnd d2 a_60840_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2533 a_44861_n5863# a_44440_n5863# a_44033_n6369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2534 a_79686_n5755# a_79316_n4429# a_78290_n3749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2535 a_8196_9109# a_9289_9771# a_9240_9961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2536 a_36395_n10437# a_36182_n10437# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2537 a_24191_9826# a_23770_9826# a_23143_9151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2538 gnd d0 a_63595_n14226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2539 vdd d0 a_20462_n10491# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2540 a_35967_12109# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2541 a_33848_7551# a_33427_7551# a_33019_7118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2542 gnd d0 a_52889_n8891# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2543 a_5333_n8839# a_4912_n8839# a_4265_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2544 gnd d3 a_17927_n6768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2545 a_63082_5217# a_63078_5394# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2546 gnd d2 a_39643_n8215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2547 a_3053_n1225# a_43280_n1602# a_43231_n1412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 a_66114_n8832# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2549 a_71547_6923# a_73043_6053# a_72998_6066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2550 a_30916_12070# a_31169_12057# a_29864_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2551 a_66900_3818# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2552 a_22313_12481# a_22934_12797# a_23142_12797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2553 gnd d1 a_8708_n5920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2554 a_73001_10554# a_74094_11216# a_74049_11229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2555 a_12014_n11877# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2556 a_14462_7548# a_14249_7548# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2557 a_63338_n13268# a_63595_n13458# a_62290_n13264# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2558 a_34897_3812# a_34476_3812# a_33849_3137# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2559 a_74307_n14888# a_74560_n14901# a_73255_n14707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2560 a_1309_n8830# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2561 a_39341_n12588# a_39433_n14223# a_39388_n14210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2562 a_51585_n11915# a_51838_n11928# a_50134_n11058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2563 vdd d0 a_74300_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2564 a_84751_5392# a_84755_4536# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2565 a_67321_3818# a_68560_4585# a_68711_6107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2566 a_78080_n9757# a_77867_n9757# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2567 a_60845_n8023# a_62341_n8893# a_62296_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2568 vdd d0 a_20204_12053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2569 gnd d2 a_17969_n5246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2570 a_19159_n4289# a_20256_n4483# a_20207_n4293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2571 a_65705_n3404# a_65705_n3660# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2572 a_64664_n1444# a_75350_n1647# a_70453_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2573 a_1262_10600# a_1049_10600# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2574 a_28415_6923# a_28672_6733# a_28377_5224# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2575 a_30915_3095# a_30911_3272# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2576 a_77607_8226# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2577 a_900_n3658# a_900_n4053# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2578 a_62029_7686# a_62286_7496# a_60586_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2579 a_76821_n5192# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2580 vdd a_19416_n4479# a_19208_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2581 vdd d0 a_41876_4523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2582 vdd a_30122_9094# a_29914_9094# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2583 gnd a_84220_n13456# a_84012_n13456# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2584 a_65705_n3404# a_74561_n3800# a_73260_n4462# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2585 a_78081_n14171# a_77868_n14171# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2586 gnd a_9496_14185# a_9288_14185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2587 a_44601_14246# a_45441_14242# a_45649_14242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2588 a_55359_n11198# a_55146_n11198# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2589 a_41879_n12591# a_41883_n13447# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2590 a_12435_n10430# a_12014_n10430# a_11606_n10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2591 a_65703_n10063# a_66324_n9747# a_66532_n9747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2592 a_639_4955# a_1260_5271# a_1468_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2593 a_63343_n5917# a_63596_n5930# a_62291_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2594 a_41622_6056# a_41618_6233# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2595 a_18900_10727# a_19997_10533# a_19952_10546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2596 a_6745_9966# a_8241_9096# a_8196_9109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2597 a_22982_n6706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2598 vdd a_52887_n14899# a_52679_n14899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2599 a_2095_3820# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2600 vdd a_7260_n14215# a_7052_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2601 vdd a_41089_n4481# a_40881_n4481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2602 a_23142_12118# a_23982_12793# a_24190_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2603 vdd a_42138_n6773# a_41930_n6773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2604 a_12177_13561# a_11756_13561# a_11348_13669# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2605 a_74044_12926# a_74048_12070# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2606 a_12017_n8836# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2607 vdd d2 a_50393_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2608 a_41623_3089# a_41876_3076# a_40571_3270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2609 a_36138_10587# a_35925_10587# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2610 a_58013_n5753# a_57643_n4427# a_56617_n5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2611 a_19161_n10474# a_20254_n9812# a_20209_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2612 a_9238_5400# a_9495_5210# a_8194_4548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2613 a_84756_12743# a_85009_12730# a_83708_12068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2614 a_75885_984# a_80510_5265# a_80586_9136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2615 a_44600_5271# a_44179_5271# a_43771_5350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2616 vdd d1 a_51841_n7440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2617 a_84752_14367# a_84756_13511# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2618 gnd d2 a_17707_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2619 a_56148_5261# a_55935_5261# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2620 a_55309_12793# a_54888_12793# a_54480_12477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2621 vdd a_20202_6724# a_19994_6724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2622 vdd a_61057_n12776# a_60849_n12776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2623 vdd d1 a_8448_12063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2624 a_22314_9514# a_22314_9259# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2625 vdd d0 a_42138_n8899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2626 a_12017_n6710# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2627 a_33280_n13036# a_33901_n12720# a_34109_n12720# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2628 a_62292_n7256# a_63389_n7450# a_63344_n7437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2629 a_72999_3099# a_74092_3761# a_74047_3774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2630 a_50098_n6749# a_50185_n5240# a_50136_n5050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2631 a_67115_11273# a_66902_11273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2632 a_68812_12115# a_68391_12115# a_68713_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2633 a_36182_n10437# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2634 a_66273_3822# a_65852_3822# a_65444_3901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2635 gnd d0 a_9755_n12773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2636 a_55570_n8836# a_56410_n8161# a_56618_n8161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2637 a_33851_9824# a_33430_9824# a_33022_9508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2638 a_20205_n11748# a_20462_n11938# a_19157_n11744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2639 a_11179_986# a_10758_986# a_5418_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2640 a_65443_8571# a_66067_9151# a_66275_9151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2641 gnd d0 a_20202_6045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2642 a_6746_6748# a_6999_6735# a_6704_5226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2643 vdd d1 a_8706_n10481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2644 vdd a_31170_9769# a_30962_9769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2645 vdd d4 a_16599_8180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2646 a_31171_n14032# a_31428_n14222# a_30127_n14884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2647 a_11608_n5761# a_11609_n6375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2648 a_23770_11273# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2649 gnd a_31170_11216# a_30962_11216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2650 a_60589_9783# a_62081_10537# a_62036_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2651 a_29869_9107# a_30962_9769# a_30913_9959# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2652 a_54886_7553# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2653 a_60848_n5233# a_61101_n5246# a_60806_n6755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2654 a_38275_n9615# a_38532_n9805# a_37930_n5744# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2655 a_49832_5403# a_49924_3768# a_49875_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2656 a_51324_9286# a_52421_9092# a_52376_9105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2657 a_17712_n5056# a_19208_n5926# a_19159_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2658 gnd a_50351_n6762# a_50143_n6762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2659 a_3586_12117# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2660 gnd d1 a_51578_7502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2661 vdd d2 a_60840_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2662 a_29864_13698# a_30961_13504# a_30916_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2663 a_68978_n5749# a_68608_n4423# a_67582_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2664 a_8196_9109# a_9289_9771# a_9244_9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2665 a_18900_9280# a_19997_9086# a_19948_9276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2666 gnd d0 a_42135_n10493# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2667 a_63339_n5061# a_63596_n5251# a_62295_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2668 gnd d2 a_7261_n5240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2669 a_11756_14240# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2670 gnd d1 a_83962_9088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2671 vdd a_8708_n4473# a_8500_n4473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2672 gnd a_40830_10535# a_40622_10535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2673 a_39129_12748# a_39382_12735# a_39087_11226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2674 a_25477_n7390# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2675 a_17711_n14031# a_19207_n14901# a_19158_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2676 a_56194_n9755# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2677 a_40577_9101# a_40830_9088# a_39126_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2678 a_11606_n9672# a_11606_n10067# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2679 a_55934_6781# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2680 a_82522_n8202# a_84014_n7448# a_83965_n7258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2681 a_9499_n4287# a_9756_n4477# a_8451_n4283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2682 a_68609_n7390# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2683 a_44860_n13391# a_45700_n12716# a_45908_n12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2684 gnd d0 a_31428_n14222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2685 gnd d1 a_40828_3080# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2686 a_17450_6919# a_17707_6729# a_17412_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2687 gnd d0 a_41878_11210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 a_13065_n8161# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2689 a_45488_n3741# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2690 a_66274_14244# a_65853_14244# a_65445_13928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2691 a_67159_n11198# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2692 a_22572_n13826# a_22572_n14082# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2693 a_23141_3143# a_22720_3143# a_22314_3152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2694 a_19952_9099# a_20205_9086# a_18900_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_22571_n11510# a_23192_n11194# a_23400_n11194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2696 gnd a_9754_n11253# a_9546_n11253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2697 a_67372_n9751# a_67159_n9751# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2698 a_73254_n10293# a_73511_n10483# a_71811_n11237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2699 a_49878_6748# a_50131_6735# a_49836_5226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2700 a_45647_8234# a_45226_8234# a_44599_7559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2701 a_9502_n13439# a_9498_n13262# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2702 vdd d1 a_84221_n4481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2703 a_2944_n1225# a_2731_n1225# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2704 vdd a_85009_14177# a_84801_14177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2705 a_899_n14730# gnd gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2706 a_57643_n4427# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2707 a_23195_n7385# a_22982_n7385# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2708 gnd d2 a_50391_n11248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2709 a_33850_12791# a_34690_12787# a_34898_12787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2710 a_63080_11402# a_63084_10546# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2711 a_639_5350# a_639_4955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2712 vdd a_9496_14185# a_9288_14185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2713 a_13276_n14169# a_13063_n14169# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2714 a_62035_13517# a_63128_14179# a_63083_14192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2715 a_9497_n10295# a_9754_n10485# a_8449_n10291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2716 a_59389_n5742# a_59783_n9803# a_59738_n9790# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2717 a_23140_6789# a_22719_6789# a_22311_6868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2718 a_44031_n13824# a_44031_n14080# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2719 a_76412_n13832# a_76412_n14088# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2720 a_68821_n4423# a_68608_n4423# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2721 a_52634_n14207# a_52887_n14220# a_51586_n14882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2722 a_77035_n6712# a_76822_n6712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2723 gnd a_41876_4523# a_41668_4523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2724 a_13226_9822# a_14465_10589# a_14616_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2725 a_8193_7515# a_8446_7502# a_6746_6748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2726 a_3801_n10429# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2727 a_54739_n14086# a_55360_n14165# a_55568_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2728 a_83968_n5915# a_85061_n5253# a_85012_n5063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2729 a_76983_10592# a_77823_11267# a_78031_11267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2730 a_63342_n13445# a_63338_n13268# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2731 a_41619_3266# a_41876_3076# a_40571_3270# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2732 a_66533_n14840# a_67373_n14165# a_67581_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2733 gnd d1 a_73511_n10483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2734 a_2518_9828# a_2097_9828# a_1470_9153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2735 a_16606_n9790# a_17719_n6768# a_17670_n6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2736 a_30916_14196# a_33021_14317# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2737 a_84752_12920# a_85009_12730# a_83708_12068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2738 a_1259_7559# a_1046_7559# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2739 a_23402_n5186# a_22981_n5186# a_22573_n5107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2740 a_36396_n13404# a_36183_n13404# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2741 a_62034_3095# a_63127_3757# a_63082_3770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2742 a_56195_n12722# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2743 a_85012_n3616# a_85269_n3806# a_83968_n4468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2744 a_30910_7686# a_31167_7496# a_29862_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2745 a_63343_n5917# a_63339_n5740# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2746 a_76411_n9418# a_77035_n8838# a_77243_n8838# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2747 a_9243_14198# a_9239_14375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2748 a_51582_n13258# a_52679_n13452# a_52634_n13439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2749 a_62296_n8880# a_62549_n8893# a_60845_n8023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2750 gnd a_9497_9092# a_9289_9092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2751 a_76151_6212# a_76772_6104# a_76980_6104# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2752 a_24242_n5190# a_24029_n5190# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2753 a_77032_n11200# a_76819_n11200# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2754 a_39386_n8025# a_39643_n8215# a_39343_n6580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2755 a_22312_5604# a_22312_5348# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2756 gnd d0 a_74302_11216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2757 a_9241_6743# a_9494_6730# a_8193_6068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2758 vdd a_9754_n11932# a_9546_n11932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2759 a_58837_5267# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 a_22980_n12714# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2761 a_40833_n7258# a_41930_n7452# a_41885_n7439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2762 a_33688_n13399# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2763 a_45442_9828# a_45229_9828# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2764 a_17674_n6755# a_17761_n5246# a_17712_n5056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2765 a_36386_6101# a_35965_6101# a_36292_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2766 a_22574_n7022# a_22574_n7277# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2767 a_22933_3822# a_22720_3822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2768 a_74046_6062# a_74299_6049# a_72994_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2769 a_68649_n11876# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2770 a_25429_13560# a_25216_13560# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2771 a_54740_n5111# a_55361_n5190# a_55569_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2772 a_67162_n8157# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2773 a_79686_n5755# a_79572_n5874# a_79780_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 gnd a_62289_9090# a_62081_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2775 a_6742_6925# a_6999_6735# a_6704_5226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2776 a_51587_n5907# a_51840_n5920# a_50136_n5050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2777 vdd d0 a_20202_6045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2778 a_84750_8359# a_84754_7503# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2779 a_2307_6787# a_2094_6787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2780 a_52636_n6752# a_52632_n6575# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2781 a_83702_7684# a_84799_7490# a_84750_7680# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2782 a_55099_6785# a_54886_6785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2783 a_27222_n5738# a_27479_n5928# a_27321_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2784 a_54741_n7281# a_54741_n7822# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2785 a_56617_n5194# a_56196_n5194# a_55569_n5869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2786 a_11607_n13034# a_11607_n13289# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2787 a_63341_n9799# a_63337_n9622# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2788 a_19164_n7433# a_20257_n6771# a_20208_n6581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2789 vdd a_31170_11216# a_30962_11216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2790 a_23194_n3739# a_22981_n3739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2791 a_51583_n5730# a_52680_n5924# a_52631_n5734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2792 a_10971_986# a_10758_986# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2793 a_55100_3818# a_54887_3818# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2794 a_2357_n8155# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2795 a_83964_n5738# a_85061_n5932# a_85016_n5919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2796 a_12229_n5869# a_12016_n5869# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2797 a_30124_n4285# a_30381_n4475# a_28681_n5229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2798 a_34108_n10432# a_34948_n9757# a_35156_n9757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2799 a_901_n8072# a_901_n8467# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2800 a_55310_9147# a_54889_9147# a_54478_8567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2801 a_31173_n6577# a_31430_n6767# a_30129_n7429# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2802 vdd a_32426_n1647# a_32218_n1647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2803 a_23769_12793# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2804 a_18900_9280# a_19997_9086# a_19952_9099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2805 a_55362_n7389# a_55149_n7389# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2806 a_12228_n14844# a_12015_n14844# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2807 a_74307_n14209# a_74303_n14032# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2808 a_60588_12750# a_62080_13504# a_62031_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2809 a_76152_4692# a_76773_4584# a_76981_4584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2810 a_84757_9097# a_85010_9084# a_83705_9278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2811 a_12436_n13397# a_12015_n13397# a_11607_n13830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2812 a_8456_n8874# a_9549_n8212# a_9504_n8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2813 a_52631_n5055# a_52635_n5911# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2814 vdd d0 a_20464_n3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2815 a_20208_n8707# a_20465_n8897# a_19160_n8703# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2816 vdd d8 a_43488_n1602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2817 a_33428_3816# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2818 a_51324_9286# a_51581_9096# a_49877_9966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2819 a_11349_9905# a_11970_9826# a_12178_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2820 a_55309_14240# a_54888_14240# a_54480_14319# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2821 vdd a_40830_10535# a_40622_10535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2822 a_66064_6110# a_65851_6110# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2823 a_39125_12925# a_39382_12735# a_39087_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2824 a_84756_13511# a_84752_13688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2825 a_22314_11356# a_22935_11277# a_23143_11277# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2826 vdd d1 a_30382_n8889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2827 a_25584_6226# a_25214_7552# a_24188_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2828 a_50141_n8194# a_51633_n7440# a_51588_n7427# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2829 vdd a_52886_n11253# a_52678_n11253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2830 a_50092_n12580# a_50349_n12770# a_49026_n9607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2831 a_45486_n11196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2832 gnd a_42136_n14228# a_41928_n14228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2833 a_56409_n3747# a_56196_n3747# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2834 a_13063_n14169# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2835 vdd d1 a_40828_3080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2836 a_66066_13565# a_65853_13565# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2837 vdd d0 a_41878_11210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2838 a_1262_9153# a_1049_9153# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2839 a_33642_14238# a_33429_14238# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2840 a_19948_9276# a_20205_9086# a_18900_9280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2841 a_76981_3816# a_77821_3812# a_78029_3812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2842 a_49874_6925# a_50131_6735# a_49836_5226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2843 a_62289_n10297# a_62546_n10487# a_60846_n11241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2844 a_79780_n5874# a_79359_n5874# a_79686_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2845 a_85012_n4295# a_85016_n5240# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2846 a_28678_n8019# a_30174_n8889# a_30125_n8699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2847 a_46935_n4421# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2848 vdd d0 a_63335_5204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2849 a_11609_n8078# a_12230_n8157# a_12438_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2850 a_41879_n13270# a_42136_n13460# a_40831_n13266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2851 gnd d0 a_9497_10539# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2852 a_12175_6785# a_11754_6785# a_11346_6864# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2853 a_44030_n10061# a_44651_n9745# a_44859_n9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2854 a_37033_9136# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2855 a_47137_6109# a_47997_9144# a_48205_9144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2856 gnd a_74300_5208# a_74092_5208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 a_62035_12070# a_62288_12057# a_60584_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2858 a_20206_n14715# a_20463_n14905# a_19158_n14711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2859 vdd a_41877_13498# a_41669_13498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2860 a_40570_7684# a_40827_7494# a_39127_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2861 a_82515_n11066# a_82772_n11256# a_82477_n12765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2862 gnd a_28933_n14217# a_28725_n14217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2863 gnd d0 a_52626_7498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2864 a_66065_4590# a_65852_4590# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2865 a_23143_11277# a_23983_11273# a_24191_11273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2866 vdd a_41876_4523# a_41668_4523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2867 a_33429_13559# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2868 a_71767_n6574# a_72024_n6764# a_70703_n9786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2869 a_11607_n13034# a_12228_n12718# a_12436_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2870 a_51587_n5907# a_52680_n5245# a_52635_n5232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2871 a_29866_6066# a_30119_6053# a_28415_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2872 a_33687_n11200# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2873 a_83706_6060# a_83959_6047# a_82255_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2874 vdd a_31428_n12775# a_31220_n12775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2875 a_59389_n5742# a_59646_n5932# a_53628_n1455# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2876 a_638_7126# a_638_6870# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2877 a_1307_n14838# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2878 a_37591_5265# a_37378_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2879 a_83709_9101# a_84802_9763# a_84753_9953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2880 a_57595_4581# a_57382_4581# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2881 gnd d0 a_85007_8169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2882 a_12438_n6710# a_12017_n6710# a_11609_n7026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2883 a_23401_n14161# a_22980_n14161# a_22572_n14477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2884 a_36289_12109# a_35925_10587# a_34899_11267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2885 a_33022_10700# a_33643_10592# a_33851_10592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2886 a_20212_n6758# a_20208_n6581# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2887 gnd a_20462_n10491# a_20254_n10491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2888 a_55146_n9751# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2889 vdd d0 a_74302_11216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2890 a_9237_6920# a_9494_6730# a_8193_6068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2891 a_47191_n5866# a_46978_n5866# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2892 a_1307_n12712# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2893 a_9500_n6575# a_9757_n6765# a_8456_n7427# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2894 a_9498_n12583# a_9502_n13439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2895 gnd a_41088_n14903# a_40880_n14903# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2896 a_44438_n11871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2897 a_54480_12477# a_55101_12793# a_55309_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2898 a_55567_n10430# a_55146_n10430# a_54738_n10863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2899 a_33021_12870# a_33021_12475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2900 a_70703_n9786# a_70956_n9799# a_70354_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2901 a_28379_11232# a_28632_11219# a_27311_8197# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2902 a_639_4955# a_639_4700# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2903 a_76154_9903# a_76775_9824# a_76983_9824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2904 a_2776_n12716# a_2355_n12716# a_1728_n12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2905 a_34477_12787# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2906 a_43773_9261# a_43770_8573# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2907 a_24448_n11198# a_24027_n11198# a_23400_n11873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2908 a_63342_n13445# a_63595_n13458# a_62290_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2909 a_41885_n7439# a_42138_n7452# a_40833_n7258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2910 vdd a_74559_n9808# a_74351_n9808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2911 a_23400_n9747# a_24240_n9751# a_24448_n9751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2912 a_19948_9955# a_19952_9099# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2913 a_33903_n8159# a_33690_n8159# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2914 a_76981_4584# a_76560_4584# a_76152_4692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2915 gnd a_20202_6045# a_19994_6045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2916 a_65705_n5757# a_66326_n5865# a_66534_n5865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2917 a_25730_n11876# a_25517_n11876# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2918 a_44654_n7383# a_44441_n7383# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2919 a_64664_n1444# a_75350_n1647# a_75301_n1457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2920 a_12178_9147# a_13018_9822# a_13226_9822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2921 a_76414_n7824# a_76414_n8080# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2922 a_72995_3276# a_74092_3082# a_74043_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2923 a_51323_13700# a_52420_13506# a_52375_13519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2924 a_84753_9274# a_85010_9084# a_83705_9278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2925 gnd a_19416_n4479# a_19208_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2926 a_638_7667# a_1259_7559# a_1467_7559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2927 gnd a_28934_n5242# a_28726_n5242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_23401_n12714# a_24241_n12718# a_24449_n12718# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 a_83963_n14713# a_85060_n14907# a_85015_n14894# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2930 a_6700_5403# a_6792_3768# a_6747_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2931 a_14614_6103# a_14250_4581# a_13224_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2932 gnd a_85270_n8899# a_85062_n8899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2933 gnd a_51578_7502# a_51370_7502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2934 a_40835_n13443# a_41928_n12781# a_41883_n12768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2935 a_3802_n13396# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2936 vdd d0 a_85267_n9814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2937 a_73258_n10470# a_74351_n9808# a_74302_n9618# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2938 a_12177_12114# a_11756_12114# a_11349_11608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2939 a_9237_8367# a_9241_7511# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2940 a_30915_3774# a_31168_3761# a_29867_3099# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2941 a_901_n6369# a_1521_n5863# a_1729_n5863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2942 a_47300_n5866# a_46936_n7388# a_45910_n6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2943 gnd d0 a_52887_n12773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2944 a_20206_n13268# a_20210_n14213# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2945 gnd a_31170_9090# a_30962_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2946 a_34950_n3749# a_34737_n3749# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2947 gnd a_83962_9088# a_83754_9088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2948 gnd a_42137_n5253# a_41929_n5253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2949 gnd d1 a_62286_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2950 gnd a_7260_n14215# a_7052_n14215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2951 a_3913_12236# a_3543_13562# a_2517_14242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2952 vdd d0 a_85009_13498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2953 gnd a_52627_3763# a_52419_3763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2954 gnd d2 a_50393_n5240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2955 a_77608_5259# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2956 a_73001_10554# a_73254_10541# a_71554_9787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2957 a_8192_9286# a_9289_9092# a_9240_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2958 a_34111_n8838# a_33690_n8838# a_33279_n9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2959 a_44861_n5184# a_44440_n5184# a_44032_n5500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2960 a_12177_13561# a_13017_14236# a_13225_14236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2961 a_76774_13559# a_76561_13559# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2962 a_22311_8571# a_22311_8315# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2963 gnd d2 a_71804_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2964 a_14510_n13402# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2965 gnd d0 a_41877_14177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2966 a_39390_n8202# a_40882_n7448# a_40837_n7435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2967 gnd a_40828_3080# a_40620_3080# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2968 a_84750_7680# a_85007_7490# a_83702_7684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2969 vdd a_9755_n14899# a_9547_n14899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2970 a_27571_n9786# a_28684_n6764# a_28639_n6751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2971 a_11607_n12639# a_11607_n13034# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2972 gnd d0 a_52889_n8212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2973 gnd d1 a_51841_n7440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2974 a_8195_12076# a_9288_12738# a_9243_12751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2975 a_71814_n8196# a_72067_n8209# a_71767_n6574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2976 a_66114_n8153# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2977 vdd d1 a_62289_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2978 gnd a_61057_n12776# a_60849_n12776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2979 gnd a_17968_n14221# a_17760_n14221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2980 a_66273_3143# a_67113_3818# a_67321_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2981 a_30915_3774# a_30911_3951# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2982 a_22314_11612# a_22934_12118# a_23142_12118# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2983 gnd d0 a_63334_6724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2984 a_62292_n7256# a_63389_n7450# a_63340_n7260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2985 a_34111_n6712# a_33690_n6712# a_33282_n6633# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2986 vdd a_52629_10539# a_52421_10539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2987 a_12014_n11198# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2988 a_45907_n9749# a_45486_n9749# a_44859_n10424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2989 a_33281_n3410# a_42137_n3806# a_40836_n4468# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2990 a_54886_6106# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2991 a_57637_6103# a_57424_6103# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2992 a_19946_4715# a_19950_3770# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2993 a_29862_6243# a_30119_6053# a_28415_6923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2994 a_20209_n11925# a_20462_n11938# a_19157_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2995 a_38275_n9615# a_39390_n12778# a_39345_n12765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2996 a_74307_n14209# a_74560_n14222# a_73259_n14884# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2997 a_43772_13134# a_43772_12878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2998 a_1309_n8151# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2999 a_56355_8228# a_55934_8228# a_55307_7553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3000 a_44653_n3737# a_44440_n3737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 a_33279_n10069# a_33900_n9753# a_34108_n9753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3002 a_41622_6735# a_41618_6912# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3003 a_13225_12789# a_12804_12789# a_12177_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3004 a_83709_9101# a_84802_9763# a_84757_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3005 a_67322_12793# a_66901_12793# a_66274_12118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3006 a_24030_n6710# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3007 vdd a_85270_n8220# a_85062_n8220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3008 a_39128_3773# a_40620_4527# a_40575_4540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3009 vdd a_42137_n5932# a_41929_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3010 a_70223_5271# a_75776_984# a_64849_973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3011 a_74303_n13264# a_74307_n14209# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3012 a_5898_n9784# a_7011_n6762# a_6966_n6749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3013 a_74043_3272# a_65446_3152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3014 a_73255_n13260# a_74352_n13454# a_74307_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3015 vdd a_17970_n8213# a_17762_n8213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3016 a_2356_n3741# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3017 a_641_10708# a_1262_10600# a_1470_10600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3018 a_44033_n6625# a_44033_n7020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3019 a_28419_6746# a_29911_7500# a_29862_7690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3020 a_2096_12795# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3021 a_18904_9103# a_19157_9090# a_17453_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3022 gnd d3 a_82470_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3023 a_82256_3950# a_83752_3080# a_83703_3270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3024 a_74309_n7433# a_74305_n7256# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3025 a_48205_9144# a_48342_5273# a_48550_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3026 a_12017_n8157# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3027 a_1047_4592# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3028 vdd d2 a_28935_n8209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3029 a_54887_4586# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3030 a_23983_9826# a_23770_9826# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3031 a_63084_9778# a_63337_9765# a_62036_9103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3032 a_9503_n4464# a_9756_n4477# a_8451_n4283# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3033 a_11080_986# a_15705_5267# a_15781_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3034 vdd a_52889_n8891# a_52681_n8891# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3035 a_71769_n12759# a_71856_n11250# a_71811_n11237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3036 a_84756_12064# a_85009_12051# a_83704_12245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3037 gnd d1 a_8447_3088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3038 a_23192_n10426# a_22979_n10426# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3039 a_22720_3822# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3040 a_33849_5263# a_33428_5263# a_33020_5342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3041 a_36440_n5874# a_36227_n5874# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3042 a_2515_8234# a_3754_7554# a_3911_6228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3043 gnd d3 a_28630_5211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3044 gnd d1 a_30121_12061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3045 vdd a_20202_6045# a_19994_6045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3046 a_2094_6787# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3047 a_79057_10587# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3048 a_65446_9514# a_66067_9830# a_66275_9830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3049 a_72995_3276# a_74092_3082# a_74047_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3050 a_19159_n4289# a_20256_n4483# a_20211_n4470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3051 a_68347_4585# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3052 a_18904_10550# a_19157_10537# a_17457_9783# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3053 a_48780_n5913# a_48730_n5926# a_48465_n8839# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3054 vdd a_51840_n5920# a_51632_n5920# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3055 a_66273_3143# a_65852_3143# a_65444_3251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3056 a_20205_n11069# a_20462_n11259# a_19161_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3057 a_12437_n5869# a_13277_n5194# a_13485_n5194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3058 a_33851_9145# a_33430_9145# a_33019_8565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3059 vdd d1 a_73254_9094# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3060 a_33427_8230# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3061 a_55935_3814# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3062 a_30911_3951# a_31168_3761# a_29867_3099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3063 vdd d0 a_52628_12738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3064 a_76412_n12641# a_77033_n12720# a_77241_n12720# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3065 a_68391_12115# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3066 a_34478_9820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3067 a_9501_n10472# a_9754_n10485# a_8449_n10291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3068 vdd a_62547_n14901# a_62339_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3069 a_13486_n8161# a_14725_n7394# a_14876_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3070 a_76153_14317# a_76774_14238# a_76982_14238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3071 a_33903_n7391# a_33690_n7391# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3072 a_49880_12756# a_50133_12743# a_49838_11234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3073 vdd a_52627_3763# a_52419_3763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3074 gnd d0 a_74560_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3075 a_54479_4153# a_55100_4586# a_55308_4586# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3076 a_54888_12793# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3077 a_45649_12795# a_46888_13562# a_47045_12236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3078 a_72997_10731# a_73254_10541# a_71554_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3079 a_1046_8238# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3080 vdd d2 a_71804_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3081 a_36549_n5874# a_36185_n7396# a_35159_n6716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3082 vdd a_40828_3080# a_40620_3080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3083 a_74044_12247# a_74049_11229# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3084 a_65704_n12379# a_66324_n11873# a_66532_n11873# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3085 gnd d1 a_51579_3088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3086 a_13485_n3747# a_13064_n3747# a_12437_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3087 vdd d1 a_19154_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3088 a_55568_n13397# a_55147_n13397# a_54739_n13830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3089 a_39390_n8202# a_39643_n8215# a_39343_n6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3090 vdd d0 a_63334_6724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3091 a_25581_12115# a_25217_10593# a_24191_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3092 vdd a_63335_5204# a_63127_5204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3093 a_25678_6107# a_26538_9142# a_26746_9142# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3094 a_67581_n12718# a_68820_n13398# a_68971_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3095 a_1468_4592# a_1047_4592# a_639_4700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3096 gnd d1 a_8448_13510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3097 vdd a_83959_7494# a_83751_7494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3098 a_33019_7659# a_33019_7118# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3099 vdd d0 a_9755_n12773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3100 a_77243_n8159# a_78083_n8163# a_78291_n8163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3101 a_76982_14238# a_77822_14234# a_78030_14234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3102 a_9241_7511# a_9237_7688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3103 a_74309_n8880# a_74562_n8893# a_73257_n8699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3104 gnd a_27824_n9799# a_27616_n9799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3105 a_27006_n8841# a_27479_n5928# a_27321_n5915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3106 gnd a_52628_13506# a_52420_13506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3107 a_56149_14236# a_55936_14236# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3108 gnd a_85010_11210# a_84802_11210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3109 a_17457_9783# a_17710_9770# a_17410_11405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3110 a_44392_4592# a_44179_4592# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3111 a_30128_n4462# a_30381_n4475# a_28681_n5229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3112 vdd a_50351_n6762# a_50143_n6762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3113 a_31177_n6754# a_31430_n6767# a_30129_n7429# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3114 a_66534_n5186# a_67374_n5190# a_67582_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3115 a_41879_n13270# a_41883_n14215# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3116 a_1519_n10424# a_1306_n10424# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3117 a_54740_n4855# a_54740_n5111# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3118 a_11608_n3664# a_11608_n4059# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3119 gnd a_32426_n1647# a_32218_n1647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3120 a_83704_13692# a_84801_13498# a_84756_13511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3121 a_78289_n12724# a_77868_n12724# a_77241_n13399# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3122 a_54481_11352# a_55102_11273# a_55310_11273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3123 a_55567_n11877# a_56407_n11202# a_56615_n11202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3124 a_23140_6110# a_22719_6110# a_22311_6218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3125 gnd a_9497_11218# a_9289_11218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3126 a_57382_4581# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3127 a_62036_10550# a_63129_11212# a_63080_11402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3128 gnd a_85007_8169# a_84799_8169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3129 a_33902_n3745# a_33689_n3745# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3130 a_12804_14236# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3131 a_66066_12118# a_65853_12118# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3132 a_36552_n11763# a_36182_n10437# a_35156_n11204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3133 a_82256_3950# a_83752_3080# a_83707_3093# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3134 a_9243_14198# a_11348_14319# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3135 a_1730_n7383# a_1309_n7383# a_901_n7816# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3136 a_33022_10159# a_33022_9903# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3137 gnd a_31427_n9808# a_31219_n9808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3138 a_40576_13515# a_41669_14177# a_41620_14367# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3139 vdd d0 a_20462_n11938# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3140 a_51325_7515# a_52418_8177# a_52373_8190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3141 a_33640_7551# a_33427_7551# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3142 a_1729_n5863# a_2569_n5188# a_2777_n5188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3143 gnd d1 a_30382_n8889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3144 a_12178_10594# a_11757_10594# a_11349_10702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3145 a_54739_n13034# a_55360_n12718# a_55568_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3146 a_50141_n8194# a_51633_n7440# a_51584_n7250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3147 a_76152_3245# a_76154_3146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3148 a_63080_9955# a_63337_9765# a_62036_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3149 a_50096_n12757# a_50349_n12770# a_49026_n9607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3150 a_77032_n11879# a_76819_n11879# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3151 a_84752_12241# a_85009_12051# a_83704_12245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3152 a_71551_6746# a_73043_7500# a_72998_7513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3153 gnd d0 a_63336_13500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3154 vdd d0 a_31428_n14222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3155 a_62030_3272# a_63127_3078# a_63082_3091# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3156 a_2778_n8155# a_4017_n7388# a_4168_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3157 a_44032_n5755# a_44653_n5863# a_44861_n5863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3158 a_1467_8238# a_1046_8238# a_638_7922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3159 a_76414_n8475# a_77035_n8159# a_77243_n8159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3160 vdd d3 a_28630_5211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3161 a_79315_n13404# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3162 a_18902_4542# a_19995_5204# a_19946_5394# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3163 a_67322_14240# a_66901_14240# a_66274_14244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3164 vdd d1 a_30121_12061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3165 gnd a_28674_12741# a_28466_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3166 vdd a_9754_n11253# a_9546_n11253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3167 a_62293_n10474# a_62546_n10487# a_60846_n11241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3168 a_9241_6064# a_9494_6051# a_8189_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3169 gnd a_7262_n8207# a_7054_n8207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3170 a_41623_4536# a_41619_4713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3171 a_78291_n8163# a_77870_n8163# a_77243_n8159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3172 vdd d0 a_74300_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3173 a_39388_n14210# a_40880_n13456# a_40835_n13443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3174 vdd d0 a_20204_13500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3175 a_33687_n9753# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3176 a_22933_3143# a_22720_3143# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3177 a_41883_n13447# a_42136_n13460# a_40831_n13266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3178 gnd a_63594_n10491# a_63386_n10491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3179 a_79316_n4429# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3180 a_62034_3095# a_62287_3082# a_60583_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3181 a_25579_6107# a_25215_4585# a_24189_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3182 a_74045_9280# a_74302_9090# a_72997_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3183 vdd a_19416_n5926# a_19208_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3184 a_65443_8315# a_65443_7920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3185 a_901_n8722# a_898_n9410# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3186 a_44391_8238# a_44178_8238# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3187 gnd a_84220_n14903# a_84012_n14903# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3188 a_74305_n8024# a_74562_n8214# a_73261_n8876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3189 a_82519_n11243# a_82772_n11256# a_82477_n12765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3190 a_67161_n5190# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3191 a_66113_n4418# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3192 a_899_n12633# a_899_n13028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3193 a_47399_n5866# a_48257_n8839# a_48465_n8839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3194 a_44602_11279# a_44181_11279# a_43773_11358# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3195 a_41885_n7439# a_41881_n7262# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3196 a_71771_n6751# a_72024_n6764# a_70703_n9786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3197 a_4173_n5747# a_3803_n4421# a_2777_n3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3198 a_17668_n12586# a_17925_n12776# a_16602_n9613# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3199 a_51587_n5907# a_52680_n5245# a_52631_n5055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3200 a_19950_5217# a_20203_5204# a_18902_4542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3201 a_55100_3139# a_54887_3139# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3202 a_49876_12933# a_50133_12743# a_49838_11234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3203 a_54738_n9672# a_55359_n9751# a_55567_n9751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3204 a_54478_6469# a_54478_6214# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3205 a_83968_n5915# a_85061_n5253# a_85016_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3206 a_22719_8236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3207 vdd a_41089_n5928# a_40881_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3208 gnd a_31428_n12775# a_31220_n12775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3209 a_76411_n10865# a_77032_n10432# a_77240_n10432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3210 a_22932_6789# a_22719_6789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3211 a_6744_12933# a_8240_12063# a_8191_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3212 a_44393_12120# a_44180_12120# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3213 a_30123_n14707# a_30380_n14897# a_28676_n14027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3214 vdd a_84222_n7448# a_84014_n7448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3215 a_12228_n14165# a_12015_n14165# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3216 vdd d1 a_73511_n10483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3217 a_12176_3818# a_11755_3818# a_11347_3502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3218 a_41623_4536# a_41876_4523# a_40571_4717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3219 a_28635_n6574# a_28727_n8209# a_28682_n8196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3220 a_52631_n3608# a_52888_n3798# a_51587_n4460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3221 a_33428_3137# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3222 a_11349_9255# a_11970_9147# a_12178_9147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3223 a_68862_n11876# a_68649_n11876# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3224 a_65704_n13826# a_65704_n14082# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3225 a_56357_14236# a_57596_13556# a_57753_12230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3226 a_33279_n10865# a_33279_n11121# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3227 a_77607_6779# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3228 a_73000_13521# a_73253_13508# a_71553_12754# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3229 a_75776_984# a_75563_984# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3230 gnd a_71804_6733# a_71596_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3231 a_52634_n13439# a_52630_n13262# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3232 a_3757_10595# a_3544_10595# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3233 a_66272_8236# a_67112_8232# a_67320_8232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3234 a_9504_n6752# a_9757_n6765# a_8456_n7427# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3235 a_20209_n10478# a_20205_n10301# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3236 vdd d1 a_8448_13510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3237 a_14881_n5753# a_14511_n4427# a_13485_n5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3238 a_54740_n3408# a_63339_n3614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3239 a_29862_7690# a_30959_7496# a_30914_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3240 gnd d3 a_6957_5213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3241 vdd a_63596_n3804# a_63388_n3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3242 a_41624_12743# a_41877_12730# a_40576_12068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3243 a_23193_n13393# a_22980_n13393# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3244 a_79269_13554# a_79056_13554# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3245 a_13226_11269# a_12805_11269# a_12178_10594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3246 a_22722_10598# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3247 gnd a_63334_6724# a_63126_6724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3248 vdd d1 a_8706_n11928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3249 a_54738_n10863# a_54738_n11119# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3250 a_15781_9138# a_15360_9138# a_14713_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3251 a_19164_n7433# a_20257_n6771# a_20212_n6758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3252 vdd d6 a_10753_n1645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3253 vdd a_9757_n8891# a_9549_n8891# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3254 vdd d3 a_39600_n6770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3255 a_57424_6103# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3256 a_12175_6106# a_11754_6106# a_11346_6214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3257 vdd a_85010_11210# a_84802_11210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3258 a_17453_9960# a_17710_9770# a_17410_11405# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3259 a_56616_n12722# a_56195_n12722# a_55568_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3260 a_14512_n7394# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3261 a_11608_n5506# a_12229_n5190# a_12437_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3262 a_66274_12118# a_67114_12793# a_67322_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3263 a_76561_14238# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3264 a_14879_n11761# a_14509_n10435# a_13483_n9755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3265 a_62036_10550# a_63129_11212# a_63084_11225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3266 a_46675_13562# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3267 a_45441_12795# a_45228_12795# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3268 a_14251_13556# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3269 a_23401_n14840# a_22980_n14840# a_21274_n15026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3270 a_25690_n7390# a_25477_n7390# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3271 a_62289_n10297# a_63386_n10491# a_63337_n10301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3272 gnd d0 a_85267_n9814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3273 vdd a_8708_n5920# a_8500_n5920# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3274 a_65445_12481# a_65445_12226# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3275 a_33643_10592# a_33430_10592# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3276 a_1307_n14159# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3277 a_2515_8234# a_2094_8234# a_1467_8238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3278 a_83705_9278# a_84802_9084# a_84753_9274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3279 vdd d0 a_85270_n8899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3280 a_640_13675# a_1261_13567# a_1469_13567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3281 vdd d0 a_9496_12738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3282 a_30912_13694# a_31169_13504# a_29864_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3283 a_82518_n8025# a_84014_n8895# a_83965_n8705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3284 a_9499_n5734# a_9756_n5924# a_8451_n5730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3285 a_67323_9826# a_66902_9826# a_66275_9151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3286 a_68559_7552# a_68346_7552# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3287 a_60587_3775# a_60840_3762# a_60540_5397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3288 a_12437_n3743# a_12016_n3743# a_11608_n3664# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3289 a_66064_7557# a_65851_7557# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3290 a_43772_13930# a_44393_14246# a_44601_14246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3291 a_1048_12799# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3292 a_23401_n12714# a_22980_n12714# a_22572_n12635# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3293 vdd a_28674_12741# a_28466_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3294 a_23770_9826# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3295 a_66535_n7385# a_66114_n7385# a_65706_n7818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3296 a_9237_6241# a_9494_6051# a_8189_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3297 a_11348_12872# a_11348_12477# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3298 a_43773_9911# a_43773_9516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3299 a_77609_14234# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3300 a_25257_6107# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3301 a_73254_n11740# a_73511_n11930# a_71807_n11060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3302 a_39390_n8202# a_40882_n7448# a_40833_n7258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3303 gnd d1 a_51580_12063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3304 a_44438_n11192# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3305 a_27571_n9786# a_28684_n6764# a_28635_n6574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3306 gnd a_8447_3088# a_8239_3088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3307 a_54481_11608# a_55101_12114# a_55309_12114# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3308 a_58006_n11880# a_57897_n11880# a_58105_n11880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3309 a_44033_n6625# a_44654_n6704# a_44862_n6704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3310 a_62030_3272# a_62287_3082# a_60583_3952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3311 vdd d1 a_84221_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3312 a_26538_9142# a_26325_9142# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3313 vref a_640_14325# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3314 a_23195_n8832# a_22982_n8832# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3315 a_57594_7548# a_57381_7548# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3316 a_78029_3812# a_77608_3812# a_76981_3137# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3317 a_78082_n5196# a_77869_n5196# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3318 a_33281_n5763# a_33902_n5871# a_34110_n5871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3319 a_28679_n11237# a_30171_n10483# a_30122_n10293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3320 a_641_9516# a_641_9261# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3321 a_76154_9253# a_76775_9145# a_76983_9145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3322 a_55148_n4422# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3323 a_41620_13688# a_41624_12743# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3324 a_56197_n6714# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3325 a_1260_5271# a_1047_5271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3326 a_76414_n7283# a_77035_n7391# a_77243_n7391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3327 a_11967_6785# a_11754_6785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3328 a_45907_n11196# a_45486_n11196# a_44859_n11192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3329 a_85014_n11248# a_85010_n11071# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3330 a_44600_3824# a_45440_3820# a_45648_3820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3331 a_13484_n14169# a_13063_n14169# a_12436_n14844# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3332 a_67112_6785# a_66899_6785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3333 a_9500_n6575# a_9504_n7431# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3334 a_54889_11273# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3335 a_38275_n9615# a_39390_n12778# a_39341_n12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3336 vdd a_73254_9094# a_73046_9094# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3337 a_14507_12111# a_14294_12111# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3338 a_40831_n13266# a_41088_n13456# a_39388_n14210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3339 a_13224_3814# a_12803_3814# a_12176_3818# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3340 gnd a_83962_10535# a_83754_10535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3341 a_65705_n5107# a_66326_n5186# a_66534_n5186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3342 a_6744_12933# a_8240_12063# a_8195_12076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3343 gnd a_51580_12063# a_51372_12063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3344 vdd d1 a_62546_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3345 a_41619_4713# a_41876_4523# a_40571_4717# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3346 a_2310_9828# a_2097_9828# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3347 gnd a_31170_9769# a_30962_9769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3348 a_44651_n11871# a_44438_n11871# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3349 a_36648_n5874# a_37506_n8847# a_37714_n8847# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3350 a_60589_9783# a_62081_10537# a_62032_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3351 a_11346_7916# a_11967_8232# a_12175_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3352 vdd d0 a_42136_n13460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3353 gnd a_85270_n8220# a_85062_n8220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3354 a_21816_973# a_21395_973# a_21717_973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3355 a_80586_9136# a_80165_9136# a_79520_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3356 vdd a_74561_n4479# a_74353_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3357 a_30915_3095# a_31168_3082# a_29863_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3358 a_3804_n7388# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3359 a_900_n5500# a_1521_n5184# a_1729_n5184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3360 vdd a_43488_n1602# a_43280_n1602# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3361 a_73255_n13260# a_74352_n13454# a_74303_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3362 vdd d5 a_5806_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3363 a_21395_973# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3364 vdd d0 a_20463_n14905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3365 vdd a_71804_6733# a_71596_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3366 vdd a_30382_n8889# a_30174_n8889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3367 a_70223_5271# a_69802_5271# a_69878_9142# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3368 a_22571_n9412# a_22571_n9668# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3369 a_6743_3958# a_8239_3088# a_8194_3101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3370 vdd d3 a_6957_5213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3371 a_5638_8199# a_5891_8186# a_5319_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3372 a_41620_12920# a_41877_12730# a_40576_12068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3373 a_33019_6467# a_33640_6783# a_33848_6783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3374 vdd a_19154_6049# a_18946_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3375 a_1520_n12712# a_1307_n12712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3376 a_33688_n14846# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3377 gnd a_52627_3084# a_52419_3084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3378 a_47040_12117# a_46676_10595# a_45650_9828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3379 a_66067_10598# a_65854_10598# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3380 a_24191_9826# a_25430_10593# a_25581_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3381 gnd d1 a_30119_6053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3382 a_34111_n8159# a_33690_n8159# a_33282_n8475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3383 a_66534_n3739# a_66113_n3739# a_65705_n4055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3384 vdd a_63334_6724# a_63126_6724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3385 a_1728_n14838# a_1307_n14838# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3386 vdd d0 a_20202_7492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3387 a_71769_n12759# a_71856_n11250# a_71807_n11060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3388 a_4059_n5866# a_3846_n5866# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3389 gnd d4 a_59991_n9803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3390 a_34110_n5871# a_33689_n5871# a_33281_n5763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3391 a_41881_n6583# a_41885_n7439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3392 vdd a_50392_n14215# a_50184_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3393 a_8191_12253# a_9288_12059# a_9243_12072# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3394 a_17454_6742# a_17707_6729# a_17412_5220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3395 a_41881_n7262# a_42138_n7452# a_40833_n7258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3396 a_76983_9824# a_76562_9824# a_76154_9508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3397 a_1729_n3737# a_1308_n3737# a_900_n3658# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3398 a_24030_n8157# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3399 a_33850_12791# a_33429_12791# a_33021_12475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3400 a_76413_n3666# a_77034_n3745# a_77242_n3745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3401 gnd d0 a_63334_6045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3402 a_66114_n6706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3403 a_48780_n5913# a_48730_n5926# a_48681_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3404 a_65852_3822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3405 a_1728_n12712# a_1307_n12712# a_899_n12633# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3406 gnd a_51840_n5920# a_51632_n5920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3407 a_55362_n8836# a_55149_n8836# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3408 gnd a_85009_14177# a_84801_14177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3409 a_19948_9276# a_19949_8184# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3410 a_20209_n11246# a_20462_n11259# a_19161_n11921# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3411 vdd a_28934_n5242# a_28726_n5242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3412 a_10758_986# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3413 a_12436_n14844# a_12015_n14844# a_10566_n15020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3414 a_56358_9822# a_55937_9822# a_55310_9147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3415 a_76983_11271# a_76562_11271# a_76154_11350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3416 a_34108_n11879# a_34948_n11204# a_35156_n11204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3417 a_83705_9278# a_84802_9084# a_84757_9097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3418 a_62035_13517# a_63128_14179# a_63079_14369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3419 vdd d0 a_52887_n12773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3420 a_52630_n12583# a_52634_n13439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3421 a_71769_n12759# a_72022_n12772# a_70699_n9609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3422 a_13483_n11202# a_14722_n10435# a_14879_n11761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3423 a_57899_n5872# a_57686_n5872# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3424 a_85015_n12768# a_85268_n12781# a_83967_n13443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3425 a_60583_3952# a_60840_3762# a_60540_5397# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3426 vdd d1 a_40828_4527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3427 vdd a_42137_n5253# a_41929_n5253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3428 a_22572_n12635# a_23193_n12714# a_23401_n12714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3429 a_60586_6742# a_62078_7496# a_62029_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3430 vdd d1 a_8709_n8887# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3431 a_29869_9107# a_30122_9094# a_28418_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3432 a_76772_6783# a_76559_6783# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3433 a_19157_n10297# a_20254_n10491# a_20209_n10478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3434 a_33281_n4857# a_33902_n4424# a_34110_n4424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3435 gnd d3 a_17665_5207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3436 a_83709_9101# a_83962_9088# a_82258_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3437 a_41882_n10480# a_41878_n10303# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3438 vdd d1 a_51580_12063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3439 a_62289_n11744# a_62546_n11934# a_60842_n11064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3440 a_62034_3095# a_63127_3757# a_63078_3947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3441 a_22934_13565# a_22721_13565# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3442 a_13275_n9755# a_13062_n9755# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3443 a_10595_n1632# a_10545_n1645# a_5648_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3444 vdd a_74559_n10487# a_74351_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3445 a_639_5606# a_639_5350# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3446 a_63084_9099# a_63337_9086# a_62032_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3447 a_63341_n9799# a_63594_n9812# a_62293_n10474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3448 vdd a_52889_n8212# a_52681_n8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3449 a_12016_n5190# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3450 gnd a_20464_n4483# a_20256_n4483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3451 a_66901_12793# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3452 a_40575_3093# a_40828_3080# a_39124_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3453 vdd a_17968_n14221# a_17760_n14221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3454 gnd d0 a_52627_5210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3455 a_74046_8188# a_74042_8365# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3456 a_22720_3143# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3457 a_44651_n10424# a_44438_n10424# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3458 a_22312_3901# a_22933_3822# a_23141_3822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3459 vdd d1 a_8707_n14895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3460 vdd a_83962_10535# a_83754_10535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3461 gnd a_50394_n8207# a_50186_n8207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3462 a_74303_n14032# a_74560_n14222# a_73259_n14884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3463 a_63338_n13268# a_63342_n14213# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3464 vdd a_51580_12063# a_51372_12063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3465 a_14874_n11880# a_14510_n13402# a_13484_n12722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3466 a_44441_n7383# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3467 a_34948_n11204# a_34735_n11204# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3468 a_50092_n12580# a_50184_n14215# a_50139_n14202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3469 a_30911_3272# a_31168_3082# a_29863_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3470 vdd d0 a_52628_12059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3471 a_9240_11408# a_9497_11218# a_8196_10556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3472 a_65443_7665# a_66064_7557# a_66272_7557# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3473 a_33640_6104# a_33427_6104# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3474 a_36292_6220# a_35922_7546# a_34896_6779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3475 vdd a_20462_n9812# a_20254_n9812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3476 a_5634_8376# a_5891_8186# a_5319_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3477 a_52635_n5232# a_52631_n5055# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3478 a_47397_n11874# a_46976_n11874# a_47303_n11755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3479 vdd a_52627_3084# a_52419_3084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3480 gnd d0 a_20462_n11938# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3481 gnd d0 a_74560_n14222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3482 a_3908_12117# a_3544_10595# a_2518_11275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3483 a_74042_7686# a_74299_7496# a_72994_7690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3484 a_24449_n14165# a_25688_n13398# a_25839_n11876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3485 a_54888_12114# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3486 a_56355_8228# a_57594_7548# a_57751_6222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3487 a_45700_n14163# a_45487_n14163# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3488 a_1049_9832# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3489 vdd d1 a_30119_6053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3490 a_48129_5273# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3491 a_63083_12745# a_63336_12732# a_62035_12070# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3492 a_11606_n11769# a_11607_n12383# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3493 a_75563_984# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3494 a_33689_n5871# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3495 a_17453_9960# a_18949_9090# a_18900_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3496 a_65703_n11510# a_66324_n11194# a_66532_n11194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3497 a_66275_11277# a_67115_11273# a_67323_11273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3498 gnd a_6957_5213# a_6749_5213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3499 a_34691_11267# a_34478_11267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3500 a_73255_n14707# a_73512_n14897# a_71808_n14027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3501 a_79518_6101# a_79097_6101# a_79424_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3502 vdd d2 a_39383_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3503 a_57847_12111# a_58705_9138# a_58913_9138# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3504 a_63342_n14892# a_63595_n14905# a_62290_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3505 a_15918_5267# a_15705_5267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3506 vdd d0 a_63334_6045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3507 a_45442_11275# a_45229_11275# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3508 vdd d0 a_74562_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3509 a_35965_6101# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3510 a_39388_n14210# a_40880_n13456# a_40831_n13266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3511 a_3911_6228# a_3541_7554# a_2515_6787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3512 a_33641_4584# a_33428_4584# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3513 a_35157_n12724# a_34736_n12724# a_34109_n12720# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3514 a_19946_5394# a_19950_4538# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3515 a_3911_6228# a_3797_6109# a_4005_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3516 gnd a_19416_n5926# a_19208_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3517 vdd d0 a_63597_n8897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3518 a_34110_n5192# a_34950_n5196# a_35158_n5196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3519 a_76154_10700# a_76775_10592# a_76983_10592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3520 a_25688_n13398# a_25475_n13398# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3521 a_2567_n9749# a_2354_n9749# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3522 a_74309_n8201# a_74562_n8214# a_73261_n8876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3523 a_48681_n5736# a_49075_n9797# a_49030_n9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3524 a_45487_n12716# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3525 a_77243_n7391# a_78083_n6716# a_78291_n6716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3526 a_17408_5397# a_17500_3762# a_17451_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3527 a_5073_9144# a_4652_9144# a_4005_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3528 gnd d2 a_71806_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3529 a_44440_n3737# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3530 a_55102_10594# a_54889_10594# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3531 a_17672_n12763# a_17925_n12776# a_16602_n9613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3532 a_1049_11279# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3533 gnd d2 a_82513_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3534 a_54481_9905# a_55102_9826# a_55310_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3535 gnd a_41089_n5928# a_40881_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3536 gnd a_71762_5211# a_71554_5211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3537 a_11349_10161# a_11349_9905# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3538 gnd a_84222_n7448# a_84014_n7448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3539 a_9499_n5734# a_9504_n6752# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3540 gnd a_85010_9763# a_84802_9763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3541 vdd a_20463_n13458# a_20255_n13458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3542 a_51585_n10468# a_52678_n9806# a_52633_n9793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3543 a_19160_n7256# a_19417_n7446# a_17717_n8200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3544 vdd d0 a_20462_n11259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3545 a_85017_n7439# a_85270_n7452# a_83965_n7258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3546 a_35158_n3749# a_34737_n3749# a_34110_n4424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3547 a_51322_3278# a_51579_3088# a_49875_3958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3548 a_33850_14238# a_33429_14238# a_33021_14317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3549 a_76820_n13399# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3550 a_22314_10706# a_22314_10165# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3551 vdd d2 a_61099_n11254# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3552 a_29867_4546# a_30960_5208# a_30911_5398# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3553 a_63080_9276# a_63337_9086# a_62032_9280# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3554 a_23980_8232# a_23767_8232# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3555 a_30125_n7252# a_31222_n7446# a_31177_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3556 a_63077_8361# a_63081_7505# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3557 a_40571_3270# a_40828_3080# a_39124_3950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3558 a_62031_13694# a_62288_13504# a_60588_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3559 vdd d0 a_52627_5210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3560 a_40575_4540# a_41668_5202# a_41623_5215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3561 a_44601_14246# a_44180_14246# a_43772_13930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3562 a_57748_12111# a_57639_12111# a_57847_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3563 a_22574_n7818# a_23195_n7385# a_23403_n7385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3564 a_44032_n5105# a_44653_n5184# a_44861_n5184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3565 a_62292_n8703# a_63389_n8897# a_63340_n8707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3566 a_26325_9142# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3567 a_33430_11271# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3568 a_57381_7548# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3569 a_55307_6785# a_54886_6785# a_54478_6864# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3570 a_63338_n14036# a_63595_n14226# a_62294_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3571 a_29862_7690# a_30119_7500# a_28419_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3572 a_85017_n8886# a_85013_n8709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3573 a_23142_12797# a_22721_12797# a_22313_12876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3574 vdd a_63336_14179# a_63128_14179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3575 a_20211_n5238# a_20207_n5061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3576 a_83702_7684# a_83959_7494# a_82259_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3577 gnd d1 a_8706_n11928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3578 vdd d0 a_41875_8169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3579 a_19163_n5913# a_20256_n5251# a_20207_n5061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3580 a_9244_9784# a_9240_9961# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3581 a_11754_6785# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3582 gnd d6 a_10753_n1645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3583 a_76151_8565# a_76151_8309# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3584 gnd d3 a_39600_n6770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3585 a_12177_12793# a_13017_12789# a_13225_12789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3586 a_44394_9832# a_44181_9832# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3587 a_52373_7511# a_52626_7498# a_51321_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3588 vdd d1 a_41087_n10489# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3589 a_41880_n5742# a_41885_n6760# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3590 gnd d0 a_9754_n9806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3591 a_18903_12070# a_19996_12732# a_19947_12922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3592 a_7005_n8017# a_8501_n8887# a_8456_n8874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3593 a_33281_n5508# a_33281_n5763# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3594 a_34898_14234# a_34477_14234# a_33850_14238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3595 a_1259_6791# a_1046_6791# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3596 a_33689_n4424# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3597 a_71811_n11237# a_73303_n10483# a_73254_n10293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3598 gnd a_8708_n5920# a_8500_n5920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3599 a_6700_5403# a_6792_3768# a_6743_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3600 a_9243_14198# a_9496_14185# a_8195_13523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3601 a_45649_14242# a_45228_14242# a_44601_13567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3602 a_2310_11275# a_2097_11275# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3603 a_13484_n14169# a_14723_n13402# a_14874_n11880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3604 a_48550_5273# a_48129_5273# a_48205_9144# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3605 a_11347_5344# a_11347_4949# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3606 a_22932_6110# a_22719_6110# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3607 a_63079_12922# a_63336_12732# a_62035_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3608 a_12176_3139# a_11755_3139# a_11349_3148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3609 vdd d1 a_19417_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3610 a_45650_9828# a_46889_10595# a_47040_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3611 a_9503_n5911# a_9756_n5924# a_8451_n5730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3612 vdd a_6957_5213# a_6749_5213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3613 a_54740_n4314# a_55361_n4422# a_55569_n4422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3614 gnd d1 a_8447_4535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3615 a_24190_12793# a_25429_13560# a_25586_12234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3616 a_12227_n9751# a_12014_n9751# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3617 a_49877_9966# a_51373_9096# a_51324_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3618 a_45910_n8155# a_45489_n8155# a_44862_n8151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3619 a_79359_n5874# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3620 a_55309_13561# a_54888_13561# a_54480_13128# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3621 vdd a_20202_7492# a_19994_7492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3622 a_33690_n6712# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3623 a_73258_n11917# a_73511_n11930# a_71807_n11060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3624 gnd a_20465_n6771# a_20257_n6771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3625 a_22573_n4055# a_23194_n3739# a_23402_n3739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3626 a_62296_n8880# a_63389_n8218# a_63344_n8205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3627 a_72995_4723# a_74092_4529# a_74047_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3628 vdd a_74301_12057# a_74093_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3629 gnd d1 a_84221_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3630 a_19159_n5736# a_20256_n5930# a_20211_n5917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3631 a_41624_12064# a_41877_12051# a_40572_12245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3632 a_2516_5267# a_2095_5267# a_1468_4592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3633 vdd d1 a_51839_n13448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3634 a_44652_n13391# a_44439_n13391# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3635 a_8195_12076# a_9288_12738# a_9239_12928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3636 a_8452_n7250# a_8709_n7440# a_7009_n8194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3637 a_11609_n6375# a_12229_n5869# a_12437_n5869# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3638 vdd d2 a_61101_n5246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3639 a_34737_n3749# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3640 a_30911_3951# a_30915_3095# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3641 gnd a_63334_6045# a_63126_6045# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3642 gnd d1 a_62289_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3643 a_17408_5397# a_17500_3762# a_17455_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3644 a_40576_13515# a_40829_13502# a_39129_12748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3645 vdd d2 a_71806_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3646 a_35925_10587# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3647 a_8452_n7250# a_9549_n7444# a_9504_n7431# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3648 a_9501_n11919# a_9754_n11932# a_8449_n11738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3649 vdd a_9757_n8212# a_9549_n8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3650 a_22313_14323# a_22313_13928# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3651 a_901_n6625# a_901_n7020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3652 a_65443_6218# a_65444_5604# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3653 gnd a_52629_10539# a_52421_10539# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3654 vdd d2 a_82513_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3655 a_40835_n13443# a_41088_n13456# a_39388_n14210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3656 a_79679_n11882# a_79315_n13404# a_78289_n14171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3657 a_57746_6103# a_57382_4581# a_56356_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3658 vdd a_71762_5211# a_71554_5211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3659 a_54740_n5506# a_54740_n5761# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3660 a_34949_n14171# a_34736_n14171# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3661 a_78291_n6716# a_79530_n7396# a_79681_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3662 a_45440_5267# a_45227_5267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3663 vdd a_85010_9763# a_84802_9763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3664 a_41618_6912# a_41622_6056# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3665 gnd d1 a_62546_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3666 a_55569_n3743# a_56409_n3747# a_56617_n3747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3667 a_74043_5398# a_74300_5208# a_72999_4546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3668 vdd d0 a_20203_3757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3669 a_65445_13132# a_66066_13565# a_66274_13565# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3670 a_39127_6740# a_40619_7494# a_40570_7684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3671 a_13275_n11202# a_13062_n11202# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3672 gnd d0 a_42136_n13460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3673 a_30914_7509# a_30910_7686# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3674 a_44860_n14838# a_44439_n14838# a_44031_n14730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3675 vdd a_40828_4527# a_40620_4527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3676 gnd a_74561_n4479# a_74353_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3677 gnd d1 a_51579_4535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3678 a_66902_11273# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3679 a_39128_3773# a_40620_4527# a_40571_4717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3680 gnd d5 a_5806_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3681 a_51582_n14705# a_52679_n14899# a_52630_n14709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3682 a_14975_n5872# a_14554_n5872# a_14881_n5753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3683 a_11968_3818# a_11755_3818# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3684 a_67113_3818# a_66900_3818# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3685 a_55568_n14844# a_55147_n14844# a_53698_n15020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3686 a_27006_n8841# a_26585_n8841# a_25940_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3687 a_44393_13567# a_44180_13567# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3688 vdd d0 a_9496_12059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3689 gnd a_30382_n8889# a_30174_n8889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3690 a_12015_n12718# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3691 a_9499_n5055# a_9756_n5245# a_8455_n5907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3692 a_71813_n5229# a_73305_n4475# a_73260_n4462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3693 vdd d1 a_19157_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3694 a_40833_n8705# a_41930_n8899# a_41881_n8709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3695 gnd d3 a_60799_11215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3696 gnd a_83960_3080# a_83752_3080# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3697 a_34689_5259# a_34476_5259# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3698 gnd d0 a_63337_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3699 a_1048_12120# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3700 a_66272_8236# a_65851_8236# a_65443_7920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3701 a_71551_6746# a_71804_6733# a_71509_5224# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3702 a_1261_12799# a_1048_12799# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3703 a_20206_n14715# a_21274_n15026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3704 a_23143_9830# a_23983_9826# a_24191_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3705 a_40574_6060# a_41667_6722# a_41618_6912# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3706 gnd d0 a_52626_6730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3707 a_66324_n9747# a_66111_n9747# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3708 a_76562_10592# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3709 a_85014_n11927# a_85010_n11750# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3710 a_11347_5344# a_11968_5265# a_12176_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3711 a_44178_6112# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3712 a_2517_14242# a_2096_14242# a_1469_14246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3713 gnd a_50392_n14215# a_50184_n14215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3714 a_67583_n6710# a_67162_n6710# a_66535_n6706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3715 a_43771_4159# a_43771_3903# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3716 a_23195_n8153# a_22982_n8153# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3717 a_898_n11763# a_899_n12377# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3718 a_44032_n5105# a_44032_n5500# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3719 a_36185_n7396# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3720 a_33281_n5113# a_33902_n5192# a_34110_n5192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3721 a_33687_n10432# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3722 a_65444_3901# a_65444_3506# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3723 a_14765_n11880# a_14552_n11880# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3724 a_1519_n9745# a_1306_n9745# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3725 a_30128_n5909# a_30381_n5922# a_28677_n5052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3726 a_18903_12070# a_19996_12732# a_19951_12745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3727 a_13064_n3747# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3728 a_66532_n10426# a_67372_n9751# a_67580_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3729 a_33020_3895# a_33641_3816# a_33849_3816# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3730 a_11967_6106# a_11754_6106# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3731 a_22721_14244# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3732 a_54478_7120# a_54478_6864# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3733 a_44030_n10857# a_44030_n11113# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3734 a_76411_n10865# a_76411_n11121# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3735 a_9239_14375# a_9496_14185# a_8195_13523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3736 a_82260_3773# a_83752_4527# a_83707_4540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3737 a_76151_6862# a_76151_6467# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3738 a_24188_6785# a_23767_6785# a_23140_6789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3739 a_73260_n4462# a_74353_n3800# a_65705_n3404# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3740 gnd d0 a_52628_12738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3741 a_63341_n10478# a_63337_n10301# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3742 a_44651_n11192# a_44438_n11192# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3743 a_11349_10702# a_11970_10594# a_12178_10594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3744 a_2309_12795# a_2096_12795# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3745 a_52372_11408# a_52629_11218# a_51328_10556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3746 a_84752_13688# a_85009_13498# a_83704_13692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3747 vdd d1 a_8447_4535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3748 a_41624_14190# a_43772_14325# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3749 a_33279_n11516# a_33279_n11771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3750 gnd d1 a_8709_n8887# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3751 a_22934_12118# a_22721_12118# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3752 a_22982_n7385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3753 a_44599_6112# a_45439_6787# a_45647_6787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3754 a_44179_4592# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3755 a_51586_n14882# a_52679_n14220# a_52634_n14207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3756 a_56150_11269# a_55937_11269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3757 a_8192_9286# a_8449_9096# a_6745_9966# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3758 vdd d1 a_30121_13508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3759 a_85011_n14038# a_85015_n14894# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3760 a_62293_n11921# a_62546_n11934# a_60842_n11064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3761 a_36388_12109# a_37246_9136# a_37454_9136# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3762 a_77243_n8838# a_76822_n8838# a_76414_n8730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3763 a_41620_12241# a_41877_12051# a_40572_12245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3764 a_40837_n8882# a_41930_n8220# a_41885_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3765 a_54479_4949# a_54479_4694# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3766 a_33688_n14167# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3767 a_33020_5598# a_33640_6104# a_33848_6104# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3768 a_3544_10595# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3769 a_45701_n5188# a_45488_n5188# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3770 a_41883_n14894# a_42136_n14907# a_40831_n14713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3771 a_10595_n1632# a_10545_n1645# a_10496_n1455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3772 a_83707_4540# a_84800_5202# a_84751_5392# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3773 gnd d1 a_19154_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3774 gnd a_74559_n10487# a_74351_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3775 a_24029_n3743# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3776 a_15705_5267# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3777 a_12804_12789# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3778 a_1728_n14159# a_1307_n14159# a_899_n14475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3779 vdd a_63334_6045# a_63126_6045# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3780 a_28679_n11237# a_30171_n10483# a_30126_n10470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3781 a_10496_n1455# a_16306_n5932# a_16257_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3782 a_54738_n11514# a_54738_n11769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3783 a_34110_n5192# a_33689_n5192# a_33281_n5113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3784 a_43771_4955# a_44392_5271# a_44600_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3785 a_66113_n5865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3786 a_55099_7553# a_54886_7553# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3787 a_76773_3816# a_76560_3816# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3788 a_28377_5224# a_28630_5211# a_27307_8374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3789 a_45227_3820# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3790 a_11606_n10067# a_11606_n10322# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3791 a_74309_n8880# a_74305_n8703# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3792 a_39343_n6580# a_39600_n6770# a_38279_n9792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3793 a_76983_9145# a_76562_9145# a_76151_8565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3794 a_55937_11269# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3795 a_33019_6467# a_33019_6212# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3796 a_55310_10594# a_54889_10594# a_54481_10702# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3797 a_80846_n8847# a_80425_n8847# a_79780_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3798 a_65852_3143# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3799 a_6748_12756# a_8240_13510# a_8191_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3800 vdd d1 a_73511_n11930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3801 a_55362_n8157# a_55149_n8157# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3802 a_22573_n3404# a_22573_n3660# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3803 a_13016_3814# a_12803_3814# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3804 a_12436_n14165# a_12015_n14165# a_11607_n14481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3805 vdd d7 a_64921_n1634# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3806 a_46676_10595# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3807 gnd a_82513_3760# a_82305_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3808 a_50092_n12580# a_50184_n14215# a_50135_n14025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3809 a_33428_4584# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3810 vdd d1 a_51579_4535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3811 a_65445_13132# a_65445_12876# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3812 a_24449_n14165# a_24028_n14165# a_23401_n14161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3813 a_37930_n5744# a_38187_n5934# a_32169_n1457# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3814 a_52372_9282# a_52629_9092# a_51324_9286# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3815 a_67320_8232# a_66899_8232# a_66272_8236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3816 vdd d3 a_60799_11215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3817 vdd a_83960_3080# a_83752_3080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3818 a_23143_11277# a_22722_11277# a_22314_10961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3819 vdd d0 a_63337_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3820 a_12176_4586# a_13016_5261# a_13224_5261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3821 a_22981_n3739# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3822 a_51328_10556# a_51581_10543# a_49881_9789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3823 a_45909_n5188# a_47148_n4421# a_47305_n5747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3824 a_76772_6104# a_76559_6104# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3825 a_79424_6220# a_79054_7546# a_78028_8226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3826 a_71547_6923# a_71804_6733# a_71509_5224# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3827 gnd d2 a_28673_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3828 a_51325_7515# a_52418_8177# a_52369_8367# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3829 a_40574_6060# a_41667_6722# a_41622_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3830 vdd d0 a_52626_6730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3831 a_42947_n15028# a_44652_n14838# a_44860_n14838# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3832 a_76413_n5763# a_76414_n6377# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3833 a_22719_6789# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3834 a_54739_n14086# a_54739_n14481# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3835 a_12016_n5869# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3836 a_12014_n10430# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3837 gnd d1 a_19156_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3838 vdd d4 a_49283_n9797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3839 vdd a_42135_n9814# a_41927_n9814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3840 a_62030_3272# a_63127_3078# a_63078_3268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3841 a_41879_n14038# a_42136_n14228# a_40835_n14890# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3842 a_33849_3137# a_34689_3812# a_34897_3812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3843 vdd a_59991_n9803# a_59783_n9803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3844 vdd d1 a_41090_n8895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3845 vdd a_63595_n13458# a_63387_n13458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3846 a_60849_n8200# a_62341_n7446# a_62296_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3847 a_41620_14367# a_41624_13511# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3848 a_55568_n12718# a_56408_n12722# a_56616_n12722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3849 gnd d0 a_74562_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3850 vdd a_41875_8169# a_41667_8169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3851 a_33901_n12720# a_33688_n12720# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3852 a_2568_n14163# a_2355_n14163# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3853 gnd d0 a_74300_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3854 a_22312_3251# a_22933_3143# a_23141_3143# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3855 a_64849_973# a_64740_973# a_43150_941# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3856 a_44181_9832# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3857 a_56357_14236# a_55936_14236# a_55309_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3858 a_76411_n9674# a_76411_n10069# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3859 vdd d4 a_70956_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3860 a_65853_13565# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3861 gnd a_50131_6735# a_49923_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3862 a_49838_11234# a_50091_11221# a_48770_8199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3863 a_52635_n5911# a_52631_n5734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3864 a_11970_9826# a_11757_9826# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3865 a_71765_n12582# a_72022_n12772# a_70699_n9609# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3866 a_58006_n11880# a_57642_n13402# a_56616_n14169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3867 a_34951_n8163# a_34738_n8163# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3868 a_34690_14234# a_34477_14234# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3869 a_85011_n12591# a_85268_n12781# a_83967_n13443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3870 a_77035_n7391# a_76822_n7391# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3871 a_17457_9783# a_18949_10537# a_18904_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3872 a_22311_6473# a_22932_6789# a_23140_6789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3873 a_33279_n11516# a_33900_n11200# a_34108_n11200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3874 a_9237_7688# a_9494_7498# a_8189_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3875 a_66535_n8832# a_66114_n8832# a_65703_n9412# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3876 gnd a_20463_n13458# a_20255_n13458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3877 a_52375_14198# a_52628_14185# a_51327_13523# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3878 vdd a_50391_n11248# a_50183_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3879 a_39386_n8025# a_40882_n8895# a_40833_n8705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3880 a_19164_n7433# a_19417_n7446# a_17717_n8200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3881 gnd a_8447_4535# a_8239_4535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3882 gnd d1 a_51580_13510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3883 gnd d0 a_20462_n11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3884 a_62030_4719# a_62287_4529# a_60587_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3885 a_25216_13560# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3886 a_30912_12926# a_30916_12070# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3887 a_18899_12247# a_19156_12057# a_17452_12927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3888 a_1049_9153# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3889 a_77821_3812# a_77608_3812# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3890 gnd d2 a_61099_n11254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3891 a_41879_n14717# a_42947_n15028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3892 a_63083_12066# a_63336_12053# a_62031_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3893 a_11970_11273# a_11757_11273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3894 a_76411_n11771# a_77032_n11879# a_77240_n11879# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3895 a_52633_n9793# a_52629_n9616# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3896 a_30125_n7252# a_31222_n7446# a_31173_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3897 a_79312_12109# a_79099_12109# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3898 a_33689_n5192# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3899 vdd a_20464_n4483# a_20256_n4483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3900 a_45700_n12716# a_45487_n12716# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3901 a_28373_5401# a_28630_5211# a_27307_8374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3902 gnd a_7001_12743# a_6793_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3903 a_2515_6787# a_2094_6787# a_1467_6112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3904 gnd d3 a_72022_n12772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3905 a_47300_n5866# a_47191_n5866# a_47399_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3906 gnd d0 a_85268_n12781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3907 a_22980_n13393# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3908 gnd a_74301_12736# a_74093_12736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3909 a_63342_n14213# a_63595_n14226# a_62294_n14888# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3910 a_57384_10589# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3911 a_22571_n9668# a_23192_n9747# a_23400_n9747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3912 gnd d0 a_74561_n3800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3913 a_76152_4692# a_76152_4151# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3914 vdd d0 a_31429_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3915 a_43772_12878# a_44393_12799# a_44601_12799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3916 a_77241_n14846# a_78081_n14171# a_78289_n14171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3917 a_44654_n8151# a_44441_n8151# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3918 a_36397_n4429# a_36184_n4429# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3919 a_6748_12756# a_8240_13510# a_8195_13523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3920 vdd d1 a_40830_9088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3921 gnd a_51580_13510# a_51372_13510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3922 vdd d1 a_62546_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3923 a_24448_n9751# a_24027_n9751# a_23400_n10426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3924 vdd a_82513_3760# a_82305_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3925 a_81411_n9792# a_81664_n9805# a_81062_n5744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3926 a_63082_5217# a_63335_5204# a_62034_4542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3927 a_23981_5265# a_23768_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3928 a_11757_10594# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3929 vdd a_74561_n5926# a_74353_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3930 gnd d1 a_41087_n10489# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3931 a_62290_n13264# a_63387_n13458# a_63342_n13445# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3932 a_7005_n8017# a_8501_n8887# a_8452_n8697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3933 a_73255_n14707# a_74352_n14901# a_74303_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3934 gnd d2 a_17708_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3935 a_55308_3818# a_54887_3818# a_54479_3502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3936 vdd a_20203_3757# a_19995_3757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3937 a_20205_n10301# a_20209_n11246# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3938 a_52375_13519# a_52371_13696# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3939 a_1309_n7383# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3940 a_1262_11279# a_1049_11279# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3941 a_51324_10733# a_51581_10543# a_49881_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3942 a_54481_9255# a_55102_9147# a_55310_9147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3943 a_47149_n7388# a_46936_n7388# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3944 a_84755_3768# a_85008_3755# a_83707_3093# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3945 a_65444_4953# a_66065_5269# a_66273_5269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3946 a_77034_n3745# a_76821_n3745# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3947 a_66111_n11873# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3948 vdd d2 a_28673_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3949 vdd d0 a_74560_n14222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3950 vdd a_31429_n3800# a_31221_n3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3951 a_21717_973# a_32431_984# a_32753_984# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3952 a_11755_3818# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3953 gnd a_52627_4531# a_52419_4531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3954 a_66275_10598# a_65854_10598# a_65446_10165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3955 gnd a_85010_9084# a_84802_9084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3956 a_45439_6787# a_45226_6787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3957 vdd a_51581_9096# a_51373_9096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3958 gnd d0 a_9496_12738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3959 a_34688_6779# a_34475_6779# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3960 a_12227_n10430# a_12014_n10430# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3961 a_37246_9136# a_37033_9136# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3962 a_34476_5259# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3963 a_58008_n5872# a_57644_n7394# a_56618_n6714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3964 a_53890_986# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3965 a_22935_10598# a_22722_10598# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3966 a_39083_11403# a_39175_9768# a_39130_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3967 a_30128_n4462# a_31221_n3800# a_31172_n3610# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3968 a_5073_9144# a_5210_5273# a_5418_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3969 a_11346_6864# a_11967_6785# a_12175_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3970 a_20211_n5917# a_20207_n5740# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3971 gnd d0 a_31168_5208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3972 a_24189_3818# a_25428_4585# a_25579_6107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3973 a_6704_5226# a_6957_5213# a_5634_8376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3974 a_15833_n8845# a_15620_n8845# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3975 a_59474_8370# a_60589_5207# a_60544_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3976 a_62296_n8880# a_63389_n8218# a_63340_n8028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3977 a_23400_n9747# a_22979_n9747# a_22571_n9668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3978 a_19159_n5736# a_20256_n5930# a_20207_n5740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3979 a_58913_9138# a_58492_9138# a_57845_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3980 a_1521_n4416# a_1308_n4416# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3981 gnd d1 a_51839_n13448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3982 a_55307_6106# a_54886_6106# a_54478_6214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3983 a_2570_n6708# a_2357_n6708# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3984 vdd a_17709_12737# a_17501_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3985 vdd a_50131_6735# a_49923_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3986 a_8456_n7427# a_8709_n7440# a_7009_n8194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3987 gnd d2 a_61101_n5246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3988 a_44180_14246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3989 a_23142_12118# a_22721_12118# a_22313_12226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3990 a_56150_9822# a_55937_9822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3991 vdd d4 a_38532_n9805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3992 a_43231_n1412# a_64713_n1634# a_53727_n1632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3993 a_24240_n9751# a_24027_n9751# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3994 a_49834_11411# a_50091_11221# a_48770_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3995 a_4007_12117# a_3586_12117# a_3908_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3996 a_11754_6106# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3997 gnd a_63337_11212# a_63129_11212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3998 a_8452_n7250# a_9549_n7444# a_9500_n7254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3999 a_4005_6109# a_3584_6109# a_3906_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4000 a_9504_n6752# a_9500_n6575# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4001 a_68561_13560# a_68348_13560# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4002 a_33021_12870# a_33642_12791# a_33850_12791# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4003 a_65445_12226# a_66066_12118# a_66274_12118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4004 a_60800_n12586# a_61057_n12776# a_59734_n9613# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4005 a_44394_9153# a_44181_9153# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4006 a_56194_n11202# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4007 a_48766_8376# a_49881_5213# a_49832_5403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4008 a_20209_n9799# a_20205_n9622# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4009 a_34109_n12720# a_33688_n12720# a_33280_n12641# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4010 vdd d1 a_73512_n14897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4011 a_18899_12247# a_19996_12053# a_19947_12243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4012 a_4865_9144# a_4652_9144# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4013 a_59478_8193# a_59731_8180# a_59159_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4014 a_19157_n11744# a_20254_n11938# a_20209_n11925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4015 a_44439_n12712# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4016 a_1259_6112# a_1046_6112# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4017 a_25841_n5868# a_25477_n7390# a_24451_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4018 a_52372_10729# a_52376_9784# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4019 a_56615_n9755# a_56194_n9755# a_55567_n10430# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4020 a_1308_n3737# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4021 a_52371_14375# a_52628_14185# a_51327_13523# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4022 vdd d1 a_51580_13510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4023 vdd a_8447_4535# a_8239_4535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4024 a_9499_n5055# a_9503_n5911# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4025 a_25472_12115# a_25259_12115# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4026 a_85013_n7262# a_85270_n7452# a_83965_n7258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4027 a_17456_12750# a_18948_13504# a_18899_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4028 a_45909_n3741# a_45488_n3741# a_44861_n3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4029 a_13486_n8161# a_13065_n8161# a_12438_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4030 a_12438_n7389# a_12017_n7389# a_11609_n7281# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4031 a_55361_n3743# a_55148_n3743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4032 a_32753_984# a_37378_5265# a_37454_9136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4033 a_63079_12243# a_63336_12053# a_62031_12247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4034 a_42828_941# d8 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4035 vdd a_74559_n11934# a_74351_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4036 a_45908_n12716# a_45487_n12716# a_44860_n13391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4037 a_84755_5215# a_84751_5392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4038 a_41624_13511# a_41620_13688# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4039 a_66902_9826# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4040 a_45228_14242# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4041 a_9503_n5232# a_9756_n5245# a_8455_n5907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4042 a_71813_n5229# a_73305_n4475# a_73256_n4285# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4043 vdd a_7001_12743# a_6793_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4044 a_68389_6107# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4045 a_31175_n13441# a_31171_n13264# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4046 a_23141_3822# a_22720_3822# a_22312_3901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4047 vdd a_74301_12736# a_74093_12736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4048 gnd a_19154_6049# a_18946_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4049 a_76559_6783# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4050 a_28418_9964# a_29914_9094# a_29869_9107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4051 a_70354_n5738# a_70748_n9799# a_70703_n9786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4052 a_25689_n4423# a_25476_n4423# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4053 a_1469_14246# a_1048_14246# a_640_13930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4054 vdd a_51580_13510# a_51372_13510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4055 a_76560_3816# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4056 gnd d4 a_27564_8184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4057 a_19163_n5913# a_20256_n5251# a_20211_n5238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4058 a_85017_n6760# a_85013_n6583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4059 a_8191_12253# a_9288_12059# a_9239_12249# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4060 a_12229_n4422# a_12016_n4422# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4061 a_22572_n12379# a_22572_n12635# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4062 a_30911_4719# a_31168_4529# a_29863_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4063 vdd d2 a_17708_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4064 a_8455_n4460# a_9548_n3798# a_9499_n3608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4065 gnd a_20204_13500# a_19996_13500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4066 a_9501_n11240# a_9754_n11253# a_8453_n11915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4067 a_12803_3814# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4068 a_71811_n11237# a_73303_n10483# a_73258_n10470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4069 a_41880_n5063# a_41884_n5919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4070 a_84751_3945# a_85008_3755# a_83707_3093# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4071 a_54478_7916# a_55099_8232# a_55307_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4072 vdd a_52627_4531# a_52419_4531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4073 a_47303_n11755# a_47189_n11874# a_47397_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4074 vdd a_85010_9084# a_84802_9084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4075 vdd d1 a_30119_7500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4076 vdd d0 a_20203_3078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4077 a_13224_3814# a_14463_4581# a_14614_6103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4078 a_82261_12748# a_82514_12735# a_82219_11226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4079 a_30123_n14707# a_31220_n14901# a_31175_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4080 a_44860_n14159# a_44439_n14159# a_44031_n14080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4081 a_11347_3247# a_11349_3148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4082 a_8449_n10291# a_9546_n10485# a_9501_n10472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4083 gnd d1 a_40828_4527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4084 a_76151_6467# a_76772_6783# a_76980_6783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4085 a_78030_12787# a_79269_13554# a_79426_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4086 a_51586_n14882# a_52679_n14220# a_52630_n14030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4087 a_11968_3139# a_11755_3139# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4088 a_46978_n5866# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4089 a_55568_n14165# a_55147_n14165# a_54739_n14481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4090 gnd d1 a_73251_6053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4091 a_28682_n8196# a_30174_n7442# a_30125_n7252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4092 a_67583_n8157# a_67162_n8157# a_66535_n8832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4093 a_6700_5403# a_6957_5213# a_5634_8376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4094 vdd a_52628_12738# a_52420_12738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4095 a_63078_3947# a_63082_3091# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4096 vdd d0 a_63334_7492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4097 a_22979_n9747# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4098 a_40837_n8882# a_41930_n8220# a_41881_n8030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4099 vdd a_20465_n6771# a_20257_n6771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4100 a_39384_n14033# a_40880_n14903# a_40831_n14713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4101 a_43770_7667# a_44391_7559# a_44599_7559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4102 a_57596_13556# a_57383_13556# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4103 a_24189_3818# a_23768_3818# a_23141_3143# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4104 a_66275_9830# a_65854_9830# a_65446_9514# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4105 a_1261_12120# a_1048_12120# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4106 gnd a_74299_7496# a_74091_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4107 a_34109_n12720# a_34949_n12724# a_35157_n12724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4108 gnd d0 a_52626_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4109 a_40570_6237# a_41667_6043# a_41618_6233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4110 a_2778_n8155# a_2357_n8155# a_1730_n8151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4111 a_36289_12109# a_36180_12109# a_36388_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4112 a_33429_12112# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4113 vdd a_63337_11212# a_63129_11212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4114 a_37700_5265# a_38064_8178# a_38019_8191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4115 vdd d0 a_31430_n6767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4116 a_11969_13561# a_11756_13561# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4117 a_48766_8376# a_49881_5213# a_49836_5226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4118 a_9497_n11742# a_9754_n11932# a_8449_n11738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4119 a_47045_12236# a_46931_12117# a_47139_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4120 a_39347_n6757# a_39600_n6770# a_38279_n9792# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4121 a_55310_9826# a_54889_9826# a_54481_9905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4122 vdd d0 a_20465_n8897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4123 a_57856_n4427# a_57643_n4427# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4124 a_18899_12247# a_19996_12053# a_19951_12066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4125 a_74045_10727# a_74302_10537# a_72997_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4126 a_14881_n5753# a_14767_n5872# a_14975_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4127 a_66326_n4418# a_66113_n4418# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4128 a_40573_10725# a_41670_10531# a_41621_10721# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4129 a_33020_3245# a_33641_3137# a_33849_3137# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4130 a_59474_8370# a_59731_8180# a_59159_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4131 a_67375_n6710# a_67162_n6710# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4132 a_22313_12226# a_22314_11612# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4133 a_25940_n5868# a_26798_n8841# a_27006_n8841# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4134 a_41878_n10303# a_41882_n11248# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4135 gnd d1 a_73511_n11930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4136 gnd a_84222_n8895# a_84014_n8895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4137 a_76821_n5871# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4138 a_49875_3958# a_50132_3768# a_49832_5403# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4139 a_33282_n7824# a_33282_n8080# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4140 a_44653_n4416# a_44440_n4416# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4141 gnd d7 a_64921_n1634# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4142 a_57897_n11880# a_57684_n11880# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4143 a_81147_8368# a_82262_5205# a_82217_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4144 a_41618_6233# a_41623_5215# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4145 a_1730_n8151# a_1309_n8151# a_901_n8467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4146 gnd d0 a_52628_12059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4147 a_9244_11231# a_9497_11218# a_8196_10556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4148 a_73001_9107# a_73254_9094# a_71550_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4149 gnd d2 a_50134_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4150 a_76820_n14846# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4151 a_37714_n8847# a_38187_n5934# a_32169_n1457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4152 a_55569_n5190# a_55148_n5190# a_54740_n5111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4153 a_40571_4717# a_40828_4527# a_39128_3773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4154 a_1262_9832# a_1049_9832# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4155 a_13277_n5194# a_13064_n5194# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4156 gnd d0 a_52888_n3798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4157 a_22571_n9412# a_23195_n8832# a_23403_n8832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4158 gnd d2 a_6999_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4159 vdd a_61059_n6768# a_60851_n6768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4160 a_12228_n13397# a_12015_n13397# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4161 a_17412_5220# a_17665_5207# a_16342_8370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4162 a_55936_14236# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4163 a_63084_11225# a_63080_11402# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4164 gnd a_28675_9774# a_28467_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4165 a_57751_6222# a_57637_6103# a_57845_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4166 a_33021_13922# a_33642_14238# a_33850_14238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4167 a_77243_n8159# a_76822_n8159# a_76414_n8080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4168 a_14614_6103# a_14505_6103# a_14713_6103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4169 vdd d4 a_27564_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4170 a_54481_9510# a_54481_9255# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4171 a_23400_n11194# a_24240_n11198# a_24448_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4172 gnd a_42135_n9814# a_41927_n9814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4173 a_33020_5342# a_33020_4947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4174 a_14616_12111# a_14507_12111# a_14715_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4175 a_41883_n14215# a_42136_n14228# a_40835_n14890# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4176 vdd d3 a_72024_n6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4177 gnd d0 a_85008_5202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4178 a_1522_n6704# a_1309_n6704# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4179 gnd d2 a_39383_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4180 gnd a_63595_n13458# a_63387_n13458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4181 a_60849_n8200# a_62341_n7446# a_62292_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4182 a_65853_12118# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4183 a_39123_6917# a_39380_6727# a_39085_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4184 a_67321_5265# a_66900_5265# a_66273_4590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4185 a_52374_5223# a_52627_5210# a_51326_4548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4186 a_17668_n12586# a_17760_n14221# a_17711_n14031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4187 a_60584_12927# a_62080_12057# a_62035_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4188 a_30124_n5732# a_30381_n5922# a_28677_n5052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4189 a_66113_n5186# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4190 vdd d1 a_41087_n11936# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4191 a_44030_n10316# a_44651_n10424# a_44859_n10424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4192 a_5418_5273# a_10971_986# a_11179_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4193 a_638_6220# a_1259_6112# a_1467_6112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4194 a_76773_3137# a_76560_3137# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4195 a_44178_7559# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4196 a_79419_6101# a_79055_4579# a_78029_3812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4197 a_23980_6785# a_23767_6785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4198 a_60846_n11241# a_62338_n10487# a_62293_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4199 a_37293_n8847# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4200 a_78290_n3749# a_77869_n3749# a_77242_n4424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4201 vdd a_73512_n13450# a_73304_n13450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4202 a_65704_n12635# a_66325_n12714# a_66533_n12714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4203 a_82517_n5058# a_82774_n5248# a_82479_n6757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4204 gnd a_52887_n13452# a_52679_n13452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4205 a_76412_n13832# a_77033_n13399# a_77241_n13399# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4206 a_19158_n14711# a_20255_n14905# a_20210_n14892# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4207 a_82257_12925# a_82514_12735# a_82219_11226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4208 gnd a_40829_12055# a_40621_12055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4209 a_82477_n12765# a_82564_n11256# a_82519_n11243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4210 a_65446_10165# a_66067_10598# a_66275_10598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4211 a_76559_8230# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4212 a_45647_8234# a_46886_7554# a_47043_6228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4213 a_22574_n7277# a_22574_n7818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4214 a_6749_9789# a_7002_9776# a_6702_11411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4215 a_35922_7546# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4216 a_63338_n14715# a_64406_n15026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4217 a_76774_12112# a_76561_12112# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4218 a_12436_n12718# a_12015_n12718# a_11607_n12639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4219 a_58107_n5872# a_58965_n8845# a_59173_n8845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4220 vdd d1 a_73251_6053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4221 a_45226_6787# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4222 a_54739_n14736# a_53698_n15020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4223 a_4173_n5747# a_4059_n5866# a_4267_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4224 a_3908_12117# a_3799_12117# a_4007_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4225 a_44394_10600# a_44181_10600# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4226 a_34475_6779# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4227 a_12436_n13397# a_13276_n12722# a_13484_n12722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4228 a_31171_n12585# a_31428_n12775# a_30127_n13437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4229 gnd a_50391_n11248# a_50183_n11248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4230 a_34898_12787# a_34477_12787# a_33850_12112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4231 a_639_4700# a_1260_4592# a_1468_4592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4232 a_23193_n14161# a_22980_n14161# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4233 gnd d0 a_42138_n7452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4234 gnd a_31168_5208# a_30960_5208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4235 vdd d0 a_52626_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4236 a_23140_7557# a_23980_8232# a_24188_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4237 a_44031_n14475# a_44652_n14159# a_44860_n14159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4238 a_40570_6237# a_41667_6043# a_41622_6056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4239 a_44860_n13391# a_44439_n13391# a_44031_n13824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4240 a_45650_11275# a_45229_11275# a_44602_11279# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4241 a_10496_n1455# a_16306_n5932# a_16041_n8845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4242 a_78030_14234# a_77609_14234# a_76982_14238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4243 a_63339_n3614# a_63596_n3804# a_62295_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4244 a_76821_n4424# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4245 a_20209_n10478# a_20462_n10491# a_19157_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4246 a_44862_n8830# a_45702_n8155# a_45910_n8155# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4247 a_44032_n4849# a_44032_n5105# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4248 a_2569_n5188# a_2356_n5188# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4249 a_22571_n11765# a_23192_n11873# a_23400_n11873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4250 a_73257_n8699# a_73514_n8889# a_71810_n8019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4251 a_40835_n14890# a_41088_n14903# a_39384_n14033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4252 a_55359_n10430# a_55146_n10430# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4253 a_40573_10725# a_41670_10531# a_41625_10544# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4254 gnd d0 a_31429_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4255 a_44600_4592# a_44179_4592# a_43771_4159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4256 gnd a_63336_14179# a_63128_14179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4257 a_40577_9101# a_41670_9763# a_41621_9953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4258 gnd d0 a_52629_9771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4259 vdd d1 a_8449_9096# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4260 gnd d1 a_62546_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4261 gnd d0 a_41875_8169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4262 a_54478_6864# a_54478_6469# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4263 a_76411_n11516# a_76411_n11771# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4264 a_1468_3824# a_2308_3820# a_2516_3820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4265 a_44181_9153# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4266 a_2568_n12716# a_2355_n12716# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4267 a_12177_12793# a_11756_12793# a_11348_12872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4268 gnd d0 a_42136_n14907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4269 a_77033_n12720# a_76820_n12720# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4270 gnd a_74561_n5926# a_74353_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4271 a_74048_13517# a_74301_13504# a_72996_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4272 vdd d2 a_50134_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4273 a_43770_7922# a_43770_7667# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4274 a_60584_12927# a_60841_12737# a_60546_11228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4275 a_4652_9144# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4276 a_62290_n13264# a_63387_n13458# a_63338_n13268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4277 a_77822_12787# a_77609_12787# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4278 gnd a_17710_9770# a_17502_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4279 a_76981_5263# a_76560_5263# a_76152_4947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4280 gnd d1 a_73254_10541# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4281 a_33280_n12385# a_33900_n11879# a_34108_n11879# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4282 a_11970_9147# a_11757_9147# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4283 a_12435_n10430# a_13275_n9755# a_13483_n9755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4284 vdd d2 a_6999_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4285 vdd a_10753_n1645# a_10545_n1645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4286 a_76153_14317# a_76153_13922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4287 a_85013_n8709# a_85014_n9801# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4288 a_22312_5604# a_22932_6110# a_23140_6110# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4289 vdd a_52889_n7444# a_52681_n7444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4290 a_34951_n6716# a_34738_n6716# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4291 vdd a_28675_9774# a_28467_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4292 a_31170_n9618# a_31427_n9808# a_30126_n10470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4293 gnd d2 a_72067_n8209# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4294 a_24191_9826# a_23770_9826# a_23143_9830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4295 a_66535_n8153# a_66114_n8153# a_65706_n8469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4296 a_9239_12928# a_9243_12072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4297 a_23402_n5865# a_22981_n5865# a_22574_n6371# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4298 a_56356_5261# a_55935_5261# a_55308_4586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4299 a_83708_13515# a_83961_13502# a_82261_12748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4300 a_35967_12109# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4301 a_78031_9820# a_77610_9820# a_76983_9824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4302 a_33848_7551# a_33427_7551# a_33019_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4303 a_52634_n12760# a_52887_n12773# a_51586_n13435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4304 a_76413_n3666# a_76413_n4061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4305 a_6706_11234# a_6793_12743# a_6744_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4306 gnd d0 a_42137_n3806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4307 a_76411_n11121# a_77032_n11200# a_77240_n11200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4308 a_41885_n8886# a_42138_n8899# a_40833_n8705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4309 a_52370_5400# a_52627_5210# a_51326_4548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4310 a_46718_12117# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4311 a_55149_n6710# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4312 gnd a_27564_8184# a_27356_8184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4313 a_68820_n13398# a_68607_n13398# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4314 a_44654_n8830# a_44441_n8830# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4315 a_14554_n5872# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4316 a_54886_6785# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4317 a_7005_n8017# a_7262_n8207# a_6962_n6572# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4318 a_34897_3812# a_34476_3812# a_33849_3816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4319 a_72995_4723# a_74092_4529# a_74043_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4320 gnd a_74301_12057# a_74093_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4321 a_26585_n8841# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4322 a_33019_7118# a_33019_6862# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4323 a_9498_n14709# a_9755_n14899# a_8450_n14705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4324 a_77243_n7391# a_76822_n7391# a_76414_n7824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4325 a_43231_n1412# a_64713_n1634# a_64664_n1444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4326 a_41618_8359# a_41875_8169# a_40574_7507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4327 vdd a_62547_n13454# a_62339_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4328 a_77242_n5871# a_78082_n5196# a_78290_n5196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4329 a_66327_n6706# a_66114_n6706# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4330 vout a_2731_n1225# a_3058_n1106# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4331 vdd d1 a_62286_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4332 vdd a_40829_12055# a_40621_12055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4333 a_60804_n12763# a_61057_n12776# a_59734_n9613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4334 a_44599_8238# a_44178_8238# a_43770_7922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4335 a_2777_n3741# a_2356_n3741# a_1729_n4416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4336 a_6745_9966# a_7002_9776# a_6702_11411# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4337 a_44654_n6704# a_44441_n6704# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4338 a_65445_12876# a_65445_12481# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4339 vdd d0 a_42136_n14228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4340 a_2517_12795# a_2096_12795# a_1469_12120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4341 a_44601_13567# a_45441_14242# a_45649_14242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4342 vdd a_74561_n5247# a_74353_n5247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4343 a_44032_n3402# a_52631_n3608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4344 a_22982_n8832# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4345 a_23403_n6706# a_24243_n6710# a_24451_n6710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4346 a_57639_12111# a_57426_12111# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4347 a_19157_n11744# a_20254_n11938# a_20205_n11748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4348 a_73259_n14884# a_74352_n14222# a_74303_n14032# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4349 a_54740_n4314# a_54740_n4855# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4350 a_55308_3139# a_54887_3139# a_54481_3148# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4351 vdd a_20203_3078# a_19995_3078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4352 a_44859_n9745# a_44438_n9745# a_44030_n9666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4353 gnd d0 a_20203_3757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4354 a_84755_3089# a_85008_3076# a_83703_3270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4355 a_41620_13688# a_41877_13498# a_40572_13692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4356 a_22721_12797# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4357 a_66111_n11194# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4358 gnd a_40828_4527# a_40620_4527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4359 a_33020_4947# a_33020_4692# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4360 a_900_n5105# a_900_n5500# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4361 a_11755_3139# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4362 a_22571_n10859# a_23192_n10426# a_23400_n10426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4363 gnd a_74559_n11934# a_74351_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4364 a_70703_n9786# a_71816_n6764# a_71771_n6751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4365 gnd d0 a_9496_12059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4366 vdd a_63334_7492# a_63126_7492# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4367 a_28675_n11060# a_30171_n11930# a_30126_n11917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4368 a_30912_12247# a_30917_11229# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4369 a_79421_12109# a_79057_10587# a_78031_9820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4370 a_19952_10546# a_19948_10723# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4371 gnd d1 a_19157_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4372 vdd d3 a_72022_n12772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4373 vdd d2 a_28933_n14217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4374 vdd a_85269_n4485# a_85061_n4485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4375 a_67580_n11198# a_67159_n11198# a_66532_n11194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4376 vdd d0 a_85268_n12781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4377 a_1727_n10424# a_2567_n9749# a_2775_n9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4378 a_41881_n8030# a_42138_n8220# a_40837_n8882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4379 vdd a_49283_n9797# a_49075_n9797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4380 a_13223_8228# a_12802_8228# a_12175_7553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4381 a_40577_9101# a_41670_9763# a_41625_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4382 vdd d0 a_52629_9771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4383 a_67115_11273# a_66902_11273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4384 a_68812_12115# a_68391_12115# a_68718_12234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4385 gnd a_42136_n12781# a_41928_n12781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4386 a_1047_5271# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4387 vdd d1 a_84219_n10489# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4388 a_33851_9824# a_33430_9824# a_33022_9903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4389 a_44031_n13283# a_44652_n13391# a_44860_n13391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4390 gnd d2 a_39641_n14223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4391 a_33642_12791# a_33429_12791# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4392 a_77242_n3745# a_76821_n3745# a_76413_n4061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4393 a_79570_n11882# a_79357_n11882# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4394 a_65854_10598# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4395 gnd d2 a_50133_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4396 a_14715_12111# a_15573_9138# a_15781_9138# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4397 vdd a_17710_9770# a_17502_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4398 vdd d0 a_9756_n3798# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4399 vdd d1 a_73254_10541# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4400 a_58752_n8845# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4401 vdd d0 a_63335_3757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4402 a_11609_n8473# a_11609_n8728# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4403 a_3586_12117# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4404 gnd d1 a_30382_n7442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4405 vdd a_83960_4527# a_83752_4527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4406 gnd d3 a_39338_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4407 a_82260_3773# a_83752_4527# a_83703_4717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4408 gnd d3 a_17667_11215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4409 gnd a_50134_9776# a_49926_9776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4410 vdd d5 a_81319_n5934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4411 a_19161_n11921# a_20254_n11259# a_20209_n11246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4412 a_77032_n10432# a_76819_n10432# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4413 a_32644_984# a_32431_984# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4414 a_80425_n8847# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4415 a_52376_11231# a_52629_11218# a_51328_10556# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4416 a_9497_n10295# a_9501_n11240# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4417 a_18897_7686# a_19994_7492# a_19945_7682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4418 a_62290_n14711# a_62547_n14901# a_60843_n14031# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4419 a_8449_n10291# a_9546_n10485# a_9497_n10295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4420 a_6706_11234# a_6793_12743# a_6748_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4421 gnd a_16599_8180# a_16391_8180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4422 a_33279_n10324# a_33279_n10865# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4423 a_45489_n8155# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4424 a_62030_4719# a_63127_4525# a_63078_4715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4425 gnd d1 a_83959_7494# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4426 vdd a_74559_n11255# a_74351_n11255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4427 a_76775_10592# a_76562_10592# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4428 a_69072_n5868# a_68651_n5868# a_68978_n5749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4429 a_28681_n5229# a_28934_n5242# a_28639_n6751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4430 a_83706_6060# a_84799_6722# a_84750_6912# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4431 a_24448_n9751# a_25687_n10431# a_25844_n11757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4432 gnd a_20464_n5251# a_20256_n5251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4433 a_54479_5344# a_55100_5265# a_55308_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4434 vdd a_27564_8184# a_27356_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4435 gnd d0 a_74562_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4436 a_66274_14244# a_65853_14244# a_65445_14323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4437 a_11969_12114# a_11756_12114# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4438 a_23141_3143# a_22720_3143# a_22312_3251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4439 a_54479_4694# a_54479_4153# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4440 a_65851_8236# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4441 a_11608_n3408# a_20207_n3614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4442 gnd a_85008_5202# a_84800_5202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4443 vdd d3 a_71764_11219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4444 a_52373_6743# a_52626_6730# a_51325_6068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4445 a_67320_6785# a_66899_6785# a_66272_6110# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4446 a_66273_4590# a_65852_4590# a_65444_4698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4447 a_66532_n11873# a_66111_n11873# a_65703_n11765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4448 a_44033_n7816# a_44654_n7383# a_44862_n7383# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4449 a_45647_8234# a_45226_8234# a_44599_8238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4450 a_31176_n4466# a_31172_n4289# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4451 a_63337_n10301# a_63341_n11246# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4452 gnd d0 a_31430_n6767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4453 a_76560_3137# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4454 a_76152_3895# a_76773_3816# a_76981_3816# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4455 a_54738_n10322# a_54738_n10863# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4456 a_19949_7505# a_20202_7492# a_18897_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4457 a_50141_n8194# a_50394_n8207# a_50094_n6572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4458 a_44441_n8151# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4459 gnd a_51838_n10481# a_51630_n10481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4460 a_33903_n8838# a_33690_n8838# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4461 a_1468_5271# a_1047_5271# a_639_4955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4462 a_44861_n3737# a_45701_n3741# a_45909_n3741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4463 a_19951_14192# a_19947_14369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4464 a_11608_n3408# a_20464_n3804# a_19163_n4466# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4465 a_66066_12797# a_65853_12797# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4466 a_71767_n6574# a_71859_n8209# a_71810_n8019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4467 a_84751_3266# a_85008_3076# a_83703_3270# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4468 gnd a_20463_n14905# a_20255_n14905# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4469 gnd a_61102_n8213# a_60894_n8213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4470 a_73000_12074# a_73253_12061# a_71549_12931# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4471 a_23767_6785# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4472 a_55360_n12718# a_55147_n12718# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4473 a_11606_n10067# a_12227_n9751# a_12435_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4474 a_19164_n8880# a_19417_n8893# a_17713_n8023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4475 a_2518_9828# a_2097_9828# a_1470_9832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4476 vdd d1 a_19154_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4477 a_35159_n8163# a_34738_n8163# a_34111_n8838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4478 a_33903_n6712# a_33690_n6712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4479 a_56357_12789# a_55936_12789# a_55309_12114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4480 a_80723_5265# a_80510_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4481 a_44392_5271# a_44179_5271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4482 a_30125_n8699# a_31222_n8893# a_31173_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4483 a_65706_n6371# a_65706_n6627# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4484 a_40836_n4468# a_41929_n3806# a_41880_n3616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4485 vdd a_20464_n5930# a_20256_n5930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4486 a_3755_4587# a_3542_4587# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4487 vdd d3 a_61057_n12776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4488 a_22311_8315# a_22311_7920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4489 a_56615_n11202# a_56194_n11202# a_55567_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4490 a_76152_5598# a_76772_6104# a_76980_6104# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4491 a_74305_n8703# a_74306_n9795# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4492 gnd a_61059_n6768# a_60851_n6768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4493 a_84755_3089# a_84751_3266# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4494 a_22980_n14840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4495 a_79686_n5755# a_79316_n4429# a_78290_n5196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4496 a_13017_12789# a_12804_12789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4497 a_58837_5267# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4498 a_36395_n10437# a_36182_n10437# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4499 a_1520_n13391# a_1307_n13391# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4500 a_24450_n5190# a_24029_n5190# a_23402_n5865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4501 vdd a_52628_12059# a_52420_12059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4502 a_51582_n13258# a_51839_n13448# a_50139_n14202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4503 a_66065_3822# a_65852_3822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4504 a_45442_9828# a_45229_9828# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4505 vdd d0 a_74562_n8214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4506 vdd a_9757_n7444# a_9549_n7444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4507 vdd d0 a_31429_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4508 a_22933_3822# a_22720_3822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4509 a_12178_11273# a_11757_11273# a_11349_10957# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4510 a_55568_n12718# a_55147_n12718# a_54739_n12639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4511 a_67582_n5190# a_67161_n5190# a_66534_n5186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4512 a_66534_n4418# a_66113_n4418# a_65705_n4310# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4513 a_77869_n5196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4514 a_66275_9151# a_65854_9151# a_65443_8571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4515 gnd d3 a_72024_n6764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4516 a_77823_11267# a_77610_11267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4517 vdd d2 a_50133_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4518 a_11346_8567# a_11346_8311# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4519 a_68718_12234# a_68348_13560# a_67322_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4520 a_79317_n7396# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4521 gnd d1 a_41087_n11936# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4522 gnd a_41875_8169# a_41667_8169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4523 a_12014_n11877# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4524 a_55100_3818# a_54887_3818# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4525 a_9497_n11063# a_9754_n11253# a_8453_n11915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4526 a_60846_n11241# a_62338_n10487# a_62289_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4527 a_56196_n3747# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4528 a_68810_6107# a_68389_6107# a_68711_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4529 a_55310_9147# a_54889_9147# a_54481_9255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4530 a_69070_n11876# a_68649_n11876# a_68976_n11757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4531 a_78080_n9757# a_77867_n9757# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4532 a_52632_n8701# a_52889_n8891# a_51584_n8697# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4533 vdd d3 a_17667_11215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4534 vdd a_50134_9776# a_49926_9776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4535 a_1730_n8830# a_1309_n8830# a_898_n9410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4536 gnd a_73512_n13450# a_73304_n13450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4537 a_640_12228# a_1261_12120# a_1469_12120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4538 a_68349_10593# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4539 a_82521_n5235# a_82774_n5248# a_82479_n6757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4540 a_76980_6783# a_76559_6783# a_76151_6467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4541 a_52372_11408# a_52376_10552# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4542 a_76821_n5192# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4543 gnd d1 a_73253_13508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4544 a_74307_n13441# a_74303_n13264# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4545 a_55569_n5869# a_55148_n5869# a_54740_n5761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4546 vdd a_73513_n4475# a_73305_n4475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4547 a_11349_9510# a_11970_9826# a_12178_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4548 a_69670_9142# a_69457_9142# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4549 a_67374_n3743# a_67161_n3743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4550 a_82477_n12765# a_82564_n11256# a_82515_n11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4551 a_71548_3956# a_73044_3086# a_72995_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4552 vdd a_20463_n14226# a_20255_n14226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4553 a_52636_n8199# a_52632_n8022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4554 a_22314_10961# a_22935_11277# a_23143_11277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4555 vdd a_16599_8180# a_16391_8180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4556 a_62030_4719# a_63127_4525# a_63082_4538# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4557 a_17457_9783# a_18949_10537# a_18900_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4558 a_16602_n9613# a_17717_n12776# a_17672_n12763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4559 a_76820_n14167# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4560 vdd a_63597_n8897# a_63389_n8897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4561 a_65703_n9668# a_66324_n9747# a_66532_n9747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4562 a_56355_6781# a_55934_6781# a_55307_6106# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4563 gnd a_9755_n13452# a_9547_n13452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4564 a_22572_n13826# a_23193_n13393# a_23401_n13393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4565 a_30129_n8876# a_31222_n8214# a_31177_n8201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4566 a_28682_n8196# a_30174_n7442# a_30129_n7429# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4567 a_1730_n6704# a_1309_n6704# a_901_n6625# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4568 a_83706_6060# a_84799_6722# a_84754_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4569 a_74048_13517# a_74044_13694# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4570 a_1262_9153# a_1049_9153# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4571 a_31175_n12762# a_31428_n12775# a_30127_n13437# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4572 a_33642_14238# a_33429_14238# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4573 a_28676_n14027# a_30172_n14897# a_30127_n14884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4574 a_22574_n8469# a_23195_n8153# a_23403_n8153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4575 a_30913_9280# a_31170_9090# a_29865_9284# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4576 a_28420_3779# a_28673_3766# a_28373_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4577 a_52369_6920# a_52626_6730# a_51325_6068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4578 a_65704_n12379# a_65704_n12635# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4579 a_63078_3268# a_54481_3148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4580 a_76981_3137# a_77821_3812# a_78029_3812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4581 a_62034_4542# a_62287_4529# a_60587_3775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4582 gnd d1 a_51839_n14895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4583 a_898_n10061# a_1519_n9745# a_1727_n9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4584 a_18903_12070# a_19156_12057# a_17452_12927# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4585 a_14876_n5872# a_14512_n7394# a_13486_n6714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4586 a_76982_14238# a_76561_14238# a_76153_13922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4587 a_34738_n8163# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4588 a_67160_n12718# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4589 vdd d0 a_63595_n12779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4590 a_8452_n8697# a_9549_n8891# a_9500_n8701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4591 gnd a_39340_11213# a_39132_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4592 a_17717_n8200# a_17970_n8213# a_17670_n6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4593 a_73261_n8876# a_73514_n8889# a_71810_n8019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4594 a_22572_n13030# a_22572_n13285# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4595 a_70138_n8841# a_69717_n8841# a_69072_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4596 a_14621_12230# a_14251_13556# a_13225_12789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4597 a_4014_n10429# a_3801_n10429# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4598 a_23143_10598# a_23983_11273# a_24191_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4599 a_76152_3500# a_76152_3245# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4600 a_33429_13559# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4601 a_16346_8193# a_17459_11215# a_17410_11405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4602 a_1469_12120# a_2309_12795# a_2517_12795# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4603 a_55570_n8157# a_56410_n8161# a_56618_n8161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4604 gnd a_20205_10533# a_19997_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4605 a_23141_5269# a_23981_5265# a_24189_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4606 a_52369_6920# a_52373_6064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4607 a_3058_n1106# a_42828_941# a_21816_973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4608 a_72996_12251# a_73253_12061# a_71549_12931# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4609 a_44861_n4416# a_44440_n4416# a_44032_n4849# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4610 a_56408_n12722# a_56195_n12722# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4611 a_12438_n8836# a_12017_n8836# a_11609_n8728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4612 a_32644_984# a_32431_984# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4613 a_63079_13690# a_63336_13500# a_62031_13694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4614 a_44180_12799# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4615 a_14552_n11880# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4616 a_44031_n13028# a_44031_n13283# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4617 gnd a_20203_3757# a_19995_3757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4618 a_14722_n10435# a_14509_n10435# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4619 a_71809_n5052# a_73305_n5922# a_73256_n5732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4620 a_33848_6104# a_33427_6104# a_33020_5598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4621 gnd a_10753_n1645# a_10545_n1645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4622 a_27571_n9786# a_27824_n9799# a_27222_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4623 a_34691_9820# a_34478_9820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4624 a_54741_n6631# a_55362_n6710# a_55570_n6710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4625 a_24190_12793# a_23769_12793# a_23142_12797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4626 gnd a_52889_n7444# a_52681_n7444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4627 a_78031_9820# a_79270_10587# a_79421_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4628 gnd a_16514_n5932# a_16306_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4629 a_36178_6101# a_35965_6101# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4630 a_70443_8197# a_71556_11219# a_71511_11232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4631 a_23193_n14840# a_22980_n14840# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4632 a_54481_11352# a_54481_10957# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4633 a_74045_10727# a_74049_9782# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4634 a_31172_n3610# a_31176_n4466# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4635 a_56618_n6714# a_56197_n6714# a_55570_n7389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4636 a_35157_n12724# a_36396_n13404# a_36547_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4637 a_76153_12870# a_76774_12791# a_76982_12791# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4638 a_57597_10589# a_57384_10589# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4639 a_76154_9508# a_76775_9824# a_76983_9824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4640 a_39083_11403# a_39175_9768# a_39126_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4641 a_17668_n12586# a_17760_n14221# a_17715_n14208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4642 a_55101_12793# a_54888_12793# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4643 a_1046_6791# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4644 a_23193_n12714# a_22980_n12714# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4645 a_13065_n8161# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4646 a_68973_n5868# a_68609_n7390# a_67583_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4647 a_45488_n3741# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4648 vdd d1 a_83962_9088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4649 gnd a_8449_10543# a_8241_10543# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4650 a_45228_12795# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4651 a_22571_n11115# a_23192_n11194# a_23400_n11194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4652 gnd d3 a_60797_5207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4653 a_71807_n11060# a_73303_n11930# a_73258_n11917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4654 gnd a_17709_12737# a_17501_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4655 a_58105_n11880# a_57684_n11880# a_58011_n11761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4656 a_40573_9278# a_40830_9088# a_39126_9958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4657 gnd a_62547_n13454# a_62339_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4658 a_40573_9278# a_41670_9084# a_41621_9274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4659 gnd d0 a_52629_9092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4660 a_12014_n9751# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4661 a_2944_n1225# a_2731_n1225# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4662 a_33849_4584# a_33428_4584# a_33020_4151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4663 gnd d0 a_41878_9763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4664 a_23195_n7385# a_22982_n7385# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4665 a_57643_n4427# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4666 a_638_7126# a_1259_7559# a_1467_7559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4667 vdd a_52887_n13452# a_52679_n13452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4668 vdd a_63335_3757# a_63127_3757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4669 a_11608_n3408# a_11608_n3664# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4670 a_71548_3956# a_73044_3086# a_72999_3099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4671 a_25427_7552# a_25214_7552# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4672 a_12177_12114# a_11756_12114# a_11348_12222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4673 a_30917_11229# a_31170_11216# a_29869_10554# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4674 gnd d0 a_42136_n14228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4675 a_45699_n11196# a_45486_n11196# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4676 a_13276_n14169# a_13063_n14169# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4677 gnd a_74561_n5247# a_74353_n5247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4678 a_44440_n4416# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4679 gnd a_39338_5205# a_39130_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4680 a_17455_3775# a_17708_3762# a_17408_5397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4681 gnd a_82773_n14223# a_82565_n14223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4682 a_54887_3818# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4683 a_50098_n6749# a_50351_n6762# a_49030_n9784# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4684 a_68821_n4423# a_68608_n4423# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4685 a_3801_n10429# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4686 a_28416_3956# a_28673_3766# a_28373_5401# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4687 a_47043_6228# a_46929_6109# a_47137_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4688 a_9503_n5232# a_9499_n5055# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4689 a_66533_n14161# a_67373_n14165# a_67581_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4690 a_77608_5259# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4691 gnd a_52888_n3798# a_52680_n3798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4692 gnd a_6959_11221# a_6751_11221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4693 a_76774_13559# a_76561_13559# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4694 a_1467_6112# a_2307_6787# a_2515_6787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4695 vdd d0 a_42138_n7452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4696 a_70703_n9786# a_71816_n6764# a_71767_n6574# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4697 a_4016_n4421# a_3803_n4421# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4698 a_54478_6864# a_55099_6785# a_55307_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4699 a_23402_n5186# a_22981_n5186# a_22573_n5502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4700 a_28675_n11060# a_30171_n11930# a_30122_n11740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4701 a_48205_9144# a_47784_9144# a_47137_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4702 a_56195_n12722# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4703 a_54480_13669# a_54480_13128# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4704 a_76414_n8730# a_77035_n8838# a_77243_n8838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4705 gnd d2 a_28933_n14217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4706 gnd a_85269_n4485# a_85061_n4485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4707 vdd a_39340_11213# a_39132_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4708 a_66535_n6706# a_66114_n6706# a_65706_n6627# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4709 a_41885_n8207# a_42138_n8220# a_40837_n8882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4710 a_76980_8230# a_76559_8230# a_76151_8309# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4711 a_31172_n4289# a_31429_n4479# a_30124_n4285# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4712 a_66067_11277# a_65854_11277# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4713 a_33688_n13399# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4714 a_18899_13694# a_19996_13500# a_19951_13513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4715 a_16346_8193# a_17459_11215# a_17414_11228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4716 a_65446_10706# a_65446_10165# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4717 a_52376_10552# a_52372_10729# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4718 a_54886_6106# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4719 vdd a_20205_10533# a_19997_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4720 a_68649_n11876# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4721 gnd d1 a_84219_n10489# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4722 vdd d0 a_31428_n12775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4723 a_55148_n3743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4724 a_65443_6218# a_66064_6110# a_66272_6110# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4725 a_1467_6791# a_1046_6791# a_638_6475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4726 a_44653_n5863# a_44440_n5863# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4727 gnd d1 a_51578_6055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4728 a_76414_n7028# a_77035_n6712# a_77243_n6712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4729 a_56355_8228# a_55934_8228# a_55307_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4730 a_36137_13554# a_35924_13554# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4731 a_30915_4542# a_31168_4529# a_29863_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4732 a_23194_n3739# a_22981_n3739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4733 a_5125_n8839# a_4912_n8839# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4734 vdd d2 a_7259_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4735 a_641_10708# a_641_10167# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4736 gnd d0 a_20462_n10491# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4737 a_2357_n8155# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4738 a_13018_11269# a_12805_11269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4739 a_55309_12114# a_56149_12789# a_56357_12789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4740 a_34108_n9753# a_34948_n9757# a_35156_n9757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4741 a_12229_n5869# a_12016_n5869# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4742 a_85016_n5240# a_85012_n5063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4743 vdd a_19154_7496# a_18946_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4744 a_22982_n8153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4745 gnd d5 a_81319_n5934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4746 a_44391_6791# a_44178_6791# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4747 a_19161_n11921# a_20254_n11259# a_20205_n11069# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4748 a_12228_n14844# a_12015_n14844# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4749 a_55362_n7389# a_55149_n7389# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4750 a_80510_5265# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4751 a_52632_n7254# a_52636_n8199# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4752 a_23402_n4418# a_24242_n3743# a_24450_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4753 a_67114_14240# a_66901_14240# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4754 gnd d0 a_20203_3078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4755 a_76153_12220# a_76154_11606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4756 gnd d1 a_62289_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4757 vdd d3 a_39598_n12778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4758 a_35156_n11204# a_34735_n11204# a_34108_n11200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4759 a_48451_5273# a_48342_5273# a_48550_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4760 a_33022_9508# a_33022_9253# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4761 a_52630_n12583# a_52887_n12773# a_51586_n13435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4762 a_8191_13700# a_9288_13506# a_9243_13519# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4763 a_9239_12249# a_9244_11231# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4764 a_83968_n4468# a_85061_n3806# a_76413_n3410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4765 a_23983_9826# a_23770_9826# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4766 gnd a_74559_n11255# a_74351_n11255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4767 a_45486_n11196# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4768 gnd a_63595_n14905# a_63387_n14905# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4769 a_60845_n8023# a_62341_n8893# a_62292_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4770 a_65444_4698# a_66065_4590# a_66273_4590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4771 a_35158_n5196# a_36397_n4429# a_36554_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4772 a_22720_3822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4773 gnd a_52628_12738# a_52420_12738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4774 vdd a_8449_10543# a_8241_10543# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4775 a_2515_6787# a_3754_7554# a_3911_6228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4776 a_44032_n5500# a_44032_n5755# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4777 a_33690_n7391# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4778 a_43041_941# a_42828_941# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4779 a_13226_9822# a_12805_9822# a_12178_9147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4780 a_60842_n11064# a_62338_n11934# a_62293_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4781 a_79780_n5874# a_79359_n5874# a_79681_n5874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4782 vdd d0 a_41878_9763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4783 a_40573_9278# a_41670_9084# a_41625_9097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4784 a_77241_n12720# a_76820_n12720# a_76412_n12641# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4785 a_56356_5261# a_57595_4581# a_57746_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4786 a_4015_n13396# a_3802_n13396# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4787 a_74302_n10297# a_74559_n10487# a_73254_n10293# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4788 a_37700_5265# a_38064_8178# a_38015_8368# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4789 a_38279_n9792# a_39392_n6770# a_39347_n6757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4790 a_8193_6068# a_8446_6055# a_6742_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4791 a_33851_9145# a_33430_9145# a_33022_9253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4792 a_31175_n14888# a_31171_n14711# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4793 a_44030_n9666# a_44651_n9745# a_44859_n9745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4794 a_27321_n5915# a_27271_n5928# a_27006_n8841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4795 a_55935_3814# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4796 a_60582_6919# a_62078_6049# a_62033_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4797 a_30913_11406# a_31170_11216# a_29869_10554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4798 a_75371_n15022# a_77033_n14846# a_77241_n14846# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4799 a_33640_6783# a_33427_6783# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4800 a_17451_3952# a_17708_3762# a_17408_5397# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4801 a_60802_n6578# a_60894_n8213# a_60849_n8200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4802 a_74049_10550# a_74302_10537# a_72997_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4803 a_44862_n6704# a_44441_n6704# a_44033_n7020# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4804 a_76153_13922# a_76774_14238# a_76982_14238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4805 vdd d1 a_73251_7500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4806 a_73259_n14884# a_74352_n14222# a_74307_n14209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4807 a_19161_n10474# a_20254_n9812# a_20205_n9622# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4808 a_76414_n7028# a_76414_n7283# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4809 gnd d0 a_63336_12732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4810 a_54481_10957# a_54481_10702# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4811 vdd d0 a_63335_3078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4812 a_49879_3781# a_50132_3768# a_49832_5403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4813 gnd a_8706_n10481# a_8498_n10481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4814 a_45648_5267# a_45227_5267# a_44600_4592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4815 a_14723_n13402# a_14510_n13402# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4816 vdd a_6959_11221# a_6751_11221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4817 vdd a_74300_5208# a_74092_5208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4818 a_55101_14240# a_54888_14240# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4819 a_76561_12791# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4820 a_30913_9959# a_30917_9103# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4821 a_1046_8238# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4822 a_85015_n14894# a_85011_n14717# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4823 vdd d0 a_52626_7498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4824 a_40570_7684# a_41667_7490# a_41622_7503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4825 a_22719_7557# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4826 gnd a_20464_n5930# a_20256_n5930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4827 a_40575_4540# a_40828_4527# a_39128_3773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4828 gnd d3 a_61057_n12776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4829 a_83709_10548# a_83962_10535# a_82262_9781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4830 gnd d2 a_17968_n14221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4831 a_12015_n13397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4832 a_31173_n8024# a_31177_n8880# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4833 a_47189_n11874# a_46976_n11874# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4834 vdd a_63595_n14226# a_63387_n14226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4835 a_1470_11279# a_2310_11275# a_2518_11275# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4836 a_51586_n13435# a_51839_n13448# a_50139_n14202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4837 a_640_14325# a_640_13930# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4838 a_83702_6237# a_84799_6043# a_84750_6233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4839 gnd d0 a_74299_8175# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4840 a_33021_13922# a_33021_13667# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4841 a_44438_n11871# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4842 gnd d0 a_74562_n8214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4843 gnd a_9757_n7444# a_9549_n7444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4844 a_23768_3818# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4845 gnd d0 a_31429_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4846 a_65854_9830# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4847 a_54481_9255# a_54478_8567# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4848 vdd a_42136_n12781# a_41928_n12781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4849 a_20210_n14213# a_20206_n14036# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4850 a_76982_13559# a_77822_14234# a_78030_14234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4851 a_67323_11273# a_68562_10593# a_68713_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4852 vdd d2 a_39641_n14223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4853 vdd d1 a_51578_6055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4854 a_52373_6064# a_52626_6051# a_51321_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4855 a_84757_11223# a_84753_11400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4856 a_13015_8228# a_12802_8228# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4857 a_44441_n8830# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4858 a_66532_n11194# a_66111_n11194# a_65703_n11115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4859 vdd a_6151_n9797# a_5943_n9797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4860 a_39127_6740# a_39380_6727# a_39085_5218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4861 a_71808_n14027# a_73304_n14897# a_73259_n14884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4862 vdd d0 a_52628_13506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4863 a_11348_12872# a_11969_12793# a_12177_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4864 a_76152_3245# a_76773_3137# a_76981_3137# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4865 a_60584_12927# a_62080_12057# a_62031_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4866 a_62290_n14711# a_63387_n14905# a_63338_n14715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4867 a_23140_6789# a_23980_6785# a_24188_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4868 a_46889_10595# a_46676_10595# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4869 a_56149_14236# a_55936_14236# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4870 a_20208_n7260# a_20465_n7450# a_19160_n7256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4871 a_33280_n14483# a_33280_n14738# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4872 a_9242_3776# a_9495_3763# a_8194_3101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4873 a_24191_11273# a_23770_11273# a_23143_10598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4874 a_78030_12787# a_77609_12787# a_76982_12112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4875 a_33903_n8159# a_33690_n8159# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4876 vdd d1 a_30382_n7442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4877 a_82219_11226# a_82472_11213# a_81151_8191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4878 a_55146_n11877# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4879 a_34736_n12724# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4880 gnd d0 a_85270_n7452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4881 vdd d1 a_19417_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4882 a_54481_10957# a_55102_11273# a_55310_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4883 a_44441_n6704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4884 a_33902_n5871# a_33689_n5871# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4885 a_32431_984# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4886 gnd a_73513_n4475# a_73305_n4475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4887 a_66066_12118# a_65853_12118# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4888 vdd a_60841_12737# a_60633_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4889 a_2308_3820# a_2095_3820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4890 gnd a_20463_n14226# a_20255_n14226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4891 a_3802_n13396# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4892 vdd d4 a_81664_n9805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4893 a_84755_3768# a_84751_3945# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4894 a_30911_4719# a_30915_3774# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4895 a_12230_n6710# a_12017_n6710# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4896 a_900_n4849# a_900_n5105# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4897 a_47300_n5866# a_46936_n7388# a_45910_n8155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4898 a_900_n5755# a_1521_n5863# a_1729_n5863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4899 a_33848_8230# a_34688_8226# a_34896_8226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4900 a_16602_n9613# a_17717_n12776# a_17668_n12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4901 a_54739_n14481# a_54739_n14736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4902 a_30129_n8876# a_31222_n8214# a_31173_n8024# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4903 a_1467_8238# a_1046_8238# a_638_8317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4904 a_35159_n6716# a_34738_n6716# a_34111_n6712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4905 a_28677_n5052# a_28934_n5242# a_28639_n6751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4906 vdd a_20464_n5251# a_20256_n5251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4907 a_60544_5220# a_60631_6729# a_60586_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4908 a_65444_3506# a_65444_3251# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4909 a_41618_7680# a_41622_6735# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4910 a_11608_n4855# a_12229_n4422# a_12437_n4422# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4911 gnd a_83961_13502# a_83753_13502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4912 a_7006_n11235# a_8498_n10481# a_8449_n10291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4913 gnd a_85270_n6773# a_85062_n6773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4914 a_22980_n14161# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4915 a_20206_n13268# a_20463_n13458# a_19158_n13264# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4916 a_57854_n10435# a_57641_n10435# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4917 a_66065_3143# a_65852_3143# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4918 a_59389_n5742# a_59783_n9803# a_59734_n9613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4919 gnd a_9756_n3798# a_9548_n3798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4920 vdd d0 a_31429_n5247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4921 a_22933_3143# a_22720_3143# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4922 a_8189_6245# a_8446_6055# a_6742_6925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4923 a_43772_13675# a_44393_13567# a_44601_13567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4924 vdd a_83962_9088# a_83754_9088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4925 gnd d0 a_63595_n12779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4926 vdd a_40829_13502# a_40621_13502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4927 a_44391_8238# a_44178_8238# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4928 vdd d1 a_62547_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4929 a_66900_5265# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4930 gnd a_60797_5207# a_60589_5207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4931 a_22313_14323# a_22934_14244# a_23142_14244# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4932 vdd a_51838_n10481# a_51630_n10481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4933 gnd a_28630_5211# a_28422_5211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4934 gnd a_41878_9763# a_41670_9763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4935 a_62294_n14888# a_63387_n14226# a_63342_n14213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4936 a_12014_n11198# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4937 a_55100_3139# a_54887_3139# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4938 vdd d0 a_63336_12732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4939 a_52629_n10295# a_52633_n11240# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4940 a_58008_n5872# a_57899_n5872# a_58107_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4941 a_25214_7552# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4942 a_1309_n8151# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4943 a_24027_n11198# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4944 a_44030_n10316# a_44030_n10857# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4945 a_66064_6789# a_65851_6789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4946 a_76411_n10324# a_76411_n10865# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4947 a_19951_12066# a_19947_12243# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4948 a_52632_n8022# a_52889_n8212# a_51588_n8874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4949 a_33279_n9674# a_33900_n9753# a_34108_n9753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4950 a_84755_4536# a_85008_4523# a_83703_4717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4951 vdd a_72064_n11250# a_71856_n11250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4952 gnd d0 a_85269_n3806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4953 a_43770_7667# a_43770_7126# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4954 a_85017_n8886# a_85270_n8899# a_83965_n8705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4955 a_12176_3818# a_11755_3818# a_11347_3897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4956 gnd a_30382_n7442# a_30174_n7442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4957 a_60588_12750# a_60841_12737# a_60546_11228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4958 a_77820_8226# a_77607_8226# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4959 a_25584_6226# a_25470_6107# a_25678_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4960 a_19947_14369# a_20204_14179# a_18903_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4961 a_11346_8567# a_11970_9147# a_12178_9147# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4962 a_44438_n10424# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4963 a_56357_12789# a_57596_13556# a_57753_12230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4964 a_83705_10725# a_83962_10535# a_82262_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4965 a_77607_6779# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4966 a_19950_5217# a_19946_5394# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4967 a_56409_n5194# a_56196_n5194# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4968 vdd a_72067_n8209# a_71859_n8209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4969 a_66272_7557# a_67112_8232# a_67320_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4970 a_11346_7661# a_11967_7553# a_12175_7553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4971 a_83702_6237# a_84799_6043# a_84754_6056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4972 vdd d0 a_74299_8175# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4973 a_23142_14244# a_23982_14240# a_24190_14240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4974 a_44601_12799# a_45441_12795# a_45649_12795# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4975 a_65703_n9668# a_65703_n10063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4976 a_22311_6218# a_22312_5604# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4977 a_13226_11269# a_12805_11269# a_12178_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4978 a_52369_6241# a_52626_6051# a_51321_6245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4979 vdd d1 a_84219_n11936# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4980 vdd a_42137_n3806# a_41929_n3806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4981 a_74042_6918# a_74046_6062# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4982 a_65705_n4310# a_66326_n4418# a_66534_n4418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4983 vdd d2 a_82775_n8215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4984 a_46936_n7388# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4985 a_66535_n6706# a_67375_n6710# a_67583_n6710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4986 vdd d5 a_48938_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4987 a_15781_9138# a_15360_9138# a_14715_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4988 a_52374_5223# a_52370_5400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4989 a_55310_11273# a_56150_11269# a_56358_11269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4990 a_83963_n13266# a_85060_n13460# a_85015_n13447# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4991 a_8456_n8874# a_9549_n8212# a_9500_n8022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4992 gnd d8 a_43488_n1602# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4993 a_9238_3953# a_9495_3763# a_8194_3101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4994 a_76561_14238# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4995 gnd a_51578_6055# a_51370_6055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4996 a_71807_n11060# a_73303_n11930# a_73254_n11740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4997 a_62291_n4289# a_62548_n4479# a_60848_n5233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4998 a_82215_11403# a_82472_11213# a_81151_8191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X4999 vdd d0 a_52889_n6765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5000 a_22314_10961# a_22314_10706# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5001 a_41622_8182# a_41875_8169# a_40574_7507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5002 a_63081_8184# a_63077_8361# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5003 a_14251_13556# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5004 vdd d1 a_8447_3088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5005 gnd d1 a_62286_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5006 a_12437_n5190# a_13277_n5194# a_13485_n5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5007 a_55570_n7389# a_56410_n6714# a_56618_n6714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5008 a_8449_n11738# a_9546_n11932# a_9497_n11742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5009 a_74303_n12585# a_74560_n12775# a_73259_n13437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5010 a_85013_n8030# a_85270_n8220# a_83969_n8882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5011 a_12438_n8157# a_12017_n8157# a_11609_n8078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5012 a_640_13134# a_1261_13567# a_1469_13567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5013 a_54740_n4059# a_54740_n4314# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5014 a_79528_n13404# a_79315_n13404# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5015 a_13486_n6714# a_14725_n7394# a_14876_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5016 a_65706_n7022# a_65706_n7277# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5017 a_67323_9826# a_66902_9826# a_66275_9830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5018 vdd a_9755_n13452# a_9547_n13452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5019 gnd a_20203_3078# a_19995_3078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5020 a_68559_7552# a_68346_7552# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5021 vdd a_74560_n14901# a_74352_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5022 a_76983_10592# a_76562_10592# a_76154_10159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5023 a_1470_10600# a_1049_10600# a_641_10167# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5024 a_22312_3901# a_22312_3506# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5025 vdd a_74301_13504# a_74093_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5026 a_31174_n10474# a_31170_n10297# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5027 a_68560_4585# a_68347_4585# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5028 a_30914_6062# a_30910_6239# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5029 a_11348_13924# a_11969_14240# a_12177_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5030 a_23770_9826# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5031 a_77609_14234# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5032 a_76559_7551# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5033 a_44652_n14838# a_44439_n14838# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5034 a_36549_n5874# a_36185_n7396# a_35159_n8163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5035 a_25257_6107# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5036 a_44030_n9410# a_44654_n8830# a_44862_n8830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5037 a_54740_n4059# a_55361_n3743# a_55569_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5038 a_44178_6791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5039 a_65703_n11765# a_66324_n11873# a_66532_n11873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5040 a_33281_n5763# a_33282_n6377# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5041 a_25940_n5868# a_25519_n5868# a_25846_n5749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5042 a_29865_9284# a_30962_9090# a_30917_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5043 a_13485_n3747# a_13064_n3747# a_12437_n4422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5044 a_11756_12793# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5045 gnd d0 a_9494_7498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5046 a_41883_n14215# a_41879_n14038# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5047 a_78029_3812# a_77608_3812# a_76981_3816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5048 a_76151_8565# a_76775_9145# a_76983_9145# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5049 a_31176_n4466# a_31429_n4479# a_30124_n4285# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5050 vdd a_82730_n12778# a_82522_n12778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5051 a_1260_5271# a_1047_5271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5052 vdd a_28630_5211# a_28422_5211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5053 vdd a_41878_9763# a_41670_9763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5054 a_39123_6917# a_40619_6047# a_40574_6060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5055 a_82521_n5235# a_84013_n4481# a_83964_n4291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5056 a_54889_11273# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5057 a_73257_n8699# a_74354_n8893# a_74309_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5058 gnd d0 a_31428_n12775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5059 a_66112_n12714# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5060 vdd d1 a_51579_3088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5061 gnd d2 a_71805_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5062 vdd a_52626_8177# a_52418_8177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5063 a_13065_n6714# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5064 a_84751_4713# a_85008_4523# a_83703_4717# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5065 a_66274_12797# a_65853_12797# a_65445_12481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5066 a_81062_n5744# a_81456_n9805# a_81411_n9792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5067 a_33279_n9674# a_33279_n10069# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5068 gnd d1 a_19155_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5069 gnd d0 a_41878_9084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5070 a_23401_n14840# a_24241_n14165# a_24449_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5071 gnd d1 a_30379_n10483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5072 a_43773_10167# a_44394_10600# a_44602_10600# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5073 a_52369_6241# a_52374_5223# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5074 gnd d2 a_7259_n11248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5075 vdd a_63335_3078# a_63127_3078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5076 a_28415_6923# a_29911_6053# a_29862_6243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5077 vdd d0 a_9496_13506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5078 a_45647_6787# a_45226_6787# a_44599_6112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5079 a_67581_n12718# a_67160_n12718# a_66533_n13393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5080 a_9503_n5911# a_9499_n5734# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5081 gnd d0 a_63335_3757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5082 a_22934_12797# a_22721_12797# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5083 a_11609_n7281# a_11609_n7822# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5084 a_71809_n5052# a_73305_n5922# a_73260_n5909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5085 vdd a_74299_6728# a_74091_6728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5086 a_13063_n12722# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5087 gnd a_83960_4527# a_83752_4527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5088 a_23140_8236# a_22719_8236# a_22311_7920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5089 a_34950_n5196# a_34737_n5196# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5090 a_54887_3139# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5091 a_12016_n4422# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5092 vdd a_16514_n5932# a_16306_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5093 a_33900_n11200# a_33687_n11200# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5094 gnd d3 a_39598_n12778# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5095 a_1729_n5184# a_2569_n5188# a_2777_n5188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5096 a_65704_n13030# a_65704_n13285# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5097 a_66534_n5865# a_66113_n5865# a_65705_n5757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5098 a_33279_n10069# a_33279_n10324# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5099 a_25517_n11876# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5100 a_77032_n11879# a_76819_n11879# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5101 vdd d5 a_27479_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5102 a_66533_n13393# a_67373_n12718# a_67581_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5103 a_57855_n13402# a_57642_n13402# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5104 a_9501_n9793# a_9497_n9616# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5105 a_2778_n6708# a_4017_n7388# a_4168_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5106 a_14973_n11880# a_14552_n11880# a_14874_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5107 a_76414_n8080# a_77035_n8159# a_77243_n8159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5108 a_25430_10593# a_25217_10593# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5109 a_76983_9824# a_76562_9824# a_76154_9903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5110 vdd a_51578_6055# a_51370_6055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5111 a_12802_8228# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5112 a_60842_n11064# a_62338_n11934# a_62289_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5113 a_76414_n6377# a_77034_n5871# a_77242_n5871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5114 a_57686_n5872# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5115 gnd d3 a_71764_11219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5116 a_69717_n8841# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5117 a_78291_n8163# a_77870_n8163# a_77243_n8838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5118 a_76152_4151# a_76152_3895# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5119 gnd a_73512_n14897# a_73304_n14897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5120 a_74306_n10474# a_74559_n10487# a_73254_n10293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5121 a_33687_n9753# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5122 a_38279_n9792# a_39392_n6770# a_39343_n6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5123 a_79426_12228# a_79312_12109# a_79520_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5124 a_27321_n5915# a_27271_n5928# a_27222_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5125 a_56358_9822# a_55937_9822# a_55310_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5126 a_44653_n5184# a_44440_n5184# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5127 a_2307_8234# a_2094_8234# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5128 a_85016_n5919# a_85012_n5742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5129 a_71552_3779# a_73044_4533# a_72995_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5130 a_72997_10731# a_74094_10537# a_74049_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5131 a_84757_11223# a_85010_11210# a_83709_10548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5132 a_2516_5267# a_3755_4587# a_3906_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5133 vdd a_82773_n14223# a_82565_n14223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5134 a_50094_n6572# a_50351_n6762# a_49030_n9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5135 a_4173_n5747# a_3803_n4421# a_2777_n5188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5136 a_65703_n10859# a_66324_n10426# a_66532_n10426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5137 a_21274_n15026# a_23193_n14840# a_23401_n14840# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5138 a_6966_n6749# a_7053_n5240# a_7008_n5227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5139 a_2095_3820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5140 a_55310_11273# a_54889_11273# a_54481_10957# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5141 a_23769_14240# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5142 a_44439_n13391# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5143 a_12229_n5190# a_12016_n5190# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5144 a_76411_n10324# a_77032_n10432# a_77240_n10432# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5145 a_1308_n4416# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5146 gnd a_59731_8180# a_59523_8180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5147 a_2357_n6708# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5148 a_12228_n14165# a_12015_n14165# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5149 a_78083_n6716# a_77870_n6716# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5150 a_45699_n9749# a_45486_n9749# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5151 a_79056_13554# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5152 a_31172_n4289# a_31176_n5234# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5153 a_80586_9136# a_80723_5265# a_75885_984# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5154 a_33428_5263# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5155 a_74045_11406# a_74049_10550# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5156 a_85014_n9801# a_85010_n9624# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5157 a_82475_n6580# a_82567_n8215# a_82522_n8202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5158 a_33641_3816# a_33428_3816# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5159 a_638_8317# a_638_7922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5160 a_77868_n12724# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5161 a_20205_n11069# a_20209_n11925# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5162 gnd a_63595_n14226# a_63387_n14226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5163 a_63344_n7437# a_63340_n7260# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5164 a_47997_9144# a_47784_9144# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5165 a_65706_n6627# a_66327_n6706# a_66535_n6706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5166 gnd a_30122_10541# a_29914_10541# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5167 a_22720_3143# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5168 a_33850_13559# a_33429_13559# a_33021_13126# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5169 gnd a_52628_12059# a_52420_12059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5170 a_22312_3506# a_22933_3822# a_23141_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5171 gnd d0 a_63596_n3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5172 vdd d2 a_71805_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5173 a_65852_4590# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5174 a_43773_10708# a_43773_10167# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5175 a_63081_7505# a_63334_7492# a_62029_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5176 vdd d1 a_41088_n14903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5177 a_47038_6109# a_46674_4587# a_45648_5267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5178 a_72996_13698# a_73253_13508# a_71553_12754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5179 vdd d1 a_19155_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5180 vdd d0 a_41878_9084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5181 gnd a_17970_n8213# a_17762_n8213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5182 a_12175_8232# a_11754_8232# a_11346_7916# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5183 a_80378_9136# a_80165_9136# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5184 a_28415_6923# a_29911_6053# a_29866_6066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5185 a_56616_n12722# a_56195_n12722# a_55568_n13397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5186 a_20212_n7437# a_20465_n7450# a_19160_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5187 a_67320_8232# a_68559_7552# a_68716_6226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5188 a_14512_n7394# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5189 a_76412_n14483# a_77033_n14167# a_77241_n14167# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5190 a_21532_n1444# a_21789_n1634# a_21631_n1621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5191 a_82215_11403# a_82307_9768# a_82262_9781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5192 a_65443_7124# a_66064_7557# a_66272_7557# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5193 vdd d0 a_9754_n10485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5194 a_33640_6104# a_33427_6104# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5195 a_36292_6220# a_35922_7546# a_34896_8226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5196 a_81062_n5744# a_81319_n5934# a_75301_n1457# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5197 a_66899_6785# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5198 a_14879_n11761# a_14509_n10435# a_13483_n11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5199 gnd d1 a_19417_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5200 a_25586_12234# a_25216_13560# a_24190_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5201 vdd d1 a_19156_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5202 gnd a_52889_n8891# a_52681_n8891# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5203 a_11756_14240# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5204 gnd d0 a_63336_12053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5205 a_44032_n4308# a_44653_n4416# a_44861_n4416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5206 a_56355_6781# a_57594_7548# a_57751_6222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5207 a_1049_9832# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5208 a_60585_9960# a_62081_9090# a_62032_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5209 a_51587_n4460# a_52680_n3798# a_44032_n3402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5210 a_48129_5273# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5211 gnd d0 a_31167_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5212 a_57642_n13402# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5213 vdd d2 a_50392_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5214 gnd d1 a_62288_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5215 a_57748_12111# a_57384_10589# a_56358_9822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5216 a_65705_n4055# a_65705_n4310# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5217 a_66275_10598# a_67115_11273# a_67323_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5218 a_54481_9905# a_54481_9510# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5219 a_12437_n3743# a_12016_n3743# a_11608_n4059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5220 a_57845_6103# a_58705_9138# a_58913_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5221 a_34108_n11200# a_33687_n11200# a_33279_n11121# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5222 a_20210_n13445# a_20463_n13458# a_19158_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5223 a_14294_12111# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5224 a_82519_n11243# a_84011_n10489# a_83966_n10476# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5225 a_45442_11275# a_45229_11275# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5226 a_22574_n7818# a_22574_n8074# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5227 a_54480_14319# a_55101_14240# a_55309_14240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5228 a_65446_9259# a_65443_8571# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5229 a_44438_n11192# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5230 a_3911_6228# a_3541_7554# a_2515_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5231 gnd a_62547_n14901# a_62339_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5232 gnd d0 a_31429_n5247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5233 a_9501_n9793# a_9754_n9806# a_8453_n10468# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5234 a_65854_9151# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5235 a_3906_6109# a_3797_6109# a_4005_6109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5236 a_23195_n8832# a_22982_n8832# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5237 a_13018_9822# a_12805_9822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5238 a_67583_n6710# a_68822_n7390# a_68973_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5239 a_71552_3779# a_73044_4533# a_72999_4546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5240 a_84753_11400# a_85010_11210# a_83709_10548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5241 a_11607_n13830# a_11607_n14086# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5242 vdd d0 a_9497_9092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5243 a_30123_n13260# a_30380_n13450# a_28680_n14204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5244 a_44440_n5863# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5245 a_5073_9144# a_4652_9144# a_4007_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5246 a_45907_n11196# a_45486_n11196# a_44859_n11871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5247 a_62294_n14888# a_63387_n14226# a_63338_n14036# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5248 a_77035_n8838# a_76822_n8838# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5249 vdd a_31430_n8893# a_31222_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5250 a_1049_11279# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5251 vdd a_8447_3088# a_8239_3088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5252 a_9242_3097# a_9495_3084# a_8190_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5253 a_54481_9510# a_55102_9826# a_55310_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5254 a_83965_n8705# a_84222_n8895# a_82518_n8025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5255 a_72996_13698# a_74093_13504# a_74044_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5256 a_78289_n14171# a_77868_n14171# a_77241_n14167# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5257 vdd a_8706_n10481# a_8498_n10481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5258 vdd a_59731_8180# a_59523_8180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5259 a_55146_n11198# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5260 gnd a_72064_n11250# a_71856_n11250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5261 a_33902_n5192# a_33689_n5192# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5262 a_43772_14325# a_43772_13930# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5263 a_18899_13694# a_19156_13504# a_17456_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5264 a_30913_9280# a_30914_8188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5265 a_52375_12072# a_52371_12249# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5266 vdd d2 a_17968_n14221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5267 a_3804_n7388# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5268 a_900_n5105# a_1521_n5184# a_1729_n5184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5269 a_85015_n12768# a_85011_n12591# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5270 a_64740_973# a_64527_973# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5271 a_33851_9824# a_34691_9820# a_34899_9820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5272 gnd a_85269_n5932# a_85061_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5273 a_44601_14246# a_44180_14246# a_43772_14325# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5274 vdd a_30122_10541# a_29914_10541# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5275 a_31172_n5736# a_31429_n5926# a_30124_n5732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5276 a_70443_8197# a_71556_11219# a_71507_11409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5277 a_74307_n14888# a_74303_n14711# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5278 vdd a_19414_n10487# a_19206_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5279 a_72998_7513# a_74091_8175# a_74042_8365# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5280 a_33688_n14846# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5281 a_34948_n9757# a_34735_n9757# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5282 a_33430_11271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5283 gnd a_9494_7498# a_9286_7498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5284 gnd d1 a_84219_n11936# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5285 a_640_12228# a_641_11614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5286 a_44033_n7816# a_44033_n8072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5287 a_32169_n1457# a_37979_n5934# a_37714_n8847# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5288 gnd d2 a_82775_n8215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5289 gnd d5 a_48938_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5290 a_34110_n5871# a_33689_n5871# a_33282_n6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5291 a_1522_n7383# a_1309_n7383# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5292 a_22935_11277# a_22722_11277# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5293 a_65445_12481# a_66066_12797# a_66274_12797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5294 a_83963_n13266# a_85060_n13460# a_85011_n13270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5295 a_44394_9832# a_44181_9832# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5296 gnd a_71805_3766# a_71597_3766# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5297 a_19951_12745# a_19947_12922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5298 gnd a_62286_7496# a_62078_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5299 vdd a_39380_6727# a_39172_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5300 gnd d1 a_51840_n4473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5301 a_1729_n3737# a_1308_n3737# a_900_n4053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5302 a_66273_5269# a_67113_5265# a_67321_5265# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5303 a_1309_n8830# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5304 a_62295_n4466# a_62548_n4479# a_60848_n5233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5305 gnd d0 a_52889_n6765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5306 a_9502_n14207# a_9498_n14030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5307 a_71813_n5229# a_72066_n5242# a_71771_n6751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5308 gnd a_19155_3082# a_18947_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5309 gnd a_41878_9084# a_41670_9084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5310 a_44393_12799# a_44180_12799# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5311 a_52629_n9616# a_52633_n10472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5312 vdd d0 a_85270_n7452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5313 a_3756_13562# a_3543_13562# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5314 a_30123_n13260# a_31220_n13454# a_31175_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5315 vdd d0 a_63336_12053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5316 a_54481_11608# a_54481_11352# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5317 a_74049_10550# a_74045_10727# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5318 a_55362_n8836# a_55149_n8836# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5319 a_62291_n4289# a_63388_n4483# a_63339_n4293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5320 a_42828_941# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5321 a_51327_12076# a_51580_12063# a_49876_12933# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5322 a_44181_10600# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5323 gnd a_63335_3757# a_63127_3757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5324 a_45649_14242# a_45228_14242# a_44601_14246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5325 a_55307_6106# a_56147_6781# a_56355_6781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5326 a_65704_n13826# a_66325_n13393# a_66533_n13393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5327 gnd d0 a_20203_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5328 vdd a_31170_10537# a_30962_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5329 a_66064_6110# a_65851_6110# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5330 a_22572_n14477# a_22572_n14732# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5331 a_13225_14236# a_12804_14236# a_12177_13561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5332 a_22721_13565# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5333 a_74307_n12762# a_74560_n12775# a_73259_n13437# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5334 a_85017_n8207# a_85270_n8220# a_83969_n8882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5335 a_12176_3139# a_11755_3139# a_11347_3247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5336 a_77823_9820# a_77610_9820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5337 a_1309_n6704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5338 a_74304_n4289# a_74561_n4479# a_73256_n4285# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5339 a_63340_n6581# a_63344_n7437# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5340 a_13483_n9755# a_14722_n10435# a_14879_n11761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5341 a_43770_6220# a_44391_6112# a_44599_6112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5342 a_74047_5221# a_74043_5398# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5343 a_19952_11225# a_20205_11212# a_18904_10550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5344 a_63342_n14213# a_63338_n14036# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5345 a_55362_n6710# a_55149_n6710# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5346 a_48465_n8839# a_48044_n8839# a_47399_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5347 a_34896_8226# a_34475_8226# a_33848_7551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5348 a_33281_n4316# a_33902_n4424# a_34110_n4424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5349 vdd a_85270_n6773# a_85062_n6773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5350 a_34111_n6712# a_34951_n6716# a_35159_n6716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5351 vdd d0 a_74302_9769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5352 a_7006_n11235# a_8498_n10481# a_8453_n10468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5353 a_55309_13561# a_54888_13561# a_54480_13669# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5354 a_55567_n9751# a_55146_n9751# a_54738_n9672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5355 a_44031_n14475# a_44031_n14730# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5356 a_76412_n14483# a_76412_n14738# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5357 a_2516_5267# a_2095_5267# a_1468_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5358 a_74302_n11744# a_74559_n11934# a_73254_n11740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5359 a_62293_n10474# a_63386_n9812# a_63341_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5360 a_49878_6748# a_51370_7502# a_51321_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5361 a_13275_n9755# a_13062_n9755# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5362 a_54480_12477# a_54480_12222# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5363 gnd a_82730_n12778# a_82522_n12778# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5364 gnd a_39641_n14223# a_39433_n14223# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5365 vdd d2 a_39642_n5248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5366 vdd d3 a_17665_5207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5367 a_33280_n12641# a_33901_n12720# a_34109_n12720# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5368 a_1521_n3737# a_1308_n3737# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5369 a_83705_9278# a_83962_9088# a_82258_9958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5370 a_76411_n9418# a_76411_n9674# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5371 a_44651_n10424# a_44438_n10424# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5372 a_66534_n4418# a_67374_n3743# a_67582_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5373 a_9238_3274# a_9495_3084# a_8190_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5374 a_17452_12927# a_18948_12057# a_18903_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5375 a_2094_8234# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5376 gnd d2 a_82514_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5377 a_43771_4700# a_44392_4592# a_44600_4592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5378 a_45440_5267# a_45227_5267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5379 a_54741_n8078# a_54741_n8473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5380 a_44179_3824# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5381 a_41625_9776# a_41878_9763# a_40577_9101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5382 vdd d0 a_20463_n13458# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5383 a_79778_n11882# a_80638_n8847# a_80846_n8847# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5384 a_14724_n4427# a_14511_n4427# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5385 vdd a_30382_n7442# a_30174_n7442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5386 vdd a_85267_n10493# a_85059_n10493# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5387 a_66111_n9747# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5388 a_65705_n3660# a_65705_n4055# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5389 a_77033_n13399# a_76820_n13399# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5390 a_30911_5398# a_30915_4542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5391 a_66902_11273# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5392 a_30914_6741# a_30910_6918# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5393 a_900_n5500# a_900_n5755# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5394 a_58913_9138# a_59050_5267# a_54212_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5395 a_82255_6917# a_82512_6727# a_82217_5218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5396 a_62033_7509# a_63126_8171# a_63077_8361# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5397 a_11968_3818# a_11755_3818# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5398 a_8453_n11915# a_9546_n11253# a_9497_n11063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5399 a_67113_3818# a_66900_3818# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5400 a_33427_6783# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5401 a_12015_n14844# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5402 a_34110_n4424# a_33689_n4424# a_33281_n4316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5403 a_47397_n11874# a_46976_n11874# a_47298_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5404 a_51586_n14882# a_51839_n14895# a_50135_n14025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5405 a_72998_7513# a_74091_8175# a_74046_8188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5406 a_11608_n4855# a_11608_n5111# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5407 a_54888_14240# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5408 gnd a_9757_n8891# a_9549_n8891# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5409 a_24449_n12718# a_25688_n13398# a_25839_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5410 a_24240_n11198# a_24027_n11198# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5411 a_33022_9253# a_33019_8565# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5412 a_66272_8236# a_65851_8236# a_65443_8315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5413 gnd d0 a_85007_7490# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5414 a_23143_9151# a_23983_9826# a_24191_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5415 vdd d1 a_51578_7502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5416 a_1727_n11871# a_2567_n11196# a_2775_n11196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5417 a_11347_4949# a_11968_5265# a_12176_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5418 a_44652_n14159# a_44439_n14159# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5419 a_33022_11350# a_33022_10955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5420 a_47784_9144# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5421 a_44033_n8467# a_44654_n8151# a_44862_n8151# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5422 gnd d5 a_27479_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5423 a_33429_12791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5424 a_68609_n7390# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5425 a_65703_n11115# a_66324_n11194# a_66532_n11194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5426 a_44178_6112# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5427 gnd a_17667_11215# a_17459_11215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5428 vdd d0 a_74302_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5429 vdd a_71805_3766# a_71597_3766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5430 a_74042_6239# a_74047_5221# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5431 a_56197_n8161# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5432 a_44032_n4308# a_44032_n4849# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5433 a_55149_n7389# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5434 gnd d0 a_31169_14183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5435 a_52374_3097# a_52370_3274# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5436 vdd a_19155_3082# a_18947_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5437 vdd a_41878_9084# a_41670_9084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5438 a_33020_3500# a_33641_3816# a_33849_3816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5439 a_80165_9136# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5440 a_35157_n12724# a_34736_n12724# a_34109_n13399# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5441 gnd d1 a_30120_3086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5442 a_51323_12253# a_51580_12063# a_49876_12933# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5443 a_12435_n11877# a_13275_n11202# a_13483_n11202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5444 gnd a_73513_n5922# a_73305_n5922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5445 a_57857_n7394# a_57644_n7394# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5446 vdd d0 a_20203_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5447 a_47045_12236# a_46675_13562# a_45649_12795# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5448 a_66327_n7385# a_66114_n7385# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5449 a_60582_6919# a_62078_6049# a_62029_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5450 a_2567_n9749# a_2354_n9749# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5451 vdd d1 a_8709_n7440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5452 a_63081_6058# a_63077_6235# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5453 a_8449_n11738# a_9546_n11932# a_9501_n11919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5454 vdd a_71764_11219# a_71556_11219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5455 a_83963_n14713# a_84220_n14903# a_82516_n14033# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5456 a_76982_12791# a_77822_12787# a_78030_12787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5457 gnd d1 a_40829_13502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5458 a_6966_n6749# a_7053_n5240# a_7004_n5050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5459 a_19948_11402# a_20205_11212# a_18904_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5460 a_33900_n11879# a_33687_n11879# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5461 a_899_n13824# a_899_n14080# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5462 gnd d0 a_63335_3078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5463 gnd a_31169_13504# a_30961_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5464 a_22934_12118# a_22721_12118# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5465 vdd a_74299_6049# a_74091_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5466 a_56358_9822# a_57597_10589# a_57748_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5467 a_23143_9830# a_22722_9830# a_22314_9514# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5468 a_56149_12789# a_55936_12789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5469 a_68606_n10431# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5470 gnd a_31167_7496# a_30959_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5471 a_36183_n13404# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5472 vdd d0 a_52886_n10485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5473 a_36386_6101# a_37246_9136# a_37454_9136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5474 a_82475_n6580# a_82567_n8215# a_82518_n8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5475 a_28675_n11060# a_28932_n11250# a_28637_n12759# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5476 vdd d1 a_8707_n13448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5477 a_31171_n14711# a_32239_n15022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5478 a_43773_9911# a_44394_9832# a_44602_9832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5479 a_8189_7692# a_8446_7502# a_6746_6748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5480 a_66534_n5186# a_66113_n5186# a_65705_n5107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5481 a_8189_7692# a_9286_7498# a_9237_7688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5482 a_76820_n13399# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5483 a_65853_12797# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5484 gnd a_7219_n6762# a_7011_n6762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5485 a_24242_n5190# a_24029_n5190# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5486 a_77032_n11200# a_76819_n11200# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5487 vdd d0 a_74560_n12775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5488 a_33281_n3666# a_33281_n4061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5489 vdd a_51838_n11928# a_51630_n11928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5490 a_37714_n8847# a_37293_n8847# a_36648_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5491 a_50140_n5227# a_51632_n4473# a_51583_n4283# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5492 a_899_n12377# a_1519_n11871# a_1727_n11871# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5493 a_55099_7553# a_54886_7553# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5494 a_638_6475# a_1259_6791# a_1467_6791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5495 a_22574_n7277# a_23195_n7385# a_23403_n7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5496 a_76773_3816# a_76560_3816# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5497 a_33021_13667# a_33021_13126# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5498 a_82521_n5235# a_84013_n4481# a_83968_n4468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5499 a_12805_9822# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5500 a_76983_9145# a_76562_9145# a_76154_9253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5501 a_55100_4586# a_54887_4586# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5502 a_76413_n5508# a_77034_n5192# a_77242_n5192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5503 vdd d2 a_82514_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5504 a_11347_3502# a_11347_3247# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5505 a_41621_9953# a_41878_9763# a_40577_9101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5506 vdd a_9497_9092# a_9289_9092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5507 gnd a_43488_n1602# a_43280_n1602# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5508 a_22314_11612# a_22314_11356# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5509 a_29867_4546# a_30960_5208# a_30915_5221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5510 a_48770_8199# a_49023_8186# a_48451_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5511 a_33279_n10865# a_33900_n10432# a_34108_n10432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5512 a_76980_7551# a_76559_7551# a_76151_7118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5513 vdd d1 a_30379_n10483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5514 a_9498_n13262# a_9502_n14207# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5515 a_78291_n6716# a_77870_n6716# a_77243_n6712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5516 a_62296_n7433# a_63389_n6771# a_63340_n6581# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5517 a_10595_n1632# a_21789_n1634# a_21631_n1621# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5518 a_14252_10589# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5519 a_66326_n3739# a_66113_n3739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5520 a_62033_7509# a_63126_8171# a_63081_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5521 a_74306_n10474# a_74302_n10297# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5522 gnd d0 a_9754_n10485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5523 a_33280_n13291# a_33280_n13832# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5524 a_80846_n8847# a_81319_n5934# a_75301_n1457# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5525 a_76774_12791# a_76561_12791# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5526 a_56147_6781# a_55934_6781# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5527 vdd d3 a_82730_n12778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5528 vdd a_62289_9090# a_62081_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5529 gnd a_70696_8184# a_70488_8184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5530 a_77240_n10432# a_78080_n9757# a_78288_n9757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5531 a_33689_n4424# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5532 vdd a_62549_n8893# a_62341_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5533 a_74305_n6577# a_74562_n6767# a_73261_n7429# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5534 vdd a_75558_n1647# a_75350_n1647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5535 a_641_10167# a_1262_10600# a_1470_10600# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5536 a_900_n3402# a_9499_n3608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5537 a_83702_7684# a_84799_7490# a_84754_7503# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5538 a_22572_n14477# a_23193_n14161# a_23401_n14161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5539 a_54741_n6375# a_54741_n6631# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5540 a_23143_11277# a_22722_11277# a_22314_11356# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5541 a_73255_n13260# a_73512_n13450# a_71812_n14204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5542 gnd a_60841_12737# a_60633_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5543 a_66533_n12714# a_66112_n12714# a_65704_n13030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5544 a_84751_3945# a_84755_3089# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5545 a_22932_8236# a_22719_8236# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5546 gnd d0 a_41876_5202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5547 a_63340_n8707# a_63597_n8897# a_62292_n8703# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5548 vdd a_16859_n9803# a_16651_n9803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5549 a_52369_7688# a_52626_7498# a_51321_7692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5550 a_33282_n6633# a_33903_n6712# a_34111_n6712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5551 a_24450_n5190# a_25689_n4423# a_25846_n5749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5552 gnd d2 a_50392_n14215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5553 a_65446_11356# a_66067_11277# a_66275_11277# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5554 vdd d1 a_73514_n8889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5555 a_76414_n8475# a_76414_n8730# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5556 vdd a_17667_11215# a_17459_11215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5557 a_18901_7509# a_19154_7496# a_17454_6742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5558 a_54739_n13289# a_54739_n13830# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5559 a_22313_12481# a_22313_12226# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5560 a_33641_3137# a_33428_3137# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5561 vdd d0 a_52629_11218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5562 a_12228_n12718# a_12015_n12718# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5563 a_36287_6101# a_35923_4579# a_34897_3812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5564 a_60588_12750# a_62080_13504# a_62035_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5565 vdd a_60839_6729# a_60631_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5566 a_12227_n9751# a_12014_n9751# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5567 vdd d0 a_63597_n7450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5568 a_60544_5220# a_60631_6729# a_60582_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5569 vdd d4 a_27824_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5570 vdd d0 a_31169_14183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5571 a_44394_11279# a_44181_11279# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5572 a_13484_n12722# a_13063_n12722# a_12436_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5573 a_82519_n11243# a_84011_n10489# a_83962_n10299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5574 a_79359_n5874# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5575 a_63339_n5740# a_63344_n6758# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5576 a_45910_n8155# a_45489_n8155# a_44862_n8830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5577 a_62291_n5736# a_62548_n5926# a_60844_n5056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5578 vdd d2 a_7000_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5579 a_22571_n10063# a_22571_n10318# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5580 a_22573_n3660# a_23194_n3739# a_23402_n3739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5581 a_22314_3152# a_22933_3143# a_23141_3143# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5582 a_4265_n11874# a_5125_n8839# a_5333_n8839# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5583 vdd d1 a_30120_3086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5584 gnd d0 a_74301_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5585 a_44181_9832# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5586 a_66272_6789# a_67112_6785# a_67320_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5587 a_44652_n13391# a_44439_n13391# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5588 a_33427_8230# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5589 gnd a_52887_n14899# a_52679_n14899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5590 a_30915_4542# a_30911_4719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5591 a_11608_n5761# a_12229_n5869# a_12437_n5869# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5592 a_6964_n12757# a_7051_n11248# a_7006_n11235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5593 a_34737_n3749# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5594 a_50094_n6572# a_50186_n8207# a_50141_n8194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5595 a_19157_n10297# a_20254_n10491# a_20205_n10301# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5596 a_25938_n11876# a_25517_n11876# a_25844_n11757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5597 a_71507_11409# a_71599_9774# a_71550_9964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5598 a_30127_n13437# a_30380_n13450# a_28680_n14204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5599 a_4166_n11874# a_4057_n11874# a_4265_n11874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5600 a_33281_n3410# a_41880_n3616# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5601 a_66274_14244# a_67114_14240# a_67322_14240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5602 vdd d0 a_31427_n9808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5603 a_44180_13567# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5604 a_84752_12920# a_84756_12064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5605 a_34690_14234# a_34477_14234# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5606 a_19163_n4466# a_20256_n3804# a_11608_n3408# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5607 gnd a_20203_4525# a_19995_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5608 a_44030_n10061# a_44030_n10316# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5609 a_41622_7503# a_41618_7680# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5610 a_76411_n10069# a_76411_n10324# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5611 a_45702_n6708# a_45489_n6708# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5612 a_3906_6109# a_3542_4587# a_2516_3820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5613 a_77610_9820# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5614 a_45441_14242# a_45228_14242# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5615 gnd a_52889_n8212# a_52681_n8212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5616 a_76980_8230# a_77820_8226# a_78028_8226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5617 a_79097_6101# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5618 a_33022_10955# a_33022_10700# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5619 a_55360_n13397# a_55147_n13397# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5620 a_43770_6475# a_43770_6220# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5621 gnd d0 a_42138_n8899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5622 a_17710_n11064# a_17967_n11254# a_17672_n12763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5623 a_19951_14192# a_20204_14179# a_18903_13517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5624 a_44860_n14838# a_44439_n14838# a_42947_n15028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5625 vdd a_62289_10537# a_62081_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5626 gnd d0 a_9495_5210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5627 a_1049_9153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5628 a_14874_n11880# a_14765_n11880# a_14973_n11880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5629 a_14975_n5872# a_14554_n5872# a_14876_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5630 vdd d2 a_7262_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5631 a_11970_11273# a_11757_11273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5632 vdd a_74302_9769# a_74094_9769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5633 a_34108_n11879# a_33687_n11879# a_33279_n11771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5634 a_27006_n8841# a_26585_n8841# a_25938_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5635 a_65446_9909# a_65446_9514# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5636 a_31176_n5913# a_31429_n5926# a_30124_n5732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5637 a_638_6220# a_639_5606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5638 a_29868_13521# a_30961_14183# a_30912_14373# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5639 gnd a_19414_n10487# a_19206_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5640 a_45907_n11196# a_47146_n10429# a_47303_n11755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5641 a_55101_13561# a_54888_13561# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5642 a_1048_14246# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5643 a_24028_n12718# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5644 a_44860_n12712# a_44439_n12712# a_44031_n12633# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5645 a_38279_n9792# a_38532_n9805# a_37930_n5744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5646 a_54479_4153# a_54479_3897# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5647 a_25841_n5868# a_25732_n5868# a_25940_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5648 a_56617_n5194# a_57856_n4427# a_58013_n5753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5649 a_74044_12247# a_74301_12057# a_72996_12251# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5650 a_32169_n1457# a_37979_n5934# a_37930_n5744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5651 gnd d0 a_74302_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5652 a_51586_n13435# a_52679_n12773# a_52630_n12583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5653 a_48766_8376# a_49023_8186# a_48451_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5654 a_76152_3895# a_76152_3500# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5655 a_7009_n8194# a_8501_n7440# a_8456_n7427# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5656 gnd a_20462_n9812# a_20254_n9812# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5657 a_23195_n8153# a_22982_n8153# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5658 a_39389_n5235# a_40881_n4481# a_40832_n4291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5659 a_77609_12787# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5660 a_78081_n12724# a_77868_n12724# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5661 a_46887_4587# a_46674_4587# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5662 a_23981_5265# a_23768_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5663 a_40837_n7435# a_41930_n6773# a_41881_n6583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5664 a_39129_12748# a_40621_13502# a_40572_13692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5665 vdd a_52887_n14220# a_52679_n14220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5666 a_68346_7552# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5667 a_45487_n14163# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5668 a_50138_n11235# a_51630_n10481# a_51581_n10291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5669 a_1519_n9745# a_1306_n9745# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5670 a_77240_n11200# a_78080_n11204# a_78288_n11204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5671 a_75776_984# a_75563_984# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5672 a_11967_8232# a_11754_8232# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5673 a_44440_n5184# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5674 a_67112_8232# a_66899_8232# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5675 a_66532_n9747# a_67372_n9751# a_67580_n9751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5676 vdd a_70696_8184# a_70488_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5677 a_77035_n8159# a_76822_n8159# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5678 a_55308_3818# a_54887_3818# a_54479_3897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5679 a_30123_n13260# a_31220_n13454# a_31171_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5680 a_8450_n14705# a_9547_n14899# a_9502_n14886# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5681 a_13224_5261# a_12803_5261# a_12176_4586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5682 a_68716_6226# a_68602_6107# a_68810_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5683 a_79267_7546# a_79054_7546# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5684 a_52375_12751# a_52371_12928# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5685 a_1262_11279# a_1049_11279# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5686 a_62290_n13264# a_62547_n13454# a_60847_n14208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5687 a_15620_n8845# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5688 a_54478_8567# a_55102_9147# a_55310_9147# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5689 a_11755_3818# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5690 a_63337_n11069# a_63341_n11925# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5691 a_74308_n4466# a_74561_n4479# a_73256_n4285# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5692 a_55309_12114# a_54888_12114# a_54481_11608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5693 a_69878_9142# a_69457_9142# a_68810_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5694 a_41625_9097# a_41621_9274# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5695 vdd d0 a_42138_n8220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5696 a_54478_7661# a_55099_7553# a_55307_7553# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5697 a_35158_n5196# a_34737_n5196# a_34110_n5192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5698 a_31173_n6577# a_31177_n7433# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5699 a_37246_9136# a_37033_9136# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5700 a_22982_n7385# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5701 gnd a_85007_7490# a_84799_7490# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5702 a_5319_5273# a_5210_5273# a_5418_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5703 gnd a_85269_n5253# a_85061_n5253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5704 vdd a_51578_7502# a_51370_7502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5705 a_31172_n5057# a_31429_n5247# a_30128_n5909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5706 a_40576_12068# a_40829_12055# a_39125_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5707 a_33019_8309# a_33640_8230# a_33848_8230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5708 a_55308_3818# a_56148_3814# a_56356_3814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5709 gnd a_20204_12732# a_19996_12732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5710 a_79679_n11882# a_79570_n11882# a_79778_n11882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5711 a_77243_n8838# a_76822_n8838# a_76411_n9418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5712 vdd a_31170_9090# a_30962_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5713 a_58913_9138# a_58492_9138# a_57847_12111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5714 vdd a_51839_n14895# a_51631_n14895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5715 a_21816_973# a_21395_973# a_11179_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5716 a_33688_n14167# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5717 a_74306_n11921# a_74559_n11934# a_73254_n11740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5718 vdd d1 a_62286_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5719 vdd d0 a_9757_n8891# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5720 a_71507_11409# a_71599_9774# a_71554_9787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5721 a_30914_8188# a_31167_8175# a_29866_7513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5722 gnd d2 a_39642_n5248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5723 a_4007_12117# a_3586_12117# a_3913_12236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5724 a_67372_n11198# a_67159_n11198# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5725 a_34110_n5192# a_33689_n5192# a_33281_n5508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5726 a_4005_6109# a_3584_6109# a_3911_6228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5727 a_8192_9286# a_9289_9092# a_9244_9105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5728 a_66113_n5865# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5729 a_39123_6917# a_40619_6047# a_40570_6237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5730 a_65446_11612# a_66066_12118# a_66274_12118# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5731 a_44394_9153# a_44181_9153# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5732 a_67580_n9751# a_67159_n9751# a_66532_n9747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5733 a_51584_n8697# a_51841_n8887# a_50137_n8017# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5734 a_77243_n6712# a_76822_n6712# a_76414_n6633# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5735 a_47146_n10429# a_46933_n10429# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5736 a_77867_n9757# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5737 vdd a_20203_4525# a_19995_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5738 a_76413_n3410# a_85269_n3806# a_83968_n4468# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5739 gnd d2 a_60842_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5740 a_41883_n12768# a_42136_n12781# a_40835_n13443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5741 a_41880_n4295# a_42137_n4485# a_40832_n4291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5742 gnd a_52626_8177# a_52418_8177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5743 a_83966_n10476# a_85059_n9814# a_85014_n9801# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5744 a_80846_n8847# a_80425_n8847# a_79778_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5745 a_4865_9144# a_4652_9144# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5746 gnd d0 a_20463_n13458# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5747 a_44393_12120# a_44180_12120# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5748 a_1308_n5863# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5749 a_76411_n10069# a_77032_n9753# a_77240_n9753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5750 a_55362_n8157# a_55149_n8157# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5751 a_70124_5271# a_70488_8184# a_70439_8374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5752 a_25476_n4423# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5753 a_65854_11277# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5754 gnd a_63335_3078# a_63127_3078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5755 vdd d0 a_9495_5210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5756 a_25472_12115# a_25259_12115# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5757 a_24449_n14165# a_24028_n14165# a_23401_n14840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5758 a_51328_10556# a_52421_11218# a_52376_11231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5759 a_43772_12228# a_43773_11614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5760 gnd a_74299_6728# a_74091_6728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5761 a_9504_n8199# a_9500_n8022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5762 vdd a_85269_n5932# a_85061_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5763 a_66902_9826# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5764 vdd a_31427_n10487# a_31219_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5765 a_27222_n5738# a_27616_n9799# a_27571_n9786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5766 a_29868_13521# a_30961_14183# a_30916_14196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5767 vdd d4 a_38272_8178# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5768 a_68389_6107# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5769 a_35924_13554# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5770 a_54741_n7822# a_55362_n7389# a_55570_n7389# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5771 a_76772_8230# a_76559_8230# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5772 gnd a_62288_13504# a_62080_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5773 a_11969_12793# a_11756_12793# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5774 a_34899_9820# a_34478_9820# a_33851_9145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5775 a_22981_n3739# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5776 a_4912_n8839# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5777 a_45909_n3741# a_47148_n4421# a_47305_n5747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5778 a_44031_n14730# a_44652_n14838# a_44860_n14838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5779 a_12016_n5869# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5780 a_1469_14246# a_1048_14246# a_640_14325# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5781 a_52631_n3608# a_52635_n4464# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5782 a_60843_n14031# a_62339_n14901# a_62294_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5783 a_76560_3816# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5784 vdd d1 a_19155_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5785 a_74302_n11065# a_74559_n11255# a_73258_n11917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5786 a_76775_11271# a_76562_11271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5787 gnd d0 a_20464_n3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5788 a_28419_6746# a_29911_7500# a_29866_7513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5789 a_18900_9280# a_19157_9090# a_17453_9960# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5790 a_20212_n8884# a_20465_n8897# a_19160_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5791 a_52632_n7254# a_52889_n7444# a_51584_n7250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5792 vdd d3 a_82470_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5793 a_66901_14240# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5794 a_33021_13667# a_33642_13559# a_33850_13559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5795 a_54741_n8728# a_54738_n9416# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5796 vdd d1 a_51840_n4473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5797 a_71809_n5052# a_72066_n5242# a_71771_n6751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5798 gnd d1 a_73253_12061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5799 a_44031_n13028# a_44652_n12712# a_44860_n12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5800 gnd d1 a_19417_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5801 a_55569_n4422# a_55148_n4422# a_54740_n4314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5802 a_71552_3779# a_71805_3766# a_71505_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5803 a_66273_5269# a_65852_5269# a_65444_4953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5804 a_66324_n11873# a_66111_n11873# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5805 gnd d0 a_52627_3763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5806 a_62291_n4289# a_63388_n4483# a_63343_n4470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5807 a_40575_3093# a_41668_3755# a_41619_3945# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5808 gnd d1 a_8709_n7440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5809 a_44179_3145# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5810 vdd d1 a_83959_6047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5811 a_41625_9097# a_41878_9084# a_40573_9278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5812 a_41885_n8207# a_41881_n8030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5813 a_55569_n5869# a_56409_n5194# a_56617_n5194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5814 a_72997_10731# a_74094_10537# a_74045_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5815 vdd a_9497_10539# a_9289_10539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5816 a_33022_9903# a_33022_9508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5817 a_77035_n7391# a_76822_n7391# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5818 a_11968_3139# a_11755_3139# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5819 gnd a_41876_5202# a_41668_5202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5820 a_40830_n10299# a_41927_n10493# a_41882_n10480# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5821 a_23141_4590# a_22720_4590# a_22312_4698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5822 a_12015_n14165# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5823 a_20210_n14892# a_20463_n14905# a_19158_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5824 a_82515_n11066# a_84011_n11936# a_83966_n11923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5825 gnd d0 a_52886_n10485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5826 a_25519_n5868# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5827 a_74047_3095# a_74043_3272# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5828 a_40572_12245# a_40829_12055# a_39125_12925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5829 a_73001_9107# a_74094_9769# a_74049_9782# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5830 vdd a_20204_12732# a_19996_12732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5831 a_76413_n3410# a_76413_n3666# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5832 a_43770_7126# a_44391_7559# a_44599_7559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5833 a_28679_n11237# a_28932_n11250# a_28637_n12759# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5834 a_55099_6106# a_54886_6106# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5835 a_24189_3818# a_23768_3818# a_23141_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5836 gnd d1 a_8707_n13448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5837 gnd a_9757_n8212# a_9549_n8212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5838 a_30916_13517# a_30912_13694# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5839 a_79681_n5874# a_79317_n7396# a_78291_n6716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5840 a_11349_11352# a_11349_10957# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5841 a_73261_n7429# a_73514_n7442# a_71814_n8196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5842 a_45908_n14163# a_47147_n13396# a_47298_n11874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5843 a_52634_n14207# a_52630_n14030# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5844 a_52374_3776# a_52370_3953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5845 a_56617_n3747# a_56196_n3747# a_55569_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5846 a_55934_8228# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5847 a_30910_8365# a_31167_8175# a_29866_7513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5848 a_20209_n11246# a_20205_n11069# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5849 gnd d0 a_74560_n12775# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5850 a_33429_12112# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5851 gnd a_51838_n11928# a_51630_n11928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5852 a_56407_n11202# a_56194_n11202# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5853 vdd a_39641_n14223# a_39433_n14223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5854 a_44600_3145# a_45440_3820# a_45648_3820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5855 a_11348_13669# a_11969_13561# a_12177_13561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5856 a_47305_n5747# a_47191_n5866# a_47399_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5857 a_47040_12117# a_46931_12117# a_47139_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5858 a_49834_11411# a_49926_9776# a_49877_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5859 a_22980_n13393# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5860 a_65704_n14477# a_65704_n14732# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5861 a_20208_n8028# a_20465_n8218# a_19164_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5862 vdd d2 a_60842_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5863 a_13064_n5194# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5864 a_9242_4544# a_9495_4531# a_8190_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5865 a_63081_6737# a_63077_6914# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5866 a_33022_3146# a_33641_3137# a_33849_3137# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5867 vdd a_8706_n11928# a_8498_n11928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5868 a_36397_n4429# a_36184_n4429# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5869 a_77241_n14167# a_78081_n14171# a_78289_n14171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5870 a_70124_5271# a_70488_8184# a_70443_8197# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5871 a_3543_13562# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5872 a_71765_n12582# a_71857_n14217# a_71812_n14204# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5873 a_23194_n4418# a_22981_n4418# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5874 a_82215_11403# a_82307_9768# a_82258_9958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5875 a_639_3903# a_1260_3824# a_1468_3824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5876 vdd a_39383_9768# a_39175_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5877 vdd a_17927_n6768# a_17719_n6768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5878 gnd d3 a_82730_n12778# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5879 a_8453_n11915# a_9546_n11253# a_9501_n11240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5880 gnd d4 a_59731_8180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5881 a_74309_n6754# a_74562_n6767# a_73261_n7429# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5882 gnd a_75558_n1647# a_75350_n1647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5883 gnd d1 a_19156_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5884 gnd d0 a_9494_6730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5885 vdd a_52628_13506# a_52420_13506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5886 vdd a_19414_n11934# a_19206_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5887 a_73259_n13437# a_73512_n13450# a_71812_n14204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5888 a_1520_n14838# a_1307_n14838# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5889 a_47149_n7388# a_46936_n7388# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5890 a_72998_7513# a_73251_7500# a_71551_6746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5891 a_77034_n3745# a_76821_n3745# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5892 gnd a_9495_5210# a_9287_5210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5893 a_23143_9151# a_22722_9151# a_22311_8571# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5894 a_51327_13523# a_52420_14185# a_52371_14375# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5895 a_44599_6791# a_44178_6791# a_43770_6475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5896 a_66111_n11873# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5897 vdd d1 a_41090_n7448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5898 vdd d3 a_28892_n6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5899 a_55936_14236# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5900 gnd a_74559_n9808# a_74351_n9808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5901 a_57746_6103# a_57637_6103# a_57845_6103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5902 a_20206_n14036# a_20463_n14226# a_19162_n14888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5903 gnd d1 a_73514_n8889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5904 a_44600_3824# a_44179_3824# a_43771_3508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5905 a_30913_10727# a_30917_9782# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5906 vdd a_74562_n8893# a_74354_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5907 vdd d2 a_50394_n8207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5908 a_24029_n5190# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5909 a_56148_3814# a_55935_3814# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5910 a_43773_9261# a_44394_9153# a_44602_9153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5911 a_9237_6920# a_9241_6064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5912 a_1522_n8830# a_1309_n8830# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5913 a_74047_3774# a_74300_3761# a_72999_3099# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5914 a_54480_13128# a_54480_12872# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5915 a_74048_12070# a_74044_12247# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5916 gnd d0 a_63597_n7450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5917 a_9502_n13439# a_9755_n13452# a_8450_n13258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5918 a_83963_n14713# a_85060_n14907# a_85011_n14717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5919 a_58008_n5872# a_57644_n7394# a_56618_n8161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5920 a_11348_13669# a_11348_13128# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5921 a_6748_12756# a_7001_12743# a_6706_11234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5922 a_65853_12118# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5923 a_67321_5265# a_66900_5265# a_66273_5269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5924 gnd a_74302_9090# a_74094_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5925 vdd a_81664_n9805# a_81456_n9805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5926 a_74048_12749# a_74301_12736# a_73000_12074# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5927 a_62295_n5913# a_62548_n5926# a_60844_n5056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5928 vdd d1 a_73253_12061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5929 a_31172_n5736# a_31177_n6754# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5930 a_898_n11508# a_1519_n11192# a_1727_n11192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5931 a_76773_3137# a_76560_3137# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5932 a_639_5606# a_1259_6112# a_1467_6112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5933 a_39385_n5058# a_39642_n5248# a_39347_n6757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5934 a_79419_6101# a_79055_4579# a_78029_5259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5935 a_23400_n9747# a_22979_n9747# a_22571_n10063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5936 a_71548_3956# a_71805_3766# a_71505_5401# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5937 a_55307_8232# a_54886_8232# a_54478_7916# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5938 vdd d0 a_52627_3763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5939 a_40575_3093# a_41668_3755# a_41623_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5940 a_46674_4587# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5941 a_23142_14244# a_22721_14244# a_22313_13928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5942 vdd d0 a_63336_13500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5943 a_44601_12799# a_44180_12799# a_43772_12483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5944 a_76819_n9753# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5945 a_51327_13523# a_51580_13510# a_49880_12756# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5946 vdd a_73513_n5922# a_73305_n5922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5947 a_6964_n12757# a_7051_n11248# a_7002_n11058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5948 a_41621_9274# a_41878_9084# a_40573_9278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5949 a_47147_n13396# a_46934_n13396# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5950 a_24240_n9751# a_24027_n9751# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5951 a_68864_n5868# a_68651_n5868# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5952 a_18902_4542# a_19995_5204# a_19950_5217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5953 a_64406_n15026# a_66325_n14840# a_66533_n14840# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5954 a_11754_8232# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5955 vdd d0 a_31168_5208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5956 a_67161_n5190# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5957 a_63338_n12589# a_63595_n12779# a_62294_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5958 a_13223_6781# a_12802_6781# a_12175_6106# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5959 a_12176_4586# a_11755_4586# a_11347_4694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5960 a_74304_n5736# a_74561_n5926# a_73256_n5732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5961 vdd a_41877_14177# a_41669_14177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5962 gnd a_85267_n11261# a_85059_n11261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5963 a_79054_7546# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5964 a_45647_6787# a_46886_7554# a_47043_6228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5965 a_33848_6783# a_33427_6783# a_33019_6862# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5966 gnd a_9755_n14899# a_9547_n14899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5967 a_35922_7546# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5968 a_44862_n7383# a_44441_n7383# a_44033_n7275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5969 a_76774_12112# a_76561_12112# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5970 a_901_n7816# a_901_n8072# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5971 a_2356_n5188# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5972 a_19945_8361# a_19949_7505# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5973 a_7002_n11058# a_8498_n11928# a_8453_n11915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5974 a_17714_n11241# a_17967_n11254# a_17672_n12763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5975 a_11608_n5506# a_11608_n5761# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5976 gnd a_9496_13506# a_9288_13506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5977 a_22935_9830# a_22722_9830# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5978 a_62031_13694# a_63128_13500# a_63079_13690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5979 a_9500_n7254# a_9504_n8199# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5980 a_19946_5394# a_20203_5204# a_18902_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5981 a_13486_n8161# a_13065_n8161# a_12438_n8836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5982 a_12438_n7389# a_12017_n7389# a_11609_n7822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5983 a_45909_n3741# a_45488_n3741# a_44861_n4416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5984 vdd a_7219_n6762# a_7011_n6762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5985 a_45649_12795# a_45228_12795# a_44601_12120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5986 vdd d1 a_84220_n14903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5987 a_50140_n5227# a_51632_n4473# a_51587_n4460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5988 a_49834_11411# a_49926_9776# a_49881_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5989 a_55102_9826# a_54889_9826# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5990 a_55147_n12718# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5991 a_83967_n14890# a_85060_n14228# a_85015_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5992 a_9238_4721# a_9495_4531# a_8190_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5993 a_68976_n11757# a_68606_n10431# a_67580_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5994 a_36547_n11882# a_36183_n13404# a_35157_n14171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5995 gnd d0 a_31170_11216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5996 a_7009_n8194# a_8501_n7440# a_8452_n7250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5997 a_45910_n6708# a_45489_n6708# a_44862_n6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5998 a_44181_9153# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5999 gnd d3 a_50351_n6762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6000 vdd a_85267_n11940# a_85059_n11940# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6001 gnd a_52887_n14220# a_52679_n14220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6002 a_12229_n4422# a_12016_n4422# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6003 a_19947_12922# a_19951_12066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6004 a_30917_9103# a_30913_9280# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6005 a_77033_n14846# a_76820_n14846# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6006 a_11608_n5111# a_12229_n5190# a_12437_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6007 vdd d3 a_82732_n6770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6008 a_62296_n7433# a_63389_n6771# a_63344_n6758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6009 a_13278_n6714# a_13065_n6714# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6010 gnd a_60842_9770# a_60634_9770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6011 gnd a_39380_6727# a_39172_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6012 a_66111_n10426# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6013 vdd d5 a_70611_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6014 a_4652_9144# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6015 a_48451_5273# a_48815_8186# a_48766_8376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6016 a_57644_n7394# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6017 a_43771_5350# a_43771_4955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6018 vdd d4 a_59731_8180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6019 gnd d2 a_28935_n8209# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6020 a_76981_5263# a_76560_5263# a_76152_5342# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6021 a_44859_n11871# a_44438_n11871# a_44030_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6022 a_74303_n14711# a_75371_n15022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6023 gnd d1 a_40830_10535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6024 vdd d0 a_9494_6730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6025 vdd a_82775_n8215# a_82567_n8215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6026 a_62294_n13441# a_62547_n13454# a_60847_n14208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6027 vdd a_9755_n14220# a_9547_n14220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6028 a_41881_n7262# a_41885_n8207# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6029 vdd a_9495_5210# a_9287_5210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6030 a_25690_n7390# a_25477_n7390# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6031 a_33282_n7028# a_33282_n7283# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6032 a_44861_n3737# a_44440_n3737# a_44032_n3658# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6033 a_51327_13523# a_52420_14185# a_52375_14198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6034 a_11349_10957# a_11349_10702# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6035 a_57383_13556# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6036 gnd a_31170_10537# a_30962_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6037 gnd a_59991_n9803# a_59783_n9803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6038 a_68822_n7390# a_68609_n7390# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6039 a_76983_9824# a_77823_9820# a_78031_9820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6040 a_54478_8311# a_54478_7916# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6041 a_22572_n13285# a_22572_n13826# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6042 a_14713_6103# a_14292_6103# a_14614_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6043 vdd a_38272_8178# a_38064_8178# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6044 a_45701_n3741# a_45488_n3741# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6045 a_56356_5261# a_55935_5261# a_55308_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6046 a_77240_n11200# a_76819_n11200# a_76411_n11121# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6047 gnd d0 a_42138_n8220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6048 a_12230_n7389# a_12017_n7389# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6049 a_84751_3266# a_76154_3146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6050 a_44860_n14159# a_44439_n14159# a_44031_n14475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6051 a_74043_3951# a_74300_3761# a_72999_3099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6052 a_82520_n14210# a_82773_n14223# a_82473_n12588# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6053 a_11756_13561# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6054 a_6744_12933# a_7001_12743# a_6706_11234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6055 a_46978_n5866# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6056 a_46718_12117# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6057 a_41882_n11248# a_41878_n11071# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6058 a_63082_4538# a_63078_4715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6059 a_74044_12926# a_74301_12736# a_73000_12074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6060 a_55149_n8836# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6061 vdd d0 a_85009_14177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6062 a_17454_6742# a_18946_7496# a_18897_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6063 gnd d0 a_74302_9769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6064 a_31176_n5234# a_31429_n5247# a_30128_n5909# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6065 vdd a_19155_4529# a_18947_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6066 a_60582_6919# a_60839_6729# a_60544_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6067 a_58011_n11761# a_57897_n11880# a_58105_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6068 a_52630_n13262# a_52634_n14207# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6069 a_44031_n13283# a_44031_n13824# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6070 a_63339_n5061# a_63343_n5917# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6071 a_9499_n3608# a_9756_n3798# a_8455_n4460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6072 a_1261_14246# a_1048_14246# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6073 vdd d1 a_73512_n13450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6074 a_76412_n13291# a_76412_n13832# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6075 gnd d1 a_30120_4533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6076 a_51323_13700# a_51580_13510# a_49880_12756# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6077 a_28377_5224# a_28464_6733# a_28415_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6078 a_84750_8359# a_85007_8169# a_83706_7507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6079 gnd d0 a_41878_10531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6080 a_66327_n8832# a_66114_n8832# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6081 a_2778_n8155# a_2357_n8155# a_1730_n8830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6082 a_66274_13565# a_65853_13565# a_65445_13132# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6083 a_41625_11223# a_41621_11400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6084 a_66272_6789# a_65851_6789# a_65443_6473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6085 vdd a_8707_n14895# a_8499_n14895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6086 a_44599_8238# a_44178_8238# a_43770_8317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6087 a_51588_n8874# a_51841_n8887# a_50137_n8017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6088 a_17452_12927# a_18948_12057# a_18899_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6089 a_18901_6062# a_19994_6724# a_19945_6914# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6090 a_41884_n4472# a_42137_n4485# a_40832_n4291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6091 gnd d0 a_63335_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6092 a_83966_n10476# a_85059_n9814# a_85010_n9624# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6093 a_23195_n6706# a_22982_n6706# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6094 a_57639_12111# a_57426_12111# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6095 a_84752_12241# a_84757_11223# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6096 a_41625_9776# a_41621_9953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6097 a_55308_3139# a_54887_3139# a_54479_3247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6098 a_22719_6110# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6099 a_54741_n7026# a_54741_n7281# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6100 a_83965_n8705# a_85062_n8899# a_85017_n8886# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6101 a_24188_8232# a_23767_8232# a_23140_7557# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6102 a_11755_3139# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6103 a_82259_6740# a_82512_6727# a_82217_5218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6104 a_900_n4308# a_900_n4849# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6105 a_8194_4548# a_9287_5210# a_9238_5400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6106 a_78028_8226# a_77607_8226# a_76980_7551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6107 a_76820_n14846# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6108 a_65703_n10063# a_65703_n10318# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6109 gnd a_31427_n10487# a_31219_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6110 a_2309_14242# a_2096_14242# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6111 a_22313_13132# a_22313_12876# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6112 a_44599_8238# a_45439_8234# a_45647_8234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6113 a_22574_n8724# a_23195_n8832# a_23403_n8832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6114 a_19949_6737# a_20202_6724# a_18901_6062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6115 a_82517_n5058# a_84013_n5928# a_83968_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6116 a_27091_5271# a_32644_984# a_21717_973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6117 a_13223_8228# a_12802_8228# a_12175_8232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6118 vdd d0 a_31170_11216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6119 a_34735_n11204# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6120 a_72997_9284# a_74094_9090# a_74045_9280# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6121 a_51586_n13435# a_52679_n12773# a_52634_n12760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6122 gnd a_20204_12053# a_19996_12053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6123 a_77243_n8159# a_76822_n8159# a_76414_n8475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6124 a_1047_5271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6125 a_2570_n8155# a_2357_n8155# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6126 a_74306_n11242# a_74559_n11255# a_73258_n11917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6127 gnd d0 a_74302_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6128 a_77242_n5871# a_76821_n5871# a_76413_n5763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6129 a_39389_n5235# a_40881_n4481# a_40836_n4468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6130 vdd d1 a_30379_n11930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6131 vdd d0 a_9757_n8212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6132 a_52636_n7431# a_52889_n7444# a_51584_n7250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6133 a_23982_12793# a_23769_12793# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6134 vdd a_60842_9770# a_60634_9770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6135 a_55146_n10430# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6136 a_40837_n7435# a_41930_n6773# a_41885_n6760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6137 a_48451_5273# a_48815_8186# a_48770_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6138 a_17408_5397# a_17665_5207# a_16342_8370# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6139 a_14713_6103# a_15573_9138# a_15781_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6140 gnd d0 a_9754_n11932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6141 a_50138_n11235# a_51630_n10481# a_51585_n10468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6142 a_66113_n5186# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6143 a_76982_12791# a_76561_12791# a_76153_12475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6144 vdd d1 a_40830_10535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6145 a_24241_n12718# a_24028_n12718# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6146 a_37378_5265# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6147 a_37293_n8847# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6148 gnd a_52629_9771# a_52421_9771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6149 a_1728_n12712# a_2568_n12716# a_2776_n12716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6150 a_1308_n5184# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6151 a_43770_7126# a_43770_6870# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6152 a_13016_5261# a_12803_5261# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6153 a_33022_11606# a_33022_11350# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6154 gnd a_71764_11219# a_71556_11219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6155 a_76412_n13291# a_77033_n13399# a_77241_n13399# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6156 gnd a_9494_6730# a_9286_6730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6157 a_39128_3773# a_39381_3760# a_39081_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6158 a_7003_n14025# a_8499_n14895# a_8454_n14882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6159 a_65446_10961# a_65446_10706# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6160 a_65443_6868# a_65443_6473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6161 a_55361_n5190# a_55148_n5190# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6162 a_45650_9828# a_45229_9828# a_44602_9153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6163 a_45908_n14163# a_45487_n14163# a_44860_n14159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6164 vdd d3 a_28632_11219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6165 gnd a_74299_6049# a_74091_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6166 a_25217_10593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6167 vdd a_85269_n5253# a_85061_n5253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6168 a_33690_n8838# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6169 a_82515_n11066# a_84011_n11936# a_83962_n11746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6170 a_8453_n10468# a_8706_n10481# a_7006_n11235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6171 a_34689_3812# a_34476_3812# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6172 a_54479_4949# a_55100_5265# a_55308_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6173 a_24449_n12718# a_24028_n12718# a_23401_n12714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6174 gnd a_8448_12063# a_8240_12063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6175 a_12436_n12718# a_13276_n12722# a_13484_n12722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6176 a_43772_12228# a_44393_12120# a_44601_12120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6177 a_22314_10706# a_22935_10598# a_23143_10598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6178 a_11969_12114# a_11756_12114# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6179 a_29869_10554# a_30962_11216# a_30913_11406# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6180 a_65851_8236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6181 a_68711_6107# a_68347_4585# a_67321_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6182 vdd d1 a_30120_4533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6183 vdd d1 a_62547_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6184 a_28377_5224# a_28464_6733# a_28419_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6185 a_22571_n9668# a_22571_n10063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6186 a_28422_9787# a_29914_10541# a_29865_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6187 vdd d0 a_41878_10531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6188 a_60586_6742# a_62078_7496# a_62033_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6189 a_44031_n14080# a_44652_n14159# a_44860_n14159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6190 vdd d0 a_20465_n7450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6191 a_29865_9284# a_30122_9094# a_28418_9964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6192 a_56407_n9755# a_56194_n9755# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6193 a_12016_n5190# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6194 a_53727_n1632# a_53677_n1645# a_48780_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6195 a_33642_13559# a_33429_13559# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6196 a_81411_n9792# a_82524_n6770# a_82479_n6757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6197 a_76560_3137# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6198 a_43771_4955# a_43771_4700# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6199 a_76152_3500# a_76773_3816# a_76981_3816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6200 a_70453_n5915# a_70403_n5928# a_70138_n8841# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6201 a_76821_n4424# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6202 gnd d3 a_82472_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6203 a_30127_n14884# a_30380_n14897# a_28676_n14027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6204 a_44862_n8151# a_45702_n8155# a_45910_n8155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6205 a_77870_n6716# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6206 gnd d1 a_73252_3086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6207 a_33021_12475# a_33021_12220# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6208 a_28635_n6574# a_28727_n8209# a_28678_n8019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6209 a_6706_11234# a_6959_11221# a_5638_8199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6210 a_20212_n8205# a_20465_n8218# a_19164_n8880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6211 a_44032_n3402# a_52888_n3798# a_51587_n4460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6212 a_18901_6062# a_19994_6724# a_19949_6737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6213 a_1468_5271# a_1047_5271# a_639_5350# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6214 a_29866_7513# a_30959_8175# a_30910_8365# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6215 vdd d0 a_63335_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6216 a_39130_9781# a_40622_10535# a_40573_10725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6217 vdd d0 a_31167_6728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6218 vdd a_85268_n14907# a_85060_n14907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6219 vdd a_31168_5208# a_30960_5208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6220 gnd a_8706_n11928# a_8498_n11928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6221 a_41879_n12591# a_42136_n12781# a_40835_n13443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6222 a_66112_n13393# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6223 a_54478_7916# a_54478_7661# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6224 a_66324_n11194# a_66111_n11194# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6225 gnd d0 a_52627_3084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6226 a_40571_3270# a_41668_3076# a_41619_3266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6227 a_22312_3506# a_22312_3251# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6228 a_55360_n14844# a_55147_n14844# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6229 a_71765_n12582# a_71857_n14217# a_71808_n14027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6230 a_44032_n5755# a_44033_n6369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6231 gnd a_63596_n3804# a_63388_n3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6232 gnd a_17927_n6768# a_17719_n6768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6233 a_8194_4548# a_9287_5210# a_9242_5223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6234 a_74047_3774# a_74043_3951# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6235 a_80723_5265# a_80510_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6236 a_44392_5271# a_44179_5271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6237 a_33279_n11771# a_33900_n11879# a_34108_n11879# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6238 a_83708_13515# a_84801_14177# a_84756_14190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6239 a_22722_9830# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6240 a_19945_6914# a_20202_6724# a_18901_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6241 gnd a_19414_n11934# a_19206_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6242 a_12435_n9751# a_13275_n9755# a_13483_n9755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6243 a_22311_8315# a_22932_8236# a_23140_8236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6244 gnd d1 a_41090_n7448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6245 gnd d3 a_28892_n6764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6246 a_20209_n11925# a_20205_n11748# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6247 gnd d0 a_42136_n12781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6248 a_9243_13519# a_9239_13696# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6249 a_34690_12787# a_34477_12787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6250 a_20210_n14213# a_20463_n14226# a_19162_n14888# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6251 a_66065_3822# a_65852_3822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6252 vdd a_20204_12053# a_19996_12053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6253 a_12178_11273# a_11757_11273# a_11349_11352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6254 a_60847_n14208# a_61100_n14221# a_60800_n12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6255 a_44030_n9666# a_44030_n10061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6256 vdd d0 a_74559_n9808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6257 a_66275_9151# a_65854_9151# a_65446_9259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6258 a_76414_n7283# a_76414_n7824# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6259 gnd d0 a_52629_11218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6260 a_34109_n14846# a_34949_n14171# a_35157_n14171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6261 a_30916_14196# a_31169_14183# a_29868_13521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6262 a_55937_9822# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6263 gnd a_60839_6729# a_60631_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6264 a_77823_11267# a_77610_11267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6265 a_39389_n5235# a_39642_n5248# a_39347_n6757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6266 gnd d2 a_7000_3768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6267 a_11606_n10863# a_11606_n11119# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6268 a_19158_n13264# a_20255_n13458# a_20210_n13445# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6269 gnd d0 a_85270_n8899# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6270 a_54741_n6631# a_54741_n7026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6271 a_17453_9960# a_18949_9090# a_18904_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6272 a_30123_n14707# a_31220_n14901# a_31171_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6273 a_68810_6107# a_68389_6107# a_68716_6226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6274 a_68562_10593# a_68349_10593# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6275 vdd a_52629_9771# a_52421_9771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6276 vdd d0 a_20204_14179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6277 a_67375_n8157# a_67162_n8157# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6278 a_40836_n4468# a_41089_n4481# a_39389_n5235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6279 a_60804_n12763# a_60891_n11254# a_60846_n11241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6280 a_77242_n5192# a_78082_n5196# a_78290_n5196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6281 a_63342_n12766# a_63595_n12779# a_62294_n13441# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6282 a_74306_n9795# a_74302_n9618# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6283 a_41885_n6760# a_42138_n6773# a_40837_n7435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6284 vdd a_50393_n5240# a_50185_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6285 vout a_2731_n1225# a_3053_n1225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6286 a_36225_n11882# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6287 vdd a_74560_n13454# a_74352_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6288 a_74308_n5913# a_74561_n5926# a_73256_n5732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6289 a_69670_9142# a_69457_9142# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6290 a_65445_13928# a_65445_13673# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6291 vdd a_9494_6730# a_9286_6730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6292 a_39124_3950# a_39381_3760# a_39081_5395# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6293 a_39126_9958# a_40622_9088# a_40573_9278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6294 gnd d1 a_51581_9096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6295 a_52636_n7431# a_52632_n7254# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6296 a_639_3253# a_1260_3145# a_1468_3145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6297 a_20206_n14036# a_20210_n14892# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6298 a_22982_n8832# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6299 a_9242_5223# a_9238_5400# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6300 a_7002_n11058# a_8498_n11928# a_8449_n11738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6301 vdd a_8448_12063# a_8240_12063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6302 a_44859_n9745# a_44438_n9745# a_44030_n10061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6303 vdd a_42138_n8899# a_41930_n8899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6304 a_71807_n11060# a_72064_n11250# a_71769_n12759# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6305 a_2354_n11196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6306 gnd d0 a_9494_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6307 a_74048_12749# a_74044_12926# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6308 a_29869_10554# a_30962_11216# a_30917_11229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6309 a_76154_10700# a_76154_10159# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6310 a_1520_n14159# a_1307_n14159# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6311 a_41623_5215# a_41876_5202# a_40575_4540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6312 a_66111_n11194# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6313 a_22933_4590# a_22720_4590# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6314 gnd a_62289_10537# a_62081_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6315 a_73257_n7252# a_73514_n7442# a_71814_n8196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6316 a_45439_8234# a_45226_8234# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6317 a_22571_n10318# a_23192_n10426# a_23400_n10426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6318 gnd d1 a_62287_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6319 a_9240_10729# a_9244_9784# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6320 a_28422_9787# a_29914_10541# a_29869_10554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6321 a_76982_14238# a_76561_14238# a_76153_14317# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6322 a_39387_n11243# a_40879_n10489# a_40834_n10476# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6323 gnd a_74302_9769# a_74094_9769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6324 a_52631_n4287# a_52635_n5232# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6325 a_44600_3145# a_44179_3145# a_43773_3154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6326 gnd a_30119_7500# a_29911_7500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6327 a_33849_3816# a_33428_3816# a_33020_3500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6328 a_45648_5267# a_46887_4587# a_47038_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6329 a_35923_4579# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6330 vdd d1 a_62548_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6331 vdd d3 a_82472_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6332 gnd d1 a_51838_n10481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6333 a_73257_n7252# a_74354_n7446# a_74309_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6334 a_1522_n8151# a_1309_n8151# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6335 vdd d1 a_73252_3086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6336 a_74047_3095# a_74300_3082# a_72995_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6337 a_67580_n11198# a_67159_n11198# a_66532_n11873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6338 a_45227_3820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6339 a_6702_11411# a_6959_11221# a_5638_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6340 a_83967_n14890# a_85060_n14228# a_85011_n14038# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6341 a_65706_n7818# a_66327_n7385# a_66535_n7385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6342 a_1727_n9745# a_2567_n9749# a_2775_n9749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6343 a_14621_12230# a_14251_13556# a_13225_14236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6344 a_39130_9781# a_40622_10535# a_40577_10548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6345 a_29866_7513# a_30959_8175# a_30914_8188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6346 gnd d0 a_41877_13498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6347 a_13062_n11202# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6348 a_74048_12070# a_74301_12057# a_72996_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6349 vdd d1 a_30380_n14897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6350 a_6746_6748# a_8238_7502# a_8189_7692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6351 gnd d0 a_20463_n14905# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6352 a_9501_n11240# a_9497_n11063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6353 vdd d0 a_85270_n8220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6354 vdd d0 a_52627_3084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6355 a_40571_3270# a_41668_3076# a_41623_3089# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6356 a_23141_4590# a_23981_5265# a_24189_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6357 a_78290_n5196# a_77869_n5196# a_77242_n5192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6358 gnd d0 a_20202_8171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6359 gnd a_85267_n11940# a_85059_n11940# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6360 a_62295_n5913# a_63388_n5251# a_63339_n5061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6361 a_65444_4698# a_65444_4157# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6362 gnd d3 a_82732_n6770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6363 vdd d2 a_17970_n8213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6364 gnd a_63335_4525# a_63127_4525# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6365 a_11607_n12383# a_12227_n11877# a_12435_n11877# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6366 a_65704_n14477# a_66325_n14161# a_66533_n14161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6367 gnd d5 a_70611_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6368 a_8455_n4460# a_8708_n4473# a_7008_n5227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6369 vdd a_51841_n8887# a_51633_n8887# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6370 a_27311_8197# a_28424_11219# a_28379_11232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6371 a_14619_6222# a_14249_7548# a_13223_6781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6372 a_74304_n5057# a_74561_n5247# a_73260_n5909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6373 a_23402_n4418# a_22981_n4418# a_22573_n4851# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6374 a_83708_12068# a_83961_12055# a_82257_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6375 vdd a_31427_n11934# a_31219_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6376 gnd a_82775_n8215# a_82567_n8215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6377 a_24451_n6710# a_24030_n6710# a_23403_n7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6378 gnd a_9755_n14220# a_9547_n14220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6379 a_33848_6104# a_33427_6104# a_33019_6212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6380 gnd a_41878_11210# a_41670_11210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6381 a_76151_7659# a_76151_7118# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6382 a_54738_n9416# a_55362_n8836# a_55570_n8836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6383 a_8193_6068# a_9286_6730# a_9237_6920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6384 a_44651_n9745# a_44438_n9745# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6385 a_63341_n11246# a_63337_n11069# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6386 a_40834_n11923# a_41927_n11261# a_41878_n11071# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6387 a_77032_n10432# a_76819_n10432# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6388 a_36178_6101# a_35965_6101# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6389 a_23983_11273# a_23770_11273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6390 a_2731_n1225# d9 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6391 a_22935_9151# a_22722_9151# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6392 a_62036_9103# a_62289_9090# a_60585_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6393 a_73259_n13437# a_74352_n12775# a_74307_n12762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6394 a_31177_n6754# a_31173_n6577# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6395 a_78082_n3749# a_77869_n3749# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6396 a_1306_n11871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6397 a_30912_14373# a_31169_14183# a_29868_13521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6398 a_45489_n8155# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6399 a_9498_n13262# a_9755_n13452# a_8450_n13258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6400 a_79270_10587# a_79057_10587# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6401 a_69072_n5868# a_68651_n5868# a_68973_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6402 a_13486_n6714# a_13065_n6714# a_12438_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6403 vdd d1 a_51840_n5920# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6404 a_9237_6241# a_9242_5223# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6405 a_20212_n7437# a_20208_n7260# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6406 a_76822_n6712# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6407 a_55102_9147# a_54889_9147# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6408 gnd d1 a_73512_n13450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6409 a_65705_n4055# a_66326_n3739# a_66534_n3739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6410 gnd d3 a_71762_5211# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6411 a_8453_n10468# a_9546_n9806# a_9501_n9793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6412 a_59173_n8845# a_58752_n8845# a_58107_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6413 a_66532_n11873# a_66111_n11873# a_65704_n12379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6414 a_44033_n7275# a_44654_n7383# a_44862_n7383# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6415 a_62291_n5736# a_63388_n5930# a_63343_n5917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6416 a_31172_n5057# a_31176_n5913# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6417 a_4267_n5866# a_3846_n5866# a_4173_n5747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6418 a_12178_9826# a_11757_9826# a_11349_9510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6419 a_49877_9966# a_51373_9096# a_51328_9109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6420 vdd d0 a_20463_n14226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6421 a_25427_7552# a_25214_7552# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6422 vdd a_85267_n11261# a_85059_n11261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6423 a_77867_n11204# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6424 a_1469_12799# a_1048_12799# a_640_12483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6425 a_77033_n14167# a_76820_n14167# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6426 a_54479_5600# a_54479_5344# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6427 a_5210_5273# a_4997_5273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6428 a_13015_6781# a_12802_6781# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6429 a_54887_3818# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6430 a_11968_4586# a_11755_4586# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6431 a_40830_n11746# a_41927_n11940# a_41882_n11927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6432 a_60845_n8023# a_61102_n8213# a_60802_n6578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6433 a_12803_5261# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6434 a_33427_7551# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6435 a_65444_3901# a_66065_3822# a_66273_3822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6436 gnd a_74302_11216# a_74094_11216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6437 a_44859_n11192# a_44438_n11192# a_44030_n11113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6438 a_17713_n8023# a_19209_n8893# a_19164_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6439 vdd d0 a_9494_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6440 a_60842_n11064# a_61099_n11254# a_60804_n12763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6441 gnd d0 a_52886_n11932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6442 a_77240_n11879# a_76819_n11879# a_76411_n11771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6443 a_47038_6109# a_46929_6109# a_47137_6109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6444 a_40572_13692# a_40829_13502# a_39129_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6445 a_11606_n9672# a_12227_n9751# a_12435_n9751# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6446 a_41882_n11927# a_41878_n11750# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6447 gnd d1 a_8707_n14895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6448 a_25216_13560# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6449 vdd d1 a_62287_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6450 a_76153_13667# a_76774_13559# a_76982_13559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6451 a_43773_11358# a_44394_11279# a_44602_11279# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6452 a_51328_10556# a_52421_11218# a_52372_11408# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6453 vdd d3 a_50349_n12770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6454 a_67373_n12718# a_67160_n12718# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6455 a_34476_3812# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6456 a_33850_12112# a_33429_12112# a_33022_11606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6457 a_48205_9144# a_47784_9144# a_47139_12117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6458 vdd a_7217_n12770# a_7009_n12770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6459 a_30913_11406# a_30917_10550# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6460 gnd d4 a_38272_8178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6461 a_76151_8309# a_76772_8230# a_76980_8230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6462 a_74043_3272# a_74300_3082# a_72995_3276# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6463 a_39127_6740# a_40619_7494# a_40574_7507# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6464 vdd d1 a_41088_n13456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6465 a_22573_n4055# a_22573_n4310# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6466 a_43150_941# a_64527_973# a_54311_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6467 a_1046_7559# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6468 a_82517_n5058# a_84013_n5928# a_83964_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6469 a_28421_12754# a_29913_13508# a_29864_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6470 a_1520_n13391# a_1307_n13391# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6471 a_55149_n8157# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6472 a_66067_11277# a_65854_11277# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6473 a_74046_8188# a_74299_8175# a_72998_7513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6474 a_33020_4151# a_33641_4584# a_33849_4584# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6475 gnd d0 a_85010_11210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6476 a_65706_n7277# a_65706_n7818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6477 a_77869_n5196# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6478 gnd d1 a_19155_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6479 gnd a_73252_3086# a_73044_3086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6480 vdd d0 a_20202_8171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6481 vdd a_20464_n3804# a_20256_n3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6482 vdd d3 a_50351_n6762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6483 gnd d1 a_30379_n11930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6484 a_84754_8182# a_84750_8359# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6485 vdd a_17925_n12776# a_17717_n12776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6486 vdd a_63335_4525# a_63127_4525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6487 vdd a_31167_6728# a_30959_6728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6488 a_36137_13554# a_35924_13554# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6489 a_14765_n11880# a_14552_n11880# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6490 a_66327_n8153# a_66114_n8153# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6491 a_23194_n5865# a_22981_n5865# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6492 a_79317_n7396# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6493 a_1729_n4416# a_1308_n4416# a_900_n4308# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6494 a_83704_12245# a_83961_12055# a_82257_12925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6495 a_19947_12243# a_19952_11225# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6496 a_2778_n6708# a_2357_n6708# a_1730_n6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6497 a_56196_n3747# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6498 a_79426_12228# a_79056_13554# a_78030_12787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6499 a_13018_11269# a_12805_11269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6500 vdd a_41878_11210# a_41670_11210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6501 a_60589_9783# a_60842_9770# a_60542_11405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6502 a_8193_6068# a_9286_6730# a_9241_6743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6503 a_18897_6239# a_19994_6045# a_19945_6235# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6504 a_41879_n14038# a_41883_n14894# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6505 a_23403_n8832# a_24243_n8157# a_24451_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6506 a_69070_n11876# a_68649_n11876# a_68971_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6507 a_73259_n14884# a_73512_n14897# a_71808_n14027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6508 a_898_n10857# a_898_n11113# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6509 vdd d0 a_52886_n9806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6510 a_85016_n4472# a_85012_n4295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6511 gnd d1 a_83959_6047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6512 gnd a_85010_10531# a_84802_10531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6513 a_80510_5265# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6514 a_68607_n13398# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6515 a_55569_n5869# a_55148_n5869# a_54741_n6375# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6516 a_19946_3947# a_19950_3091# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6517 a_67374_n3743# a_67161_n3743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6518 gnd a_8449_9096# a_8241_9096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6519 vdd a_41090_n8895# a_40882_n8895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6520 gnd a_9497_10539# a_9289_10539# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6521 a_54481_10702# a_55102_10594# a_55310_10594# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6522 a_82516_n14033# a_82773_n14223# a_82473_n12588# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6523 a_36388_12109# a_35967_12109# a_36289_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6524 a_62032_10727# a_63129_10533# a_63080_10723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6525 a_31170_n11744# a_31175_n12762# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6526 a_2775_n11196# a_4014_n10429# a_4171_n11755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6527 a_66532_n10426# a_66111_n10426# a_65703_n10318# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6528 gnd d0 a_63597_n8897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6529 a_76820_n14167# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6530 a_22572_n13285# a_23193_n13393# a_23401_n13393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6531 a_48681_n5736# a_49075_n9797# a_49026_n9607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6532 a_33900_n9753# a_33687_n9753# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6533 a_2569_n3741# a_2356_n3741# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6534 a_40572_13692# a_41669_13498# a_41620_13688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6535 vdd d1 a_73253_13508# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6536 a_73001_9107# a_74094_9769# a_74045_9959# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6537 a_76773_4584# a_76560_4584# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6538 a_22574_n8074# a_23195_n8153# a_23403_n8153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6539 a_19949_6058# a_20202_6045# a_18897_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6540 vdd d3 a_71762_5211# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6541 gnd d1 a_62547_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6542 a_13226_9822# a_12805_9822# a_12178_9826# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6543 a_898_n9666# a_1519_n9745# a_1727_n9745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6544 gnd d0 a_20465_n7450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6545 a_52370_3953# a_52374_3097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6546 a_14876_n5872# a_14512_n7394# a_13486_n8161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6547 a_1467_7559# a_1046_7559# a_638_7126# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6548 a_53727_n1632# a_53677_n1645# a_53628_n1455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6549 a_34738_n8163# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6550 a_81411_n9792# a_82524_n6770# a_82475_n6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6551 a_17670_n6578# a_17762_n8213# a_17717_n8200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6552 a_14463_4581# a_14250_4581# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6553 a_55936_12789# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6554 vdd a_31430_n7446# a_31222_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6555 a_70453_n5915# a_70403_n5928# a_70354_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6556 a_51325_7515# a_51578_7502# a_49878_6748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6557 a_11346_6214# a_11347_5600# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6558 a_67159_n9751# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6559 a_53628_n1455# a_59438_n5932# a_59389_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6560 a_85010_n11750# a_85015_n12768# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6561 a_68561_13560# a_68348_13560# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6562 a_77242_n5192# a_76821_n5192# a_76413_n5113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6563 a_33280_n13832# a_33901_n13399# a_34109_n13399# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6564 a_70138_n8841# a_69717_n8841# a_69070_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6565 a_51585_n10468# a_52678_n9806# a_52629_n9616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6566 a_65704_n13285# a_65704_n13826# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6567 gnd d0 a_9754_n11253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6568 a_63077_6914# a_63081_6058# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6569 a_4014_n10429# a_3801_n10429# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6570 a_83707_4540# a_84800_5202# a_84755_5215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6571 a_44862_n8830# a_44441_n8830# a_44033_n8722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6572 a_44439_n14838# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6573 a_36292_6220# a_36178_6101# a_36386_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6574 a_65852_5269# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6575 vdd a_74302_11216# a_74094_11216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6576 a_51584_n8697# a_52681_n8891# a_52636_n8878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6577 a_52374_3776# a_52627_3763# a_51326_3101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6578 a_44391_7559# a_44178_7559# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6579 a_23403_n6706# a_22982_n6706# a_22574_n7022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6580 a_9497_n9616# a_9501_n10472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6581 a_45648_5267# a_45227_5267# a_44600_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6582 a_11349_11608# a_11349_11352# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6583 gnd a_52629_9092# a_52421_9092# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6584 a_55361_n5869# a_55148_n5869# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6585 gnd a_39383_9768# a_39175_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6586 a_56408_n12722# a_56195_n12722# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6587 a_12438_n8836# a_12017_n8836# a_11606_n9416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6588 a_22719_7557# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6589 a_14715_12111# a_14294_12111# a_14616_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6590 vdd a_8709_n8887# a_8501_n8887# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6591 gnd a_9494_6051# a_9286_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6592 a_14722_n10435# a_14509_n10435# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6593 a_50136_n5050# a_51632_n5920# a_51587_n5907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6594 a_74045_9959# a_74049_9103# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6595 a_20208_n6581# a_20212_n7437# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6596 a_22720_4590# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6597 a_45226_8234# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6598 a_79357_n11882# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6599 vdd d0 a_63597_n8218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6600 a_1470_10600# a_2310_11275# a_2518_11275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6601 a_33690_n8159# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6602 a_74042_8365# a_74299_8175# a_72998_7513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6603 a_23768_3818# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6604 vdd d0 a_85010_11210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6605 gnd a_30379_n10483# a_30171_n10483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6606 a_12438_n6710# a_12017_n6710# a_11609_n6631# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6607 a_12014_n10430# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6608 a_34110_n4424# a_34950_n3749# a_35158_n3749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6609 vdd a_73252_3086# a_73044_3086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6610 a_44859_n11871# a_45699_n11196# a_45907_n11196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6611 a_24188_8232# a_25427_7552# a_25584_6226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6612 a_13015_8228# a_12802_8228# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6613 a_11347_3897# a_11347_3502# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6614 a_34899_11267# a_36138_10587# a_36289_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6615 vdd a_85267_n9814# a_85059_n9814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6616 a_11348_12477# a_11348_12222# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6617 a_39087_11226# a_39340_11213# a_38019_8191# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6618 a_43773_9516# a_43773_9261# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6619 vdd d0 a_9754_n11932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6620 vdd d1 a_84222_n8895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6621 a_76154_3146# a_76773_3137# a_76981_3137# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6622 a_76413_n4857# a_76413_n5113# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6623 a_33901_n12720# a_33688_n12720# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6624 a_19158_n13264# a_20255_n13458# a_20206_n13268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6625 a_41878_n9624# a_41882_n10480# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6626 a_14465_10589# a_14252_10589# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6627 a_24191_11273# a_23770_11273# a_23143_11277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6628 a_60585_9960# a_60842_9770# a_60542_11405# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6629 gnd a_20202_8171# a_19994_8171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6630 a_33279_n9418# a_33279_n9674# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6631 vdd d1 a_19156_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6632 a_2097_9828# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6633 a_18897_6239# a_19994_6045# a_19949_6058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6634 a_62294_n14888# a_62547_n14901# a_60843_n14031# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6635 a_44862_n7383# a_45702_n6708# a_45910_n6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6636 vdd d0 a_31167_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6637 vdd d1 a_62288_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6638 a_60804_n12763# a_60891_n11254# a_60842_n11064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6639 a_78288_n11204# a_79527_n10437# a_79684_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6640 vdd a_85010_10531# a_84802_10531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6641 a_12014_n9751# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6642 vdd a_63597_n7450# a_63389_n7450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6643 gnd a_50393_n5240# a_50185_n5240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6644 a_76561_13559# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6645 a_33019_8309# a_33019_7914# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6646 gnd a_74560_n13454# a_74352_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6647 a_40831_n14713# a_41928_n14907# a_41883_n14894# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6648 a_12177_14240# a_11756_14240# a_11348_13924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6649 a_55360_n14165# a_55147_n14165# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6650 a_12230_n8836# a_12017_n8836# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6651 gnd a_41877_14177# a_41669_14177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6652 a_30917_10550# a_30913_10727# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6653 a_28680_n14204# a_30172_n13450# a_30127_n13437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6654 a_45699_n11196# a_45486_n11196# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6655 a_62036_9103# a_63129_9765# a_63080_9955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6656 a_22573_n3660# a_22573_n4055# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6657 a_62032_10727# a_63129_10533# a_63084_10546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6658 a_33848_7551# a_34688_8226# a_34896_8226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6659 vdd d3 a_60797_5207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6660 a_899_n12633# a_1520_n12712# a_1728_n12712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6661 a_77822_14234# a_77609_14234# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6662 a_44032_n4053# a_44653_n3737# a_44861_n3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6663 a_22313_12876# a_22313_12481# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6664 a_33279_n11121# a_33900_n11200# a_34108_n11200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6665 a_8449_n10291# a_8706_n10481# a_7006_n11235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6666 a_55570_n6710# a_55149_n6710# a_54741_n7026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6667 a_54739_n12383# a_55359_n11877# a_55567_n11877# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6668 a_71811_n11237# a_72064_n11250# a_71769_n12759# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6669 a_22722_9151# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6670 a_19945_6235# a_20202_6045# a_18897_6239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6671 a_11608_n4314# a_11608_n4855# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6672 a_83709_10548# a_84802_11210# a_84753_11400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6673 a_66275_9830# a_65854_9830# a_65446_9909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6674 a_56410_n6714# a_56197_n6714# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6675 a_4016_n4421# a_3803_n4421# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6676 a_39387_n11243# a_40879_n10489# a_40830_n10299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6677 a_68348_13560# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6678 a_66065_3143# a_65852_3143# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6679 a_63340_n8707# a_63341_n9799# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6680 gnd d1 a_62548_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6681 a_73257_n7252# a_74354_n7446# a_74305_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6682 gnd d2 a_72066_n5242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6683 a_43772_13134# a_44393_13567# a_44601_13567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6684 a_33851_10592# a_33430_10592# a_33022_10700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6685 a_72996_12251# a_74093_12057# a_74048_12070# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6686 a_66900_5265# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6687 a_22313_13928# a_22934_14244# a_23142_14244# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6688 a_19157_n10297# a_19414_n10487# a_17714_n11241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6689 a_44602_10600# a_44181_10600# a_43773_10167# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6690 a_44033_n6369# a_44033_n6625# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6691 a_41884_n5919# a_42137_n5932# a_40832_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6692 a_640_12483# a_1261_12799# a_1469_12799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6693 a_54886_8232# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6694 a_52370_3953# a_52627_3763# a_51326_3101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6695 a_54738_n9416# a_54738_n9672# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6696 gnd d0 a_85270_n8220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6697 a_54103_986# a_53890_986# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6698 a_55308_4586# a_54887_4586# a_54479_4694# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6699 a_25214_7552# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6700 a_30127_n14884# a_31220_n14222# a_31171_n14032# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6701 vdd d0 a_74561_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6702 a_55148_n3743# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6703 a_79529_n4429# a_79316_n4429# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6704 a_44653_n5863# a_44440_n5863# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6705 a_1260_4592# a_1047_4592# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6706 a_39383_n11066# a_39640_n11256# a_39345_n12765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6707 a_12802_6781# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6708 gnd d0 a_20205_11212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6709 gnd a_51841_n8887# a_51633_n8887# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6710 a_11755_4586# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6711 a_54889_10594# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6712 a_25579_6107# a_25470_6107# a_25678_6107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6713 a_77820_8226# a_77607_8226# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6714 vdd a_28935_n8209# a_28727_n8209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6715 a_5125_n8839# a_4912_n8839# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6716 a_74308_n5234# a_74561_n5247# a_73260_n5909# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6717 a_43770_6475# a_44391_6791# a_44599_6791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6718 gnd a_31427_n11934# a_31219_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6719 vdd a_9494_6051# a_9286_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6720 a_65446_11612# a_65446_11356# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6721 a_74308_n4466# a_74304_n4289# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6722 a_22982_n8153# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6723 a_63078_5394# a_63335_5204# a_62034_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6724 a_2518_11275# a_3757_10595# a_3908_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6725 a_11346_7120# a_11967_7553# a_12175_7553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6726 vdd d0 a_42136_n12781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6727 a_2776_n14163# a_4015_n13396# a_4166_n11874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6728 a_66533_n13393# a_66112_n13393# a_65704_n13285# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6729 vdd a_74561_n3800# a_74353_n3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6730 a_23402_n3739# a_24242_n3743# a_24450_n3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6731 gnd a_38272_8178# a_38064_8178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6732 a_73259_n13437# a_74352_n12775# a_74303_n12585# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6733 a_60843_n14031# a_61100_n14221# a_60800_n12586# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6734 a_33282_n7824# a_33903_n7391# a_34111_n7391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6735 vdd a_62286_6049# a_62078_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6736 a_39385_n5058# a_40881_n5928# a_40836_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6737 a_19159_n4289# a_19416_n4479# a_17716_n5233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6738 a_39083_11403# a_39340_11213# a_38019_8191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6739 a_52636_n8878# a_52889_n8891# a_51584_n8697# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6740 a_43771_5606# a_43771_5350# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6741 a_9501_n11919# a_9497_n11742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6742 a_67160_n14165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6743 gnd d1 a_51840_n5920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6744 a_33849_3137# a_33428_3137# a_33022_3146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6745 a_35158_n3749# a_36397_n4429# a_36554_n5755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6746 gnd d0 a_85009_14177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6747 a_55310_10594# a_56150_11269# a_56358_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6748 a_17410_11405# a_17502_9770# a_17453_9960# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6749 a_50134_n11058# a_51630_n11928# a_51585_n11915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6750 a_73260_n4462# a_74353_n3800# a_74304_n3610# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6751 a_30124_n4285# a_31221_n4479# a_31176_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6752 gnd a_19155_4529# a_18947_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6753 a_33021_13126# a_33021_12870# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6754 vdd a_20202_8171# a_19994_8171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6755 a_60586_6742# a_60839_6729# a_60544_5220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6756 a_34949_n12724# a_34736_n12724# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6757 a_33690_n7391# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6758 a_12175_6106# a_13015_6781# a_13223_6781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6759 a_66532_n9747# a_66111_n9747# a_65703_n9668# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6760 a_62291_n5736# a_63388_n5930# a_63339_n5740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6761 a_22573_n4851# a_23194_n4418# a_23402_n4418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6762 a_84754_8182# a_85007_8169# a_83706_7507# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6763 a_83963_n13266# a_84220_n13456# a_82520_n14210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6764 a_40832_n4291# a_41089_n4481# a_39389_n5235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6765 gnd d0 a_20463_n14226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6766 a_4015_n13396# a_3802_n13396# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6767 a_41881_n6583# a_42138_n6773# a_40837_n7435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6768 a_33900_n10432# a_33687_n10432# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6769 gnd d2 a_61100_n14221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6770 a_76412_n14738# a_77033_n14846# a_77241_n14846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6771 a_62036_9103# a_63129_9765# a_63084_9778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6772 a_63341_n11925# a_63337_n11748# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6773 a_34109_n12720# a_33688_n12720# a_33280_n13036# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6774 a_11606_n11514# a_12227_n11198# a_12435_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6775 gnd a_85009_13498# a_84801_13498# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6776 vdd d0 a_31170_9769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6777 a_1259_8238# a_1046_8238# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6778 a_40830_n11746# a_41927_n11940# a_41878_n11750# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6779 a_41621_9953# a_41625_9097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6780 a_54311_986# a_64740_973# a_43150_941# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6781 a_57845_6103# a_57424_6103# a_57746_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6782 vdd a_31427_n11255# a_31219_n11255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6783 a_60846_n11241# a_61099_n11254# a_60804_n12763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6784 gnd a_8448_13510# a_8240_13510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6785 a_54741_n8473# a_55362_n8157# a_55570_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6786 a_83709_10548# a_84802_11210# a_84757_11223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6787 a_24450_n3743# a_24029_n3743# a_23402_n3739# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6788 a_8189_6245# a_9286_6051# a_9237_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6789 a_85010_n10303# a_85267_n10493# a_83962_n10299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6790 a_9242_3097# a_9238_3274# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6791 gnd d3 a_50349_n12770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6792 a_68604_12115# a_68391_12115# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6793 a_76559_7551# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6794 a_60583_3952# a_62079_3082# a_62030_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6795 a_25428_4585# a_25215_4585# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6796 a_56618_n8161# a_56197_n8161# a_55570_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6797 a_23400_n11873# a_22979_n11873# a_22571_n11765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6798 gnd a_7217_n12770# a_7009_n12770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6799 a_36646_n11882# a_36225_n11882# a_36552_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6800 a_33281_n4061# a_33902_n3745# a_34110_n3745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6801 a_76560_4584# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6802 vdd d1 a_51838_n10481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6803 gnd d1 a_41088_n13456# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6804 a_1306_n11192# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6805 a_33282_n8475# a_33282_n8730# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6806 a_12015_n13397# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6807 a_55568_n14844# a_56408_n14169# a_56616_n14169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6808 gnd d1 a_73252_4533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6809 a_47189_n11874# a_46976_n11874# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6810 a_17456_12750# a_18948_13504# a_18903_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6811 a_37930_n5744# a_38324_n9805# a_38279_n9792# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6812 a_11606_n11514# a_11606_n11769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6813 a_45489_n6708# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6814 a_14250_4581# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6815 a_20207_n5740# a_20212_n6758# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6816 a_66112_n14840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6817 vdd d0 a_9755_n14899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6818 a_33019_7914# a_33019_7659# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6819 a_2775_n11196# a_2354_n11196# a_1727_n11192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6820 a_1468_3145# a_2308_3820# a_2516_3820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6821 vdd d2 a_72064_n11250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6822 gnd d0 a_52627_4531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6823 a_6702_11411# a_6794_9776# a_6745_9966# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6824 a_66532_n11194# a_66111_n11194# a_65703_n11510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6825 gnd a_17925_n12776# a_17717_n12776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6826 a_63338_n14036# a_63342_n14892# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6827 a_62295_n5913# a_63388_n5251# a_63343_n5238# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6828 a_40571_4717# a_41668_4523# a_41619_4713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6829 a_15781_9138# a_15918_5267# a_11080_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6830 vdd d0 a_20205_11212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6831 a_65851_6789# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6832 a_12178_9147# a_11757_9147# a_11346_8567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6833 vdd a_62549_n7446# a_62341_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6834 a_8451_n4283# a_8708_n4473# a_7008_n5227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6835 a_78289_n14171# a_79528_n13404# a_79679_n11882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6836 a_39087_11226# a_39174_12735# a_39125_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6837 gnd a_63336_13500# a_63128_13500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6838 a_8451_n4283# a_9548_n4477# a_9503_n4464# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6839 a_41620_12920# a_41624_12064# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6840 gnd d4 a_49283_n9797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6841 a_23140_8236# a_22719_8236# a_22311_8315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6842 gnd d0 a_41875_7490# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6843 a_56615_n11202# a_57854_n10435# a_58011_n11761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6844 a_55146_n11877# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6845 a_54887_3139# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6846 a_41619_4713# a_41623_3768# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6847 a_34736_n12724# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6848 a_13483_n11202# a_13062_n11202# a_12435_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6849 gnd d1 a_41090_n8895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6850 a_33902_n5871# a_33689_n5871# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6851 a_40834_n11923# a_41927_n11261# a_41882_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6852 a_66066_14244# a_65853_14244# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6853 a_65444_3251# a_66065_3143# a_66273_3143# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6854 a_9240_10729# a_9497_10539# a_8192_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6855 gnd d0 a_52886_n11253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6856 a_22574_n8074# a_22574_n8469# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6857 a_23767_8232# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6858 vdd a_20204_13500# a_19996_13500# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6859 a_82516_n14033# a_84012_n14903# a_83967_n14890# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6860 a_71771_n6751# a_71858_n5242# a_71809_n5052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6861 a_63081_6737# a_63334_6724# a_62033_6062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6862 a_9240_11408# a_9244_10552# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6863 a_84752_14367# a_85009_14177# a_83708_13515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6864 a_15573_9138# a_15360_9138# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6865 gnd d4 a_70956_n9799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6866 gnd d3 a_28632_11219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6867 a_52633_n11240# a_52629_n11063# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6868 a_17410_11405# a_17502_9770# a_17457_9783# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6869 a_11607_n14086# a_11607_n14481# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6870 a_13017_14236# a_12804_14236# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6871 vdd d2 a_82515_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6872 a_12802_8228# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6873 a_11608_n4314# a_12229_n4422# a_12437_n4422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6874 a_52629_n10295# a_52886_n10485# a_51581_n10291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6875 a_65443_6473# a_66064_6789# a_66272_6789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6876 a_22980_n14161# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6877 a_12438_n6710# a_13278_n6714# a_13486_n6714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6878 a_900_n5755# a_901_n6369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6879 a_28637_n12759# a_28724_n11250# a_28679_n11237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6880 a_57854_n10435# a_57641_n10435# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6881 a_14616_12111# a_14252_10589# a_13226_11269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6882 a_68713_12115# a_68349_10593# a_67323_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6883 a_36227_n5874# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6884 gnd a_31430_n7446# a_31222_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6885 a_44180_12120# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6886 a_34896_8226# a_36135_7546# a_36292_6220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6887 a_5894_n9607# a_6151_n9797# a_5549_n5736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6888 a_79421_12109# a_79312_12109# a_79520_12109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6889 vdd a_31169_12057# a_30961_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6890 a_2307_8234# a_2094_8234# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6891 vdd d0 a_74562_n6767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6892 a_3542_4587# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6893 a_1727_n11871# a_1306_n11871# a_898_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6894 gnd a_73511_n10483# a_73303_n10483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6895 vdd a_31167_6049# a_30959_6049# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6896 a_85013_n8030# a_85017_n8886# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6897 a_23194_n5186# a_22981_n5186# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6898 a_74304_n3610# a_74308_n4466# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6899 gnd d0 a_31167_6728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6900 a_67115_9826# a_66902_9826# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6901 a_82217_5218# a_82470_5205# a_81147_8368# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6902 vdd a_74299_7496# a_74091_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6903 a_60540_5397# a_60632_3762# a_60583_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6904 a_55100_5265# a_54887_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6905 a_22314_10165# a_22314_9909# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6906 a_58013_n5753# a_57899_n5872# a_58107_n5872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6907 a_639_3508# a_639_3253# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6908 a_55310_11273# a_54889_11273# a_54481_11352# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6909 vdd a_8448_13510# a_8240_13510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6910 a_39343_n6580# a_39435_n8215# a_39390_n8202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6911 vdd d0 a_52886_n11932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6912 a_24027_n11198# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6913 a_898_n9666# a_898_n10061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6914 a_8189_6245# a_9286_6051# a_9241_6064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6915 a_76819_n11200# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6916 a_34108_n10432# a_33687_n10432# a_33279_n10324# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6917 vdd a_60797_5207# a_60589_5207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6918 vdd a_19415_n14901# a_19207_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6919 a_8194_3101# a_8447_3088# a_6743_3958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6920 a_79056_13554# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6921 a_60583_3952# a_62079_3082# a_62034_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6922 a_74043_3951# a_74047_3095# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6923 a_80832_5265# a_80723_5265# a_75885_984# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6924 a_33428_5263# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6925 a_55569_n5190# a_55148_n5190# a_54740_n5506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6926 a_39383_n11066# a_40879_n11936# a_40834_n11923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6927 a_44438_n10424# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6928 gnd a_8709_n8887# a_8501_n8887# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6929 a_33641_3816# a_33428_3816# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6930 vdd d1 a_62548_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6931 a_50136_n5050# a_51632_n5920# a_51583_n5730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6932 a_78080_n11204# a_77867_n11204# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6933 a_83708_13515# a_84801_14177# a_84752_14367# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6934 vdd d1 a_73252_4533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6935 gnd d0 a_63597_n8218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6936 a_56409_n5194# a_56196_n5194# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6937 a_641_11358# a_1262_11279# a_1470_11279# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6938 vdd a_20463_n12779# a_20255_n12779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6939 a_65703_n9412# a_66327_n8832# a_66535_n8832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6940 vdd d0 a_52888_n4477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6941 a_47997_9144# a_47784_9144# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6942 a_71812_n14204# a_73304_n13450# a_73259_n13437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6943 a_22981_n4418# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6944 a_85017_n6760# a_85270_n6773# a_83969_n7435# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6945 a_33022_9903# a_33643_9824# a_33851_9824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6946 a_72997_9284# a_73254_9094# a_71550_9964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6947 a_66325_n12714# a_66112_n12714# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6948 a_33850_13559# a_33429_13559# a_33021_13667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6949 a_28681_n5229# a_30173_n4475# a_30128_n4462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6950 a_50135_n14025# a_51631_n14895# a_51586_n14882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6951 a_35156_n9757# a_34735_n9757# a_34108_n9753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6952 a_30129_n7429# a_31222_n6767# a_31177_n6754# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6953 a_32169_n1457# a_32426_n1647# a_21532_n1444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6954 a_74046_7509# a_74042_7686# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6955 vdd d0 a_52627_4531# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6956 a_6702_11411# a_6794_9776# a_6749_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6957 a_40571_4717# a_41668_4523# a_41623_4536# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6958 a_44601_13567# a_44180_13567# a_43772_13134# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6959 a_73000_12074# a_74093_12736# a_74044_12926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6960 gnd a_85267_n9814# a_85059_n9814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6961 a_46936_n7388# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6962 a_22574_n7022# a_23195_n6706# a_23403_n6706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6963 a_19160_n8703# a_20257_n8897# a_20212_n8884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6964 a_33902_n4424# a_33689_n4424# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6965 a_12175_8232# a_11754_8232# a_11346_8311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6966 gnd a_31429_n3800# a_31221_n3800# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6967 a_33430_10592# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6968 a_80378_9136# a_80165_9136# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6969 a_39087_11226# a_39174_12735# a_39129_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6970 vdd a_9496_12738# a_9288_12738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6971 a_67320_6785# a_68559_7552# a_68716_6226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6972 a_13276_n12722# a_13063_n12722# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6973 a_84754_6056# a_84750_6233# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6974 a_34738_n6716# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6975 gnd d0 a_74300_5208# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6976 a_900_n4308# a_1521_n4416# a_1729_n4416# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6977 gnd d0 a_20204_14179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6978 a_1730_n6704# a_2570_n6708# a_2778_n6708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6979 a_44862_n8151# a_44441_n8151# a_44033_n8072# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6980 vdd d0 a_85008_5202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6981 a_44439_n14159# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6982 gnd a_63597_n7450# a_63389_n7450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6983 a_5319_5273# a_5683_8186# a_5634_8376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6984 a_1469_14246# a_2309_14242# a_2517_14242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6985 a_18897_6239# a_19154_6049# a_17450_6919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6986 a_51588_n8874# a_52681_n8212# a_52636_n8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6987 a_52374_3097# a_52627_3084# a_51322_3278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6988 a_65445_13673# a_65445_13132# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6989 gnd a_40830_9088# a_40622_9088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6990 a_28680_n14204# a_30172_n13450# a_30123_n13260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6991 a_63077_6914# a_63334_6724# a_62033_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6992 a_4265_n11874# a_3844_n11874# a_4171_n11755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6993 a_67322_14240# a_68561_13560# a_68718_12234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6994 a_79572_n5874# a_79359_n5874# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6995 gnd a_83961_12055# a_83753_12055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6996 a_54740_n5111# a_54740_n5506# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6997 a_33689_n3745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6998 a_12438_n8157# a_12017_n8157# a_11609_n8473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6999 a_19946_3268# a_11349_3148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7000 gnd d4 a_38532_n9805# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7001 vdd d0 a_74301_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7002 a_9243_13519# a_9496_13506# a_8191_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7003 a_46888_13562# a_46675_13562# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7004 a_76775_9824# a_76562_9824# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7005 a_31170_n11065# a_31174_n11921# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7006 vdd d0 a_9757_n7444# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7007 a_22312_4157# a_22933_4590# a_23141_4590# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7008 a_24190_14240# a_23769_14240# a_23142_13565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7009 a_9237_8367# a_9494_8177# a_8193_7515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7010 a_14294_12111# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7011 gnd d1 a_73512_n14897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7012 a_25586_12234# a_25472_12115# a_25680_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7013 a_17672_n12763# a_17759_n11254# a_17714_n11241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7014 a_44652_n14838# a_44439_n14838# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7015 a_54740_n3664# a_55361_n3743# a_55569_n3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7016 a_60802_n6578# a_60894_n8213# a_60845_n8023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7017 a_25940_n5868# a_25519_n5868# a_25841_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7018 a_65854_9151# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7019 a_68971_n11876# a_68607_n13398# a_67581_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7020 a_13018_9822# a_12805_9822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7021 a_9499_n3608# a_9503_n4464# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7022 a_52370_3274# a_43773_3154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7023 a_33849_5263# a_34689_5259# a_34897_5259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7024 a_53628_n1455# a_59438_n5932# a_59173_n8845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7025 a_19161_n10474# a_19414_n10487# a_17714_n11241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7026 a_47303_n11755# a_46933_n10429# a_45907_n9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7027 a_16041_n8845# a_15620_n8845# a_14975_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7028 a_33020_5598# a_33020_5342# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7029 vdd d4 a_81404_8178# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7030 vdd d0 a_9754_n11253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7031 vdd a_5806_n5926# a_5598_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7032 a_36138_10587# a_35925_10587# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7033 a_85010_n11071# a_85014_n11927# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7034 a_60540_5397# a_60632_3762# a_60587_3775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7035 a_2355_n12716# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7036 a_60848_n5233# a_62340_n4479# a_62295_n4466# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7037 a_44652_n12712# a_44439_n12712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7038 gnd d0 a_74561_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7039 a_63077_6235# a_63082_5217# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7040 vdd d0 a_9494_7498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7041 a_82258_9958# a_83754_9088# a_83705_9278# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7042 a_74302_n11744# a_74307_n12762# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7043 a_39387_n11243# a_39640_n11256# a_39345_n12765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7044 gnd d2 a_28675_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7045 a_8456_n7427# a_9549_n6765# a_9504_n6752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7046 a_9244_10552# a_9240_10729# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7047 a_55309_12793# a_54888_12793# a_54480_12872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7048 a_56616_n14169# a_57855_n13402# a_58006_n11880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7049 a_23401_n14161# a_24241_n14165# a_24449_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7050 vdd d1 a_62287_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7051 a_11346_6214# a_11967_6106# a_12175_6106# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7052 a_70354_n5738# a_70748_n9799# a_70699_n9609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7053 vdd a_52886_n9806# a_52678_n9806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7054 a_27311_8197# a_28424_11219# a_28375_11409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7055 a_78288_n11204# a_77867_n11204# a_77240_n11879# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7056 a_12230_n8157# a_12017_n8157# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7057 a_62032_9280# a_63129_9086# a_63080_9276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7058 a_13063_n12722# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7059 a_74043_4719# a_74300_4529# a_72995_4723# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7060 a_34950_n5196# a_34737_n5196# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7061 a_76151_6467# a_76151_6212# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7062 gnd d0 a_31170_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7063 a_55567_n10430# a_56407_n9755# a_56615_n9755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7064 a_12016_n4422# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7065 a_60847_n14208# a_62339_n13454# a_62294_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7066 a_25215_4585# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7067 vdd a_82732_n6770# a_82524_n6770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7068 a_74044_13694# a_74301_13504# a_72996_13698# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7069 a_74045_9280# a_74046_8188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7070 a_54738_n11514# a_55359_n11198# a_55567_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7071 gnd a_73251_7500# a_73043_7500# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7072 a_74302_n9618# a_74559_n9808# a_73258_n10470# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7073 vdd a_30379_n10483# a_30171_n10483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7074 a_41880_n3616# a_41884_n4472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7075 a_33279_n11121# a_33279_n11516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7076 a_66534_n5865# a_66113_n5865# a_65706_n6371# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7077 a_33281_n3410# a_33281_n3666# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7078 a_33021_12220# a_33642_12112# a_33850_12112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7079 a_1467_8238# a_2307_8234# a_2515_8234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7080 a_52636_n8878# a_52632_n8701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7081 a_77821_5259# a_77608_5259# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7082 a_73000_12074# a_74093_12736# a_74048_12749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7083 gnd a_73252_4533# a_73044_4533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7084 a_25517_n11876# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7085 a_39385_n5058# a_40881_n5928# a_40832_n5738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7086 a_19163_n4466# a_19416_n4479# a_17716_n5233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7087 a_43771_3903# a_44392_3824# a_44600_3824# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7088 a_50134_n11058# a_51630_n11928# a_51581_n11738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7089 a_22935_11277# a_22722_11277# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7090 vdd d0 a_42137_n4485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7091 gnd a_74300_3761# a_74092_3761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7092 a_30124_n4285# a_31221_n4479# a_31172_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7093 a_66272_7557# a_65851_7557# a_65443_7124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7094 a_1729_n5863# a_1308_n5863# a_900_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7095 a_83704_13692# a_83961_13502# a_82261_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7096 a_36135_7546# a_35922_7546# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7097 a_66273_4590# a_67113_5265# a_67321_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7098 a_16602_n9613# a_16859_n9803# a_16257_n5742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7099 a_11347_4694# a_11968_4586# a_12176_4586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7100 a_76413_n5763# a_77034_n5871# a_77242_n5871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7101 a_57686_n5872# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7102 gnd d0 a_63334_8171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7103 a_25846_n5749# a_25476_n4423# a_24450_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7104 a_31176_n5234# a_31172_n5057# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7105 a_79778_n11882# a_79357_n11882# a_79684_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7106 a_69717_n8841# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7107 a_83967_n13443# a_84220_n13456# a_82520_n14210# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7108 a_5319_5273# a_5683_8186# a_5638_8199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7109 a_41884_n5240# a_42137_n5253# a_40836_n5915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7110 a_641_11614# a_1261_12120# a_1469_12120# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7111 a_3756_13562# a_3543_13562# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7112 a_54738_n11119# a_54738_n11514# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7113 a_52370_3274# a_52627_3084# a_51322_3278# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7114 a_26746_9142# a_26325_9142# a_25678_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7115 a_57751_6222# a_57381_7548# a_56355_6781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7116 a_44653_n5184# a_44440_n5184# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7117 a_71554_9787# a_73046_10541# a_72997_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7118 a_74305_n8024# a_74309_n8880# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7119 a_13225_14236# a_12804_14236# a_12177_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7120 vdd a_83961_12055# a_83753_12055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7121 gnd a_41875_7490# a_41667_7490# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7122 gnd d0 a_85007_6722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7123 a_22721_13565# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7124 a_7003_n14025# a_7260_n14215# a_6960_n12580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7125 vdd d0 a_52887_n14899# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7126 a_13062_n9755# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7127 a_33019_6212# a_33020_5598# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7128 a_76559_6104# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7129 gnd a_51579_3088# a_51371_3088# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7130 gnd a_31427_n11255# a_31219_n11255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7131 a_65703_n10318# a_66324_n10426# a_66532_n10426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7132 a_43771_5606# a_44391_6112# a_44599_6112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7133 a_12176_3818# a_13016_3814# a_13224_3814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7134 a_55309_14240# a_56149_14236# a_56357_14236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7135 a_44439_n13391# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7136 a_34896_8226# a_34475_8226# a_33848_8230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7137 gnd d1 a_62547_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7138 a_15360_9138# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7139 a_52372_10729# a_52629_10539# a_51324_10733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7140 a_45699_n9749# a_45486_n9749# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7141 a_33850_12112# a_34690_12787# a_34898_12787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7142 a_3754_7554# a_3541_7554# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7143 gnd d0 a_20465_n8897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7144 a_74048_14196# a_76153_14317# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7145 a_22982_n6706# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7146 a_79520_12109# a_80378_9136# a_80586_9136# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7147 a_77868_n12724# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7148 vdd d2 a_72066_n5242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7149 vdd a_82515_9768# a_82307_9768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7150 a_31170_n10297# a_31427_n10487# a_30122_n10293# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7151 a_34108_n9753# a_33687_n9753# a_33279_n9674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7152 a_38015_8368# a_39130_5205# a_39081_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7153 a_67114_12793# a_66901_12793# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7154 a_66535_n8832# a_67375_n8157# a_67583_n8157# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7155 a_52636_n8199# a_52889_n8212# a_51588_n8874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7156 a_11348_13128# a_11348_12872# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7157 gnd d2 a_39382_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7158 a_32239_n15022# a_33901_n14846# a_34109_n14846# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7159 a_69878_9142# a_70015_5271# a_70223_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7160 a_55147_n13397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7161 a_41880_n5742# a_42137_n5932# a_40832_n5738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7162 a_71509_5224# a_71762_5211# a_70439_8374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7163 gnd d2 a_72064_n11250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7164 a_2094_8234# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7165 a_30127_n14884# a_31220_n14222# a_31175_n14209# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7166 a_24027_n9751# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7167 gnd a_31169_12736# a_30961_12736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7168 a_44179_3824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7169 a_79520_12109# a_79099_12109# a_79421_12109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7170 vdd d2 a_28675_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7171 a_11757_9826# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7172 gnd a_31167_6728# a_30959_6728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7173 a_901_n6625# a_1522_n6704# a_1730_n6704# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7174 gnd a_62549_n7446# a_62341_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7175 a_55935_5261# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7176 vdd a_62288_12057# a_62080_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7177 a_20206_n12589# a_20210_n13445# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7178 a_76412_n14088# a_77033_n14167# a_77241_n14167# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7179 a_33640_8230# a_33427_8230# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7180 a_59159_5267# a_59050_5267# a_54212_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7181 a_62032_9280# a_63129_9086# a_63084_9099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7182 a_8451_n4283# a_9548_n4477# a_9499_n4287# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7183 a_9242_3776# a_9238_3953# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7184 vdd d1 a_19414_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7185 a_34691_9820# a_34478_9820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7186 gnd d1 a_73514_n7442# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7187 a_55099_6785# a_54886_6785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7188 a_77608_3812# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7189 vdd a_74562_n7446# a_74354_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7190 a_36549_n5874# a_36440_n5874# a_36648_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7191 vdd a_73252_4533# a_73044_4533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7192 gnd d0 a_41877_12730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7193 a_76413_n4857# a_77034_n4424# a_77242_n4424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7194 a_65705_n5107# a_65705_n5502# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7195 a_28416_3956# a_29912_3086# a_29863_3276# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7196 a_47784_9144# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7197 a_2354_n9749# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7198 a_23143_10598# a_22722_10598# a_22314_10165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7199 vdd d0 a_20465_n8218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7200 vdd d3 a_39338_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7201 a_23400_n11194# a_22979_n11194# a_22571_n11115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7202 a_13485_n5194# a_13064_n5194# a_12437_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7203 vdd a_74300_3761# a_74092_3761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7204 a_76152_4151# a_76773_4584# a_76981_4584# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7205 a_23141_5269# a_22720_5269# a_22312_4953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7206 gnd a_71806_12741# a_71598_12741# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7207 a_51321_7692# a_52418_7498# a_52369_7688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7208 a_19158_n14711# a_20255_n14905# a_20206_n14715# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7209 a_52633_n10472# a_52886_n10485# a_51581_n10291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7210 vdd d0 a_63334_8171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7211 a_30916_12070# a_30912_12247# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7212 a_18897_7686# a_19994_7492# a_19949_7505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7213 a_28637_n12759# a_28724_n11250# a_28675_n11060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7214 a_44033_n7020# a_44033_n7275# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7215 a_47298_n11874# a_46934_n13396# a_45908_n12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7216 vdd a_28632_11219# a_28424_11219# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7217 a_80165_9136# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7218 vdd d1 a_83959_7494# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7219 a_66112_n14161# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7220 vdd a_63595_n12779# a_63387_n12779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7221 a_71554_9787# a_73046_10541# a_73001_10554# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7222 gnd a_74560_n14901# a_74352_n14901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7223 a_47045_12236# a_46675_13562# a_45649_14242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7224 vdd d2 a_61100_n14221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7225 gnd d0 a_74562_n6767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7226 vdd d0 a_85007_6722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7227 a_36398_n7396# a_36185_n7396# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7228 vdd a_85008_5202# a_84800_5202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7229 a_44440_n5863# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7230 a_21631_n1621# a_21581_n1634# a_10595_n1632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7231 a_77035_n8838# a_76822_n8838# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7232 a_75301_n1457# a_81111_n5934# a_80846_n8847# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7233 a_13277_n3747# a_13064_n3747# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7234 a_67581_n14165# a_67160_n14165# a_66533_n14161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7235 a_22574_n8724# a_22571_n9412# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7236 a_39343_n6580# a_39435_n8215# a_39386_n8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7237 a_8449_n11738# a_8706_n11928# a_7002_n11058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7238 a_54740_n3408# a_63596_n3804# a_62295_n4466# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7239 a_78289_n14171# a_77868_n14171# a_77241_n14846# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7240 a_19945_7682# a_20202_7492# a_18897_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7241 a_55146_n11198# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7242 a_41621_9274# a_41622_8182# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7243 a_33902_n5192# a_33689_n5192# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7244 a_52633_n11919# a_52629_n11742# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7245 vdd d1 a_84220_n13456# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7246 a_11607_n14736# a_10566_n15020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7247 vdd d1 a_30381_n4475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7248 gnd d2 a_7001_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7249 a_2308_5267# a_2095_5267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7250 a_39383_n11066# a_40879_n11936# a_40830_n11746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7251 a_19947_13690# a_19951_12745# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7252 a_77035_n6712# a_76822_n6712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7253 gnd d0 a_74301_12736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7254 a_76562_9824# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7255 a_43773_9516# a_44394_9832# a_44602_9832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7256 gnd d1 a_62548_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7257 a_73257_n8699# a_74354_n8893# a_74305_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7258 a_40832_n4291# a_41929_n4485# a_41884_n4472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7259 a_63081_6058# a_63334_6045# a_62029_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7260 vdd a_9754_n9806# a_9546_n9806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7261 gnd a_20463_n12779# a_20255_n12779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7262 gnd d0 a_52888_n4477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7263 a_52375_13519# a_52628_13506# a_51323_13700# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7264 vdd d2 a_39382_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7265 a_22980_n14840# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7266 a_19157_n11744# a_19414_n11934# a_17710_n11064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7267 a_71812_n14204# a_73304_n13450# a_73255_n13260# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7268 a_33848_6783# a_34688_6779# a_34896_6779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7269 a_34948_n9757# a_34735_n9757# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7270 a_28681_n5229# a_30173_n4475# a_30124_n4285# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7271 a_57595_4581# a_57382_4581# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7272 a_71505_5401# a_71762_5211# a_70439_8374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7273 a_12805_9822# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7274 a_30129_n7429# a_31222_n6767# a_31173_n6577# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7275 a_67582_n5190# a_67161_n5190# a_66534_n5865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7276 a_11970_10594# a_11757_10594# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7277 a_27321_n5915# a_32426_n1647# a_21532_n1444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7278 a_76153_12870# a_76153_12475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7279 a_19162_n14888# a_20255_n14226# a_20210_n14213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7280 vdd a_31169_12736# a_30961_12736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7281 a_65444_5604# a_66064_6110# a_66272_6110# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7282 vdd d0 a_74561_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7283 a_33022_10159# a_33643_10592# a_33851_10592# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7284 vdd d0 a_85267_n10493# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7285 a_20207_n5061# a_20211_n5917# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7286 vdd a_81404_8178# a_81196_8178# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7287 a_22980_n12714# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7288 a_8450_n13258# a_9547_n13452# a_9498_n13262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7289 a_1522_n7383# a_1309_n7383# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7290 a_31174_n9795# a_31427_n9808# a_30126_n10470# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7291 a_79424_6220# a_79310_6101# a_79518_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7292 a_76980_7551# a_76559_7551# a_76151_7659# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7293 vdd a_19417_n8893# a_19209_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7294 a_2777_n5188# a_2356_n5188# a_1729_n5184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7295 vdd a_9494_7498# a_9286_7498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7296 a_1727_n11192# a_1306_n11192# a_898_n11113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7297 vdd d0 a_31429_n3800# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7298 a_31173_n8703# a_31430_n8893# a_30125_n8699# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7299 a_50136_n5050# a_50393_n5240# a_50098_n6749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7300 a_76819_n11879# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7301 gnd d0 a_31167_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7302 a_4168_n5866# a_3804_n7388# a_2778_n6708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7303 gnd d1 a_62288_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7304 a_22313_12876# a_22934_12797# a_23142_12797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7305 a_11346_7661# a_11346_7120# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7306 gnd a_50089_5213# a_49881_5213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7307 a_34477_12787# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7308 a_44860_n12712# a_45700_n12716# a_45908_n12716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7309 a_67114_14240# a_66901_14240# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7310 a_41620_12241# a_41625_11223# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7311 a_49026_n9607# a_50141_n12770# a_50096_n12757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7312 a_66533_n14840# a_66112_n14840# a_65704_n14732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7313 a_66064_8236# a_65851_8236# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7314 vdd d0 a_52886_n11253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7315 a_28421_12754# a_28674_12741# a_28379_11232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7316 a_65704_n13285# a_66325_n13393# a_66533_n13393# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7317 a_22932_8236# a_22719_8236# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7318 a_62294_n13441# a_63387_n12779# a_63342_n12766# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7319 a_7009_n8194# a_7262_n8207# a_6962_n6572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7320 vdd d0 a_41877_12730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7321 a_78083_n8163# a_77870_n8163# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7322 a_12176_5265# a_11755_5265# a_11347_4949# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7323 a_85014_n11248# a_85267_n11261# a_83966_n11923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7324 a_71771_n6751# a_71858_n5242# a_71813_n5229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7325 a_28416_3956# a_29912_3086# a_29867_3099# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7326 a_67321_5265# a_68560_4585# a_68711_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7327 a_65446_10961# a_66067_11277# a_66275_11277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7328 a_9502_n14886# a_9755_n14899# a_8450_n14705# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7329 a_19159_n5736# a_19416_n5926# a_17712_n5056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7330 gnd a_39381_3760# a_39173_3760# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7331 a_901_n6369# a_901_n6625# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7332 vdd d2 a_39380_6727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7333 a_33641_3137# a_33428_3137# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7334 a_36287_6101# a_35923_4579# a_34897_5259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7335 vdd a_71806_12741# a_71598_12741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7336 a_44602_9832# a_45442_9828# a_45650_9828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7337 a_73261_n8876# a_74354_n8214# a_74309_n8201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7338 a_77820_6779# a_77607_6779# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7339 gnd d0 a_9757_n7444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7340 a_30124_n5732# a_31221_n5926# a_31176_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7341 a_48465_n8839# a_48044_n8839# a_47397_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7342 a_11608_n4059# a_11608_n4314# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7343 a_44394_11279# a_44181_11279# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7344 a_17672_n12763# a_17759_n11254# a_17710_n11064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7345 a_65706_n8469# a_66327_n8153# a_66535_n8153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7346 a_22574_n6371# a_23194_n5865# a_23402_n5865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7347 a_33022_9253# a_33643_9145# a_33851_9145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7348 a_55567_n9751# a_55146_n9751# a_54738_n10067# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7349 a_84754_6735# a_84750_6912# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7350 a_30910_7686# a_30914_6741# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7351 a_40832_n5738# a_41089_n5928# a_39385_n5058# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7352 a_23142_12797# a_23982_12793# a_24190_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7353 a_83965_n7258# a_84222_n7448# a_82522_n8202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7354 a_72996_12251# a_74093_12057# a_74044_12247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7355 gnd a_63334_8171# a_63126_8171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7356 vdd a_73511_n10483# a_73303_n10483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7357 gnd a_5806_n5926# a_5598_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7358 a_1521_n3737# a_1308_n3737# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7359 a_60848_n5233# a_62340_n4479# a_62291_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7360 a_57753_12230# a_57383_13556# a_56357_12789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7361 a_44180_13567# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7362 vdd a_9496_12059# a_9288_12059# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7363 a_66534_n3739# a_67374_n3743# a_67582_n3743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7364 a_68819_n10431# a_68606_n10431# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7365 a_71553_12754# a_73045_13508# a_72996_13698# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7366 a_36396_n13404# a_36183_n13404# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7367 a_33851_11271# a_34691_11267# a_34899_11267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7368 vdd a_19157_10537# a_18949_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7369 vdd a_31428_n14901# a_31220_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7370 a_20210_n14892# a_20206_n14715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7371 gnd a_85007_6722# a_84799_6722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7372 gnd a_63337_10533# a_63129_10533# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7373 a_8456_n7427# a_9549_n6765# a_9500_n6575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7374 a_41619_5392# a_41623_4536# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7375 a_37454_9136# a_37033_9136# a_36386_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7376 a_14724_n4427# a_14511_n4427# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7377 a_79780_n5874# a_80638_n8847# a_80846_n8847# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7378 a_45441_14242# a_45228_14242# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7379 a_30913_10727# a_31170_10537# a_29865_10731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7380 a_76980_7551# a_77820_8226# a_78028_8226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7381 a_85010_n11750# a_85267_n11940# a_83962_n11746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7382 gnd a_49283_n9797# a_49075_n9797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7383 a_79097_6101# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7384 vdd d2 a_7001_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7385 a_40576_12068# a_41669_12730# a_41620_12920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7386 a_24243_n6710# a_24030_n6710# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7387 a_1729_n4416# a_2569_n3741# a_2777_n3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7388 a_66111_n9747# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7389 a_77033_n13399# a_76820_n13399# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7390 vdd d0 a_74301_12736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7391 a_63077_6235# a_63334_6045# a_62029_6239# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7392 a_27091_5271# a_26670_5271# a_26992_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7393 vdd d1 a_51838_n11928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7394 a_899_n13028# a_899_n13283# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7395 gnd d1 a_41088_n14903# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7396 a_12015_n14844# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7397 a_27307_8374# a_28422_5211# a_28373_5401# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7398 a_60847_n14208# a_62339_n13454# a_62290_n13264# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7399 a_9498_n14030# a_9755_n14220# a_8454_n14882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7400 a_9500_n8701# a_9757_n8891# a_8452_n8697# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7401 a_1306_n9745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7402 gnd a_82732_n6770# a_82524_n6770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7403 a_34110_n4424# a_33689_n4424# a_33281_n4857# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7404 a_12437_n5190# a_12016_n5190# a_11608_n5111# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7405 a_67322_12793# a_66901_12793# a_66274_12797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7406 a_85013_n6583# a_85270_n6773# a_83969_n7435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7407 a_55101_13561# a_54888_13561# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7408 a_76775_9145# a_76562_9145# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7409 gnd a_59646_n5932# a_59438_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7410 a_1048_14246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7411 a_65854_9830# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7412 gnd d0 a_9756_n3798# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7413 a_24240_n11198# a_24027_n11198# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7414 a_17670_n6578# a_17927_n6768# a_16606_n9790# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7415 gnd a_62286_6049# a_62078_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7416 a_1727_n11192# a_2567_n11196# a_2775_n11196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7417 a_44652_n14159# a_44439_n14159# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7418 a_82473_n12588# a_82565_n14223# a_82516_n14033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7419 a_44033_n8072# a_44654_n8151# a_44862_n8151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7420 a_25470_6107# a_25257_6107# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7421 a_63082_3091# a_63078_3268# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7422 a_82260_3773# a_82513_3760# a_82213_5395# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7423 gnd d0 a_42137_n4485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7424 a_19949_8184# a_19945_8361# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7425 a_8451_n5730# a_8708_n5920# a_7004_n5050# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7426 a_2096_12795# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7427 a_68346_7552# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7428 a_56197_n8161# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7429 a_55149_n7389# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7430 a_1469_13567# a_1048_13567# a_640_13134# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7431 a_44861_n5863# a_45701_n5188# a_45909_n5188# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7432 a_74304_n4289# a_74308_n5234# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7433 a_22721_12118# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7434 a_11967_8232# a_11754_8232# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7435 a_58105_n11880# a_57684_n11880# a_58006_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7436 a_48044_n8839# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7437 a_8451_n5730# a_9548_n5924# a_9503_n5911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7438 a_72999_4546# a_74092_5208# a_74043_5398# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7439 a_67112_8232# a_66899_8232# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7440 a_55934_6781# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7441 a_54887_4586# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7442 a_12229_n3743# a_12016_n3743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7443 vdd a_50089_5213# a_49881_5213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7444 a_13224_5261# a_12803_5261# a_12176_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7445 a_68711_6107# a_68602_6107# a_68810_6107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7446 a_79267_7546# a_79054_7546# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7447 a_28417_12931# a_28674_12741# a_28379_11232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7448 a_57857_n7394# a_57644_n7394# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7449 a_66327_n7385# a_66114_n7385# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7450 a_76152_5342# a_76152_4947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7451 a_7007_n14202# a_7260_n14215# a_6960_n12580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7452 a_8450_n14705# a_8707_n14895# a_7003_n14025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7453 a_52373_8190# a_52369_8367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7454 a_17450_6919# a_18946_6049# a_18901_6062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7455 a_55309_12114# a_54888_12114# a_54480_12222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7456 a_69878_9142# a_69457_9142# a_68812_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7457 vdd a_39381_3760# a_39173_3760# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7458 gnd d0 a_31170_9769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7459 a_54478_7120# a_55099_7553# a_55307_7553# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7460 a_79057_10587# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7461 vdd d0 a_52629_9092# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7462 a_33900_n11879# a_33687_n11879# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7463 a_22934_14244# a_22721_14244# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7464 a_23401_n13393# a_24241_n12718# a_24449_n12718# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7465 a_49874_6925# a_51370_6055# a_51321_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7466 a_68606_n10431# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7467 a_33642_12112# a_33429_12112# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7468 vdd a_39338_5205# a_39130_5205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7469 a_41620_14367# a_41877_14177# a_40576_13515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7470 a_55308_3139# a_56148_3814# a_56356_3814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7471 a_23140_6789# a_22719_6789# a_22311_6473# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7472 vdd a_52888_n4477# a_52680_n4477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7473 gnd a_31430_n8893# a_31222_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7474 a_13226_11269# a_14465_10589# a_14616_12111# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7475 a_66534_n5186# a_66113_n5186# a_65705_n5502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7476 a_11607_n12639# a_12228_n12718# a_12436_n12718# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7477 a_31174_n10474# a_31427_n10487# a_30122_n10293# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7478 vdd a_63334_8171# a_63126_8171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7479 a_31176_n5913# a_31172_n5736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7480 a_46976_n11874# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7481 a_33282_n7283# a_33282_n7824# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7482 a_43771_3253# a_44392_3145# a_44600_3145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7483 a_37714_n8847# a_37293_n8847# a_36646_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7484 a_898_n11763# a_1519_n11871# a_1727_n11871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7485 a_80832_5265# a_81196_8178# a_81151_8191# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7486 gnd a_74300_3082# a_74092_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7487 a_34897_5259# a_34476_5259# a_33849_4584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7488 a_79314_n10437# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7489 a_22311_6868# a_22311_6473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7490 a_11606_n10322# a_11606_n10863# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7491 a_1729_n5184# a_1308_n5184# a_900_n5105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7492 a_43231_n1412# a_43488_n1602# a_3053_n1225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7493 vdd d0 a_63594_n10491# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7494 a_76413_n5113# a_77034_n5192# a_77242_n5192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7495 vdd a_63337_10533# a_63129_10533# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7496 vdd a_85007_6722# a_84799_6722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7497 a_30125_n8699# a_30382_n8889# a_28678_n8019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7498 a_8189_7692# a_9286_7498# a_9241_7511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7499 a_40576_12068# a_41669_12730# a_41624_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7500 a_33279_n10324# a_33900_n10432# a_34108_n10432# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7501 a_8194_4548# a_8447_4535# a_6747_3781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7502 a_60587_3775# a_62079_4529# a_62034_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7503 a_25581_12115# a_25217_10593# a_24191_11273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7504 a_74302_n11065# a_74306_n11921# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7505 a_1307_n12712# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7506 a_31174_n9795# a_31170_n9618# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7507 a_65854_11277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7508 a_10971_986# a_10758_986# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7509 a_66326_n3739# a_66113_n3739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7510 gnd a_19156_13504# a_18948_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7511 vdd d3 a_61059_n6768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7512 gnd d0 a_85007_6043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7513 gnd d1 a_19414_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7514 a_65706_n7818# a_65706_n8074# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7515 a_27307_8374# a_28422_5211# a_28377_5224# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7516 a_13223_8228# a_14462_7548# a_14619_6222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7517 a_2307_6787# a_2094_6787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7518 a_9504_n7431# a_9500_n7254# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7519 a_18902_3095# a_19995_3757# a_19950_3770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7520 a_77240_n9753# a_78080_n9757# a_78288_n9757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7521 vdd d0 a_52888_n5924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7522 a_2095_5267# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7523 a_35924_13554# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7524 a_22572_n14082# a_23193_n14161# a_23401_n14161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7525 gnd a_74562_n7446# a_74354_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7526 a_23142_13565# a_23982_14240# a_24190_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7527 a_2776_n12716# a_2355_n12716# a_1728_n13391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7528 a_22981_n5865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7529 a_84755_4536# a_84751_4713# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7530 a_9244_10552# a_9497_10539# a_8192_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7531 a_76154_10159# a_76154_9903# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7532 a_34111_n8838# a_34951_n8163# a_35159_n8163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7533 a_60544_5220# a_60797_5207# a_59474_8370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7534 vdd a_70956_n9799# a_70748_n9799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7535 a_24450_n3743# a_25689_n4423# a_25846_n5749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7536 a_23769_12793# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7537 gnd d0 a_20465_n8218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7538 a_84756_14190# a_85009_14177# a_83708_13515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7539 a_82256_3950# a_82513_3760# a_82213_5395# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7540 a_62034_4542# a_63127_5204# a_63078_5394# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7541 a_57382_4581# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7542 a_9499_n4287# a_9503_n5232# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7543 a_76775_11271# a_76562_11271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7544 vdd a_31430_n8214# a_31222_n8214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7545 a_78290_n5196# a_79529_n4429# a_79686_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7546 a_33021_13126# a_33642_13559# a_33850_13559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7547 a_32753_984# a_32644_984# a_21717_973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7548 gnd d2 a_82515_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7549 vdd d1 a_62289_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7550 a_13484_n12722# a_13063_n12722# a_12436_n13397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7551 a_22571_n11115# a_22571_n11510# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7552 a_33280_n14483# a_33901_n14167# a_34109_n14167# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7553 a_19946_3947# a_20203_3757# a_18902_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7554 a_76822_n7391# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7555 a_34478_11267# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7556 a_77241_n12720# a_76820_n12720# a_76412_n13036# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7557 a_4267_n5866# a_5125_n8839# a_5333_n8839# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7558 a_41880_n5063# a_42137_n5253# a_40836_n5915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7559 gnd d1 a_40829_12055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7560 gnd a_63597_n8897# a_63389_n8897# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7561 a_66273_5269# a_65852_5269# a_65444_5348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7562 gnd a_63595_n12779# a_63387_n12779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7563 a_52374_4544# a_52627_4531# a_51322_4725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7564 gnd d0 a_20205_9765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7565 gnd a_31169_12057# a_30961_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7566 a_41883_n14894# a_41879_n14717# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7567 a_44179_3145# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7568 a_65444_4157# a_65444_3901# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7569 a_41618_8359# a_41622_7503# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7570 a_28676_n14027# a_30172_n14897# a_30123_n14707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7571 a_11757_9147# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7572 a_25938_n11876# a_25517_n11876# a_25839_n11876# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7573 a_21631_n1621# a_21581_n1634# a_21532_n1444# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7574 gnd a_31167_6049# a_30959_6049# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7575 a_4171_n11755# a_4057_n11874# a_4265_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7576 gnd a_60840_3762# a_60632_3762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7577 a_75301_n1457# a_81111_n5934# a_81062_n5744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7578 a_85017_n7439# a_85013_n7262# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7579 a_85011_n14717# a_85268_n14907# a_83963_n14713# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7580 gnd a_30121_13508# a_29913_13508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7581 a_44030_n11113# a_44030_n11508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7582 a_14510_n13402# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7583 a_639_3253# a_641_3154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7584 a_76411_n11121# a_76411_n11516# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7585 a_5418_5273# a_4997_5273# a_5319_5273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7586 a_8453_n11915# a_8706_n11928# a_7002_n11058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7587 a_49874_6925# a_51370_6055# a_51325_6068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7588 a_66899_8232# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7589 a_41622_7503# a_41875_7490# a_40570_7684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7590 a_12175_6785# a_11754_6785# a_11346_6469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7591 a_62293_n10474# a_63386_n9812# a_63337_n9622# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7592 a_20211_n4470# a_20464_n4483# a_19159_n4289# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7593 a_25579_6107# a_25215_4585# a_24189_5265# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7594 a_1470_10600# a_1049_10600# a_641_10708# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7595 a_5634_8376# a_6749_5213# a_6700_5403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7596 a_76151_7118# a_76151_6862# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7597 gnd a_52887_n12773# a_52679_n12773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7598 gnd d1 a_84220_n13456# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7599 gnd d1 a_30381_n4475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7600 a_58705_9138# a_58492_9138# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7601 a_55360_n13397# a_55147_n13397# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7602 a_898_n10857# a_1519_n10424# a_1727_n10424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7603 a_55099_6106# a_54886_6106# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7604 a_41880_n4295# a_41884_n5240# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7605 a_34111_n6712# a_33690_n6712# a_33282_n7028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7606 a_36184_n4429# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7607 a_30916_12749# a_30912_12926# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7608 a_40832_n4291# a_41929_n4485# a_41880_n4295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7609 gnd d0 a_41877_12051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7610 a_55934_8228# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7611 a_48342_5273# a_48129_5273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7612 a_34108_n11879# a_33687_n11879# a_33280_n12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7613 a_3797_6109# a_3584_6109# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7614 vdd d2 a_7260_n14215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7615 a_19161_n11921# a_19414_n11934# a_17710_n11064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7616 a_45488_n5188# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7617 a_52371_13696# a_52375_12751# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7618 a_9243_12072# a_9239_12249# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7619 vdd a_74300_3082# a_74092_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7620 a_11348_13128# a_11969_13561# a_12177_13561# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7621 a_45907_n9749# a_47146_n10429# a_47303_n11755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7622 a_8196_10556# a_9289_11218# a_9244_11231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7623 gnd a_85267_n10493# a_85059_n10493# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7624 a_76980_6104# a_76559_6104# a_76152_5598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7625 a_78028_8226# a_79267_7546# a_79424_6220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7626 gnd d0 a_42138_n6773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7627 a_60844_n5056# a_62340_n5926# a_62295_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7628 a_36289_12109# a_35925_10587# a_34899_9820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7629 a_19162_n14888# a_20255_n14226# a_20206_n14036# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7630 gnd d0 a_74561_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7631 a_25846_n5749# a_25732_n5868# a_25940_n5868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7632 a_11606_n10863# a_12227_n10430# a_12435_n10430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7633 a_56617_n3747# a_57856_n4427# a_58013_n5753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7634 a_59159_5267# a_59523_8180# a_59474_8370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7635 a_76152_4947# a_76152_4692# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7636 a_20205_n9622# a_20462_n9812# a_19161_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7637 gnd a_85009_12730# a_84801_12730# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7638 a_76821_n3745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7639 a_35157_n14171# a_34736_n14171# a_34109_n14167# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7640 a_8190_4725# a_8447_4535# a_6747_3781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7641 vdd a_63597_n8218# a_63389_n8218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7642 a_3757_10595# a_3544_10595# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7643 a_14973_n11880# a_15833_n8845# a_16041_n8845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7644 a_78081_n12724# a_77868_n12724# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7645 a_39341_n12588# a_39598_n12778# a_38275_n9615# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7646 gnd a_74560_n14222# a_74352_n14222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7647 a_3543_13562# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7648 gnd a_9496_12738# a_9288_12738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7649 a_54480_12872# a_55101_12793# a_55309_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7650 a_45487_n14163# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7651 a_62035_12070# a_63128_12732# a_63079_12922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7652 a_11179_986# a_21608_973# a_21816_973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7653 vdd d0 a_31427_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7654 a_639_3508# a_1260_3824# a_1468_3824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7655 vdd d0 a_85007_6043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7656 a_63340_n7260# a_63597_n7450# a_62292_n7256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7657 a_50140_n5227# a_50393_n5240# a_50098_n6749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7658 a_44440_n5184# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7659 a_67323_11273# a_66902_11273# a_66275_10598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7660 a_68718_12234# a_68604_12115# a_68812_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7661 a_84753_10721# a_84757_9776# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7662 gnd a_5891_8186# a_5683_8186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7663 a_77035_n8159# a_76822_n8159# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7664 a_22722_10598# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7665 vdd d1 a_73514_n7442# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7666 a_18901_6062# a_19154_6049# a_17450_6919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7667 a_49026_n9607# a_50141_n12770# a_50092_n12580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7668 a_15620_n8845# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7669 a_77034_n5871# a_76821_n5871# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7670 a_23143_9151# a_22722_9151# a_22314_9259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7671 a_62294_n13441# a_63387_n12779# a_63338_n12589# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7672 vdd a_30379_n11930# a_30171_n11930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7673 a_22979_n11873# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7674 a_46931_12117# a_46718_12117# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7675 a_76981_4584# a_76560_4584# a_76152_4151# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7676 gnd d0 a_85010_9763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7677 vdd a_38532_n9805# a_38324_n9805# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7678 a_44600_3824# a_44179_3824# a_43771_3903# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7679 a_19163_n5913# a_19416_n5926# a_17712_n5056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7680 a_56195_n14169# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7681 a_2097_11275# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7682 a_35158_n5196# a_34737_n5196# a_34110_n5871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7683 gnd d0 a_74301_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7684 a_63084_10546# a_63080_10723# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7685 a_76562_9145# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7686 a_56148_3814# a_55935_3814# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7687 a_43770_8573# a_44394_9153# a_44602_9153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7688 a_73261_n8876# a_74354_n8214# a_74305_n8024# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7689 vdd a_52889_n6765# a_52681_n6765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7690 a_22312_4698# a_22312_4157# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7691 a_31174_n11242# a_31170_n11065# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7692 a_30124_n5732# a_31221_n5926# a_31172_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7693 a_14614_6103# a_14250_4581# a_13224_3814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7694 a_9241_8190# a_9494_8177# a_8193_7515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7695 a_33643_10592# a_33430_10592# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7696 vdd d1 a_40829_12055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7697 a_83967_n14890# a_84220_n14903# a_82516_n14033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7698 a_22933_5269# a_22720_5269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7699 a_55307_8232# a_54886_8232# a_54478_8311# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7700 a_79684_n11763# a_79570_n11882# a_79778_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7701 a_63338_n12589# a_63342_n13445# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7702 a_40836_n5915# a_41089_n5928# a_39385_n5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7703 gnd a_39382_12735# a_39174_12735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7704 a_52370_4721# a_52627_4531# a_51322_4725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7705 vdd d0 a_20205_9765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7706 a_23142_14244# a_22721_14244# a_22313_14323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7707 a_79315_n13404# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7708 a_83969_n7435# a_84222_n7448# a_82522_n8202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7709 vdd d0 a_74561_n5247# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7710 vdd a_9756_n4477# a_9548_n4477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7711 a_11754_8232# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7712 a_59738_n9790# a_60851_n6768# a_60806_n6755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7713 vdd a_83961_13502# a_83753_13502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7714 a_67372_n11198# a_67159_n11198# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7715 vdd a_60840_3762# a_60632_3762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7716 a_65445_14323# a_66066_14244# a_66274_14244# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7717 gnd d4 a_81404_8178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7718 a_17717_n8200# a_19209_n7446# a_19164_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7719 a_83965_n7258# a_85062_n7452# a_85013_n7262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7720 a_77240_n10432# a_76819_n10432# a_76411_n10324# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7721 a_79054_7546# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7722 a_67580_n9751# a_67159_n9751# a_66532_n10426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7723 a_47146_n10429# a_46933_n10429# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7724 a_77867_n9757# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7725 gnd a_51579_4535# a_51371_4535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7726 a_23769_14240# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7727 a_76153_12220# a_76774_12112# a_76982_12112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7728 vdd a_61099_n11254# a_60891_n11254# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7729 a_5634_8376# a_6749_5213# a_6704_5226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7730 a_44393_14246# a_44180_14246# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7731 a_22574_n6627# a_22574_n7022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7732 a_23403_n7385# a_22982_n7385# a_22574_n7277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7733 a_1308_n5863# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7734 a_85014_n11927# a_85267_n11940# a_83962_n11746# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7735 a_898_n10316# a_898_n10857# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7736 a_44599_7559# a_44178_7559# a_43770_7126# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7737 a_76411_n9674# a_77032_n9753# a_77240_n9753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7738 gnd d1 a_62287_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7739 a_66067_9830# a_65854_9830# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7740 a_25476_n4423# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7741 a_12435_n11877# a_12014_n11877# a_11606_n11769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7742 a_66533_n14161# a_66112_n14161# a_65704_n14082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7743 vdd d0 a_85269_n4485# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7744 a_55101_12114# a_54888_12114# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7745 a_11609_n8078# a_11609_n8473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7746 a_1046_6112# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7747 a_63079_14369# a_63336_14179# a_62035_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7748 a_28417_12931# a_29913_12061# a_29864_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7749 vdd d0 a_41877_12051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7750 gnd d1 a_51838_n11928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7751 a_59734_n9613# a_59991_n9803# a_59389_n5742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7752 a_31170_n11744# a_31427_n11934# a_30122_n11740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7753 a_65705_n4851# a_65705_n5107# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7754 a_74047_4542# a_74300_4529# a_72995_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7755 a_9502_n14207# a_9755_n14220# a_8454_n14882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7756 a_13225_12789# a_12804_12789# a_12177_12114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7757 a_74302_n9618# a_74306_n10474# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7758 a_54741_n7281# a_55362_n7389# a_55570_n7389# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7759 a_55102_9826# a_54889_9826# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7760 a_55147_n14844# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7761 a_30128_n5909# a_31221_n5247# a_31176_n5234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7762 a_39125_12925# a_40621_12055# a_40572_12245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7763 a_4912_n8839# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7764 a_17674_n6755# a_17927_n6768# a_16606_n9790# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7765 a_76981_5263# a_77821_5259# a_78029_5259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7766 a_59159_5267# a_59523_8180# a_59478_8193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7767 vdd a_85009_12730# a_84801_12730# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7768 a_22573_n5502# a_23194_n5186# a_23402_n5186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7769 a_34896_6779# a_34475_6779# a_33848_6104# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7770 vdd a_85269_n3806# a_85061_n3806# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7771 gnd d3 a_28890_n12772# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7772 a_55567_n11198# a_56407_n11202# a_56615_n11202# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7773 gnd a_62549_n8893# a_62341_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7774 a_8455_n5907# a_8708_n5920# a_7004_n5050# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7775 a_8195_13523# a_9288_14185# a_9239_14375# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7776 a_8450_n13258# a_9547_n13452# a_9502_n13439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7777 a_85013_n6583# a_85017_n7439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7778 vdd d2 a_61102_n8213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7779 vdd a_39643_n8215# a_39435_n8215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7780 a_34737_n5196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7781 a_62035_12070# a_63128_12732# a_63083_12745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7782 a_71550_9964# a_73046_9094# a_72997_9284# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7783 vdd a_42135_n10493# a_41927_n10493# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7784 a_33901_n13399# a_33688_n13399# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7785 a_47040_12117# a_46676_10595# a_45650_11275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7786 a_54311_986# a_53890_986# a_48550_5273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7787 a_8451_n5730# a_9548_n5924# a_9499_n5734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7788 a_63083_14192# a_63079_14369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7789 vdd a_5891_8186# a_5683_8186# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7790 gnd a_16859_n9803# a_16651_n9803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7791 a_1047_4592# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7792 vdd d1 a_19414_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7793 a_54739_n12639# a_55360_n12718# a_55568_n12718# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7794 a_83968_n4468# a_85061_n3806# a_85012_n3616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7795 a_55569_n4422# a_55148_n4422# a_54740_n4855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7796 a_25586_12234# a_25216_13560# a_24190_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7797 a_74049_9103# a_74045_9280# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7798 a_66324_n11873# a_66111_n11873# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7799 a_54478_6214# a_55099_6106# a_55307_6106# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7800 a_52370_4721# a_52374_3776# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7801 a_16342_8370# a_17457_5207# a_17408_5397# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7802 a_45702_n8155# a_45489_n8155# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7803 a_28422_9787# a_28675_9774# a_28375_11409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7804 a_77240_n9753# a_76819_n9753# a_76411_n9674# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7805 gnd a_85007_6043# a_84799_6043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7806 a_57383_13556# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7807 vdd a_27479_n5928# a_27271_n5928# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7808 a_52632_n8701# a_52633_n9793# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7809 a_55569_n5190# a_56409_n5194# a_56617_n5194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7810 a_20212_n6758# a_20465_n6771# a_19164_n7433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7811 a_23402_n3739# a_22981_n3739# a_22573_n3660# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7812 a_14713_6103# a_14292_6103# a_14619_6222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7813 vdd d0 a_85010_9763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7814 a_85010_n11071# a_85267_n11261# a_83966_n11923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7815 a_2094_6787# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7816 a_40572_12245# a_41669_12051# a_41620_12241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7817 a_33850_12791# a_33429_12791# a_33021_12870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7818 a_28420_3779# a_29912_4533# a_29863_4723# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7819 a_19947_14369# a_19951_13513# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7820 a_68347_4585# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7821 vdd a_51839_n13448# a_51631_n13448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7822 a_12437_n5869# a_12016_n5869# a_11608_n5761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7823 a_29867_3099# a_30960_3761# a_30911_3951# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7824 a_63077_7682# a_63081_6737# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7825 a_899_n13824# a_1520_n13391# a_1728_n13391# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7826 a_24242_n3743# a_24029_n3743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7827 a_11968_5265# a_11755_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7828 a_39085_5218# a_39172_6727# a_39127_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7829 a_51326_4548# a_52419_5210# a_52370_5400# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7830 a_67113_5265# a_66900_5265# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7831 a_11756_13561# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7832 a_45229_9828# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7833 a_55570_n7389# a_55149_n7389# a_54741_n7281# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7834 a_12015_n14165# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7835 a_1467_6112# a_1046_6112# a_639_5606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7836 a_52633_n11919# a_52886_n11932# a_51581_n11738# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7837 a_44030_n9410# a_44030_n9666# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7838 a_9500_n8022# a_9757_n8212# a_8456_n8874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7839 a_63082_3770# a_63078_3947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7840 a_79268_4579# a_79055_4579# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7841 vdd a_20465_n8897# a_20257_n8897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7842 a_25519_n5868# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7843 a_52376_10552# a_52629_10539# a_51324_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7844 a_66113_n4418# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7845 a_54480_13924# a_55101_14240# a_55309_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7846 a_24028_n14165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7847 a_44033_n8722# a_44654_n8830# a_44862_n8830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7848 gnd a_52888_n4477# a_52680_n4477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7849 vdd a_39382_12735# a_39174_12735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7850 a_67162_n6710# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7851 gnd d1 a_83960_3080# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7852 vdd a_72065_n14217# a_71857_n14217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7853 a_79681_n5874# a_79317_n7396# a_78291_n8163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7854 a_1261_14246# a_1048_14246# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7855 a_45908_n12716# a_47147_n13396# a_47298_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7856 a_51584_n7250# a_51841_n7440# a_50141_n8194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7857 a_37454_9136# a_37591_5265# a_32753_984# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7858 a_6960_n12580# a_7217_n12770# a_5894_n9607# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7859 gnd a_82515_9768# a_82307_9768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7860 a_63344_n8205# a_63340_n8028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7861 a_56617_n3747# a_56196_n3747# a_55569_n4422# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7862 a_54479_4694# a_55100_4586# a_55308_4586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7863 a_54888_12793# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7864 gnd d0 a_85267_n11261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7865 a_66274_13565# a_65853_13565# a_65445_13673# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7866 a_51584_n7250# a_52681_n7444# a_52636_n7431# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7867 a_65851_7557# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7868 a_44391_6112# a_44178_6112# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7869 a_47043_6228# a_46673_7554# a_45647_6787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7870 a_76413_n4316# a_76413_n4857# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7871 vdd a_51579_4535# a_51371_4535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7872 gnd a_20205_9765# a_19997_9765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7873 a_44033_n7020# a_44654_n6704# a_44862_n6704# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7874 a_14767_n5872# a_14554_n5872# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7875 a_33281_n4857# a_33281_n5113# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7876 a_55361_n4422# a_55148_n4422# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7877 a_18903_13517# a_19996_14179# a_19951_14192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7878 a_26798_n8841# a_26585_n8841# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7879 a_13064_n5194# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7880 a_33020_5342# a_33641_5263# a_33849_5263# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7881 a_30129_n8876# a_30382_n8889# a_28678_n8019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7882 a_8455_n5907# a_9548_n5245# a_9503_n5232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7883 a_640_12878# a_640_12483# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7884 a_56197_n6714# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7885 a_25474_n10431# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7886 a_1468_4592# a_1047_4592# a_639_4159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7887 a_20210_n12766# a_20206_n12589# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7888 gnd a_62288_12057# a_62080_12057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7889 gnd d3 a_61059_n6768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7890 a_30915_5221# a_31168_5208# a_29867_4546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7891 a_24188_8232# a_23767_8232# a_23140_8236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7892 gnd d0 a_52628_14185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7893 a_28417_12931# a_29913_12061# a_29868_12074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7894 a_9238_3953# a_9242_3097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7895 a_33851_9145# a_34691_9820# a_34899_9820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7896 a_78028_8226# a_77607_8226# a_76980_8230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7897 vdd a_30380_n14897# a_30172_n14897# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7898 vdd a_72024_n6764# a_71816_n6764# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7899 a_9502_n14886# a_9498_n14709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7900 a_2309_14242# a_2096_14242# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7901 a_58492_9138# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7902 a_67375_n6710# a_67162_n6710# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7903 gnd a_6151_n9797# a_5943_n9797# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7904 gnd d0 a_52888_n5924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7905 a_68812_12115# a_69670_9142# a_69878_9142# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7906 a_901_n7020# a_901_n7275# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7907 a_71808_n14027# a_73304_n14897# a_73255_n14707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7908 a_33900_n11200# a_33687_n11200# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7909 a_44599_7559# a_45439_8234# a_45647_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7910 a_1520_n14838# a_1307_n14838# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7911 a_26883_5271# a_26670_5271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7912 vdd a_59646_n5932# a_59438_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7913 a_39125_12925# a_40621_12055# a_40576_12068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7914 a_28677_n5052# a_30173_n5922# a_30124_n5732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7915 a_44392_4592# a_44179_4592# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7916 a_60546_11228# a_60799_11215# a_59478_8193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7917 a_3584_6109# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7918 a_79530_n7396# a_79317_n7396# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7919 a_11609_n6631# a_12230_n6710# a_12438_n6710# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7920 a_11609_n6375# a_11609_n6631# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7921 a_2516_3820# a_2095_3820# a_1468_3145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7922 vdd d0 a_85267_n11940# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7923 a_30910_8365# a_30914_7509# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7924 a_82473_n12588# a_82565_n14223# a_82520_n14210# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7925 a_8195_13523# a_9288_14185# a_9243_14198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7926 a_4171_n11755# a_3801_n10429# a_2775_n9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7927 a_41625_11223# a_41878_11210# a_40577_10548# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7928 a_66324_n10426# a_66111_n10426# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7929 gnd a_31430_n8214# a_31222_n8214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7930 a_20208_n8707# a_20209_n9799# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7931 a_59050_5267# a_58837_5267# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7932 a_65853_14244# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7933 a_63342_n14892# a_63338_n14715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7934 a_1520_n12712# a_1307_n12712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7935 gnd d4 a_81664_n9805# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7936 vdd a_9757_n6765# a_9549_n6765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7937 a_12178_10594# a_11757_10594# a_11349_10161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7938 a_76773_5263# a_76560_5263# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7939 a_898_n11113# a_1519_n11192# a_1727_n11192# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7940 a_19949_6058# a_19945_6235# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7941 a_76561_12112# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7942 a_54889_9826# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7943 gnd a_28632_11219# a_28424_11219# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7944 a_45440_3820# a_45227_3820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7945 a_37378_5265# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7946 a_44181_10600# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7947 a_76819_n9753# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7948 a_28418_9964# a_28675_9774# a_28375_11409# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7949 vdd a_85007_6043# a_84799_6043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7950 a_47147_n13396# a_46934_n13396# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7951 a_68864_n5868# a_68651_n5868# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7952 a_83967_n13443# a_85060_n12781# a_85011_n12591# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7953 a_23401_n12714# a_22980_n12714# a_22572_n13030# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7954 a_13016_5261# a_12803_5261# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7955 a_40572_12245# a_41669_12051# a_41624_12064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7956 a_77823_9820# a_77610_9820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7957 gnd a_42138_n7452# a_41930_n7452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7958 a_28420_3779# a_29912_4533# a_29867_4546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7959 a_34109_n13399# a_33688_n13399# a_33280_n13291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7960 a_54738_n10863# a_55359_n10430# a_55567_n10430# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7961 a_22574_n8469# a_22574_n8724# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7962 a_29867_3099# a_30960_3761# a_30915_3774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7963 a_22572_n14732# a_23193_n14840# a_23401_n14840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7964 a_58965_n8845# a_58752_n8845# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7965 a_33641_4584# a_33428_4584# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7966 a_51326_4548# a_52419_5210# a_52374_5223# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7967 a_45650_9828# a_45229_9828# a_44602_9832# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7968 a_44862_n7383# a_44441_n7383# a_44033_n7816# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7969 a_52373_6064# a_52369_6241# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7970 a_2356_n5188# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7971 a_76154_10159# a_76775_10592# a_76983_10592# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7972 gnd d0 a_9757_n8891# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7973 vdd d0 a_9497_11218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7974 a_27311_8197# a_27564_8184# a_26992_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7975 a_18898_3272# a_19995_3078# a_19950_3091# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7976 a_11607_n14481# a_11607_n14736# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7977 a_34689_3812# a_34476_3812# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7978 vdd d0 a_52888_n5245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7979 a_22981_n5186# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7980 vdd d1 a_83960_3080# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7981 a_11348_12222# a_11969_12114# a_12177_12114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7982 gnd d3 a_39340_11213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7983 a_45910_n8155# a_47149_n7388# a_47300_n5866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7984 vdd d0 a_52626_8177# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7985 a_55102_10594# a_54889_10594# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7986 a_40574_7507# a_41667_8169# a_41622_8182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7987 a_80638_n8847# a_80425_n8847# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7988 gnd a_9755_n12773# a_9547_n12773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7989 a_22572_n13030# a_23193_n12714# a_23401_n12714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7990 gnd d2 a_7260_n14215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7991 a_33642_13559# a_33429_13559# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7992 a_22932_6789# a_22719_6789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7993 a_1470_9832# a_1049_9832# a_641_9516# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7994 vdd a_73511_n11930# a_73303_n11930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7995 a_22720_5269# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7996 a_22573_n3404# a_31172_n3610# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7997 vdd a_20205_9765# a_19997_9765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7998 a_60844_n5056# a_62340_n5926# a_62291_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7999 gnd a_73254_10541# a_73046_10541# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8000 a_76982_13559# a_76561_13559# a_76153_13126# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8001 a_79099_12109# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8002 a_30126_n10470# a_30379_n10483# a_28679_n11237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8003 a_68976_n11757# a_68606_n10431# a_67580_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8004 a_19946_3268# a_20203_3078# a_18898_3272# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8005 a_28635_n6574# a_28892_n6764# a_27571_n9786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8006 gnd a_81404_8178# a_81196_8178# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8007 a_9239_12928# a_9496_12738# a_8195_12076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8008 gnd a_63597_n8218# a_63389_n8218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8009 a_74305_n6577# a_74309_n7433# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8010 a_54479_5344# a_54479_4949# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8011 a_639_3903# a_639_3508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8012 a_49881_9789# a_51373_10543# a_51324_10733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8013 gnd a_72067_n8209# a_71859_n8209# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8014 a_47305_n5747# a_46935_n4421# a_45909_n3741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8015 a_19951_13513# a_19947_13690# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8016 a_39345_n12765# a_39598_n12778# a_38275_n9615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8017 gnd d0 a_20205_9086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8018 vdd d0 a_52628_14185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8019 a_77033_n14846# a_76820_n14846# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8020 gnd d2 a_50131_6735# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8021 gnd d0 a_31427_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8022 a_72998_6066# a_73251_6053# a_71547_6923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8023 a_66111_n10426# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8024 a_63344_n7437# a_63597_n7450# a_62292_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8025 a_63077_7682# a_63334_7492# a_62029_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8026 a_57644_n7394# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8027 a_44033_n8467# a_44033_n8722# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8028 a_85012_n5742# a_85017_n6760# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8029 gnd a_42137_n3806# a_41929_n3806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8030 a_14249_7548# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8031 a_44859_n11871# a_44438_n11871# a_44031_n12377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8032 a_41878_n9624# a_42135_n9814# a_40834_n10476# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8033 a_60843_n14031# a_62339_n14901# a_62290_n14711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8034 a_79684_n11763# a_79314_n10437# a_78288_n9757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8035 a_44861_n3737# a_44440_n3737# a_44032_n4053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8036 a_11346_6469# a_11346_6214# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8037 a_54888_14240# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8038 a_22311_7920# a_22932_8236# a_23140_8236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8039 gnd a_30379_n11930# a_30171_n11930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8040 a_12177_12114# a_13017_12789# a_13225_12789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8041 gnd a_28672_6733# a_28464_6733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8042 a_34948_n11204# a_34735_n11204# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8043 a_66274_12797# a_67114_12793# a_67322_12793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8044 a_60542_11405# a_60799_11215# a_59478_8193# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8045 vdd d2 a_82772_n11256# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8046 gnd d1 a_8446_7502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8047 a_33688_n12720# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8048 a_9243_12751# a_9239_12928# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8049 a_45701_n3741# a_45488_n3741# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8050 a_12230_n7389# a_12017_n7389# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8051 gnd d1 a_8449_10543# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8052 a_41621_11400# a_41878_11210# a_40577_10548# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8053 a_66114_n6706# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8054 a_45441_12795# a_45228_12795# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8055 gnd d2 a_39380_6727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8056 gnd a_52889_n6765# a_52681_n6765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8057 a_1728_n12712# a_1307_n12712# a_899_n13028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8058 gnd d0 a_42137_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8059 a_76980_6783# a_77820_6779# a_78028_6779# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8060 a_55937_9822# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8061 a_34108_n11200# a_33687_n11200# a_33279_n11516# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8062 a_638_8573# a_638_8317# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8063 a_55567_n11877# a_55146_n11877# a_54738_n11769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8064 a_55149_n8836# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8065 gnd d0 a_9495_3763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8066 a_60585_9960# a_62081_9090# a_62036_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8067 a_43150_941# a_43041_941# a_3058_n1106# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8068 vdd d0 a_31167_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8069 a_34108_n11200# a_34948_n11204# a_35156_n11204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8070 gnd a_74301_14183# a_74093_14183# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8071 a_57426_12111# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8072 a_84750_6912# a_84754_6056# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8073 vdd d1 a_62288_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8074 a_63340_n7260# a_63344_n8205# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8075 a_21717_973# a_32431_984# a_27091_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8076 a_49881_9789# a_50134_9776# a_49834_11411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8077 gnd d0 a_74561_n5247# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8078 gnd a_9756_n4477# a_9548_n4477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8079 a_76154_9508# a_76154_9253# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8080 gnd a_85009_12051# a_84801_12051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8081 a_33851_11271# a_33430_11271# a_33022_10955# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8082 a_1048_12799# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8083 a_66327_n8832# a_66114_n8832# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8084 a_59738_n9790# a_60851_n6768# a_60802_n6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8085 a_40830_n10299# a_41927_n10493# a_41878_n10303# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8086 a_17717_n8200# a_19209_n7446# a_19160_n7256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8087 a_55149_n6710# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8088 a_17714_n11241# a_19206_n10487# a_19161_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8089 a_19948_10723# a_19952_9778# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8090 a_41883_n12768# a_41879_n12591# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8091 vdd a_17969_n5246# a_17761_n5246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8092 gnd a_84221_n4481# a_84013_n4481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8093 gnd a_9496_12059# a_9288_12059# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8094 a_62031_12247# a_63128_12053# a_63079_12243# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8095 gnd d3 a_6959_11221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8096 a_641_3154# a_1260_3145# a_1468_3145# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8097 gnd a_61099_n11254# a_60891_n11254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8098 a_23143_9830# a_22722_9830# a_22314_9909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8099 a_20207_n4293# a_20464_n4483# a_19159_n4289# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8100 gnd a_19157_10537# a_18949_10537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8101 gnd a_82470_5205# a_82262_5205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8102 a_55308_5265# a_54887_5265# a_54479_4949# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8103 a_27307_8374# a_27564_8184# a_26992_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8104 vdd a_52887_n12773# a_52679_n12773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8105 a_45487_n12716# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8106 a_47399_n5866# a_46978_n5866# a_47305_n5747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8107 a_30917_10550# a_31170_10537# a_29865_10731# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8108 a_84755_5215# a_85008_5202# a_83707_4540# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8109 a_11967_6785# a_11754_6785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8110 a_39345_n12765# a_39432_n11256# a_39387_n11243# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8111 a_12017_n6710# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8112 a_77034_n5192# a_76821_n5192# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8113 gnd d0 a_85269_n4485# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8114 vdd d1 a_19416_n4479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8115 vdd d3 a_39340_11213# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8116 a_51325_6068# a_52418_6730# a_52369_6920# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8117 a_67112_6785# a_66899_6785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8118 a_31174_n11921# a_31170_n11744# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8119 a_35925_10587# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8120 a_66065_4590# a_65852_4590# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8121 a_11755_5265# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8122 vdd a_52888_n5924# a_52680_n5924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8123 a_22979_n11194# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8124 a_45439_8234# a_45226_8234# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8125 a_65703_n11115# a_65703_n11510# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8126 a_36547_n11882# a_36438_n11882# a_36646_n11882# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8127 a_65446_10165# a_65446_9909# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8128 a_31174_n11921# a_31427_n11934# a_30122_n11740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8129 gnd d0 a_85010_9084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8130 gnd d0 a_9496_14185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8131 a_72996_13698# a_74093_13504# a_74048_13517# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8132 a_23403_n7385# a_24243_n6710# a_24451_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8133 a_79055_4579# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8134 a_44600_3145# a_44179_3145# a_43771_3253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8135 a_33849_3816# a_33428_3816# a_33020_3895# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8136 a_35923_4579# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8137 gnd a_50133_12743# a_49925_12743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8138 a_81062_n5744# a_81456_n9805# a_81407_n9615# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8139 vdd d0 a_85268_n14907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8140 a_22314_9259# a_22311_8571# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8141 a_14874_n11880# a_14510_n13402# a_13484_n14169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8142 a_30128_n5909# a_31221_n5247# a_31172_n5057# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8143 vdd a_73254_10541# a_73046_10541# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8144 a_4166_n11874# a_3802_n13396# a_2776_n12716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8145 vdd d0 a_42138_n6773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8146 a_9244_9784# a_9497_9771# a_8196_9109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8147 a_66325_n13393# a_66112_n13393# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8148 a_22571_n10859# a_22571_n11115# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8149 a_35159_n8163# a_36398_n7396# a_36549_n5874# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8150 a_641_10167# a_641_9911# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8151 vdd d0 a_63594_n11938# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8152 a_12437_n4422# a_13277_n3747# a_13485_n3747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8153 a_49881_9789# a_51373_10543# a_51328_10556# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8154 a_44859_n10424# a_44438_n10424# a_44030_n10316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8155 a_2570_n8155# a_2357_n8155# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8156 vdd d0 a_20205_9086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8157 a_9501_n10472# a_9497_n10295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8158 gnd a_39643_n8215# a_39435_n8215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8159 a_31172_n3610# a_31429_n3800# a_30128_n4462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8160 a_77242_n5871# a_76821_n5871# a_76414_n6377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8161 a_33019_6862# a_33640_6783# a_33848_6783# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8162 a_72994_6243# a_73251_6053# a_71547_6923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8163 a_66067_10598# a_65854_10598# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8164 vdd d2 a_50131_6735# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8165 vdd a_74560_n14222# a_74352_n14222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8166 a_24191_11273# a_25430_10593# a_25581_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8167 gnd d1 a_19414_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8168 a_14619_6222# a_14249_7548# a_13223_8228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8169 a_76562_10592# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8170 a_11609_n8728# a_11606_n9416# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8171 a_31171_n14032# a_31175_n14888# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8172 a_82520_n14210# a_84012_n13456# a_83967_n13443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8173 gnd a_74562_n8893# a_74354_n8893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8174 vdd a_28672_6733# a_28464_6733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8175 gnd a_27479_n5928# a_27271_n5928# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8176 a_11756_12114# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8177 vdd a_62286_7496# a_62078_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8178 a_33279_n9418# a_33903_n8838# a_34111_n8838# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8179 a_1308_n5184# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8180 a_23192_n9747# a_22979_n9747# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8181 a_17450_6919# a_18946_6049# a_18897_6239# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8182 a_66067_9151# a_65854_9151# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8183 vdd d1 a_8449_10543# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8184 a_65443_7920# a_65443_7665# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8185 a_12435_n11198# a_12014_n11198# a_11606_n11119# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8186 a_17452_12927# a_17709_12737# a_17414_11228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8187 a_23983_11273# a_23770_11273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8188 a_22935_9151# a_22722_9151# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8189 gnd a_51839_n13448# a_51631_n13448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8190 a_26670_5271# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8191 a_45908_n14163# a_45487_n14163# a_44860_n14838# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8192 vdd a_7261_n5240# a_7053_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8193 a_3799_12117# a_3586_12117# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8194 a_31170_n11065# a_31427_n11255# a_30126_n11917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8195 a_63084_11225# a_63337_11212# a_62036_10550# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8196 vdd d0 a_9495_3763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8197 a_33690_n8838# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8198 a_66274_12118# a_65853_12118# a_65446_11612# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8199 a_52371_14375# a_52375_13519# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8200 a_11969_14240# a_11756_14240# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8201 vdd a_74301_14183# a_74093_14183# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8202 a_41624_14190# a_41877_14177# a_40576_13515# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8203 vdd a_8707_n13448# a_8499_n13448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8204 a_77243_n6712# a_78083_n6716# a_78291_n6716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8205 a_68602_6107# a_68389_6107# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8206 a_83962_n10299# a_85059_n10493# a_85014_n10480# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8207 a_55102_9147# a_54889_9147# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8208 gnd a_72065_n14217# a_71857_n14217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8209 a_55147_n14165# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8210 a_11349_10161# a_11970_10594# a_12178_10594# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8211 a_49877_9966# a_50134_9776# a_49834_11411# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8212 a_51588_n7427# a_51841_n7440# a_50141_n8194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8213 a_23192_n11873# a_22979_n11873# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8214 a_6964_n12757# a_7217_n12770# a_5894_n9607# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8215 a_899_n14475# a_899_n14730# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8216 a_74043_4719# a_74047_3774# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8217 vdd a_85009_12051# a_84801_12051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8218 a_76772_6783# a_76559_6783# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8219 a_36438_n11882# a_36225_n11882# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8220 a_56407_n9755# a_56194_n9755# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8221 a_44179_4592# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8222 a_76560_5263# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8223 a_12178_9826# a_11757_9826# a_11349_9905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8224 a_31177_n8201# a_31173_n8024# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8225 a_51584_n7250# a_52681_n7444# a_52632_n7254# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8226 a_33690_n6712# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8227 a_638_6870# a_638_6475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8228 a_56616_n14169# a_56195_n14169# a_55568_n14165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8229 a_83965_n7258# a_85062_n7452# a_85017_n7439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8230 vdd d2 a_82774_n5248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8231 a_66274_13565# a_67114_14240# a_67322_14240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8232 a_80832_5265# a_81196_8178# a_81147_8368# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8233 a_13278_n8161# a_13065_n8161# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8234 a_62031_12247# a_63128_12053# a_63083_12066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8235 vdd d3 a_6959_11221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8236 a_5210_5273# a_4997_5273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8237 a_3544_10595# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8238 a_49878_6748# a_51370_7502# a_51325_7515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8239 vdd a_19415_n13454# a_19207_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8240 a_8455_n5907# a_9548_n5245# a_9499_n5055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8241 a_84753_11400# a_84757_10544# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8242 a_66112_n13393# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8243 a_2567_n11196# a_2354_n11196# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8244 a_12803_5261# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8245 a_77610_9820# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8246 a_12804_12789# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8247 a_66901_12793# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8248 a_33427_7551# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8249 a_65444_3506# a_66065_3822# a_66273_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8250 a_66324_n11194# a_66111_n11194# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8251 a_28373_5401# a_28465_3766# a_28416_3956# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8252 gnd d1 a_84220_n14903# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8253 gnd d1 a_30381_n5922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8254 a_51325_6068# a_52418_6730# a_52373_6743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8255 a_11080_986# a_10971_986# a_11179_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8256 a_52372_9282# a_52373_8190# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8257 a_74306_n11242# a_74302_n11065# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8258 a_55360_n14844# a_55147_n14844# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8259 a_33280_n14088# a_33280_n14483# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8260 a_60587_3775# a_62079_4529# a_62030_4719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8261 vdd a_74562_n8214# a_74354_n8214# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8262 a_21608_973# a_21395_973# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8263 a_43773_10963# a_44394_11279# a_44602_11279# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8264 a_79679_n11882# a_79315_n13404# a_78289_n12724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8265 a_76153_13126# a_76774_13559# a_76982_13559# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8266 gnd a_72024_n6764# a_71816_n6764# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8267 a_74304_n5736# a_74309_n6754# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8268 vdd d0 a_9496_14185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8269 vdd d0 a_85010_9084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8270 a_40832_n5738# a_41929_n5932# a_41880_n5742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8271 a_2777_n5188# a_4016_n4421# a_4173_n5747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8272 a_34476_3812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8273 a_33850_12112# a_33429_12112# a_33021_12220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8274 vdd a_50133_12743# a_49925_12743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8275 a_77610_11267# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8276 a_18902_3095# a_19995_3757# a_19946_3947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8277 a_58011_n11761# a_57641_n10435# a_56615_n9755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8278 a_29863_3276# a_30960_3082# a_30911_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8279 gnd d0 a_31168_3761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8280 a_1046_7559# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8281 a_13275_n11202# a_13062_n11202# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8282 a_36648_n5874# a_36227_n5874# a_36554_n5755# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8283 vdd a_74300_4529# a_74092_4529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8284 a_9240_9961# a_9497_9771# a_8196_9109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8285 a_77242_n4424# a_76821_n4424# a_76413_n4316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8286 a_44601_12120# a_44180_12120# a_43773_11614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8287 vdd d4 a_6151_n9797# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8288 a_19951_13513# a_20204_13500# a_18899_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8289 a_52633_n11240# a_52886_n11253# a_51585_n11915# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8290 a_28678_n8019# a_28935_n8209# a_28635_n6574# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8291 gnd d0 a_85267_n11940# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8292 a_44178_8238# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8293 a_24189_5265# a_23768_5265# a_23141_4590# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8294 a_12015_n12718# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8295 vdd d3 a_28890_n12772# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8296 gnd a_73253_13508# a_73045_13508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8297 a_34109_n14167# a_34949_n14171# a_35157_n14171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8298 a_78029_5259# a_77608_5259# a_76981_4584# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8299 a_67161_n3743# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8300 gnd d0 a_74299_7496# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8301 a_3908_12117# a_3544_10595# a_2518_9828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8302 gnd a_9757_n6765# a_9549_n6765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8303 a_13484_n12722# a_14723_n13402# a_14874_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8304 vdd d0 a_85007_7490# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8305 vdd a_17707_6729# a_17499_6729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8306 vdd d0 a_31427_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8307 a_51587_n4460# a_52680_n3798# a_52631_n3608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8308 a_82219_11226# a_82306_12735# a_82257_12925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8309 a_5638_8199# a_6751_11221# a_6702_11411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8310 a_19950_3770# a_20203_3757# a_18902_3095# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8311 a_44600_5271# a_45440_5267# a_45648_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8312 a_54480_14319# a_54480_13924# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8313 a_74044_13694# a_74048_12749# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8314 vdd d2 a_60841_12737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8315 a_51581_n10291# a_52678_n10485# a_52633_n10472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8316 a_22719_6789# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8317 a_79426_12228# a_79056_13554# a_78030_14234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8318 a_12178_11273# a_13018_11269# a_13226_11269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8319 gnd a_20205_9086# a_19997_9086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8320 a_7007_n14202# a_8499_n13448# a_8454_n13435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8321 a_63083_12066# a_63079_12243# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8322 a_67375_n8157# a_67162_n8157# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8323 a_52371_12928# a_52628_12738# a_51327_12076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8324 vdd a_41087_n10489# a_40879_n10489# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8325 a_18904_10550# a_19997_11212# a_19948_11402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8326 a_20208_n6581# a_20465_n6771# a_19164_n7433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8327 a_44032_n3402# a_44032_n3658# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8328 a_52376_11231# a_52372_11408# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8329 a_1519_n11871# a_1306_n11871# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8330 a_36225_n11882# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8331 gnd d1 a_83961_13502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8332 gnd d0 a_85270_n6773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8333 a_36388_12109# a_35967_12109# a_36294_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8334 a_65705_n5502# a_65705_n5757# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8335 a_63080_11402# a_63337_11212# a_62036_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8336 gnd a_8446_7502# a_8238_7502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8337 vdd d6 a_32426_n1647# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8338 a_52629_n11742# a_52886_n11932# a_51581_n11738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8339 gnd d0 a_52888_n5245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8340 a_47139_12117# a_46718_12117# a_47040_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8341 a_33019_7914# a_33640_8230# a_33848_8230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8342 a_2354_n11196# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8343 vdd d5 a_38187_n5934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8344 a_1520_n14159# a_1307_n14159# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8345 a_19158_n14711# a_19415_n14901# a_17711_n14031# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8346 vdd d1 a_40829_13502# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8347 a_1470_9832# a_2310_9828# a_2518_9828# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8348 gnd d2 a_71807_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8349 a_39126_9958# a_40622_9088# a_40577_9101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8350 vdd a_31169_13504# a_30961_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8351 vdd a_85268_n13460# a_85060_n13460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8352 a_75885_984# a_75776_984# a_64849_973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8353 a_1467_7559# a_1046_7559# a_638_7667# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8354 a_19949_6737# a_19945_6914# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8355 a_83969_n8882# a_84222_n8895# a_82518_n8025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8356 vdd a_9756_n5924# a_9548_n5924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8357 gnd a_9495_3763# a_9287_3763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8358 a_43772_12878# a_43772_12483# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8359 a_9504_n8878# a_9500_n8701# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8360 a_63078_3947# a_63335_3757# a_62034_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8361 gnd d1 a_19157_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8362 vdd d0 a_85267_n11261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8363 gnd a_73511_n11930# a_73303_n11930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8364 vdd a_31167_7496# a_30959_7496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8365 vdd d0 a_63595_n14905# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8366 a_11608_n4059# a_12229_n3743# a_12437_n3743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8367 a_1522_n8151# a_1309_n8151# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8368 a_20206_n12589# a_20463_n12779# a_19162_n13441# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8369 a_39085_5218# a_39338_5205# a_38015_8368# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8370 a_8196_10556# a_9289_11218# a_9240_11408# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8371 a_65706_n7277# a_66327_n7385# a_66535_n7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8372 gnd d0 a_63337_9765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8373 gnd a_42135_n11261# a_41927_n11261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8374 gnd d0 a_63596_n4483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8375 a_74046_6062# a_74042_6239# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8376 a_28639_n6751# a_28892_n6764# a_27571_n9786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8377 a_36287_6101# a_36178_6101# a_36386_6101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8378 a_54889_9147# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8379 a_46886_7554# a_46673_7554# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8380 a_65852_5269# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8381 a_28373_5401# a_28465_3766# a_28420_3779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8382 a_47137_6109# a_46716_6109# a_47038_6109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8383 a_44391_7559# a_44178_7559# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8384 a_24241_n14165# a_24028_n14165# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8385 a_23403_n8832# a_22982_n8832# a_22574_n8724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8386 a_22313_13673# a_22934_13565# a_23142_13565# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8387 a_60802_n6578# a_61059_n6768# a_59738_n9790# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8388 a_78290_n5196# a_77869_n5196# a_77242_n5871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8389 a_52370_5400# a_52374_4544# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8390 a_52373_6743# a_52369_6920# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8391 a_1728_n14838# a_2568_n14163# a_2776_n14163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8392 a_901_n7816# a_1522_n7383# a_1730_n7383# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8393 a_2515_6787# a_2094_6787# a_1467_6791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8394 a_55307_6785# a_54886_6785# a_54478_6469# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8395 a_11606_n11769# a_12227_n11877# a_12435_n11877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8396 a_65704_n14082# a_66325_n14161# a_66533_n14161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8397 vdd d3 a_7217_n12770# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8398 vdd d0 a_41877_13498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8399 a_23142_12797# a_22721_12797# a_22313_12481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8400 a_57384_10589# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8401 a_41882_n9801# a_42135_n9814# a_40834_n10476# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8402 a_14715_12111# a_14294_12111# a_14621_12230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8403 a_4997_5273# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8404 gnd d3 a_50091_11221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8405 a_33848_8230# a_33427_8230# a_33019_7914# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8406 a_11754_6785# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8407 a_29863_3276# a_30960_3082# a_30915_3095# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8408 a_9238_3274# a_641_3154# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8409 vdd d0 a_31168_3761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8410 a_43772_12483# a_44393_12799# a_44601_12799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8411 a_76772_8230# a_76559_8230# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8412 a_54741_n8728# a_55362_n8836# a_55570_n8836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8413 a_34899_9820# a_34478_9820# a_33851_9824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8414 a_45226_8234# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8415 a_44651_n9745# a_44438_n9745# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8416 a_9502_n12760# a_9498_n12583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8417 gnd d0 a_9757_n8212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8418 a_28677_n5052# a_30173_n5922# a_30128_n5909# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8419 a_11757_10594# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8420 gnd d2 a_82772_n11256# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8421 a_33280_n12385# a_33280_n12641# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8422 vdd d0 a_63594_n9812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8423 a_41885_n8886# a_41881_n8709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8424 a_3844_n11874# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8425 a_4057_n11874# a_3844_n11874# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8426 a_25844_n11757# a_25474_n10431# a_24448_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8427 a_66272_6110# a_65851_6110# a_65444_5604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8428 a_1259_6791# a_1046_6791# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8429 a_67582_n5190# a_68821_n4423# a_68978_n5749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8430 a_2731_n1225# d9 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8431 vdd d3 a_17925_n12776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8432 a_78082_n3749# a_77869_n3749# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8433 a_639_4700# a_639_4159# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8434 a_24188_6785# a_25427_7552# a_25584_6226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8435 a_1306_n11871# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8436 a_1260_3824# a_1047_3824# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8437 a_82479_n6757# a_82566_n5248# a_82521_n5235# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8438 a_66901_14240# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8439 a_54741_n7026# a_55362_n6710# a_55570_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8440 vdd a_42135_n11940# a_41927_n11940# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8441 a_5638_8199# a_6751_11221# a_6706_11234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8442 a_33901_n14846# a_33688_n14846# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8443 vdd d0 a_41876_5202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8444 a_82219_11226# a_82306_12735# a_82261_12748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8445 a_1470_9153# a_1049_9153# a_638_8573# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8446 a_84757_10544# a_84753_10721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8447 a_77870_n8163# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8448 a_22312_5348# a_22933_5269# a_23141_5269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8449 a_45650_11275# a_46889_10595# a_47040_12117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8450 a_66275_10598# a_65854_10598# a_65446_10706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8451 a_63342_n12766# a_63338_n12589# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8452 vdd a_20205_9086# a_19997_9086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8453 a_2097_9828# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8454 a_18897_7686# a_19154_7496# a_17454_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8455 a_65705_n3660# a_66326_n3739# a_66534_n3739# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8456 a_54739_n12383# a_54739_n12639# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8457 a_59173_n8845# a_58752_n8845# a_58105_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8458 a_31173_n7256# a_31177_n8201# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8459 a_4267_n5866# a_3846_n5866# a_4168_n5866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8460 a_18904_10550# a_19997_11212# a_19952_11225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8461 a_52634_n14886# a_52630_n14709# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8462 a_28676_n14027# a_28933_n14217# a_28633_n12582# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8463 a_83967_n13443# a_85060_n12781# a_85015_n12768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8464 a_9239_12249# a_9496_12059# a_8191_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8465 a_11346_6469# a_11967_6785# a_12175_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8466 a_76561_13559# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8467 a_17714_n11241# a_19206_n10487# a_19157_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8468 vdd a_42138_n7452# a_41930_n7452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8469 a_3803_n4421# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8470 a_7008_n5227# a_8500_n4473# a_8451_n4283# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8471 a_46933_n10429# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8472 a_900_n4053# a_1521_n3737# a_1729_n3737# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8473 gnd a_17969_n5246# a_17761_n5246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8474 a_33643_9824# a_33430_9824# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8475 a_77033_n14167# a_76820_n14167# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8476 vdd d0 a_74301_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8477 a_66273_4590# a_65852_4590# a_65444_4157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8478 a_77822_14234# a_77609_14234# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8479 a_50134_n11058# a_50391_n11248# a_50096_n12757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8480 a_62295_n4466# a_63388_n3804# a_54740_n3408# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8481 a_55570_n8836# a_55149_n8836# a_54741_n8728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8482 a_898_n10061# a_898_n10316# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8483 a_5549_n5736# a_5943_n9797# a_5898_n9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8484 a_44859_n11192# a_44438_n11192# a_44030_n11508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8485 gnd a_30119_6053# a_29911_6053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8486 gnd d1 a_19416_n4479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8487 a_22722_9151# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8488 a_77240_n11879# a_76819_n11879# a_76412_n12385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8489 a_39345_n12765# a_39432_n11256# a_39383_n11066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8490 a_71810_n8019# a_73306_n8889# a_73261_n8876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8491 gnd d2 a_28934_n5242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8492 gnd a_52888_n5924# a_52680_n5924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8493 a_58006_n11880# a_57642_n13402# a_56616_n12722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8494 a_33021_12475# a_33642_12791# a_33850_12791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8495 vdd d2 a_71807_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8496 a_63083_14192# a_63336_14179# a_62035_13517# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8497 a_14879_n11761# a_14765_n11880# a_14973_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8498 a_57746_6103# a_57382_4581# a_56356_3814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8499 vdd a_9755_n12773# a_9547_n12773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8500 a_11609_n7026# a_11609_n7281# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8501 vdd a_9495_3763# a_9287_3763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8502 vdd d1 a_30380_n13450# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8503 a_6742_6925# a_8238_6055# a_8189_6245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8504 gnd d0 a_9755_n13452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8505 a_54480_13924# a_54480_13669# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8506 a_22573_n5107# a_22573_n5502# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8507 gnd d0 a_42137_n5253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8508 a_24030_n6710# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8509 a_60546_11228# a_60633_12737# a_60588_12750# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8510 vdd d0 a_63337_9765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8511 a_12805_11269# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8512 a_55567_n11198# a_55146_n11198# a_54738_n11119# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8513 a_55149_n8157# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8514 gnd d0 a_9495_3084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8515 gnd d0 a_63594_n11938# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8516 a_30122_n10293# a_30379_n10483# a_28679_n11237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8517 gnd d4 a_70696_8184# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8518 vdd a_51841_n7440# a_51633_n7440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8519 a_54886_8232# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8520 vdd d0 a_74559_n10487# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8521 a_17412_5220# a_17499_6729# a_17454_6742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8522 a_13483_n9755# a_13062_n9755# a_12435_n9751# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8523 a_10496_n1455# a_10753_n1645# a_10595_n1632# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8524 a_30126_n10470# a_31219_n9808# a_31174_n9795# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8525 a_66327_n8153# a_66114_n8153# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8526 a_28421_12754# a_29913_13508# a_29868_13521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8527 a_23194_n5865# a_22981_n5865# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8528 a_54479_3247# a_54481_3148# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8529 a_82261_12748# a_83753_13502# a_83704_13692# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8530 a_1261_12799# a_1048_12799# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8531 a_76559_6783# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8532 a_898_n9410# a_898_n9666# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8533 vdd d0 a_74302_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8534 vdd d3 a_50091_11221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8535 a_82520_n14210# a_84012_n13456# a_83963_n13266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8536 a_1306_n10424# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8537 a_23403_n8153# a_24243_n8157# a_24451_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8538 a_85012_n5063# a_85016_n5919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8539 a_84756_14190# a_84752_14367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8540 a_39129_12748# a_40621_13502# a_40576_13515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8541 a_3846_n5866# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8542 a_19950_4538# a_19946_4715# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8543 a_6962_n6572# a_7054_n8207# a_7009_n8194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8544 gnd d0 a_20203_5204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8545 a_68607_n13398# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8546 gnd d1 a_40827_7494# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8547 a_22314_9909# a_22314_9514# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8548 gnd a_31168_3761# a_30960_3761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8549 a_51321_6245# a_52418_6051# a_52369_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8550 a_6960_n12580# a_7052_n14215# a_7007_n14202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8551 a_52630_n14709# a_52887_n14899# a_51582_n14705# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8552 a_23140_7557# a_22719_7557# a_22311_7124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8553 vdd a_52888_n5245# a_52680_n5245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8554 vdd d0 a_42137_n5932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8555 gnd a_7261_n5240# a_7053_n5240# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8556 a_12016_n3743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8557 a_43770_8317# a_43770_7922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8558 a_39085_5218# a_39172_6727# a_39123_6917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8559 a_2775_n9749# a_4014_n10429# a_4171_n11755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8560 a_31174_n11242# a_31427_n11255# a_30126_n11917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8561 a_66532_n10426# a_66111_n10426# a_65703_n10859# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8562 a_69930_n8841# a_69717_n8841# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8563 a_24188_6785# a_23767_6785# a_23140_6110# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8564 a_33900_n9753# a_33687_n9753# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8565 a_33849_3137# a_33428_3137# a_33020_3245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8566 a_2569_n3741# a_2356_n3741# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8567 a_8194_3101# a_9287_3763# a_9238_3953# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8568 gnd a_8707_n13448# a_8499_n13448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8569 a_78028_6779# a_77607_6779# a_76980_6104# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8570 a_2309_12795# a_2096_12795# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8571 a_52374_4544# a_52370_4721# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8572 a_9244_9105# a_9497_9092# a_8192_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8573 gnd a_63336_12732# a_63128_12732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8574 gnd d0 a_41875_6722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8575 a_44599_6791# a_45439_6787# a_45647_6787# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8576 vdd d0 a_63594_n11259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8577 vdd a_85007_7490# a_84799_7490# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8578 gnd d0 a_63597_n6771# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8579 a_84750_6233# a_84755_5215# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8580 a_30122_n10293# a_31219_n10487# a_31174_n10474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8581 a_33427_6104# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8582 a_67159_n9751# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8583 a_40572_13692# a_41669_13498# a_41624_13511# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8584 gnd d2 a_82774_n5248# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8585 a_23982_14240# a_23769_14240# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8586 a_34109_n14846# a_33688_n14846# a_33280_n14738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8587 a_77242_n5192# a_76821_n5192# a_76413_n5508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8588 a_76413_n4061# a_76413_n4316# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8589 a_63081_7505# a_63077_7682# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8590 a_33280_n13291# a_33901_n13399# a_34109_n13399# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8591 a_1521_n4416# a_1308_n4416# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8592 a_53890_986# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8593 vdd a_84221_n4481# a_84013_n4481# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8594 a_2570_n6708# a_2357_n6708# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8595 gnd a_19415_n13454# a_19207_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8596 a_18903_13517# a_19996_14179# a_19947_14369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8597 a_44439_n14838# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8598 a_1259_8238# a_1046_8238# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8599 a_24451_n8157# a_24030_n8157# a_23403_n8153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8600 a_57845_6103# a_57424_6103# a_57751_6222# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8601 vdd a_30119_6053# a_29911_6053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8602 a_85012_n4295# a_85269_n4485# a_83964_n4291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8603 a_45700_n12716# a_45487_n12716# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8604 a_84757_10544# a_85010_10531# a_83705_10725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8605 a_11346_7120# a_11346_6864# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8606 a_2775_n9749# a_2354_n9749# a_1727_n9745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8607 a_55307_8232# a_56147_8228# a_56355_8228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8608 a_49026_n9607# a_49283_n9797# a_48681_n5736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8609 gnd a_74562_n8214# a_74354_n8214# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8610 a_22935_9830# a_22722_9830# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8611 vdd d1 a_83960_4527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8612 a_55361_n5869# a_55148_n5869# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8613 a_40833_n8705# a_41090_n8895# a_39386_n8025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8614 a_68608_n4423# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8615 a_30917_9782# a_30913_9959# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8616 a_33282_n8475# a_33903_n8159# a_34111_n8159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8617 a_5549_n5736# a_5806_n5926# a_5648_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8618 a_68604_12115# a_68391_12115# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8619 a_55310_10594# a_54889_10594# a_54481_10161# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8620 a_43773_10167# a_43773_9911# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8621 a_6742_6925# a_8238_6055# a_8193_6068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8622 a_36180_12109# a_35967_12109# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8623 a_44439_n12712# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8624 vdd a_84219_n10489# a_84011_n10489# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8625 a_26746_9142# a_26883_5271# a_27091_5271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8626 a_46676_10595# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8627 gnd a_71807_9774# a_71599_9774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8628 a_79357_n11882# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8629 a_33428_4584# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8630 a_33690_n8159# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8631 gnd d2 a_17970_n8213# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8632 vdd d0 a_9495_3084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8633 vdd d4 a_70696_8184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8634 gnd a_19157_9090# a_18949_9090# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8635 a_45908_n12716# a_45487_n12716# a_44860_n12712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8636 vdd a_42136_n14907# a_41928_n14907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8637 a_52629_n9616# a_52886_n9806# a_51585_n10468# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8638 a_83707_3093# a_83960_3080# a_82256_3950# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8639 vdd a_19417_n7446# a_19209_n7446# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8640 a_34110_n3745# a_34950_n3749# a_35158_n3749# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8641 a_44859_n11192# a_45699_n11196# a_45907_n11196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8642 a_11347_4949# a_11347_4694# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8643 a_31173_n7256# a_31430_n7446# a_30125_n7252# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8644 a_16027_5267# a_15918_5267# a_11080_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8645 gnd a_63337_9765# a_63129_9765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8646 a_23192_n11194# a_22979_n11194# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8647 vdd a_62288_13504# a_62080_13504# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8648 a_76819_n10432# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8649 a_25678_6107# a_25257_6107# a_25579_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8650 gnd d0 a_31427_n11934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8651 a_76152_5342# a_76773_5263# a_76981_5263# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8652 a_12178_9147# a_11757_9147# a_11349_9255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8653 a_46673_7554# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8654 a_63344_n8884# a_63597_n8897# a_62292_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8655 a_9498_n14709# a_10566_n15020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8656 a_51581_n10291# a_52678_n10485# a_52629_n10295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8657 a_19948_11402# a_19952_10546# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8658 a_74306_n11921# a_74302_n11744# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8659 a_33280_n14738# a_32239_n15022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8660 vdd a_41090_n7448# a_40882_n7448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8661 a_7007_n14202# a_8499_n13448# a_8450_n13258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8662 a_46934_n13396# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8663 a_12175_7553# a_11754_7553# a_11346_7120# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8664 gnd a_41087_n10489# a_40879_n10489# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8665 a_28639_n6751# a_28726_n5242# a_28677_n5052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8666 a_78288_n9757# a_79527_n10437# a_79684_n11763# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8667 a_20211_n5238# a_20464_n5251# a_19163_n5913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8668 a_76983_9145# a_77823_9820# a_78031_9820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8669 gnd d4 a_27824_n9799# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8670 a_54741_n7822# a_54741_n8078# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8671 a_11609_n6631# a_11609_n7026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8672 a_65446_3152# a_66065_3143# a_66273_3143# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8673 a_66066_14244# a_65853_14244# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8674 a_63084_9099# a_63080_9276# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8675 a_51321_6245# a_52418_6051# a_52373_6064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8676 a_23767_8232# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8677 a_55360_n14165# a_55147_n14165# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8678 vdd a_31168_3761# a_30960_3761# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8679 a_12230_n8836# a_12017_n8836# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8680 a_23980_6785# a_23767_6785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8681 a_70015_5271# a_69802_5271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8682 a_65703_n10859# a_65703_n11115# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8683 a_67373_n14165# a_67160_n14165# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8684 a_15573_9138# a_15360_9138# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8685 a_40836_n5915# a_41929_n5253# a_41880_n5063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8686 gnd d6 a_32426_n1647# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8687 a_22313_13928# a_22313_13673# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8688 a_44032_n3658# a_44653_n3737# a_44861_n3737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8689 a_50094_n6572# a_50186_n8207# a_50137_n8017# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8690 a_8194_3101# a_9287_3763# a_9242_3776# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8691 gnd d0 a_9497_11218# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8692 a_54738_n11769# a_55359_n11877# a_55567_n11877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8693 a_52633_n10472# a_52629_n10295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8694 a_18898_3272# a_19995_3078# a_19946_3268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8695 gnd d5 a_38187_n5934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8696 a_11607_n13289# a_11607_n13830# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8697 a_63337_n9622# a_63341_n10478# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8698 gnd d0 a_31168_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8699 a_51325_6068# a_51578_6055# a_49874_6925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8700 a_13017_14236# a_12804_14236# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8701 vdd a_63336_12732# a_63128_12732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8702 a_51328_9109# a_52421_9771# a_52372_9961# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8703 gnd d0 a_31427_n9808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8704 a_12230_n6710# a_12017_n6710# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8705 gnd d0 a_52626_8177# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8706 a_56194_n11202# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8707 a_22571_n11510# a_22571_n11765# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8708 a_40574_7507# a_41667_8169# a_41618_8359# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8709 gnd a_85268_n13460# a_85060_n13460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8710 vdd d0 a_41875_6722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8711 a_19163_n4466# a_20256_n3804# a_20207_n3614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8712 gnd a_9756_n5924# a_9548_n5924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8713 gnd d1 a_41089_n4481# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8714 a_22311_6868# a_22932_6789# a_23140_6789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8715 vdd a_41876_5202# a_41668_5202# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8716 a_33429_14238# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8717 a_11607_n13830# a_12228_n13397# a_12436_n13397# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8718 a_901_n8467# a_901_n8722# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8719 vdd d0 a_31430_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8720 a_34896_6779# a_36135_7546# a_36292_6220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8721 a_60849_n8200# a_61102_n8213# a_60802_n6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8722 a_74303_n14032# a_74307_n14888# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8723 a_71549_12931# a_73045_12061# a_72996_12251# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8724 a_12435_n9751# a_12014_n9751# a_11606_n9672# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8725 a_20210_n12766# a_20463_n12779# a_19162_n13441# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8726 a_17713_n8023# a_19209_n8893# a_19160_n8703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8727 a_63083_12745# a_63079_12922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8728 a_17710_n11064# a_19206_n11934# a_19161_n11921# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8729 vdd a_31428_n13454# a_31220_n13454# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8730 a_54480_13669# a_55101_13561# a_55309_13561# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8731 a_34898_12787# a_34477_12787# a_33850_12791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8732 a_67115_9826# a_66902_9826# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8733 vdd d0 a_31427_n11255# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8734 a_639_4159# a_1260_4592# a_1468_4592# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8735 a_63340_n8028# a_63597_n8218# a_62296_n8880# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8736 a_19950_3091# a_20203_3078# a_18898_3272# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8737 a_20207_n5740# a_20464_n5930# a_19159_n5736# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8738 a_55100_5265# a_54887_5265# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8739 gnd d2 a_7262_n8207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8740 a_56196_n5194# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8741 a_74309_n6754# a_74305_n6577# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8742 a_33022_11350# a_33643_11271# a_33851_11271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8743 a_44030_n11508# a_44030_n11763# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8744 a_22719_6110# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8745 a_9243_12751# a_9496_12738# a_8195_12076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8746 vdd a_8709_n7440# a_8501_n7440# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8747 a_60806_n6755# a_61059_n6768# a_59738_n9790# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8748 a_84753_10721# a_85010_10531# a_83705_10725# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8749 vdd d1 a_30381_n5922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8750 a_33430_9824# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8751 a_79529_n4429# a_79316_n4429# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8752 gnd d0 a_85269_n5932# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8753 vdd d1 a_19416_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8754 a_52371_12249# a_52628_12059# a_51323_12253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8755 gnd d3 a_7217_n12770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8756 a_1307_n13391# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8757 a_44859_n10424# a_45699_n9749# a_45907_n9749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8758 a_9500_n7254# a_9757_n7444# a_8452_n7250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8759 a_40832_n5738# a_41929_n5932# a_41884_n5919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8760 a_67374_n5190# a_67161_n5190# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8761 a_66326_n4418# a_66113_n4418# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8762 a_1519_n11192# a_1306_n11192# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8763 a_57684_n11880# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8764 a_44033_n7275# a_44033_n7816# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8765 vdd a_48938_n5926# a_48730_n5926# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8766 a_44600_4592# a_44179_4592# a_43771_4700# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8767 a_74304_n5057# a_74308_n5913# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8768 vdd a_71807_9774# a_71599_9774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8769 a_641_10963# a_1262_11279# a_1470_11279# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8770 a_22572_n14082# a_22572_n14477# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8771 a_83706_7507# a_84799_8169# a_84754_8182# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8772 a_66325_n14840# a_66112_n14840# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8773 a_2776_n12716# a_4015_n13396# a_4166_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8774 a_52629_n11063# a_52886_n11253# a_51585_n11915# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8775 a_66533_n13393# a_66112_n13393# a_65704_n13826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8776 vdd d1 a_84222_n7448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8777 a_33022_9508# a_33643_9824# a_33851_9824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8778 a_83703_3270# a_83960_3080# a_82256_3950# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8779 gnd d3 a_17925_n12776# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8780 a_52369_8367# a_52626_8177# a_51325_7515# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8781 a_83966_n11923# a_85059_n11261# a_85010_n11071# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8782 gnd d1 a_30122_9094# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8783 a_33282_n7283# a_33903_n7391# a_34111_n7391# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8784 a_8450_n14705# a_9547_n14899# a_9498_n14709# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8785 a_1522_n8830# a_1309_n8830# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8786 a_24029_n5190# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8787 vdd a_63337_9765# a_63129_9765# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8788 a_74043_5398# a_74047_4542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8789 a_1469_12120# a_1048_12120# a_641_11614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8790 a_44601_13567# a_44180_13567# a_43772_13675# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8791 a_74046_6741# a_74042_6918# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8792 a_82479_n6757# a_82566_n5248# a_82517_n5058# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8793 a_72994_7690# a_73251_7500# a_71551_6746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8794 gnd a_42135_n11940# a_41927_n11940# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8795 vdd a_9756_n5245# a_9548_n5245# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8796 gnd a_9495_3084# a_9287_3084# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8797 a_72994_7690# a_74091_7496# a_74042_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8798 a_73256_n4285# a_73513_n4475# a_71813_n5229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8799 a_63078_3268# a_63335_3078# a_62030_3272# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8800 a_67160_n14165# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8801 a_638_8317# a_1259_8238# a_1467_8238# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8802 a_45439_6787# a_45226_6787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8803 a_45227_5267# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8804 a_76412_n14088# a_76412_n14483# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8805 a_44031_n14080# a_44031_n14475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8806 a_40831_n13266# a_41928_n13460# a_41883_n13447# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8807 vdd d0 a_31170_10537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8808 a_34949_n12724# a_34736_n12724# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8809 gnd d0 a_63337_9086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8810 gnd d0 a_52887_n13452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8811 a_77241_n13399# a_76820_n13399# a_76412_n13291# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8812 a_66532_n9747# a_66111_n9747# a_65703_n10063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8813 a_76154_9253# a_76151_8565# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8814 a_1522_n6704# a_1309_n6704# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8815 a_54480_12222# a_54481_11608# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8816 a_22935_10598# a_22722_10598# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8817 a_28680_n14204# a_28933_n14217# a_28633_n12582# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8818 a_65704_n14732# a_66325_n14840# a_66533_n14840# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8819 a_1469_13567# a_2309_14242# a_2517_14242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8820 a_66535_n7385# a_67375_n6710# a_67583_n6710# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8821 gnd a_62287_3082# a_62079_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8822 a_24189_5265# a_25428_4585# a_25579_6107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8823 vdd a_74302_9090# a_74094_9090# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8824 a_23403_n8153# a_22982_n8153# a_22574_n8074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8825 a_33900_n10432# a_33687_n10432# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8826 a_71553_12754# a_71806_12741# a_71511_11232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8827 a_1727_n9745# a_1306_n9745# a_898_n9666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8828 a_32431_984# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8829 gnd a_51839_n14895# a_51631_n14895# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8830 a_11606_n11119# a_12227_n11198# a_12435_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8831 a_14725_n7394# a_14512_n7394# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8832 vdd d0 a_85270_n6773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8833 a_76774_14238# a_76561_14238# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8834 a_56147_8228# a_55934_8228# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8835 a_34898_14234# a_36137_13554# a_36294_12228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8836 a_50138_n11235# a_50391_n11248# a_50096_n12757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8837 a_30127_n13437# a_31220_n12775# a_31175_n12762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8838 gnd a_20203_5204# a_19995_5204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8839 gnd a_40827_7494# a_40619_7494# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8840 a_65704_n13030# a_66325_n12714# a_66533_n12714# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8841 a_76775_9824# a_76562_9824# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8842 a_31171_n14711# a_31428_n14901# a_30123_n14707# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8843 a_17670_n6578# a_17762_n8213# a_17713_n8023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8844 vdd d0 a_31168_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8845 a_51321_6245# a_51578_6055# a_49874_6925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8846 a_46888_13562# a_46675_13562# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8847 a_43773_11614# a_44393_12120# a_44601_12120# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8848 a_71810_n8019# a_73306_n8889# a_73257_n8699# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8849 a_54741_n8078# a_55362_n8157# a_55570_n8157# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8850 a_14464_13556# a_14251_13556# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8851 a_51328_9109# a_52421_9771# a_52376_9784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8852 a_74304_n3610# a_74561_n3800# a_73260_n4462# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8853 a_83962_n11746# a_85059_n11940# a_85014_n11927# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8854 a_24450_n3743# a_24029_n3743# a_23402_n4418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8855 a_11347_3897# a_11968_3818# a_12176_3818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8856 a_25581_12115# a_25472_12115# a_25680_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8857 gnd d1 a_30380_n13450# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8858 a_34111_n7391# a_33690_n7391# a_33282_n7283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8859 a_2517_12795# a_2096_12795# a_1469_12799# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8860 vdd a_52629_11218# a_52421_11218# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8861 a_56618_n8161# a_56197_n8161# a_55570_n8836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8862 vdd a_85009_13498# a_84801_13498# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8863 a_19952_10546# a_20205_10533# a_18900_10727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8864 a_23400_n11873# a_22979_n11873# a_22572_n12379# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8865 a_641_9261# a_638_8573# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8866 a_36646_n11882# a_36225_n11882# a_36547_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8867 a_71549_12931# a_73045_12061# a_73000_12074# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8868 a_51584_n8697# a_52681_n8891# a_52632_n8701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8869 a_33281_n3666# a_33902_n3745# a_34110_n3745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8870 a_33849_4584# a_34689_5259# a_34897_5259# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8871 a_1306_n11192# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8872 a_8454_n14882# a_9547_n14220# a_9502_n14207# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8873 a_44653_n4416# a_44440_n4416# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8874 a_64849_973# a_75563_984# a_70223_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8875 a_1260_3145# a_1047_3145# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8876 a_55568_n14165# a_56408_n14169# a_56616_n14169# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8877 vdd a_9496_13506# a_9288_13506# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8878 a_62031_13694# a_63128_13500# a_63083_13513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8879 a_9241_8190# a_9237_8367# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8880 gnd a_41875_6722# a_41667_6722# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8881 a_22721_12797# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8882 vdd a_42135_n11261# a_41927_n11261# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8883 a_33901_n14167# a_33688_n14167# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8884 gnd a_51841_n7440# a_51633_n7440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8885 vdd d0 a_63596_n4483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8886 a_74044_14373# a_74048_13517# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8887 a_1049_10600# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8888 gnd d0 a_74559_n10487# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8889 a_14509_n10435# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8890 a_5648_n5913# a_10753_n1645# a_10595_n1632# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8891 a_2775_n11196# a_2354_n11196# a_1727_n11871# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8892 a_27222_n5738# a_27616_n9799# a_27567_n9609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8893 vdd d1 a_19415_n14901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8894 a_79421_12109# a_79057_10587# a_78031_11267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8895 a_16041_n8845# a_16514_n5932# a_10496_n1455# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8896 a_46929_6109# a_46716_6109# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8897 a_11347_5600# a_11967_6106# a_12175_6106# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8898 a_82259_6740# a_83751_7494# a_83702_7684# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8899 a_33643_9145# a_33430_9145# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8900 vdd d0 a_20463_n12779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8901 a_76820_n12720# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8902 a_22722_9830# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8903 vdd a_28932_n11250# a_28724_n11250# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8904 a_56615_n9755# a_57854_n10435# a_58011_n11761# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8905 a_54887_5265# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8906 gnd d1 a_83962_10535# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8907 a_33642_12791# a_33429_12791# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8908 a_68822_n7390# a_68609_n7390# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8909 a_55570_n8157# a_55149_n8157# a_54741_n8078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8910 a_8196_10556# a_8449_10543# a_6749_9789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8911 a_77240_n11200# a_76819_n11200# a_76411_n11516# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8912 a_62029_7686# a_63126_7492# a_63077_7682# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8913 a_65443_7665# a_65443_7124# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8914 a_6960_n12580# a_7052_n14215# a_7003_n14025# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8915 a_83707_3093# a_84800_3755# a_84751_3945# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8916 gnd a_52888_n5245# a_52680_n5245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8917 a_17456_12750# a_17709_12737# a_17414_11228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8918 a_33022_11606# a_33642_12112# a_33850_12112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8919 a_1467_7559# a_2307_8234# a_2515_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8920 a_56410_n8161# a_56197_n8161# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8921 a_77821_5259# a_77608_5259# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8922 a_41885_n6760# a_41881_n6583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8923 vdd a_38187_n5934# a_37979_n5934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8924 a_4017_n7388# a_3804_n7388# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8925 a_34110_n3745# a_33689_n3745# a_33281_n3666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8926 a_43771_3508# a_44392_3824# a_44600_3824# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8927 vdd a_9495_3084# a_9287_3084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8928 a_66275_9830# a_67115_9826# a_67323_9826# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8929 a_41623_5215# a_41619_5392# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8930 a_54888_13561# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8931 a_68716_6226# a_68346_7552# a_67320_6785# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8932 a_66272_7557# a_65851_7557# a_65443_7665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8933 a_13224_5261# a_14463_4581# a_14614_6103# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8934 a_36135_7546# a_35922_7546# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8935 a_85015_n13447# a_85011_n13270# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8936 vdd d0 a_63337_9086# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8937 a_49030_n9784# a_50143_n6762# a_50094_n6572# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8938 a_76151_6862# a_76772_6783# a_76980_6783# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8939 gnd d0 a_63594_n11259# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8940 a_899_n13283# a_899_n13824# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8941 a_17715_n14208# a_17968_n14221# a_17668_n12586# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8942 a_36227_n5874# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8943 vdd a_62287_3082# a_62079_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8944 a_2517_14242# a_3756_13562# a_3913_12236# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8945 vdd a_41087_n11936# a_40879_n11936# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8946 a_26746_9142# a_26325_9142# a_25680_12115# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8947 a_12436_n12718# a_12015_n12718# a_11607_n13034# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8948 a_30122_n10293# a_31219_n10487# a_31170_n10297# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8949 a_55148_n5190# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8950 a_71549_12931# a_71806_12741# a_71511_11232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8951 gnd a_30121_12061# a_29913_12061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8952 a_17454_6742# a_18946_7496# a_18901_7509# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8953 a_57751_6222# a_57381_7548# a_56355_8228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8954 a_45486_n9749# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8955 gnd d0 a_31169_13504# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8956 a_7008_n5227# a_8500_n4473# a_8455_n4460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8957 a_52634_n12760# a_52630_n12583# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8958 a_1727_n11871# a_1306_n11871# a_899_n12377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8959 a_25475_n13398# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8960 a_44031_n12377# a_44031_n12633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8961 a_23194_n5186# a_22981_n5186# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8962 a_76412_n12385# a_76412_n12641# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8963 a_67320_6785# a_66899_6785# a_66272_6789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8964 a_76559_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8965 a_85016_n4472# a_85269_n4485# a_83964_n4291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8966 a_12176_3139# a_13016_3814# a_13224_3814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8967 a_55309_13561# a_56149_14236# a_56357_14236# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8968 a_63337_n10301# a_63594_n10491# a_62289_n10297# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8969 a_23400_n10426# a_22979_n10426# a_22571_n10318# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8970 a_66327_n6706# a_66114_n6706# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8971 a_41621_10721# a_41625_9776# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8972 vdd d2 a_28934_n5242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8973 gnd d3 a_7219_n6762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8974 a_69802_5271# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8975 a_34108_n10432# a_33687_n10432# a_33279_n10865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8976 a_74047_4542# a_74043_4719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8977 a_15360_9138# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8978 a_5333_n8839# a_5806_n5926# a_5648_n5913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8979 a_3754_7554# a_3541_7554# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8980 a_33280_n13036# a_33280_n13291# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8981 a_23402_n5865# a_24242_n5190# a_24450_n5190# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8982 a_74049_11229# a_74045_11406# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8983 a_19948_10723# a_20205_10533# a_18900_10727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8984 a_63343_n4470# a_63339_n4293# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8985 a_79518_6101# a_80378_9136# a_80586_9136# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8986 gnd a_84219_n10489# a_84011_n10489# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8987 a_54478_8567# a_54478_8311# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8988 gnd a_31168_3082# a_30960_3082# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8989 vdd d0 a_9755_n13452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8990 a_34899_11267# a_34478_11267# a_33851_10592# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8991 a_24451_n8157# a_25690_n7390# a_25841_n5868# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8992 vdd d0 a_42137_n5253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8993 a_22312_4157# a_22312_3901# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8994 gnd a_74300_4529# a_74092_4529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8995 vdd a_41875_6722# a_41667_6722# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8996 a_2568_n12716# a_2355_n12716# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8997 a_29865_10731# a_30962_10537# a_30917_10550# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X8998 a_65706_n8724# a_66327_n8832# a_66535_n8832# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8999 a_70124_5271# a_70015_5271# a_70223_5271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9000 gnd a_52628_14185# a_52420_14185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9001 a_30911_3272# a_22314_3152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9002 a_8190_3278# a_8447_3088# a_6743_3958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9003 gnd a_19417_n7446# a_19209_n7446# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9004 a_900_n3402# a_900_n3658# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9005 a_8190_3278# a_9287_3084# a_9238_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9006 vdd a_7259_n11248# a_7051_n11248# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9007 a_56357_12789# a_55936_12789# a_55309_12793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9008 a_25839_n11876# a_25730_n11876# a_25938_n11876# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9009 a_76414_n8080# a_76414_n8475# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9010 a_35156_n9757# a_34735_n9757# a_34108_n10432# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9011 vdd a_19156_12057# a_18948_12057# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9012 a_52376_9105# a_52372_9282# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9013 a_54739_n13034# a_54739_n13289# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9014 gnd a_63336_12053# a_63128_12053# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9015 a_31177_n7433# a_31430_n7446# a_30125_n7252# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9016 a_79520_12109# a_79099_12109# a_79426_12228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9017 vdd a_39598_n12778# a_39390_n12778# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9018 a_898_n9410# a_1522_n8830# a_1730_n8830# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9019 gnd d0 a_41875_6043# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9020 a_11757_9826# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9021 a_55146_n10430# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9022 a_13485_n5194# a_14724_n4427# a_14881_n5753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9023 a_33902_n4424# a_33689_n4424# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9024 vdd d1 a_62549_n8893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9025 gnd d0 a_20464_n4483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9026 a_22314_9909# a_22935_9830# a_23143_9830# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9027 a_34951_n6716# a_34738_n6716# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9028 gnd a_17707_6729# a_17499_6729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9029 a_55935_5261# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9030 a_13276_n12722# a_13063_n12722# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9031 gnd a_41090_n7448# a_40882_n7448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9032 gnd d2 a_60841_12737# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9033 a_34109_n14167# a_33688_n14167# a_33280_n14088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9034 a_72997_9284# a_74094_9090# a_74049_9103# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9035 a_54212_986# a_54103_986# a_54311_986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9036 a_54739_n13830# a_55360_n13397# a_55568_n13397# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9037 a_29863_4723# a_30960_4529# a_30915_4542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9038 vdd d4 a_16859_n9803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9039 vdd a_17967_n11254# a_17759_n11254# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9040 gnd d2 a_50394_n8207# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9041 vdd d1 a_83962_10535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9042 a_44862_n8151# a_44441_n8151# a_44033_n8467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9043 a_36554_n5755# a_36184_n4429# a_35158_n3749# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9044 a_44439_n14159# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9045 a_52375_12751# a_52628_12738# a_51327_12076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9046 a_8192_10733# a_8449_10543# a_6749_9789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9047 gnd a_81664_n9805# a_81456_n9805# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9048 a_77608_3812# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9049 a_83707_3093# a_84800_3755# a_84755_3768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9050 a_55310_9826# a_56150_9822# a_56358_9822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9051 a_84756_12064# a_84752_12241# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9052 a_55361_n5190# a_55148_n5190# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9053 a_45909_n5188# a_45488_n5188# a_44861_n5184# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9054 a_4265_n11874# a_3844_n11874# a_4166_n11874# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9055 a_79572_n5874# a_79359_n5874# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9056 a_33689_n3745# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9057 vdd d0 a_74300_5208# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9058 a_65705_n4310# a_65705_n4851# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9059 a_1470_11279# a_1049_11279# a_641_10963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9060 a_22573_n4851# a_22573_n5107# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9061 a_68349_10593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9062 a_22932_7557# a_22719_7557# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9063 a_62033_7509# a_62286_7496# a_60586_6742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9064 vdd d0 a_20462_n9812# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9065 a_23141_5269# a_22720_5269# a_22312_5348# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9066 gnd a_30122_9094# a_29914_9094# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9067 a_76822_n8838# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9068 a_43770_6220# a_43771_5606# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9069 a_76980_6783# a_76559_6783# a_76151_6862# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9070 a_63083_14192# a_65445_14323# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9071 vdd a_40830_9088# a_40622_9088# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9072 a_31170_n9618# a_31174_n10474# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9073 a_65446_10706# a_66067_10598# a_66275_10598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9074 a_18902_3095# a_19155_3082# a_17451_3952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9075 a_1727_n10424# a_1306_n10424# a_898_n10316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9076 a_77241_n13399# a_78081_n12724# a_78289_n12724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9077 a_44654_n6704# a_44441_n6704# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9078 a_23768_5265# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9079 vdd d0 a_52629_10539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9080 a_65446_9514# a_65446_9259# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9081 a_19945_6914# a_19949_6058# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9082 a_45226_6787# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9083 vdd d0 a_63597_n6771# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9084 a_63082_3770# a_63335_3757# a_62034_3095# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9085 a_23981_3818# a_23768_3818# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9086 vdd a_30121_12061# a_29913_12061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9087 a_6745_9966# a_8241_9096# a_8192_9286# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9088 a_56355_6781# a_55934_6781# a_55307_6785# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9089 a_68971_n11876# a_68607_n13398# a_67581_n14165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9090 a_35156_n11204# a_36395_n10437# a_36552_n11763# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9091 a_11349_9510# a_11349_9255# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9092 a_56618_n8161# a_57857_n7394# a_58008_n5872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9093 a_17710_n11064# a_19206_n11934# a_19157_n11744# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9094 gnd a_63337_9086# a_63129_9086# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9095 gnd a_31428_n13454# a_31220_n13454# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9096 a_47303_n11755# a_46933_n10429# a_45907_n11196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9097 a_16041_n8845# a_15620_n8845# a_14973_n11880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9098 gnd d0 a_31427_n11255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9099 a_85014_n10480# a_85267_n10493# a_83962_n10299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9100 a_63084_9778# a_63080_9955# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9101 a_31171_n12585# a_31175_n13441# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9102 a_63344_n8205# a_63597_n8218# a_62296_n8880# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9103 a_44599_6112# a_44178_6112# a_43771_5606# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9104 a_20211_n5917# a_20464_n5930# a_19159_n5736# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9105 a_52631_n4287# a_52888_n4477# a_51583_n4283# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9106 a_47148_n4421# a_46935_n4421# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9107 a_82262_9781# a_83754_10535# a_83705_10725# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9108 a_12435_n10430# a_12014_n10430# a_11606_n10322# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9109 gnd a_8709_n7440# a_8501_n7440# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9110 a_34688_8226# a_34475_8226# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9111 gnd d1 a_19416_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9112 a_64664_n1444# a_64921_n1634# a_43231_n1412# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9113 a_34736_n14171# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9114 a_34735_n9757# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9115 a_2518_11275# a_2097_11275# a_1470_10600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9116 a_34897_5259# a_36136_4579# a_36287_6101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9117 a_11606_n9416# a_11606_n9672# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9118 a_9504_n7431# a_9757_n7444# a_8452_n7250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9119 a_2308_5267# a_2095_5267# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9120 a_9500_n8701# a_9501_n9793# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9121 a_76562_9824# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9122 gnd a_48938_n5926# a_48730_n5926# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9123 vdd a_31168_3082# a_30960_3082# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9124 a_12230_n8157# a_12017_n8157# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9125 a_76151_7914# a_76772_8230# a_76980_8230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9126 a_50139_n14202# a_51631_n13448# a_51586_n13435# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9127 a_22722_11277# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9128 a_85011_n12591# a_85015_n13447# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9129 a_12177_12793# a_11756_12793# a_11348_12477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9130 a_55360_n12718# a_55147_n12718# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9131 a_82258_9958# a_83754_9088# a_83709_9101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9132 a_16027_5267# a_16391_8180# a_16342_8370# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9133 a_55567_n9751# a_56407_n9755# a_56615_n9755# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9134 vdd a_52628_14185# a_52420_14185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9135 gnd d1 a_84222_n7448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9136 a_19160_n7256# a_20257_n7450# a_20212_n7437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9137 a_8190_3278# a_9287_3084# a_9242_3097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9138 a_54738_n11119# a_55359_n11198# a_55567_n11198# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9139 gnd d0 a_9495_4531# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9140 a_33848_6104# a_34688_6779# a_34896_6779# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9141 a_30122_n11740# a_30379_n11930# a_28675_n11060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9142 a_77822_12787# a_77609_12787# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9143 a_25680_12115# a_25259_12115# a_25581_12115# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9144 a_44180_12799# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9145 a_71554_9787# a_71807_9774# a_71507_11409# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9146 vdd d0 a_74559_n11934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9147 a_12438_n8836# a_13278_n8161# a_13486_n8161# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9148 a_11609_n7822# a_12230_n7389# a_12438_n7389# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9149 vdd a_63336_12053# a_63128_12053# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9150 a_81151_8191# a_82264_11213# a_82215_11403# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9151 a_51324_9286# a_52421_9092# a_52372_9282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9152 a_66532_n11873# a_67372_n11198# a_67580_n11198# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9153 vdd d0 a_41875_6043# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9154 a_29864_13698# a_30961_13504# a_30912_13694# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9155 gnd a_9756_n5245# a_9548_n5245# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9156 a_73260_n4462# a_73513_n4475# a_71813_n5229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9157 a_1048_13567# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9158 a_20212_n8205# a_20208_n8028# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9159 a_33020_3245# a_33022_3146# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9160 a_79419_6101# a_79310_6101# a_79518_6101# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9161 a_54212_986# a_58837_5267# a_59159_5267# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9162 a_82217_5218# a_82304_6727# a_82259_6740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9163 a_44438_n9745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9164 a_40831_n13266# a_41928_n13460# a_41879_n13270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9165 a_1729_n5863# a_1308_n5863# a_901_n6369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9166 a_11179_986# a_10758_986# a_11080_986# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9167 a_33643_11271# a_33430_11271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9168 a_76153_12475# a_76774_12791# a_76982_12791# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9169 a_82516_n14033# a_84012_n14903# a_83963_n14713# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9170 a_70699_n9609# a_70956_n9799# a_70354_n5738# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9171 a_76414_n6377# a_76414_n6633# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9172 a_33281_n4316# a_33281_n4857# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9173 a_25846_n5749# a_25476_n4423# a_24450_n5190# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9174 a_79778_n11882# a_79357_n11882# a_79679_n11882# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9175 a_640_14325# a_1261_14246# a_1469_14246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9176 a_28639_n6751# a_28726_n5242# a_28681_n5229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9177 a_46716_6109# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9178 a_33021_14317# a_33021_13922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9179 vdd d0 a_63336_14179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9180 a_33280_n12641# a_33280_n13036# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9181 a_20207_n5061# a_20464_n5251# a_19163_n5913# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9182 a_41881_n8709# a_41882_n9801# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9183 a_45648_3820# a_45227_3820# a_44600_3145# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9184 a_9243_12072# a_9496_12059# a_8191_12253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9185 a_12437_n4422# a_12016_n4422# a_11608_n4314# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9186 a_63339_n3614# a_63343_n4470# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9187 a_33430_9145# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9188 a_66064_8236# a_65851_8236# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9189 a_1046_6791# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9190 a_11346_6864# a_11346_6469# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9191 a_55101_12793# a_54888_12793# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9192 a_54886_6785# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9193 a_11967_7553# a_11754_7553# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9194 a_23401_n13393# a_22980_n13393# a_22572_n13285# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9195 gnd d0 a_85269_n5253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9196 a_22572_n14732# a_21274_n15026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9197 a_12176_5265# a_11755_5265# a_11347_5344# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9198 a_30127_n13437# a_31220_n12775# a_31171_n12585# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9199 a_13062_n9755# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9200 a_45228_12795# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9201 a_4007_12117# a_4865_9144# a_5073_9144# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9202 a_900_n3402# a_9756_n3798# a_8455_n4460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9203 a_40836_n5915# a_41929_n5253# a_41884_n5240# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9204 a_25477_n7390# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9205 a_33849_4584# a_33428_4584# a_33020_4692# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9206 a_44602_9153# a_45442_9828# a_45650_9828# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9207 a_77820_6779# a_77607_6779# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
C0 a_21816_973# d6 5.71fF
C1 d6 d7 119.31fF
C2 d8 d6 14.54fF
C3 d0 d1 114.29fF
C4 d2 d1 103.46fF
C5 d2 d0 8.48fF
C6 d5 d3 33.09fF
C7 vdd d1 153.81fF
C8 d5 vdd 4.76fF
C9 vdd d0 173.02fF
C10 d5 d4 130.31fF
C11 d3 d2 124.94fF
C12 d2 vdd 85.70fF
C13 d3 vdd 93.26fF
C14 a_43231_n1412# d6 5.71fF
C15 d3 d4 138.27fF
C16 d4 vdd 4.69fF
C17 d8 a_3058_n1106# 14.02fF
C18 a_85011_n14717# gnd 2.27fF
C19 a_83963_n14713# gnd 2.80fF
C20 a_75371_n15022# gnd 4.89fF
C21 a_74303_n14711# gnd 2.27fF
C22 a_73255_n14707# gnd 2.80fF
C23 a_76412_n14738# gnd 2.33fF
C24 a_64406_n15026# gnd 5.08fF
C25 a_63338_n14715# gnd 2.27fF
C26 a_62290_n14711# gnd 2.80fF
C27 a_65704_n14732# gnd 2.33fF
C28 a_53698_n15020# gnd 4.89fF
C29 a_52630_n14709# gnd 2.27fF
C30 a_51582_n14705# gnd 2.80fF
C31 a_54739_n14736# gnd 2.33fF
C32 a_42947_n15028# gnd 4.85fF
C33 a_41879_n14717# gnd 2.27fF
C34 a_40831_n14713# gnd 2.80fF
C35 a_32239_n15022# gnd 4.89fF
C36 a_31171_n14711# gnd 2.27fF
C37 a_30123_n14707# gnd 2.80fF
C38 a_44031_n14730# gnd 2.33fF
C39 a_33280_n14738# gnd 2.33fF
C40 a_21274_n15026# gnd 5.08fF
C41 a_20206_n14715# gnd 2.27fF
C42 a_19158_n14711# gnd 2.80fF
C43 a_22572_n14732# gnd 2.33fF
C44 a_10566_n15020# gnd 4.89fF
C45 a_9498_n14709# gnd 2.27fF
C46 a_8450_n14705# gnd 2.80fF
C47 a_11607_n14736# gnd 2.33fF
C48 a_899_n14730# gnd 2.73fF
C49 a_85015_n14894# gnd 3.17fF
C50 a_74307_n14888# gnd 3.17fF
C51 a_63342_n14892# gnd 3.17fF
C52 a_52634_n14886# gnd 3.17fF
C53 a_41883_n14894# gnd 3.17fF
C54 a_31175_n14888# gnd 3.17fF
C55 a_83967_n14890# gnd 3.33fF
C56 a_85011_n14038# gnd 2.33fF
C57 a_82516_n14033# gnd 4.35fF
C58 a_77241_n14846# gnd 3.33fF
C59 a_20210_n14892# gnd 3.17fF
C60 a_9502_n14886# gnd 3.17fF
C61 a_76412_n14483# gnd 3.17fF
C62 a_77241_n14167# gnd 2.80fF
C63 a_73259_n14884# gnd 3.33fF
C64 a_74303_n14032# gnd 2.33fF
C65 a_71808_n14027# gnd 4.35fF
C66 a_66533_n14840# gnd 3.33fF
C67 a_76412_n14088# gnd 2.27fF
C68 a_65704_n14477# gnd 3.17fF
C69 a_66533_n14161# gnd 2.80fF
C70 a_62294_n14888# gnd 3.33fF
C71 a_63338_n14036# gnd 2.33fF
C72 a_60843_n14031# gnd 4.35fF
C73 a_55568_n14844# gnd 3.33fF
C74 a_65704_n14082# gnd 2.27fF
C75 a_54739_n14481# gnd 3.17fF
C76 a_55568_n14165# gnd 2.80fF
C77 a_51586_n14882# gnd 3.33fF
C78 a_52630_n14030# gnd 2.33fF
C79 a_50135_n14025# gnd 4.35fF
C80 a_44860_n14838# gnd 3.33fF
C81 a_54739_n14086# gnd 2.27fF
C82 a_44031_n14475# gnd 3.17fF
C83 a_44860_n14159# gnd 2.80fF
C84 a_40835_n14890# gnd 3.33fF
C85 a_41879_n14038# gnd 2.33fF
C86 a_39384_n14033# gnd 4.35fF
C87 a_34109_n14846# gnd 3.33fF
C88 a_44031_n14080# gnd 2.27fF
C89 a_33280_n14483# gnd 3.17fF
C90 a_34109_n14167# gnd 2.80fF
C91 a_30127_n14884# gnd 3.33fF
C92 a_31171_n14032# gnd 2.33fF
C93 a_28676_n14027# gnd 4.35fF
C94 a_23401_n14840# gnd 3.33fF
C95 a_33280_n14088# gnd 2.27fF
C96 a_22572_n14477# gnd 3.17fF
C97 a_23401_n14161# gnd 2.80fF
C98 a_19162_n14888# gnd 3.33fF
C99 a_20206_n14036# gnd 2.33fF
C100 a_17711_n14031# gnd 4.35fF
C101 a_12436_n14844# gnd 3.33fF
C102 a_22572_n14082# gnd 2.27fF
C103 a_11607_n14481# gnd 3.17fF
C104 a_12436_n14165# gnd 2.80fF
C105 a_8454_n14882# gnd 3.33fF
C106 a_9498_n14030# gnd 2.33fF
C107 a_7003_n14025# gnd 4.35fF
C108 a_1728_n14838# gnd 3.40fF
C109 a_11607_n14086# gnd 2.27fF
C110 a_899_n14475# gnd 3.17fF
C111 a_1728_n14159# gnd 2.80fF
C112 a_899_n14080# gnd 2.27fF
C113 a_85015_n14215# gnd 3.43fF
C114 a_74307_n14209# gnd 3.43fF
C115 a_63342_n14213# gnd 3.43fF
C116 a_52634_n14207# gnd 3.43fF
C117 a_41883_n14215# gnd 3.43fF
C118 a_31175_n14209# gnd 3.43fF
C119 a_85011_n13270# gnd 2.27fF
C120 a_82520_n14210# gnd 3.43fF
C121 a_83963_n13266# gnd 2.80fF
C122 a_78289_n14171# gnd 3.35fF
C123 a_76412_n13832# gnd 3.43fF
C124 a_74303_n13264# gnd 2.27fF
C125 a_71812_n14204# gnd 3.43fF
C126 a_73255_n13260# gnd 2.80fF
C127 a_67581_n14165# gnd 3.35fF
C128 a_20210_n14213# gnd 3.43fF
C129 a_9502_n14207# gnd 3.43fF
C130 a_76412_n13291# gnd 2.33fF
C131 a_65704_n13826# gnd 3.43fF
C132 a_63338_n13268# gnd 2.27fF
C133 a_60847_n14208# gnd 3.43fF
C134 a_62290_n13264# gnd 2.80fF
C135 a_56616_n14169# gnd 3.35fF
C136 a_65704_n13285# gnd 2.33fF
C137 a_54739_n13830# gnd 3.43fF
C138 a_52630_n13262# gnd 2.27fF
C139 a_50139_n14202# gnd 3.43fF
C140 a_51582_n13258# gnd 2.80fF
C141 a_45908_n14163# gnd 3.35fF
C142 a_54739_n13289# gnd 2.33fF
C143 a_44031_n13824# gnd 3.43fF
C144 a_41879_n13270# gnd 2.27fF
C145 a_39388_n14210# gnd 3.43fF
C146 a_40831_n13266# gnd 2.80fF
C147 a_35157_n14171# gnd 3.35fF
C148 a_33280_n13832# gnd 3.43fF
C149 a_31171_n13264# gnd 2.27fF
C150 a_28680_n14204# gnd 3.43fF
C151 a_30123_n13260# gnd 2.80fF
C152 a_24449_n14165# gnd 3.35fF
C153 a_44031_n13283# gnd 2.33fF
C154 a_33280_n13291# gnd 2.33fF
C155 a_22572_n13826# gnd 3.43fF
C156 a_20206_n13268# gnd 2.27fF
C157 a_17715_n14208# gnd 3.43fF
C158 a_19158_n13264# gnd 2.80fF
C159 a_13484_n14169# gnd 3.35fF
C160 a_22572_n13285# gnd 2.33fF
C161 a_11607_n13830# gnd 3.43fF
C162 a_9498_n13262# gnd 2.27fF
C163 a_7007_n14202# gnd 3.43fF
C164 a_8450_n13258# gnd 2.80fF
C165 a_2776_n14163# gnd 3.35fF
C166 a_11607_n13289# gnd 2.33fF
C167 a_899_n13824# gnd 3.43fF
C168 a_899_n13283# gnd 2.33fF
C169 a_85015_n13447# gnd 3.17fF
C170 a_74307_n13441# gnd 3.17fF
C171 a_63342_n13445# gnd 3.17fF
C172 a_52634_n13439# gnd 3.17fF
C173 a_41883_n13447# gnd 3.17fF
C174 a_31175_n13441# gnd 3.17fF
C175 a_83967_n13443# gnd 3.33fF
C176 a_85011_n12591# gnd 2.33fF
C177 a_82473_n12588# gnd 3.27fF
C178 a_77241_n13399# gnd 3.33fF
C179 a_78289_n12724# gnd 3.73fF
C180 a_20210_n13445# gnd 3.17fF
C181 a_9502_n13439# gnd 3.17fF
C182 a_76412_n13036# gnd 3.17fF
C183 a_77241_n12720# gnd 2.80fF
C184 a_73259_n13437# gnd 3.33fF
C185 a_74303_n12585# gnd 2.33fF
C186 a_71765_n12582# gnd 3.27fF
C187 a_66533_n13393# gnd 3.33fF
C188 a_67581_n12718# gnd 3.73fF
C189 a_76412_n12641# gnd 2.27fF
C190 a_65704_n13030# gnd 3.17fF
C191 a_66533_n12714# gnd 2.80fF
C192 a_62294_n13441# gnd 3.33fF
C193 a_63338_n12589# gnd 2.33fF
C194 a_60800_n12586# gnd 3.27fF
C195 a_55568_n13397# gnd 3.33fF
C196 a_56616_n12722# gnd 3.73fF
C197 a_65704_n12635# gnd 2.27fF
C198 a_54739_n13034# gnd 3.17fF
C199 a_55568_n12718# gnd 2.80fF
C200 a_51586_n13435# gnd 3.33fF
C201 a_52630_n12583# gnd 2.33fF
C202 a_50092_n12580# gnd 3.27fF
C203 a_44860_n13391# gnd 3.33fF
C204 a_45908_n12716# gnd 3.73fF
C205 a_54739_n12639# gnd 2.27fF
C206 a_44031_n13028# gnd 3.17fF
C207 a_44860_n12712# gnd 2.80fF
C208 a_40835_n13443# gnd 3.33fF
C209 a_41879_n12591# gnd 2.33fF
C210 a_39341_n12588# gnd 3.27fF
C211 a_34109_n13399# gnd 3.33fF
C212 a_35157_n12724# gnd 3.73fF
C213 a_44031_n12633# gnd 2.27fF
C214 a_33280_n13036# gnd 3.17fF
C215 a_34109_n12720# gnd 2.80fF
C216 a_30127_n13437# gnd 3.33fF
C217 a_31171_n12585# gnd 2.33fF
C218 a_28633_n12582# gnd 3.27fF
C219 a_23401_n13393# gnd 3.33fF
C220 a_24449_n12718# gnd 3.73fF
C221 a_33280_n12641# gnd 2.27fF
C222 a_22572_n13030# gnd 3.17fF
C223 a_23401_n12714# gnd 2.80fF
C224 a_19162_n13441# gnd 3.33fF
C225 a_20206_n12589# gnd 2.33fF
C226 a_17668_n12586# gnd 3.27fF
C227 a_12436_n13397# gnd 3.33fF
C228 a_13484_n12722# gnd 3.73fF
C229 a_22572_n12635# gnd 2.27fF
C230 a_11607_n13034# gnd 3.17fF
C231 a_12436_n12718# gnd 2.80fF
C232 a_8454_n13435# gnd 3.33fF
C233 a_9498_n12583# gnd 2.33fF
C234 a_6960_n12580# gnd 3.27fF
C235 a_1728_n13391# gnd 3.33fF
C236 a_2776_n12716# gnd 3.73fF
C237 a_11607_n12639# gnd 2.27fF
C238 a_899_n13028# gnd 3.17fF
C239 a_1728_n12712# gnd 2.80fF
C240 a_899_n12633# gnd 2.27fF
C241 a_85015_n12768# gnd 3.52fF
C242 a_74307_n12762# gnd 3.52fF
C243 a_63342_n12766# gnd 3.52fF
C244 a_52634_n12760# gnd 3.52fF
C245 a_41883_n12768# gnd 3.52fF
C246 a_31175_n12762# gnd 3.52fF
C247 a_85010_n11750# gnd 2.27fF
C248 a_83962_n11746# gnd 2.80fF
C249 a_79679_n11882# gnd 3.19fF
C250 a_76412_n12385# gnd 3.52fF
C251 a_74302_n11744# gnd 2.27fF
C252 a_73254_n11740# gnd 2.80fF
C253 a_68971_n11876# gnd 3.19fF
C254 a_20210_n12766# gnd 3.52fF
C255 a_9502_n12760# gnd 3.52fF
C256 a_76411_n11771# gnd 2.33fF
C257 a_65704_n12379# gnd 3.52fF
C258 a_63337_n11748# gnd 2.27fF
C259 a_62289_n11744# gnd 2.80fF
C260 a_58006_n11880# gnd 3.19fF
C261 a_65703_n11765# gnd 2.33fF
C262 a_54739_n12383# gnd 3.52fF
C263 a_52629_n11742# gnd 2.27fF
C264 a_51581_n11738# gnd 2.80fF
C265 a_47298_n11874# gnd 3.19fF
C266 a_54738_n11769# gnd 2.33fF
C267 a_44031_n12377# gnd 3.52fF
C268 a_41878_n11750# gnd 2.27fF
C269 a_40830_n11746# gnd 2.80fF
C270 a_36547_n11882# gnd 3.19fF
C271 a_33280_n12385# gnd 3.52fF
C272 a_31170_n11744# gnd 2.27fF
C273 a_30122_n11740# gnd 2.80fF
C274 a_25839_n11876# gnd 3.19fF
C275 a_44030_n11763# gnd 2.33fF
C276 a_33279_n11771# gnd 2.33fF
C277 a_22572_n12379# gnd 3.52fF
C278 a_20205_n11748# gnd 2.27fF
C279 a_19157_n11744# gnd 2.80fF
C280 a_14874_n11880# gnd 3.19fF
C281 a_22571_n11765# gnd 2.33fF
C282 a_11607_n12383# gnd 3.52fF
C283 a_9497_n11742# gnd 2.27fF
C284 a_8449_n11738# gnd 2.80fF
C285 a_4166_n11874# gnd 3.19fF
C286 a_11606_n11769# gnd 2.33fF
C287 a_899_n12377# gnd 3.52fF
C288 a_898_n11763# gnd 2.33fF
C289 a_85014_n11927# gnd 3.17fF
C290 a_74306_n11921# gnd 3.17fF
C291 a_63341_n11925# gnd 3.17fF
C292 a_52633_n11919# gnd 3.17fF
C293 a_41882_n11927# gnd 3.17fF
C294 a_31174_n11921# gnd 3.17fF
C295 a_83966_n11923# gnd 3.33fF
C296 a_85010_n11071# gnd 2.33fF
C297 a_82477_n12765# gnd 3.19fF
C298 a_82515_n11066# gnd 3.65fF
C299 a_77240_n11879# gnd 3.33fF
C300 a_20209_n11925# gnd 3.17fF
C301 a_9501_n11919# gnd 3.17fF
C302 a_76411_n11516# gnd 3.17fF
C303 a_77240_n11200# gnd 2.80fF
C304 a_73258_n11917# gnd 3.33fF
C305 a_74302_n11065# gnd 2.33fF
C306 a_71769_n12759# gnd 3.19fF
C307 a_71807_n11060# gnd 3.65fF
C308 a_66532_n11873# gnd 3.33fF
C309 a_76411_n11121# gnd 2.27fF
C310 a_65703_n11510# gnd 3.17fF
C311 a_66532_n11194# gnd 2.80fF
C312 a_62293_n11921# gnd 3.33fF
C313 a_63337_n11069# gnd 2.33fF
C314 a_60804_n12763# gnd 3.19fF
C315 a_60842_n11064# gnd 3.65fF
C316 a_55567_n11877# gnd 3.33fF
C317 a_65703_n11115# gnd 2.27fF
C318 a_54738_n11514# gnd 3.17fF
C319 a_55567_n11198# gnd 2.80fF
C320 a_51585_n11915# gnd 3.33fF
C321 a_52629_n11063# gnd 2.33fF
C322 a_50096_n12757# gnd 3.19fF
C323 a_50134_n11058# gnd 3.65fF
C324 a_44859_n11871# gnd 3.33fF
C325 a_54738_n11119# gnd 2.27fF
C326 a_44030_n11508# gnd 3.17fF
C327 a_44859_n11192# gnd 2.80fF
C328 a_40834_n11923# gnd 3.33fF
C329 a_41878_n11071# gnd 2.33fF
C330 a_39345_n12765# gnd 3.19fF
C331 a_39383_n11066# gnd 3.65fF
C332 a_34108_n11879# gnd 3.33fF
C333 a_44030_n11113# gnd 2.27fF
C334 a_33279_n11516# gnd 3.17fF
C335 a_34108_n11200# gnd 2.80fF
C336 a_30126_n11917# gnd 3.33fF
C337 a_31170_n11065# gnd 2.33fF
C338 a_28637_n12759# gnd 3.19fF
C339 a_28675_n11060# gnd 3.65fF
C340 a_23400_n11873# gnd 3.33fF
C341 a_33279_n11121# gnd 2.27fF
C342 a_22571_n11510# gnd 3.17fF
C343 a_23400_n11194# gnd 2.80fF
C344 a_19161_n11921# gnd 3.33fF
C345 a_20205_n11069# gnd 2.33fF
C346 a_17672_n12763# gnd 3.19fF
C347 a_17710_n11064# gnd 3.65fF
C348 a_12435_n11877# gnd 3.33fF
C349 a_22571_n11115# gnd 2.27fF
C350 a_11606_n11514# gnd 3.17fF
C351 a_12435_n11198# gnd 2.80fF
C352 a_8453_n11915# gnd 3.33fF
C353 a_9497_n11063# gnd 2.33fF
C354 a_6964_n12757# gnd 3.19fF
C355 a_7002_n11058# gnd 3.65fF
C356 a_1727_n11871# gnd 3.33fF
C357 a_11606_n11119# gnd 2.27fF
C358 a_898_n11508# gnd 3.17fF
C359 a_1727_n11192# gnd 2.80fF
C360 a_898_n11113# gnd 2.27fF
C361 a_85014_n11248# gnd 3.43fF
C362 a_74306_n11242# gnd 3.43fF
C363 a_63341_n11246# gnd 3.43fF
C364 a_52633_n11240# gnd 3.43fF
C365 a_41882_n11248# gnd 3.43fF
C366 a_31174_n11242# gnd 3.43fF
C367 a_85010_n10303# gnd 2.27fF
C368 a_82519_n11243# gnd 3.20fF
C369 a_83962_n10299# gnd 2.80fF
C370 a_78288_n11204# gnd 3.43fF
C371 a_79684_n11763# gnd 3.27fF
C372 a_76411_n10865# gnd 3.43fF
C373 a_74302_n10297# gnd 2.27fF
C374 a_71811_n11237# gnd 3.20fF
C375 a_73254_n10293# gnd 2.80fF
C376 a_67580_n11198# gnd 3.43fF
C377 a_68976_n11757# gnd 3.27fF
C378 a_20209_n11246# gnd 3.43fF
C379 a_9501_n11240# gnd 3.43fF
C380 a_76411_n10324# gnd 2.33fF
C381 a_65703_n10859# gnd 3.43fF
C382 a_63337_n10301# gnd 2.27fF
C383 a_60846_n11241# gnd 3.20fF
C384 a_62289_n10297# gnd 2.80fF
C385 a_56615_n11202# gnd 3.43fF
C386 a_58011_n11761# gnd 3.27fF
C387 a_65703_n10318# gnd 2.33fF
C388 a_54738_n10863# gnd 3.43fF
C389 a_52629_n10295# gnd 2.27fF
C390 a_50138_n11235# gnd 3.20fF
C391 a_51581_n10291# gnd 2.80fF
C392 a_45907_n11196# gnd 3.43fF
C393 a_47303_n11755# gnd 3.27fF
C394 a_54738_n10322# gnd 2.33fF
C395 a_44030_n10857# gnd 3.43fF
C396 a_41878_n10303# gnd 2.27fF
C397 a_39387_n11243# gnd 3.20fF
C398 a_40830_n10299# gnd 2.80fF
C399 a_35156_n11204# gnd 3.43fF
C400 a_36552_n11763# gnd 3.27fF
C401 a_33279_n10865# gnd 3.43fF
C402 a_31170_n10297# gnd 2.27fF
C403 a_28679_n11237# gnd 3.20fF
C404 a_30122_n10293# gnd 2.80fF
C405 a_24448_n11198# gnd 3.43fF
C406 a_25844_n11757# gnd 3.27fF
C407 a_44030_n10316# gnd 2.33fF
C408 a_33279_n10324# gnd 2.33fF
C409 a_22571_n10859# gnd 3.43fF
C410 a_20205_n10301# gnd 2.27fF
C411 a_17714_n11241# gnd 3.20fF
C412 a_19157_n10297# gnd 2.80fF
C413 a_13483_n11202# gnd 3.43fF
C414 a_14879_n11761# gnd 3.27fF
C415 a_22571_n10318# gnd 2.33fF
C416 a_11606_n10863# gnd 3.43fF
C417 a_9497_n10295# gnd 2.27fF
C418 a_7006_n11235# gnd 3.20fF
C419 a_8449_n10291# gnd 2.80fF
C420 a_2775_n11196# gnd 3.43fF
C421 a_4171_n11755# gnd 3.27fF
C422 a_11606_n10322# gnd 2.33fF
C423 a_898_n10857# gnd 3.43fF
C424 a_898_n10316# gnd 2.33fF
C425 a_85014_n10480# gnd 3.17fF
C426 a_74306_n10474# gnd 3.17fF
C427 a_63341_n10478# gnd 3.17fF
C428 a_52633_n10472# gnd 3.17fF
C429 a_41882_n10480# gnd 3.17fF
C430 a_31174_n10474# gnd 3.17fF
C431 a_83966_n10476# gnd 3.33fF
C432 a_85010_n9624# gnd 2.33fF
C433 a_81407_n9615# gnd 7.02fF
C434 a_77240_n10432# gnd 3.33fF
C435 a_78288_n9757# gnd 4.35fF
C436 a_20209_n10478# gnd 3.17fF
C437 a_9501_n10472# gnd 3.17fF
C438 a_76411_n10069# gnd 3.17fF
C439 a_77240_n9753# gnd 2.80fF
C440 a_73258_n10470# gnd 3.33fF
C441 a_74302_n9618# gnd 2.33fF
C442 a_70699_n9609# gnd 7.02fF
C443 a_66532_n10426# gnd 3.33fF
C444 a_67580_n9751# gnd 4.35fF
C445 a_76411_n9674# gnd 2.27fF
C446 a_65703_n10063# gnd 3.17fF
C447 a_66532_n9747# gnd 2.80fF
C448 a_62293_n10474# gnd 3.33fF
C449 a_63337_n9622# gnd 2.33fF
C450 a_59734_n9613# gnd 7.02fF
C451 a_55567_n10430# gnd 3.33fF
C452 a_56615_n9755# gnd 4.35fF
C453 a_65703_n9668# gnd 2.27fF
C454 a_54738_n10067# gnd 3.17fF
C455 a_55567_n9751# gnd 2.80fF
C456 a_51585_n10468# gnd 3.33fF
C457 a_52629_n9616# gnd 2.33fF
C458 a_49026_n9607# gnd 7.02fF
C459 a_44859_n10424# gnd 3.33fF
C460 a_45907_n9749# gnd 4.35fF
C461 a_54738_n9672# gnd 2.27fF
C462 a_44030_n10061# gnd 3.17fF
C463 a_44859_n9745# gnd 2.80fF
C464 a_40834_n10476# gnd 3.33fF
C465 a_41878_n9624# gnd 2.33fF
C466 a_38275_n9615# gnd 7.02fF
C467 a_34108_n10432# gnd 3.33fF
C468 a_35156_n9757# gnd 4.35fF
C469 a_44030_n9666# gnd 2.27fF
C470 a_33279_n10069# gnd 3.17fF
C471 a_34108_n9753# gnd 2.80fF
C472 a_30126_n10470# gnd 3.33fF
C473 a_31170_n9618# gnd 2.33fF
C474 a_27567_n9609# gnd 7.02fF
C475 a_23400_n10426# gnd 3.33fF
C476 a_24448_n9751# gnd 4.35fF
C477 a_33279_n9674# gnd 2.27fF
C478 a_22571_n10063# gnd 3.17fF
C479 a_23400_n9747# gnd 2.80fF
C480 a_19161_n10474# gnd 3.33fF
C481 a_20205_n9622# gnd 2.33fF
C482 a_16602_n9613# gnd 7.02fF
C483 a_12435_n10430# gnd 3.33fF
C484 a_13483_n9755# gnd 4.35fF
C485 a_22571_n9668# gnd 2.27fF
C486 a_11606_n10067# gnd 3.17fF
C487 a_12435_n9751# gnd 2.80fF
C488 a_8453_n10468# gnd 3.33fF
C489 a_9497_n9616# gnd 2.33fF
C490 a_5894_n9607# gnd 7.02fF
C491 a_1727_n10424# gnd 3.33fF
C492 a_2775_n9749# gnd 4.35fF
C493 a_11606_n9672# gnd 2.27fF
C494 a_898_n10061# gnd 3.17fF
C495 a_1727_n9745# gnd 2.80fF
C496 a_898_n9666# gnd 2.27fF
C497 a_85014_n9801# gnd 3.62fF
C498 a_74306_n9795# gnd 3.62fF
C499 a_63341_n9799# gnd 3.62fF
C500 a_52633_n9793# gnd 3.62fF
C501 a_41882_n9801# gnd 3.62fF
C502 a_31174_n9795# gnd 3.62fF
C503 a_85013_n8709# gnd 2.27fF
C504 a_83965_n8705# gnd 2.80fF
C505 a_79778_n11882# gnd 4.90fF
C506 a_76411_n9418# gnd 3.62fF
C507 a_74305_n8703# gnd 2.27fF
C508 a_73257_n8699# gnd 2.80fF
C509 a_69070_n11876# gnd 4.90fF
C510 a_20209_n9799# gnd 3.62fF
C511 a_9501_n9793# gnd 3.62fF
C512 a_76414_n8730# gnd 2.33fF
C513 a_65703_n9412# gnd 3.62fF
C514 a_63340_n8707# gnd 2.27fF
C515 a_62292_n8703# gnd 2.80fF
C516 a_58105_n11880# gnd 4.90fF
C517 a_65706_n8724# gnd 2.33fF
C518 a_54738_n9416# gnd 3.62fF
C519 a_52632_n8701# gnd 2.27fF
C520 a_51584_n8697# gnd 2.80fF
C521 a_47397_n11874# gnd 4.90fF
C522 a_54741_n8728# gnd 2.33fF
C523 a_44030_n9410# gnd 3.62fF
C524 a_41881_n8709# gnd 2.27fF
C525 a_40833_n8705# gnd 2.80fF
C526 a_36646_n11882# gnd 4.90fF
C527 a_33279_n9418# gnd 3.62fF
C528 a_31173_n8703# gnd 2.27fF
C529 a_30125_n8699# gnd 2.80fF
C530 a_25938_n11876# gnd 4.90fF
C531 a_44033_n8722# gnd 2.33fF
C532 a_33282_n8730# gnd 2.33fF
C533 a_22571_n9412# gnd 3.62fF
C534 a_20208_n8707# gnd 2.27fF
C535 a_19160_n8703# gnd 2.80fF
C536 a_14973_n11880# gnd 4.90fF
C537 a_22574_n8724# gnd 2.33fF
C538 a_11606_n9416# gnd 3.62fF
C539 a_9500_n8701# gnd 2.27fF
C540 a_8452_n8697# gnd 2.80fF
C541 a_4265_n11874# gnd 4.90fF
C542 a_11609_n8728# gnd 2.33fF
C543 a_898_n9410# gnd 3.62fF
C544 a_901_n8722# gnd 2.33fF
C545 a_85017_n8886# gnd 3.17fF
C546 a_74309_n8880# gnd 3.17fF
C547 a_63344_n8884# gnd 3.17fF
C548 a_52636_n8878# gnd 3.17fF
C549 a_41885_n8886# gnd 3.17fF
C550 a_31177_n8880# gnd 3.17fF
C551 a_83969_n8882# gnd 3.33fF
C552 a_85013_n8030# gnd 2.33fF
C553 a_82518_n8025# gnd 4.35fF
C554 a_77243_n8838# gnd 3.33fF
C555 a_20212_n8884# gnd 3.17fF
C556 a_9504_n8878# gnd 3.17fF
C557 a_76414_n8475# gnd 3.17fF
C558 a_77243_n8159# gnd 2.80fF
C559 a_73261_n8876# gnd 3.33fF
C560 a_74305_n8024# gnd 2.33fF
C561 a_71810_n8019# gnd 4.35fF
C562 a_66535_n8832# gnd 3.33fF
C563 a_76414_n8080# gnd 2.27fF
C564 a_65706_n8469# gnd 3.17fF
C565 a_66535_n8153# gnd 2.80fF
C566 a_62296_n8880# gnd 3.33fF
C567 a_63340_n8028# gnd 2.33fF
C568 a_60845_n8023# gnd 4.35fF
C569 a_55570_n8836# gnd 3.33fF
C570 a_65706_n8074# gnd 2.27fF
C571 a_54741_n8473# gnd 3.17fF
C572 a_55570_n8157# gnd 2.80fF
C573 a_51588_n8874# gnd 3.33fF
C574 a_52632_n8022# gnd 2.33fF
C575 a_50137_n8017# gnd 4.35fF
C576 a_44862_n8830# gnd 3.33fF
C577 a_54741_n8078# gnd 2.27fF
C578 a_44033_n8467# gnd 3.17fF
C579 a_44862_n8151# gnd 2.80fF
C580 a_40837_n8882# gnd 3.33fF
C581 a_41881_n8030# gnd 2.33fF
C582 a_39386_n8025# gnd 4.35fF
C583 a_34111_n8838# gnd 3.33fF
C584 a_44033_n8072# gnd 2.27fF
C585 a_33282_n8475# gnd 3.17fF
C586 a_34111_n8159# gnd 2.80fF
C587 a_30129_n8876# gnd 3.33fF
C588 a_31173_n8024# gnd 2.33fF
C589 a_28678_n8019# gnd 4.35fF
C590 a_23403_n8832# gnd 3.33fF
C591 a_33282_n8080# gnd 2.27fF
C592 a_22574_n8469# gnd 3.17fF
C593 a_23403_n8153# gnd 2.80fF
C594 a_19164_n8880# gnd 3.33fF
C595 a_20208_n8028# gnd 2.33fF
C596 a_17713_n8023# gnd 4.35fF
C597 a_12438_n8836# gnd 3.33fF
C598 a_22574_n8074# gnd 2.27fF
C599 a_11609_n8473# gnd 3.17fF
C600 a_12438_n8157# gnd 2.80fF
C601 a_8456_n8874# gnd 3.33fF
C602 a_9500_n8022# gnd 2.33fF
C603 a_7005_n8017# gnd 4.35fF
C604 a_1730_n8830# gnd 3.33fF
C605 a_11609_n8078# gnd 2.27fF
C606 a_901_n8467# gnd 3.17fF
C607 a_1730_n8151# gnd 2.80fF
C608 a_901_n8072# gnd 2.27fF
C609 a_85017_n8207# gnd 3.43fF
C610 a_74309_n8201# gnd 3.43fF
C611 a_63344_n8205# gnd 3.43fF
C612 a_52636_n8199# gnd 3.43fF
C613 a_41885_n8207# gnd 3.43fF
C614 a_31177_n8201# gnd 3.43fF
C615 a_85013_n7262# gnd 2.27fF
C616 a_82522_n8202# gnd 3.43fF
C617 a_83965_n7258# gnd 2.80fF
C618 a_78291_n8163# gnd 3.20fF
C619 a_76414_n7824# gnd 3.43fF
C620 a_74305_n7256# gnd 2.27fF
C621 a_71814_n8196# gnd 3.43fF
C622 a_73257_n7252# gnd 2.80fF
C623 a_67583_n8157# gnd 3.20fF
C624 a_20212_n8205# gnd 3.43fF
C625 a_9504_n8199# gnd 3.43fF
C626 a_76414_n7283# gnd 2.33fF
C627 a_65706_n7818# gnd 3.43fF
C628 a_63340_n7260# gnd 2.27fF
C629 a_60849_n8200# gnd 3.43fF
C630 a_62292_n7256# gnd 2.80fF
C631 a_56618_n8161# gnd 3.20fF
C632 a_65706_n7277# gnd 2.33fF
C633 a_54741_n7822# gnd 3.43fF
C634 a_52632_n7254# gnd 2.27fF
C635 a_50141_n8194# gnd 3.43fF
C636 a_51584_n7250# gnd 2.80fF
C637 a_45910_n8155# gnd 3.20fF
C638 a_54741_n7281# gnd 2.33fF
C639 a_44033_n7816# gnd 3.43fF
C640 a_41881_n7262# gnd 2.27fF
C641 a_39390_n8202# gnd 3.43fF
C642 a_40833_n7258# gnd 2.80fF
C643 a_35159_n8163# gnd 3.20fF
C644 a_33282_n7824# gnd 3.43fF
C645 a_31173_n7256# gnd 2.27fF
C646 a_28682_n8196# gnd 3.43fF
C647 a_30125_n7252# gnd 2.80fF
C648 a_24451_n8157# gnd 3.20fF
C649 a_44033_n7275# gnd 2.33fF
C650 a_33282_n7283# gnd 2.33fF
C651 a_22574_n7818# gnd 3.43fF
C652 a_20208_n7260# gnd 2.27fF
C653 a_17717_n8200# gnd 3.43fF
C654 a_19160_n7256# gnd 2.80fF
C655 a_13486_n8161# gnd 3.20fF
C656 a_22574_n7277# gnd 2.33fF
C657 a_11609_n7822# gnd 3.43fF
C658 a_9500_n7254# gnd 2.27fF
C659 a_7009_n8194# gnd 3.43fF
C660 a_8452_n7250# gnd 2.80fF
C661 a_2778_n8155# gnd 3.20fF
C662 a_11609_n7281# gnd 2.33fF
C663 a_901_n7816# gnd 3.43fF
C664 a_901_n7275# gnd 2.33fF
C665 a_85017_n7439# gnd 3.17fF
C666 a_74309_n7433# gnd 3.17fF
C667 a_63344_n7437# gnd 3.17fF
C668 a_52636_n7431# gnd 3.17fF
C669 a_41885_n7439# gnd 3.17fF
C670 a_31177_n7433# gnd 3.17fF
C671 a_83969_n7435# gnd 3.33fF
C672 a_85013_n6583# gnd 2.33fF
C673 a_81411_n9792# gnd 4.97fF
C674 a_82475_n6580# gnd 3.27fF
C675 a_77243_n7391# gnd 3.33fF
C676 a_78291_n6716# gnd 3.65fF
C677 a_20212_n7437# gnd 3.17fF
C678 a_9504_n7431# gnd 3.17fF
C679 a_76414_n7028# gnd 3.17fF
C680 a_77243_n6712# gnd 2.80fF
C681 a_73261_n7429# gnd 3.33fF
C682 a_74305_n6577# gnd 2.33fF
C683 a_70703_n9786# gnd 4.97fF
C684 a_71767_n6574# gnd 3.27fF
C685 a_66535_n7385# gnd 3.33fF
C686 a_67583_n6710# gnd 3.65fF
C687 a_76414_n6633# gnd 2.27fF
C688 a_65706_n7022# gnd 3.17fF
C689 a_66535_n6706# gnd 2.80fF
C690 a_62296_n7433# gnd 3.33fF
C691 a_63340_n6581# gnd 2.33fF
C692 a_59738_n9790# gnd 4.97fF
C693 a_60802_n6578# gnd 3.27fF
C694 a_55570_n7389# gnd 3.33fF
C695 a_56618_n6714# gnd 3.65fF
C696 a_65706_n6627# gnd 2.27fF
C697 a_54741_n7026# gnd 3.17fF
C698 a_55570_n6710# gnd 2.80fF
C699 a_51588_n7427# gnd 3.33fF
C700 a_52632_n6575# gnd 2.33fF
C701 a_49030_n9784# gnd 4.97fF
C702 a_50094_n6572# gnd 3.27fF
C703 a_44862_n7383# gnd 3.33fF
C704 a_45910_n6708# gnd 3.65fF
C705 a_54741_n6631# gnd 2.27fF
C706 a_44033_n7020# gnd 3.17fF
C707 a_44862_n6704# gnd 2.80fF
C708 a_40837_n7435# gnd 3.33fF
C709 a_41881_n6583# gnd 2.33fF
C710 a_38279_n9792# gnd 4.97fF
C711 a_39343_n6580# gnd 3.27fF
C712 a_34111_n7391# gnd 3.33fF
C713 a_35159_n6716# gnd 3.65fF
C714 a_44033_n6625# gnd 2.27fF
C715 a_33282_n7028# gnd 3.17fF
C716 a_34111_n6712# gnd 2.80fF
C717 a_30129_n7429# gnd 3.33fF
C718 a_31173_n6577# gnd 2.33fF
C719 a_27571_n9786# gnd 4.97fF
C720 a_28635_n6574# gnd 3.27fF
C721 a_23403_n7385# gnd 3.33fF
C722 a_24451_n6710# gnd 3.65fF
C723 a_33282_n6633# gnd 2.27fF
C724 a_22574_n7022# gnd 3.17fF
C725 a_23403_n6706# gnd 2.80fF
C726 a_19164_n7433# gnd 3.33fF
C727 a_20208_n6581# gnd 2.33fF
C728 a_16606_n9790# gnd 4.97fF
C729 a_17670_n6578# gnd 3.27fF
C730 a_12438_n7389# gnd 3.33fF
C731 a_13486_n6714# gnd 3.65fF
C732 a_22574_n6627# gnd 2.27fF
C733 a_11609_n7026# gnd 3.17fF
C734 a_12438_n6710# gnd 2.80fF
C735 a_8456_n7427# gnd 3.33fF
C736 a_9500_n6575# gnd 2.33fF
C737 a_5898_n9784# gnd 4.97fF
C738 a_6962_n6572# gnd 3.27fF
C739 a_1730_n7383# gnd 3.33fF
C740 a_2778_n6708# gnd 3.65fF
C741 a_11609_n6631# gnd 2.27fF
C742 a_901_n7020# gnd 3.17fF
C743 a_1730_n6704# gnd 2.80fF
C744 a_901_n6625# gnd 2.27fF
C745 a_85017_n6760# gnd 3.52fF
C746 a_74309_n6754# gnd 3.52fF
C747 a_63344_n6758# gnd 3.52fF
C748 a_52636_n6752# gnd 3.52fF
C749 a_85012_n5742# gnd 2.27fF
C750 a_83964_n5738# gnd 2.80fF
C751 a_80846_n8847# gnd 4.30fF
C752 a_81062_n5744# gnd 4.72fF
C753 a_79681_n5874# gnd 3.19fF
C754 a_79780_n5874# gnd 7.03fF
C755 a_76414_n6377# gnd 3.52fF
C756 a_41885_n6760# gnd 3.52fF
C757 a_31177_n6754# gnd 3.52fF
C758 a_74304_n5736# gnd 2.27fF
C759 a_73256_n5732# gnd 2.80fF
C760 a_70138_n8841# gnd 4.30fF
C761 a_70354_n5738# gnd 4.72fF
C762 a_76413_n5763# gnd 2.33fF
C763 a_68973_n5868# gnd 3.19fF
C764 a_69072_n5868# gnd 7.03fF
C765 a_65706_n6371# gnd 3.52fF
C766 a_63339_n5740# gnd 2.27fF
C767 a_62291_n5736# gnd 2.80fF
C768 a_59173_n8845# gnd 4.30fF
C769 a_59389_n5742# gnd 4.72fF
C770 a_65705_n5757# gnd 2.33fF
C771 a_58008_n5872# gnd 3.19fF
C772 a_58107_n5872# gnd 7.03fF
C773 a_54741_n6375# gnd 3.52fF
C774 a_20212_n6758# gnd 3.52fF
C775 a_9504_n6752# gnd 3.52fF
C776 a_52631_n5734# gnd 2.27fF
C777 a_51583_n5730# gnd 2.80fF
C778 a_48465_n8839# gnd 4.30fF
C779 a_48681_n5736# gnd 4.72fF
C780 a_54740_n5761# gnd 2.33fF
C781 a_47300_n5866# gnd 3.19fF
C782 a_47399_n5866# gnd 7.03fF
C783 a_44033_n6369# gnd 3.52fF
C784 a_41880_n5742# gnd 2.27fF
C785 a_40832_n5738# gnd 2.80fF
C786 a_37714_n8847# gnd 4.30fF
C787 a_37930_n5744# gnd 4.72fF
C788 a_44032_n5755# gnd 2.33fF
C789 a_36549_n5874# gnd 3.19fF
C790 a_36648_n5874# gnd 7.03fF
C791 a_33282_n6377# gnd 3.52fF
C792 a_31172_n5736# gnd 2.27fF
C793 a_30124_n5732# gnd 2.80fF
C794 a_27006_n8841# gnd 4.30fF
C795 a_27222_n5738# gnd 4.72fF
C796 a_33281_n5763# gnd 2.33fF
C797 a_25841_n5868# gnd 3.19fF
C798 a_25940_n5868# gnd 7.03fF
C799 a_22574_n6371# gnd 3.52fF
C800 a_20207_n5740# gnd 2.27fF
C801 a_19159_n5736# gnd 2.80fF
C802 a_16041_n8845# gnd 4.30fF
C803 a_16257_n5742# gnd 4.72fF
C804 a_22573_n5757# gnd 2.33fF
C805 a_14876_n5872# gnd 3.19fF
C806 a_14975_n5872# gnd 7.03fF
C807 a_11609_n6375# gnd 3.52fF
C808 a_9499_n5734# gnd 2.27fF
C809 a_8451_n5730# gnd 2.80fF
C810 a_5333_n8839# gnd 4.30fF
C811 a_5549_n5736# gnd 4.72fF
C812 a_11608_n5761# gnd 2.33fF
C813 a_4168_n5866# gnd 3.19fF
C814 a_4267_n5866# gnd 7.03fF
C815 a_901_n6369# gnd 3.52fF
C816 a_900_n5755# gnd 2.33fF
C817 a_85016_n5919# gnd 3.17fF
C818 a_74308_n5913# gnd 3.17fF
C819 a_63343_n5917# gnd 3.17fF
C820 a_52635_n5911# gnd 3.17fF
C821 a_41884_n5919# gnd 3.17fF
C822 a_31176_n5913# gnd 3.17fF
C823 a_83968_n5915# gnd 3.33fF
C824 a_85012_n5063# gnd 2.33fF
C825 a_82479_n6757# gnd 3.19fF
C826 a_82517_n5058# gnd 3.64fF
C827 a_77242_n5871# gnd 3.33fF
C828 a_20211_n5917# gnd 3.17fF
C829 a_9503_n5911# gnd 3.17fF
C830 a_76413_n5508# gnd 3.17fF
C831 a_77242_n5192# gnd 2.80fF
C832 a_73260_n5909# gnd 3.33fF
C833 a_74304_n5057# gnd 2.33fF
C834 a_71771_n6751# gnd 3.19fF
C835 a_71809_n5052# gnd 3.64fF
C836 a_66534_n5865# gnd 3.33fF
C837 a_76413_n5113# gnd 2.27fF
C838 a_65705_n5502# gnd 3.17fF
C839 a_66534_n5186# gnd 2.80fF
C840 a_62295_n5913# gnd 3.33fF
C841 a_63339_n5061# gnd 2.33fF
C842 a_60806_n6755# gnd 3.19fF
C843 a_60844_n5056# gnd 3.64fF
C844 a_55569_n5869# gnd 3.33fF
C845 a_65705_n5107# gnd 2.27fF
C846 a_54740_n5506# gnd 3.17fF
C847 a_55569_n5190# gnd 2.80fF
C848 a_51587_n5907# gnd 3.33fF
C849 a_52631_n5055# gnd 2.33fF
C850 a_50098_n6749# gnd 3.19fF
C851 a_50136_n5050# gnd 3.64fF
C852 a_44861_n5863# gnd 3.33fF
C853 a_54740_n5111# gnd 2.27fF
C854 a_44032_n5500# gnd 3.17fF
C855 a_44861_n5184# gnd 2.80fF
C856 a_40836_n5915# gnd 3.33fF
C857 a_41880_n5063# gnd 2.33fF
C858 a_39347_n6757# gnd 3.19fF
C859 a_39385_n5058# gnd 3.64fF
C860 a_34110_n5871# gnd 3.33fF
C861 a_44032_n5105# gnd 2.27fF
C862 a_33281_n5508# gnd 3.17fF
C863 a_34110_n5192# gnd 2.80fF
C864 a_30128_n5909# gnd 3.33fF
C865 a_31172_n5057# gnd 2.33fF
C866 a_28639_n6751# gnd 3.19fF
C867 a_28677_n5052# gnd 3.64fF
C868 a_23402_n5865# gnd 3.33fF
C869 a_33281_n5113# gnd 2.27fF
C870 a_22573_n5502# gnd 3.17fF
C871 a_23402_n5186# gnd 2.80fF
C872 a_19163_n5913# gnd 3.33fF
C873 a_20207_n5061# gnd 2.33fF
C874 a_17674_n6755# gnd 3.19fF
C875 a_17712_n5056# gnd 3.64fF
C876 a_12437_n5869# gnd 3.33fF
C877 a_22573_n5107# gnd 2.27fF
C878 a_11608_n5506# gnd 3.17fF
C879 a_12437_n5190# gnd 2.80fF
C880 a_8455_n5907# gnd 3.33fF
C881 a_9499_n5055# gnd 2.33fF
C882 a_6966_n6749# gnd 3.19fF
C883 a_7004_n5050# gnd 3.64fF
C884 a_1729_n5863# gnd 3.33fF
C885 a_11608_n5111# gnd 2.27fF
C886 a_900_n5500# gnd 3.17fF
C887 a_1729_n5184# gnd 2.80fF
C888 a_900_n5105# gnd 2.27fF
C889 a_85016_n5240# gnd 3.43fF
C890 a_74308_n5234# gnd 3.43fF
C891 a_63343_n5238# gnd 3.43fF
C892 a_52635_n5232# gnd 3.43fF
C893 a_41884_n5240# gnd 3.43fF
C894 a_31176_n5234# gnd 3.43fF
C895 a_85012_n4295# gnd 2.27fF
C896 a_82521_n5235# gnd 3.16fF
C897 a_83964_n4291# gnd 2.80fF
C898 a_78290_n5196# gnd 3.43fF
C899 a_79686_n5755# gnd 3.27fF
C900 a_76413_n4857# gnd 3.43fF
C901 a_74304_n4289# gnd 2.27fF
C902 a_71813_n5229# gnd 3.16fF
C903 a_73256_n4285# gnd 2.80fF
C904 a_67582_n5190# gnd 3.43fF
C905 a_68978_n5749# gnd 3.27fF
C906 a_20211_n5238# gnd 3.43fF
C907 a_9503_n5232# gnd 3.43fF
C908 a_76413_n4316# gnd 2.33fF
C909 a_65705_n4851# gnd 3.43fF
C910 a_63339_n4293# gnd 2.27fF
C911 a_60848_n5233# gnd 3.16fF
C912 a_62291_n4289# gnd 2.80fF
C913 a_56617_n5194# gnd 3.43fF
C914 a_58013_n5753# gnd 3.27fF
C915 a_65705_n4310# gnd 2.33fF
C916 a_54740_n4855# gnd 3.43fF
C917 a_52631_n4287# gnd 2.27fF
C918 a_50140_n5227# gnd 3.16fF
C919 a_51583_n4283# gnd 2.80fF
C920 a_45909_n5188# gnd 3.43fF
C921 a_47305_n5747# gnd 3.27fF
C922 a_54740_n4314# gnd 2.33fF
C923 a_44032_n4849# gnd 3.43fF
C924 a_41880_n4295# gnd 2.27fF
C925 a_39389_n5235# gnd 3.16fF
C926 a_40832_n4291# gnd 2.80fF
C927 a_35158_n5196# gnd 3.43fF
C928 a_36554_n5755# gnd 3.27fF
C929 a_33281_n4857# gnd 3.43fF
C930 a_31172_n4289# gnd 2.27fF
C931 a_28681_n5229# gnd 3.16fF
C932 a_30124_n4285# gnd 2.80fF
C933 a_24450_n5190# gnd 3.43fF
C934 a_25846_n5749# gnd 3.27fF
C935 a_44032_n4308# gnd 2.33fF
C936 a_33281_n4316# gnd 2.33fF
C937 a_22573_n4851# gnd 3.43fF
C938 a_20207_n4293# gnd 2.27fF
C939 a_17716_n5233# gnd 3.16fF
C940 a_19159_n4289# gnd 2.80fF
C941 a_13485_n5194# gnd 3.43fF
C942 a_14881_n5753# gnd 3.27fF
C943 a_22573_n4310# gnd 2.33fF
C944 a_11608_n4855# gnd 3.43fF
C945 a_9499_n4287# gnd 2.27fF
C946 a_7008_n5227# gnd 3.16fF
C947 a_8451_n4283# gnd 2.80fF
C948 a_2777_n5188# gnd 3.43fF
C949 a_4173_n5747# gnd 3.27fF
C950 a_11608_n4314# gnd 2.33fF
C951 a_900_n4849# gnd 3.43fF
C952 a_900_n4308# gnd 2.33fF
C953 a_85016_n4472# gnd 3.17fF
C954 a_74308_n4466# gnd 3.17fF
C955 a_63343_n4470# gnd 3.17fF
C956 a_52635_n4464# gnd 3.17fF
C957 a_41884_n4472# gnd 3.17fF
C958 a_31176_n4466# gnd 3.17fF
C959 a_83968_n4468# gnd 3.33fF
C960 a_85012_n3616# gnd 2.28fF
C961 a_77242_n4424# gnd 3.33fF
C962 a_78290_n3749# gnd 4.37fF
C963 a_20211_n4470# gnd 3.17fF
C964 a_9503_n4464# gnd 3.17fF
C965 a_76413_n4061# gnd 3.17fF
C966 a_77242_n3745# gnd 2.80fF
C967 a_73260_n4462# gnd 3.33fF
C968 a_74304_n3610# gnd 2.28fF
C969 a_66534_n4418# gnd 3.33fF
C970 a_67582_n3743# gnd 4.37fF
C971 a_76413_n3666# gnd 2.27fF
C972 a_65705_n4055# gnd 3.17fF
C973 a_66534_n3739# gnd 2.80fF
C974 a_62295_n4466# gnd 3.33fF
C975 a_63339_n3614# gnd 2.28fF
C976 a_55569_n4422# gnd 3.33fF
C977 a_56617_n3747# gnd 4.37fF
C978 a_65705_n3660# gnd 2.27fF
C979 a_54740_n4059# gnd 3.17fF
C980 a_55569_n3743# gnd 2.80fF
C981 a_51587_n4460# gnd 3.33fF
C982 a_52631_n3608# gnd 2.28fF
C983 a_44861_n4416# gnd 3.33fF
C984 a_45909_n3741# gnd 4.37fF
C985 a_54740_n3664# gnd 2.27fF
C986 a_44032_n4053# gnd 3.17fF
C987 a_44861_n3737# gnd 2.80fF
C988 a_40836_n4468# gnd 3.33fF
C989 a_41880_n3616# gnd 2.28fF
C990 a_34110_n4424# gnd 3.33fF
C991 a_35158_n3749# gnd 4.37fF
C992 a_44032_n3658# gnd 2.27fF
C993 a_33281_n4061# gnd 3.17fF
C994 a_34110_n3745# gnd 2.80fF
C995 a_30128_n4462# gnd 3.33fF
C996 a_31172_n3610# gnd 2.28fF
C997 a_23402_n4418# gnd 3.33fF
C998 a_24450_n3743# gnd 4.37fF
C999 a_76413_n3410# gnd 17.59fF
C1000 a_65705_n3404# gnd 17.59fF
C1001 a_33281_n3666# gnd 2.27fF
C1002 a_22573_n4055# gnd 3.17fF
C1003 a_23402_n3739# gnd 2.80fF
C1004 a_19163_n4466# gnd 3.33fF
C1005 a_20207_n3614# gnd 2.28fF
C1006 a_12437_n4422# gnd 3.33fF
C1007 a_13485_n3747# gnd 4.37fF
C1008 a_22573_n3660# gnd 2.27fF
C1009 a_11608_n4059# gnd 3.17fF
C1010 a_12437_n3743# gnd 2.80fF
C1011 a_8455_n4460# gnd 3.33fF
C1012 a_9499_n3608# gnd 2.28fF
C1013 a_1729_n4416# gnd 3.33fF
C1014 a_2777_n3741# gnd 4.37fF
C1015 a_54740_n3408# gnd 17.59fF
C1016 a_44032_n3402# gnd 17.59fF
C1017 a_11608_n3664# gnd 2.27fF
C1018 a_900_n4053# gnd 3.17fF
C1019 a_1729_n3737# gnd 2.80fF
C1020 a_900_n3658# gnd 2.27fF
C1021 a_33281_n3410# gnd 17.59fF
C1022 a_22573_n3404# gnd 17.59fF
C1023 a_11608_n3408# gnd 17.59fF
C1024 a_900_n3402# gnd 17.59fF
C1025 a_70453_n5915# gnd 10.85fF
C1026 a_75301_n1457# gnd 11.63fF
C1027 a_64664_n1444# gnd 12.71fF
C1028 a_48780_n5913# gnd 10.85fF
C1029 a_53727_n1632# gnd 12.30fF
C1030 a_53628_n1455# gnd 11.63fF
C1031 a_27321_n5915# gnd 10.85fF
C1032 a_32169_n1457# gnd 11.63fF
C1033 a_21631_n1621# gnd 27.41fF
C1034 a_21532_n1444# gnd 12.71fF
C1035 a_5648_n5913# gnd 10.85fF
C1036 a_10595_n1632# gnd 12.21fF
C1037 a_10496_n1455# gnd 11.63fF
C1038 a_43231_n1412# gnd 23.98fF
C1039 a_3053_n1225# gnd 44.03fF
C1040 vout gnd 4.53fF
C1041 d9 gnd 4.15fF
C1042 a_64849_973# gnd 12.30fF
C1043 a_54311_986# gnd 12.71fF
C1044 a_43150_941# gnd 27.41fF
C1045 a_3058_n1106# gnd 46.08fF
C1046 d8 gnd 53.48fF
C1047 a_21717_973# gnd 12.30fF
C1048 a_21816_973# gnd 23.94fF
C1049 d7 gnd 104.11fF
C1050 a_11179_986# gnd 12.71fF
C1051 d6 gnd 240.69fF
C1052 a_84751_3266# gnd 2.27fF
C1053 a_83703_3270# gnd 2.80fF
C1054 a_76154_3146# gnd 17.59fF
C1055 a_74043_3272# gnd 2.27fF
C1056 a_72995_3276# gnd 2.80fF
C1057 a_76152_3245# gnd 2.28fF
C1058 a_65446_3152# gnd 17.59fF
C1059 a_63078_3268# gnd 2.27fF
C1060 a_62030_3272# gnd 2.80fF
C1061 a_65444_3251# gnd 2.28fF
C1062 a_54481_3148# gnd 17.59fF
C1063 a_52370_3274# gnd 2.27fF
C1064 a_51322_3278# gnd 2.80fF
C1065 a_54479_3247# gnd 2.28fF
C1066 a_43773_3154# gnd 17.59fF
C1067 a_41619_3266# gnd 2.27fF
C1068 a_40571_3270# gnd 2.80fF
C1069 a_33022_3146# gnd 17.59fF
C1070 a_30911_3272# gnd 2.27fF
C1071 a_29863_3276# gnd 2.80fF
C1072 a_43771_3253# gnd 2.28fF
C1073 a_33020_3245# gnd 2.28fF
C1074 a_22314_3152# gnd 17.59fF
C1075 a_19946_3268# gnd 2.27fF
C1076 a_18898_3272# gnd 2.80fF
C1077 a_22312_3251# gnd 2.28fF
C1078 a_11349_3148# gnd 17.59fF
C1079 a_9238_3274# gnd 2.27fF
C1080 a_8190_3278# gnd 2.80fF
C1081 a_11347_3247# gnd 2.28fF
C1082 a_641_3154# gnd 17.59fF
C1083 a_639_3253# gnd 2.28fF
C1084 a_84755_3089# gnd 3.17fF
C1085 a_74047_3095# gnd 3.17fF
C1086 a_63082_3091# gnd 3.17fF
C1087 a_52374_3097# gnd 3.17fF
C1088 a_41623_3089# gnd 3.17fF
C1089 a_30915_3095# gnd 3.17fF
C1090 a_83707_3093# gnd 3.33fF
C1091 a_84751_3945# gnd 2.33fF
C1092 a_82256_3950# gnd 4.37fF
C1093 a_76981_3137# gnd 3.33fF
C1094 a_19950_3091# gnd 3.17fF
C1095 a_9242_3097# gnd 3.17fF
C1096 a_76152_3500# gnd 3.17fF
C1097 a_76981_3816# gnd 2.80fF
C1098 a_72999_3099# gnd 3.33fF
C1099 a_74043_3951# gnd 2.33fF
C1100 a_71548_3956# gnd 4.37fF
C1101 a_66273_3143# gnd 3.33fF
C1102 a_76152_3895# gnd 2.27fF
C1103 a_65444_3506# gnd 3.17fF
C1104 a_66273_3822# gnd 2.80fF
C1105 a_62034_3095# gnd 3.33fF
C1106 a_63078_3947# gnd 2.33fF
C1107 a_60583_3952# gnd 4.37fF
C1108 a_55308_3139# gnd 3.33fF
C1109 a_65444_3901# gnd 2.27fF
C1110 a_54479_3502# gnd 3.17fF
C1111 a_55308_3818# gnd 2.80fF
C1112 a_51326_3101# gnd 3.33fF
C1113 a_52370_3953# gnd 2.33fF
C1114 a_49875_3958# gnd 4.37fF
C1115 a_44600_3145# gnd 3.33fF
C1116 a_54479_3897# gnd 2.27fF
C1117 a_43771_3508# gnd 3.17fF
C1118 a_44600_3824# gnd 2.80fF
C1119 a_40575_3093# gnd 3.33fF
C1120 a_41619_3945# gnd 2.33fF
C1121 a_39124_3950# gnd 4.37fF
C1122 a_33849_3137# gnd 3.33fF
C1123 a_43771_3903# gnd 2.27fF
C1124 a_33020_3500# gnd 3.17fF
C1125 a_33849_3816# gnd 2.80fF
C1126 a_29867_3099# gnd 3.33fF
C1127 a_30911_3951# gnd 2.33fF
C1128 a_28416_3956# gnd 4.37fF
C1129 a_23141_3143# gnd 3.33fF
C1130 a_33020_3895# gnd 2.27fF
C1131 a_22312_3506# gnd 3.17fF
C1132 a_23141_3822# gnd 2.80fF
C1133 a_18902_3095# gnd 3.33fF
C1134 a_19946_3947# gnd 2.33fF
C1135 a_17451_3952# gnd 4.37fF
C1136 a_12176_3139# gnd 3.33fF
C1137 a_22312_3901# gnd 2.27fF
C1138 a_11347_3502# gnd 3.17fF
C1139 a_12176_3818# gnd 2.80fF
C1140 a_8194_3101# gnd 3.33fF
C1141 a_9238_3953# gnd 2.33fF
C1142 a_6743_3958# gnd 4.37fF
C1143 a_1468_3145# gnd 3.33fF
C1144 a_11347_3897# gnd 2.27fF
C1145 a_639_3508# gnd 3.17fF
C1146 a_1468_3824# gnd 2.80fF
C1147 a_639_3903# gnd 2.27fF
C1148 a_84755_3768# gnd 3.43fF
C1149 a_74047_3774# gnd 3.43fF
C1150 a_63082_3770# gnd 3.43fF
C1151 a_52374_3776# gnd 3.43fF
C1152 a_41623_3768# gnd 3.43fF
C1153 a_30915_3774# gnd 3.43fF
C1154 a_84751_4713# gnd 2.27fF
C1155 a_82260_3773# gnd 3.43fF
C1156 a_83703_4717# gnd 2.80fF
C1157 a_78029_3812# gnd 3.16fF
C1158 a_76152_4151# gnd 3.43fF
C1159 a_74043_4719# gnd 2.27fF
C1160 a_71552_3779# gnd 3.43fF
C1161 a_72995_4723# gnd 2.80fF
C1162 a_67321_3818# gnd 3.16fF
C1163 a_19950_3770# gnd 3.43fF
C1164 a_9242_3776# gnd 3.43fF
C1165 a_76152_4692# gnd 2.33fF
C1166 a_65444_4157# gnd 3.43fF
C1167 a_63078_4715# gnd 2.27fF
C1168 a_60587_3775# gnd 3.43fF
C1169 a_62030_4719# gnd 2.80fF
C1170 a_56356_3814# gnd 3.16fF
C1171 a_65444_4698# gnd 2.33fF
C1172 a_54479_4153# gnd 3.43fF
C1173 a_52370_4721# gnd 2.27fF
C1174 a_49879_3781# gnd 3.43fF
C1175 a_51322_4725# gnd 2.80fF
C1176 a_45648_3820# gnd 3.16fF
C1177 a_54479_4694# gnd 2.33fF
C1178 a_43771_4159# gnd 3.43fF
C1179 a_41619_4713# gnd 2.27fF
C1180 a_39128_3773# gnd 3.43fF
C1181 a_40571_4717# gnd 2.80fF
C1182 a_34897_3812# gnd 3.16fF
C1183 a_33020_4151# gnd 3.43fF
C1184 a_30911_4719# gnd 2.27fF
C1185 a_28420_3779# gnd 3.43fF
C1186 a_29863_4723# gnd 2.80fF
C1187 a_24189_3818# gnd 3.16fF
C1188 a_43771_4700# gnd 2.33fF
C1189 a_33020_4692# gnd 2.33fF
C1190 a_22312_4157# gnd 3.43fF
C1191 a_19946_4715# gnd 2.27fF
C1192 a_17455_3775# gnd 3.43fF
C1193 a_18898_4719# gnd 2.80fF
C1194 a_13224_3814# gnd 3.16fF
C1195 a_22312_4698# gnd 2.33fF
C1196 a_11347_4153# gnd 3.43fF
C1197 a_9238_4721# gnd 2.27fF
C1198 a_6747_3781# gnd 3.43fF
C1199 a_8190_4725# gnd 2.80fF
C1200 a_2516_3820# gnd 3.16fF
C1201 a_11347_4694# gnd 2.33fF
C1202 a_639_4159# gnd 3.43fF
C1203 a_639_4700# gnd 2.33fF
C1204 a_84755_4536# gnd 3.17fF
C1205 a_74047_4542# gnd 3.17fF
C1206 a_63082_4538# gnd 3.17fF
C1207 a_52374_4544# gnd 3.17fF
C1208 a_41623_4536# gnd 3.17fF
C1209 a_30915_4542# gnd 3.17fF
C1210 a_83707_4540# gnd 3.33fF
C1211 a_84751_5392# gnd 2.33fF
C1212 a_82213_5395# gnd 3.27fF
C1213 a_75885_984# gnd 10.85fF
C1214 a_76981_4584# gnd 3.33fF
C1215 a_78029_5259# gnd 3.64fF
C1216 a_76152_4947# gnd 3.17fF
C1217 a_76981_5263# gnd 2.80fF
C1218 a_19950_4538# gnd 3.17fF
C1219 a_9242_4544# gnd 3.17fF
C1220 a_72999_4546# gnd 3.33fF
C1221 a_74043_5398# gnd 2.33fF
C1222 a_71505_5401# gnd 3.27fF
C1223 a_76152_5342# gnd 2.27fF
C1224 a_70223_5271# gnd 11.63fF
C1225 a_66273_4590# gnd 3.33fF
C1226 a_67321_5265# gnd 3.64fF
C1227 a_65444_4953# gnd 3.17fF
C1228 a_66273_5269# gnd 2.80fF
C1229 a_62034_4542# gnd 3.33fF
C1230 a_63078_5394# gnd 2.33fF
C1231 a_60540_5397# gnd 3.27fF
C1232 a_65444_5348# gnd 2.27fF
C1233 a_54212_986# gnd 10.85fF
C1234 a_55308_4586# gnd 3.33fF
C1235 a_56356_5261# gnd 3.64fF
C1236 a_54479_4949# gnd 3.17fF
C1237 a_55308_5265# gnd 2.80fF
C1238 a_51326_4548# gnd 3.33fF
C1239 a_52370_5400# gnd 2.33fF
C1240 a_49832_5403# gnd 3.27fF
C1241 a_54479_5344# gnd 2.27fF
C1242 a_48550_5273# gnd 11.63fF
C1243 a_44600_4592# gnd 3.33fF
C1244 a_45648_5267# gnd 3.64fF
C1245 a_43771_4955# gnd 3.17fF
C1246 a_44600_5271# gnd 2.80fF
C1247 a_40575_4540# gnd 3.33fF
C1248 a_41619_5392# gnd 2.33fF
C1249 a_39081_5395# gnd 3.27fF
C1250 a_43771_5350# gnd 2.27fF
C1251 a_32753_984# gnd 10.85fF
C1252 a_33849_4584# gnd 3.33fF
C1253 a_34897_5259# gnd 3.64fF
C1254 a_33020_4947# gnd 3.17fF
C1255 a_33849_5263# gnd 2.80fF
C1256 a_29867_4546# gnd 3.33fF
C1257 a_30911_5398# gnd 2.33fF
C1258 a_28373_5401# gnd 3.27fF
C1259 a_33020_5342# gnd 2.27fF
C1260 a_27091_5271# gnd 11.63fF
C1261 a_23141_4590# gnd 3.33fF
C1262 a_24189_5265# gnd 3.64fF
C1263 a_22312_4953# gnd 3.17fF
C1264 a_23141_5269# gnd 2.80fF
C1265 a_18902_4542# gnd 3.33fF
C1266 a_19946_5394# gnd 2.33fF
C1267 a_17408_5397# gnd 3.27fF
C1268 a_22312_5348# gnd 2.27fF
C1269 a_11080_986# gnd 10.85fF
C1270 a_12176_4586# gnd 3.33fF
C1271 a_13224_5261# gnd 3.64fF
C1272 a_11347_4949# gnd 3.17fF
C1273 a_12176_5265# gnd 2.80fF
C1274 a_8194_4548# gnd 3.33fF
C1275 a_9238_5400# gnd 2.33fF
C1276 a_6700_5403# gnd 3.27fF
C1277 a_11347_5344# gnd 2.27fF
C1278 a_5418_5273# gnd 11.63fF
C1279 a_1468_4592# gnd 3.33fF
C1280 a_2516_5267# gnd 3.64fF
C1281 d5 gnd 403.42fF
C1282 a_639_4955# gnd 3.17fF
C1283 a_1468_5271# gnd 2.80fF
C1284 a_639_5350# gnd 2.27fF
C1285 a_84755_5215# gnd 3.52fF
C1286 a_74047_5221# gnd 3.52fF
C1287 a_63082_5217# gnd 3.52fF
C1288 a_52374_5223# gnd 3.52fF
C1289 a_41623_5215# gnd 3.52fF
C1290 a_30915_5221# gnd 3.52fF
C1291 a_84750_6233# gnd 2.27fF
C1292 a_83702_6237# gnd 2.80fF
C1293 a_79419_6101# gnd 3.19fF
C1294 a_76152_5598# gnd 3.52fF
C1295 a_74042_6239# gnd 2.27fF
C1296 a_72994_6243# gnd 2.80fF
C1297 a_68711_6107# gnd 3.19fF
C1298 a_19950_5217# gnd 3.52fF
C1299 a_9242_5223# gnd 3.52fF
C1300 a_76151_6212# gnd 2.33fF
C1301 a_65444_5604# gnd 3.52fF
C1302 a_63077_6235# gnd 2.27fF
C1303 a_62029_6239# gnd 2.80fF
C1304 a_57746_6103# gnd 3.19fF
C1305 a_65443_6218# gnd 2.33fF
C1306 a_54479_5600# gnd 3.52fF
C1307 a_52369_6241# gnd 2.27fF
C1308 a_51321_6245# gnd 2.80fF
C1309 a_47038_6109# gnd 3.19fF
C1310 a_54478_6214# gnd 2.33fF
C1311 a_43771_5606# gnd 3.52fF
C1312 a_41618_6233# gnd 2.27fF
C1313 a_40570_6237# gnd 2.80fF
C1314 a_36287_6101# gnd 3.19fF
C1315 a_33020_5598# gnd 3.52fF
C1316 a_30910_6239# gnd 2.27fF
C1317 a_29862_6243# gnd 2.80fF
C1318 a_25579_6107# gnd 3.19fF
C1319 a_43770_6220# gnd 2.33fF
C1320 a_33019_6212# gnd 2.33fF
C1321 a_22312_5604# gnd 3.52fF
C1322 a_19945_6235# gnd 2.27fF
C1323 a_18897_6239# gnd 2.80fF
C1324 a_14614_6103# gnd 3.19fF
C1325 a_22311_6218# gnd 2.33fF
C1326 a_11347_5600# gnd 3.52fF
C1327 a_9237_6241# gnd 2.27fF
C1328 a_8189_6245# gnd 2.80fF
C1329 a_3906_6109# gnd 3.19fF
C1330 a_11346_6214# gnd 2.33fF
C1331 a_639_5606# gnd 3.52fF
C1332 a_638_6220# gnd 2.33fF
C1333 a_84754_6056# gnd 3.17fF
C1334 a_74046_6062# gnd 3.17fF
C1335 a_63081_6058# gnd 3.17fF
C1336 a_52373_6064# gnd 3.17fF
C1337 a_41622_6056# gnd 3.17fF
C1338 a_30914_6062# gnd 3.17fF
C1339 a_83706_6060# gnd 3.33fF
C1340 a_84750_6912# gnd 2.33fF
C1341 a_82217_5218# gnd 3.19fF
C1342 a_82255_6917# gnd 3.65fF
C1343 a_76980_6104# gnd 3.33fF
C1344 a_19949_6058# gnd 3.17fF
C1345 a_9241_6064# gnd 3.17fF
C1346 a_76151_6467# gnd 3.17fF
C1347 a_76980_6783# gnd 2.80fF
C1348 a_72998_6066# gnd 3.33fF
C1349 a_74042_6918# gnd 2.33fF
C1350 a_71509_5224# gnd 3.19fF
C1351 a_71547_6923# gnd 3.65fF
C1352 a_66272_6110# gnd 3.33fF
C1353 a_76151_6862# gnd 2.27fF
C1354 a_65443_6473# gnd 3.17fF
C1355 a_66272_6789# gnd 2.80fF
C1356 a_62033_6062# gnd 3.33fF
C1357 a_63077_6914# gnd 2.33fF
C1358 a_60544_5220# gnd 3.19fF
C1359 a_60582_6919# gnd 3.65fF
C1360 a_55307_6106# gnd 3.33fF
C1361 a_65443_6868# gnd 2.27fF
C1362 a_54478_6469# gnd 3.17fF
C1363 a_55307_6785# gnd 2.80fF
C1364 a_51325_6068# gnd 3.33fF
C1365 a_52369_6920# gnd 2.33fF
C1366 a_49836_5226# gnd 3.19fF
C1367 a_49874_6925# gnd 3.65fF
C1368 a_44599_6112# gnd 3.33fF
C1369 a_54478_6864# gnd 2.27fF
C1370 a_43770_6475# gnd 3.17fF
C1371 a_44599_6791# gnd 2.80fF
C1372 a_40574_6060# gnd 3.33fF
C1373 a_41618_6912# gnd 2.33fF
C1374 a_39085_5218# gnd 3.19fF
C1375 a_39123_6917# gnd 3.65fF
C1376 a_33848_6104# gnd 3.33fF
C1377 a_43770_6870# gnd 2.27fF
C1378 a_33019_6467# gnd 3.17fF
C1379 a_33848_6783# gnd 2.80fF
C1380 a_29866_6066# gnd 3.33fF
C1381 a_30910_6918# gnd 2.33fF
C1382 a_28377_5224# gnd 3.19fF
C1383 a_28415_6923# gnd 3.65fF
C1384 a_23140_6110# gnd 3.33fF
C1385 a_33019_6862# gnd 2.27fF
C1386 a_22311_6473# gnd 3.17fF
C1387 a_23140_6789# gnd 2.80fF
C1388 a_18901_6062# gnd 3.33fF
C1389 a_19945_6914# gnd 2.33fF
C1390 a_17412_5220# gnd 3.19fF
C1391 a_17450_6919# gnd 3.65fF
C1392 a_12175_6106# gnd 3.33fF
C1393 a_22311_6868# gnd 2.27fF
C1394 a_11346_6469# gnd 3.17fF
C1395 a_12175_6785# gnd 2.80fF
C1396 a_8193_6068# gnd 3.33fF
C1397 a_9237_6920# gnd 2.33fF
C1398 a_6704_5226# gnd 3.19fF
C1399 a_6742_6925# gnd 3.65fF
C1400 a_1467_6112# gnd 3.33fF
C1401 a_11346_6864# gnd 2.27fF
C1402 a_638_6475# gnd 3.17fF
C1403 a_1467_6791# gnd 2.80fF
C1404 a_638_6870# gnd 2.27fF
C1405 a_84754_6735# gnd 3.43fF
C1406 a_74046_6741# gnd 3.43fF
C1407 a_63081_6737# gnd 3.43fF
C1408 a_52373_6743# gnd 3.43fF
C1409 a_41622_6735# gnd 3.43fF
C1410 a_30914_6741# gnd 3.43fF
C1411 a_84750_7680# gnd 2.27fF
C1412 a_82259_6740# gnd 3.20fF
C1413 a_83702_7684# gnd 2.80fF
C1414 a_78028_6779# gnd 3.43fF
C1415 a_79424_6220# gnd 3.27fF
C1416 a_76151_7118# gnd 3.43fF
C1417 a_74042_7686# gnd 2.27fF
C1418 a_71551_6746# gnd 3.20fF
C1419 a_72994_7690# gnd 2.80fF
C1420 a_67320_6785# gnd 3.43fF
C1421 a_68716_6226# gnd 3.27fF
C1422 a_19949_6737# gnd 3.43fF
C1423 a_9241_6743# gnd 3.43fF
C1424 a_76151_7659# gnd 2.33fF
C1425 a_65443_7124# gnd 3.43fF
C1426 a_63077_7682# gnd 2.27fF
C1427 a_60586_6742# gnd 3.20fF
C1428 a_62029_7686# gnd 2.80fF
C1429 a_56355_6781# gnd 3.43fF
C1430 a_57751_6222# gnd 3.27fF
C1431 a_65443_7665# gnd 2.33fF
C1432 a_54478_7120# gnd 3.43fF
C1433 a_52369_7688# gnd 2.27fF
C1434 a_49878_6748# gnd 3.20fF
C1435 a_51321_7692# gnd 2.80fF
C1436 a_45647_6787# gnd 3.43fF
C1437 a_47043_6228# gnd 3.27fF
C1438 a_54478_7661# gnd 2.33fF
C1439 a_43770_7126# gnd 3.43fF
C1440 a_41618_7680# gnd 2.27fF
C1441 a_39127_6740# gnd 3.20fF
C1442 a_40570_7684# gnd 2.80fF
C1443 a_34896_6779# gnd 3.43fF
C1444 a_36292_6220# gnd 3.27fF
C1445 a_33019_7118# gnd 3.43fF
C1446 a_30910_7686# gnd 2.27fF
C1447 a_28419_6746# gnd 3.20fF
C1448 a_29862_7690# gnd 2.80fF
C1449 a_24188_6785# gnd 3.43fF
C1450 a_25584_6226# gnd 3.27fF
C1451 a_43770_7667# gnd 2.33fF
C1452 a_33019_7659# gnd 2.33fF
C1453 a_22311_7124# gnd 3.43fF
C1454 a_19945_7682# gnd 2.27fF
C1455 a_17454_6742# gnd 3.20fF
C1456 a_18897_7686# gnd 2.80fF
C1457 a_13223_6781# gnd 3.43fF
C1458 a_14619_6222# gnd 3.27fF
C1459 a_22311_7665# gnd 2.33fF
C1460 a_11346_7120# gnd 3.43fF
C1461 a_9237_7688# gnd 2.27fF
C1462 a_6746_6748# gnd 3.20fF
C1463 a_8189_7692# gnd 2.80fF
C1464 a_2515_6787# gnd 3.43fF
C1465 a_3911_6228# gnd 3.27fF
C1466 a_11346_7661# gnd 2.33fF
C1467 a_638_7126# gnd 3.43fF
C1468 a_638_7667# gnd 2.33fF
C1469 a_84754_7503# gnd 3.17fF
C1470 a_74046_7509# gnd 3.17fF
C1471 a_63081_7505# gnd 3.17fF
C1472 a_52373_7511# gnd 3.17fF
C1473 a_41622_7503# gnd 3.17fF
C1474 a_30914_7509# gnd 3.17fF
C1475 a_83706_7507# gnd 3.33fF
C1476 a_84750_8359# gnd 2.33fF
C1477 a_80832_5265# gnd 4.30fF
C1478 a_81147_8368# gnd 7.03fF
C1479 a_76980_7551# gnd 3.33fF
C1480 a_78028_8226# gnd 4.35fF
C1481 a_19949_7505# gnd 3.17fF
C1482 a_9241_7511# gnd 3.17fF
C1483 a_76151_7914# gnd 3.17fF
C1484 a_76980_8230# gnd 2.80fF
C1485 a_72998_7513# gnd 3.33fF
C1486 a_74042_8365# gnd 2.33fF
C1487 a_70124_5271# gnd 4.30fF
C1488 a_70439_8374# gnd 7.03fF
C1489 a_66272_7557# gnd 3.33fF
C1490 a_67320_8232# gnd 4.35fF
C1491 a_76151_8309# gnd 2.27fF
C1492 a_65443_7920# gnd 3.17fF
C1493 a_66272_8236# gnd 2.80fF
C1494 a_62033_7509# gnd 3.33fF
C1495 a_63077_8361# gnd 2.33fF
C1496 a_59159_5267# gnd 4.30fF
C1497 a_59474_8370# gnd 7.03fF
C1498 a_55307_7553# gnd 3.33fF
C1499 a_56355_8228# gnd 4.35fF
C1500 a_65443_8315# gnd 2.27fF
C1501 a_54478_7916# gnd 3.17fF
C1502 a_55307_8232# gnd 2.80fF
C1503 a_51325_7515# gnd 3.33fF
C1504 a_52369_8367# gnd 2.33fF
C1505 a_48451_5273# gnd 4.30fF
C1506 a_48766_8376# gnd 7.03fF
C1507 a_44599_7559# gnd 3.33fF
C1508 a_45647_8234# gnd 4.35fF
C1509 a_54478_8311# gnd 2.27fF
C1510 a_43770_7922# gnd 3.17fF
C1511 a_44599_8238# gnd 2.80fF
C1512 a_40574_7507# gnd 3.33fF
C1513 a_41618_8359# gnd 2.33fF
C1514 a_37700_5265# gnd 4.30fF
C1515 a_38015_8368# gnd 7.03fF
C1516 a_33848_7551# gnd 3.33fF
C1517 a_34896_8226# gnd 4.35fF
C1518 a_43770_8317# gnd 2.27fF
C1519 a_33019_7914# gnd 3.17fF
C1520 a_33848_8230# gnd 2.80fF
C1521 a_29866_7513# gnd 3.33fF
C1522 a_30910_8365# gnd 2.33fF
C1523 a_26992_5271# gnd 4.30fF
C1524 a_27307_8374# gnd 7.03fF
C1525 a_23140_7557# gnd 3.33fF
C1526 a_24188_8232# gnd 4.35fF
C1527 a_33019_8309# gnd 2.27fF
C1528 a_22311_7920# gnd 3.17fF
C1529 a_23140_8236# gnd 2.80fF
C1530 a_18901_7509# gnd 3.33fF
C1531 a_19945_8361# gnd 2.33fF
C1532 a_16027_5267# gnd 4.30fF
C1533 a_16342_8370# gnd 7.03fF
C1534 a_12175_7553# gnd 3.33fF
C1535 a_13223_8228# gnd 4.35fF
C1536 a_22311_8315# gnd 2.27fF
C1537 a_11346_7916# gnd 3.17fF
C1538 a_12175_8232# gnd 2.80fF
C1539 a_8193_7515# gnd 3.33fF
C1540 a_9237_8367# gnd 2.33fF
C1541 a_5319_5273# gnd 4.30fF
C1542 a_5634_8376# gnd 7.03fF
C1543 a_1467_7559# gnd 3.33fF
C1544 a_2515_8234# gnd 4.35fF
C1545 a_11346_8311# gnd 2.27fF
C1546 a_638_7922# gnd 3.17fF
C1547 a_1467_8238# gnd 2.80fF
C1548 a_638_8317# gnd 2.27fF
C1549 a_84754_8182# gnd 3.62fF
C1550 a_74046_8188# gnd 3.62fF
C1551 a_63081_8184# gnd 3.62fF
C1552 a_52373_8190# gnd 3.62fF
C1553 a_41622_8182# gnd 3.62fF
C1554 a_30914_8188# gnd 3.62fF
C1555 a_84753_9274# gnd 2.27fF
C1556 a_83705_9278# gnd 2.80fF
C1557 a_79518_6101# gnd 4.97fF
C1558 a_80586_9136# gnd 4.72fF
C1559 a_76151_8565# gnd 3.62fF
C1560 a_74045_9280# gnd 2.27fF
C1561 a_72997_9284# gnd 2.80fF
C1562 a_68810_6107# gnd 4.97fF
C1563 a_69878_9142# gnd 4.72fF
C1564 a_19949_8184# gnd 3.62fF
C1565 a_9241_8190# gnd 3.62fF
C1566 a_76154_9253# gnd 2.33fF
C1567 a_65443_8571# gnd 3.62fF
C1568 a_63080_9276# gnd 2.27fF
C1569 a_62032_9280# gnd 2.80fF
C1570 a_57845_6103# gnd 4.97fF
C1571 a_58913_9138# gnd 4.72fF
C1572 a_65446_9259# gnd 2.33fF
C1573 a_54478_8567# gnd 3.62fF
C1574 a_52372_9282# gnd 2.27fF
C1575 a_51324_9286# gnd 2.80fF
C1576 a_47137_6109# gnd 4.97fF
C1577 a_48205_9144# gnd 4.72fF
C1578 a_54481_9255# gnd 2.33fF
C1579 a_43770_8573# gnd 3.62fF
C1580 a_41621_9274# gnd 2.27fF
C1581 a_40573_9278# gnd 2.80fF
C1582 a_36386_6101# gnd 4.97fF
C1583 a_37454_9136# gnd 4.72fF
C1584 a_33019_8565# gnd 3.62fF
C1585 a_30913_9280# gnd 2.27fF
C1586 a_29865_9284# gnd 2.80fF
C1587 a_25678_6107# gnd 4.97fF
C1588 a_26746_9142# gnd 4.72fF
C1589 a_43773_9261# gnd 2.33fF
C1590 a_33022_9253# gnd 2.33fF
C1591 a_22311_8571# gnd 3.62fF
C1592 a_19948_9276# gnd 2.27fF
C1593 a_18900_9280# gnd 2.80fF
C1594 a_14713_6103# gnd 4.97fF
C1595 a_15781_9138# gnd 4.72fF
C1596 a_22314_9259# gnd 2.33fF
C1597 a_11346_8567# gnd 3.62fF
C1598 a_9240_9282# gnd 2.27fF
C1599 a_8192_9286# gnd 2.80fF
C1600 a_4005_6109# gnd 4.97fF
C1601 a_5073_9144# gnd 4.72fF
C1602 a_11349_9255# gnd 2.33fF
C1603 d4 gnd 489.14fF
C1604 a_638_8573# gnd 3.62fF
C1605 a_641_9261# gnd 2.33fF
C1606 a_84757_9097# gnd 3.17fF
C1607 a_74049_9103# gnd 3.17fF
C1608 a_63084_9099# gnd 3.17fF
C1609 a_52376_9105# gnd 3.17fF
C1610 a_41625_9097# gnd 3.17fF
C1611 a_30917_9103# gnd 3.17fF
C1612 a_83709_9101# gnd 3.33fF
C1613 a_84753_9953# gnd 2.33fF
C1614 a_82258_9958# gnd 4.35fF
C1615 a_76983_9145# gnd 3.33fF
C1616 a_19952_9099# gnd 3.17fF
C1617 a_9244_9105# gnd 3.17fF
C1618 a_76154_9508# gnd 3.17fF
C1619 a_76983_9824# gnd 2.80fF
C1620 a_73001_9107# gnd 3.33fF
C1621 a_74045_9959# gnd 2.33fF
C1622 a_71550_9964# gnd 4.35fF
C1623 a_66275_9151# gnd 3.33fF
C1624 a_76154_9903# gnd 2.27fF
C1625 a_65446_9514# gnd 3.17fF
C1626 a_66275_9830# gnd 2.80fF
C1627 a_62036_9103# gnd 3.33fF
C1628 a_63080_9955# gnd 2.33fF
C1629 a_60585_9960# gnd 4.35fF
C1630 a_55310_9147# gnd 3.33fF
C1631 a_65446_9909# gnd 2.27fF
C1632 a_54481_9510# gnd 3.17fF
C1633 a_55310_9826# gnd 2.80fF
C1634 a_51328_9109# gnd 3.33fF
C1635 a_52372_9961# gnd 2.33fF
C1636 a_49877_9966# gnd 4.35fF
C1637 a_44602_9153# gnd 3.33fF
C1638 a_54481_9905# gnd 2.27fF
C1639 a_43773_9516# gnd 3.17fF
C1640 a_44602_9832# gnd 2.80fF
C1641 a_40577_9101# gnd 3.33fF
C1642 a_41621_9953# gnd 2.33fF
C1643 a_39126_9958# gnd 4.35fF
C1644 a_33851_9145# gnd 3.33fF
C1645 a_43773_9911# gnd 2.27fF
C1646 a_33022_9508# gnd 3.17fF
C1647 a_33851_9824# gnd 2.80fF
C1648 a_29869_9107# gnd 3.33fF
C1649 a_30913_9959# gnd 2.33fF
C1650 a_28418_9964# gnd 4.35fF
C1651 a_23143_9151# gnd 3.33fF
C1652 a_33022_9903# gnd 2.27fF
C1653 a_22314_9514# gnd 3.17fF
C1654 a_23143_9830# gnd 2.80fF
C1655 a_18904_9103# gnd 3.33fF
C1656 a_19948_9955# gnd 2.33fF
C1657 a_17453_9960# gnd 4.35fF
C1658 a_12178_9147# gnd 3.33fF
C1659 a_22314_9909# gnd 2.27fF
C1660 a_11349_9510# gnd 3.17fF
C1661 a_12178_9826# gnd 2.80fF
C1662 a_8196_9109# gnd 3.33fF
C1663 a_9240_9961# gnd 2.33fF
C1664 a_6745_9966# gnd 4.35fF
C1665 a_1470_9153# gnd 3.33fF
C1666 a_11349_9905# gnd 2.27fF
C1667 a_641_9516# gnd 3.17fF
C1668 a_1470_9832# gnd 2.80fF
C1669 a_641_9911# gnd 2.27fF
C1670 a_84757_9776# gnd 3.43fF
C1671 a_74049_9782# gnd 3.43fF
C1672 a_63084_9778# gnd 3.43fF
C1673 a_52376_9784# gnd 3.43fF
C1674 a_41625_9776# gnd 3.43fF
C1675 a_30917_9782# gnd 3.43fF
C1676 a_84753_10721# gnd 2.27fF
C1677 a_82262_9781# gnd 3.43fF
C1678 a_83705_10725# gnd 2.80fF
C1679 a_78031_9820# gnd 3.20fF
C1680 a_76154_10159# gnd 3.43fF
C1681 a_74045_10727# gnd 2.27fF
C1682 a_71554_9787# gnd 3.43fF
C1683 a_72997_10731# gnd 2.80fF
C1684 a_67323_9826# gnd 3.20fF
C1685 a_19952_9778# gnd 3.43fF
C1686 a_9244_9784# gnd 3.43fF
C1687 a_76154_10700# gnd 2.33fF
C1688 a_65446_10165# gnd 3.43fF
C1689 a_63080_10723# gnd 2.27fF
C1690 a_60589_9783# gnd 3.43fF
C1691 a_62032_10727# gnd 2.80fF
C1692 a_56358_9822# gnd 3.20fF
C1693 a_65446_10706# gnd 2.33fF
C1694 a_54481_10161# gnd 3.43fF
C1695 a_52372_10729# gnd 2.27fF
C1696 a_49881_9789# gnd 3.43fF
C1697 a_51324_10733# gnd 2.80fF
C1698 a_45650_9828# gnd 3.20fF
C1699 a_54481_10702# gnd 2.33fF
C1700 a_43773_10167# gnd 3.43fF
C1701 a_41621_10721# gnd 2.27fF
C1702 a_39130_9781# gnd 3.43fF
C1703 a_40573_10725# gnd 2.80fF
C1704 a_34899_9820# gnd 3.20fF
C1705 a_33022_10159# gnd 3.43fF
C1706 a_30913_10727# gnd 2.27fF
C1707 a_28422_9787# gnd 3.43fF
C1708 a_29865_10731# gnd 2.80fF
C1709 a_24191_9826# gnd 3.20fF
C1710 a_43773_10708# gnd 2.33fF
C1711 a_33022_10700# gnd 2.33fF
C1712 a_22314_10165# gnd 3.43fF
C1713 a_19948_10723# gnd 2.27fF
C1714 a_17457_9783# gnd 3.43fF
C1715 a_18900_10727# gnd 2.80fF
C1716 a_13226_9822# gnd 3.20fF
C1717 a_22314_10706# gnd 2.33fF
C1718 a_11349_10161# gnd 3.43fF
C1719 a_9240_10729# gnd 2.27fF
C1720 a_6749_9789# gnd 3.43fF
C1721 a_8192_10733# gnd 2.80fF
C1722 a_2518_9828# gnd 3.20fF
C1723 a_11349_10702# gnd 2.33fF
C1724 a_641_10167# gnd 3.43fF
C1725 a_641_10708# gnd 2.33fF
C1726 a_84757_10544# gnd 3.17fF
C1727 a_74049_10550# gnd 3.17fF
C1728 a_63084_10546# gnd 3.17fF
C1729 a_52376_10552# gnd 3.17fF
C1730 a_41625_10544# gnd 3.17fF
C1731 a_30917_10550# gnd 3.17fF
C1732 a_83709_10548# gnd 3.33fF
C1733 a_84753_11400# gnd 2.33fF
C1734 a_81151_8191# gnd 4.90fF
C1735 a_82215_11403# gnd 3.27fF
C1736 a_76983_10592# gnd 3.33fF
C1737 a_78031_11267# gnd 3.65fF
C1738 a_19952_10546# gnd 3.17fF
C1739 a_9244_10552# gnd 3.17fF
C1740 a_76154_10955# gnd 3.17fF
C1741 a_76983_11271# gnd 2.80fF
C1742 a_73001_10554# gnd 3.33fF
C1743 a_74045_11406# gnd 2.33fF
C1744 a_70443_8197# gnd 4.90fF
C1745 a_71507_11409# gnd 3.27fF
C1746 a_66275_10598# gnd 3.33fF
C1747 a_67323_11273# gnd 3.65fF
C1748 a_76154_11350# gnd 2.27fF
C1749 a_65446_10961# gnd 3.17fF
C1750 a_66275_11277# gnd 2.80fF
C1751 a_62036_10550# gnd 3.33fF
C1752 a_63080_11402# gnd 2.33fF
C1753 a_59478_8193# gnd 4.90fF
C1754 a_60542_11405# gnd 3.27fF
C1755 a_55310_10594# gnd 3.33fF
C1756 a_56358_11269# gnd 3.65fF
C1757 a_65446_11356# gnd 2.27fF
C1758 a_54481_10957# gnd 3.17fF
C1759 a_55310_11273# gnd 2.80fF
C1760 a_51328_10556# gnd 3.33fF
C1761 a_52372_11408# gnd 2.33fF
C1762 a_48770_8199# gnd 4.90fF
C1763 a_49834_11411# gnd 3.27fF
C1764 a_44602_10600# gnd 3.33fF
C1765 a_45650_11275# gnd 3.65fF
C1766 a_54481_11352# gnd 2.27fF
C1767 a_43773_10963# gnd 3.17fF
C1768 a_44602_11279# gnd 2.80fF
C1769 a_40577_10548# gnd 3.33fF
C1770 a_41621_11400# gnd 2.33fF
C1771 a_38019_8191# gnd 4.90fF
C1772 a_39083_11403# gnd 3.27fF
C1773 a_33851_10592# gnd 3.33fF
C1774 a_34899_11267# gnd 3.65fF
C1775 a_43773_11358# gnd 2.27fF
C1776 a_33022_10955# gnd 3.17fF
C1777 a_33851_11271# gnd 2.80fF
C1778 a_29869_10554# gnd 3.33fF
C1779 a_30913_11406# gnd 2.33fF
C1780 a_27311_8197# gnd 4.90fF
C1781 a_28375_11409# gnd 3.27fF
C1782 a_23143_10598# gnd 3.33fF
C1783 a_24191_11273# gnd 3.65fF
C1784 a_33022_11350# gnd 2.27fF
C1785 a_22314_10961# gnd 3.17fF
C1786 a_23143_11277# gnd 2.80fF
C1787 a_18904_10550# gnd 3.33fF
C1788 a_19948_11402# gnd 2.33fF
C1789 a_16346_8193# gnd 4.90fF
C1790 a_17410_11405# gnd 3.27fF
C1791 a_12178_10594# gnd 3.33fF
C1792 a_13226_11269# gnd 3.65fF
C1793 a_22314_11356# gnd 2.27fF
C1794 a_11349_10957# gnd 3.17fF
C1795 a_12178_11273# gnd 2.80fF
C1796 a_8196_10556# gnd 3.33fF
C1797 a_9240_11408# gnd 2.33fF
C1798 a_5638_8199# gnd 4.90fF
C1799 a_6702_11411# gnd 3.27fF
C1800 a_1470_10600# gnd 3.33fF
C1801 a_2518_11275# gnd 3.65fF
C1802 a_11349_11352# gnd 2.27fF
C1803 a_641_10963# gnd 3.17fF
C1804 a_1470_11279# gnd 2.80fF
C1805 a_641_11358# gnd 2.27fF
C1806 a_84757_11223# gnd 3.52fF
C1807 a_74049_11229# gnd 3.52fF
C1808 a_63084_11225# gnd 3.52fF
C1809 a_52376_11231# gnd 3.52fF
C1810 a_41625_11223# gnd 3.52fF
C1811 a_30917_11229# gnd 3.52fF
C1812 a_84752_12241# gnd 2.27fF
C1813 a_83704_12245# gnd 2.80fF
C1814 a_79421_12109# gnd 3.19fF
C1815 a_79520_12109# gnd 7.02fF
C1816 a_76154_11606# gnd 3.52fF
C1817 a_74044_12247# gnd 2.27fF
C1818 a_72996_12251# gnd 2.80fF
C1819 a_68713_12115# gnd 3.19fF
C1820 a_68812_12115# gnd 7.02fF
C1821 a_19952_11225# gnd 3.52fF
C1822 a_9244_11231# gnd 3.52fF
C1823 a_76153_12220# gnd 2.33fF
C1824 a_65446_11612# gnd 3.52fF
C1825 a_63079_12243# gnd 2.27fF
C1826 a_62031_12247# gnd 2.80fF
C1827 a_57748_12111# gnd 3.19fF
C1828 a_57847_12111# gnd 7.02fF
C1829 a_65445_12226# gnd 2.33fF
C1830 a_54481_11608# gnd 3.52fF
C1831 a_52371_12249# gnd 2.27fF
C1832 a_51323_12253# gnd 2.80fF
C1833 a_47040_12117# gnd 3.19fF
C1834 a_47139_12117# gnd 7.02fF
C1835 a_54480_12222# gnd 2.33fF
C1836 a_43773_11614# gnd 3.52fF
C1837 a_41620_12241# gnd 2.27fF
C1838 a_40572_12245# gnd 2.80fF
C1839 a_36289_12109# gnd 3.19fF
C1840 a_36388_12109# gnd 7.02fF
C1841 a_33022_11606# gnd 3.52fF
C1842 a_30912_12247# gnd 2.27fF
C1843 a_29864_12251# gnd 2.80fF
C1844 a_25581_12115# gnd 3.19fF
C1845 a_25680_12115# gnd 7.02fF
C1846 a_43772_12228# gnd 2.33fF
C1847 a_33021_12220# gnd 2.33fF
C1848 a_22314_11612# gnd 3.52fF
C1849 a_19947_12243# gnd 2.27fF
C1850 a_18899_12247# gnd 2.80fF
C1851 a_14616_12111# gnd 3.19fF
C1852 a_14715_12111# gnd 7.02fF
C1853 a_22313_12226# gnd 2.33fF
C1854 a_11349_11608# gnd 3.52fF
C1855 a_9239_12249# gnd 2.27fF
C1856 a_8191_12253# gnd 2.80fF
C1857 a_3908_12117# gnd 3.19fF
C1858 a_4007_12117# gnd 7.02fF
C1859 a_11348_12222# gnd 2.33fF
C1860 d3 gnd 856.70fF
C1861 a_641_11614# gnd 3.52fF
C1862 a_640_12228# gnd 2.33fF
C1863 a_84756_12064# gnd 3.17fF
C1864 a_74048_12070# gnd 3.17fF
C1865 a_63083_12066# gnd 3.17fF
C1866 a_52375_12072# gnd 3.17fF
C1867 a_41624_12064# gnd 3.17fF
C1868 a_30916_12070# gnd 3.17fF
C1869 a_83708_12068# gnd 3.33fF
C1870 a_84752_12920# gnd 2.33fF
C1871 a_82219_11226# gnd 3.19fF
C1872 a_82257_12925# gnd 3.73fF
C1873 a_76982_12112# gnd 3.33fF
C1874 a_19951_12066# gnd 3.17fF
C1875 a_9243_12072# gnd 3.17fF
C1876 a_76153_12475# gnd 3.17fF
C1877 a_76982_12791# gnd 2.80fF
C1878 a_73000_12074# gnd 3.33fF
C1879 a_74044_12926# gnd 2.33fF
C1880 a_71511_11232# gnd 3.19fF
C1881 a_71549_12931# gnd 3.73fF
C1882 a_66274_12118# gnd 3.33fF
C1883 a_76153_12870# gnd 2.27fF
C1884 a_65445_12481# gnd 3.17fF
C1885 a_66274_12797# gnd 2.80fF
C1886 a_62035_12070# gnd 3.33fF
C1887 a_63079_12922# gnd 2.33fF
C1888 a_60546_11228# gnd 3.19fF
C1889 a_60584_12927# gnd 3.73fF
C1890 a_55309_12114# gnd 3.33fF
C1891 a_65445_12876# gnd 2.27fF
C1892 a_54480_12477# gnd 3.17fF
C1893 a_55309_12793# gnd 2.80fF
C1894 a_51327_12076# gnd 3.33fF
C1895 a_52371_12928# gnd 2.33fF
C1896 a_49838_11234# gnd 3.19fF
C1897 a_49876_12933# gnd 3.73fF
C1898 a_44601_12120# gnd 3.33fF
C1899 a_54480_12872# gnd 2.27fF
C1900 a_43772_12483# gnd 3.17fF
C1901 a_44601_12799# gnd 2.80fF
C1902 a_40576_12068# gnd 3.33fF
C1903 a_41620_12920# gnd 2.33fF
C1904 a_39087_11226# gnd 3.19fF
C1905 a_39125_12925# gnd 3.73fF
C1906 a_33850_12112# gnd 3.33fF
C1907 a_43772_12878# gnd 2.27fF
C1908 a_33021_12475# gnd 3.17fF
C1909 a_33850_12791# gnd 2.80fF
C1910 a_29868_12074# gnd 3.33fF
C1911 a_30912_12926# gnd 2.33fF
C1912 a_28379_11232# gnd 3.19fF
C1913 a_28417_12931# gnd 3.73fF
C1914 a_23142_12118# gnd 3.33fF
C1915 a_33021_12870# gnd 2.27fF
C1916 a_22313_12481# gnd 3.17fF
C1917 a_23142_12797# gnd 2.80fF
C1918 a_18903_12070# gnd 3.33fF
C1919 a_19947_12922# gnd 2.33fF
C1920 a_17414_11228# gnd 3.19fF
C1921 a_17452_12927# gnd 3.73fF
C1922 a_12177_12114# gnd 3.33fF
C1923 a_22313_12876# gnd 2.27fF
C1924 a_11348_12477# gnd 3.17fF
C1925 a_12177_12793# gnd 2.80fF
C1926 a_8195_12076# gnd 3.33fF
C1927 a_9239_12928# gnd 2.33fF
C1928 a_6706_11234# gnd 3.19fF
C1929 a_6744_12933# gnd 3.73fF
C1930 a_1469_12120# gnd 3.33fF
C1931 a_11348_12872# gnd 2.27fF
C1932 a_640_12483# gnd 3.17fF
C1933 a_1469_12799# gnd 2.80fF
C1934 a_640_12878# gnd 2.27fF
C1935 a_84756_12743# gnd 3.43fF
C1936 a_74048_12749# gnd 3.43fF
C1937 a_63083_12745# gnd 3.43fF
C1938 a_52375_12751# gnd 3.43fF
C1939 a_41624_12743# gnd 3.43fF
C1940 a_30916_12749# gnd 3.43fF
C1941 a_84752_13688# gnd 2.27fF
C1942 a_82261_12748# gnd 3.35fF
C1943 a_83704_13692# gnd 2.80fF
C1944 a_78030_12787# gnd 3.43fF
C1945 a_79426_12228# gnd 3.27fF
C1946 a_76153_13126# gnd 3.43fF
C1947 a_74044_13694# gnd 2.27fF
C1948 a_71553_12754# gnd 3.35fF
C1949 a_72996_13698# gnd 2.80fF
C1950 a_67322_12793# gnd 3.43fF
C1951 a_68718_12234# gnd 3.27fF
C1952 a_19951_12745# gnd 3.43fF
C1953 a_9243_12751# gnd 3.43fF
C1954 a_76153_13667# gnd 2.33fF
C1955 a_65445_13132# gnd 3.43fF
C1956 a_63079_13690# gnd 2.27fF
C1957 a_60588_12750# gnd 3.35fF
C1958 a_62031_13694# gnd 2.80fF
C1959 a_56357_12789# gnd 3.43fF
C1960 a_57753_12230# gnd 3.27fF
C1961 a_65445_13673# gnd 2.33fF
C1962 a_54480_13128# gnd 3.43fF
C1963 a_52371_13696# gnd 2.27fF
C1964 a_49880_12756# gnd 3.35fF
C1965 a_51323_13700# gnd 2.80fF
C1966 a_45649_12795# gnd 3.43fF
C1967 a_47045_12236# gnd 3.27fF
C1968 a_54480_13669# gnd 2.33fF
C1969 a_43772_13134# gnd 3.43fF
C1970 a_41620_13688# gnd 2.27fF
C1971 a_39129_12748# gnd 3.35fF
C1972 a_40572_13692# gnd 2.80fF
C1973 a_34898_12787# gnd 3.43fF
C1974 a_36294_12228# gnd 3.27fF
C1975 a_33021_13126# gnd 3.43fF
C1976 a_30912_13694# gnd 2.27fF
C1977 a_28421_12754# gnd 3.35fF
C1978 a_29864_13698# gnd 2.80fF
C1979 a_24190_12793# gnd 3.43fF
C1980 a_25586_12234# gnd 3.27fF
C1981 a_43772_13675# gnd 2.33fF
C1982 a_33021_13667# gnd 2.33fF
C1983 a_22313_13132# gnd 3.43fF
C1984 a_19947_13690# gnd 2.27fF
C1985 a_17456_12750# gnd 3.35fF
C1986 a_18899_13694# gnd 2.80fF
C1987 a_13225_12789# gnd 3.43fF
C1988 a_14621_12230# gnd 3.27fF
C1989 a_22313_13673# gnd 2.33fF
C1990 a_11348_13128# gnd 3.43fF
C1991 a_9239_13696# gnd 2.27fF
C1992 a_6748_12756# gnd 3.35fF
C1993 a_8191_13700# gnd 2.80fF
C1994 a_2517_12795# gnd 3.43fF
C1995 a_3913_12236# gnd 3.27fF
C1996 a_11348_13669# gnd 2.33fF
C1997 d2 gnd 864.08fF
C1998 a_640_13134# gnd 3.43fF
C1999 a_640_13675# gnd 2.33fF
C2000 a_84756_13511# gnd 3.17fF
C2001 a_74048_13517# gnd 3.17fF
C2002 a_63083_13513# gnd 3.17fF
C2003 a_52375_13519# gnd 3.17fF
C2004 a_41624_13511# gnd 3.17fF
C2005 a_30916_13517# gnd 3.17fF
C2006 a_84756_14190# gnd 41.87fF
C2007 a_83708_13515# gnd 3.33fF
C2008 a_84752_14367# gnd 2.33fF
C2009 a_76982_13559# gnd 3.33fF
C2010 a_78030_14234# gnd 4.35fF
C2011 a_19951_13513# gnd 3.17fF
C2012 a_9243_13519# gnd 3.17fF
C2013 a_76153_13922# gnd 3.17fF
C2014 a_76982_14238# gnd 2.80fF
C2015 a_73000_13521# gnd 3.33fF
C2016 a_74044_14373# gnd 2.33fF
C2017 a_66274_13565# gnd 3.33fF
C2018 a_67322_14240# gnd 4.35fF
C2019 a_76153_14317# gnd 2.27fF
C2020 a_65445_13928# gnd 3.17fF
C2021 a_66274_14244# gnd 2.80fF
C2022 a_62035_13517# gnd 3.33fF
C2023 a_63079_14369# gnd 2.33fF
C2024 a_55309_13561# gnd 3.33fF
C2025 a_56357_14236# gnd 4.35fF
C2026 a_65445_14323# gnd 2.27fF
C2027 a_54480_13924# gnd 3.17fF
C2028 a_55309_14240# gnd 2.80fF
C2029 a_51327_13523# gnd 3.33fF
C2030 a_52371_14375# gnd 2.33fF
C2031 a_44601_13567# gnd 3.33fF
C2032 a_45649_14242# gnd 4.35fF
C2033 a_54480_14319# gnd 2.27fF
C2034 a_43772_13930# gnd 3.17fF
C2035 a_44601_14246# gnd 2.80fF
C2036 a_40576_13515# gnd 3.33fF
C2037 a_41620_14367# gnd 2.33fF
C2038 a_33850_13559# gnd 3.33fF
C2039 a_34898_14234# gnd 4.35fF
C2040 a_43772_14325# gnd 2.27fF
C2041 a_33021_13922# gnd 3.17fF
C2042 a_33850_14238# gnd 2.80fF
C2043 a_29868_13521# gnd 3.33fF
C2044 a_30912_14373# gnd 2.33fF
C2045 a_23142_13565# gnd 3.33fF
C2046 a_24190_14240# gnd 4.35fF
C2047 a_74048_14196# gnd 4.89fF
C2048 a_63083_14192# gnd 5.08fF
C2049 a_33021_14317# gnd 2.27fF
C2050 a_22313_13928# gnd 3.17fF
C2051 a_23142_14244# gnd 2.80fF
C2052 a_18903_13517# gnd 3.33fF
C2053 a_19947_14369# gnd 2.33fF
C2054 a_12177_13561# gnd 3.33fF
C2055 a_13225_14236# gnd 4.35fF
C2056 a_22313_14323# gnd 2.27fF
C2057 a_11348_13924# gnd 3.17fF
C2058 a_12177_14240# gnd 2.80fF
C2059 a_8195_13523# gnd 3.33fF
C2060 a_9239_14375# gnd 2.33fF
C2061 a_1469_13567# gnd 3.33fF
C2062 a_2517_14242# gnd 4.35fF
C2063 a_52375_14198# gnd 4.89fF
C2064 a_41624_14190# gnd 4.85fF
C2065 a_11348_14319# gnd 2.27fF
C2066 d1 gnd 1003.49fF
C2067 a_640_13930# gnd 3.17fF
C2068 a_1469_14246# gnd 2.80fF
C2069 d0 gnd 1239.36fF
C2070 a_640_14325# gnd 2.27fF
C2071 a_30916_14196# gnd 4.89fF
C2072 a_19951_14192# gnd 5.08fF
C2073 a_9243_14198# gnd 4.89fF
C2074 vdd gnd 5237.13fF
