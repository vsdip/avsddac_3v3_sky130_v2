* SPICE3 file created from switchfinal.ext - technology: sky130A

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_308_n101# a_95_n101# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 a_95_n101# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2 vrefl a_308_n101# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3 vrefh a_308_n101# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_95_n101# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5 vout a_95_n101# vrefh vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6 vout a_95_n101# vrefl gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7 a_308_n101# a_95_n101# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5

Vdd vdd 0 dc 1.8
Vin1 vrefh 0 dc 0.5
Vin2 vrefl 0 dc 0.2
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)

.tran 0.1ns 20ns
.control
run
plot V(vout) V(d0)
.endc
.end
